`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dHLKy/nz06UYVZQugnMYVzoizdQga5eiPviTNijLVrfka0e4n10maZroENH+i/d3D4nP+6rCehwJ
Pg9u9lMPEA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FU+YgOMEW7wHhcRbjPDmbCo7UM2CGV7VwVVl4gjrfWCjnM9rBXIcGtwrCocUfVrUK5yAzNllJcbk
RkDirhqVsH3Dq1TEQbXSZIdRul0B5/DsmxVfyk6xwHMQT4GRVIhAj9IY2BPlyuQe+uiGABvn7SO9
708Iw6IfcBM3Akln2XQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sCyiVB27tH4McbS42COLF49X2klsN9rEOOt6PRuLABV0U4bnrzrPA7cgvCNRl5ervASr1Eq8O0E/
6sNkTJ0CNnexp9PRJnvCTuVEqf5rDmOexlkysQSuvCf5I9IjBWrob+rfkQE29AHt4/iWieHDAA03
fAnUI5CoEWnbH6V5/BSBkNIB/STwgBz+UXKuJnqAumwRextGnYVz1D3Vlf7gpOMaqMaG+OYUB6Db
3wK0S+kLVMhec5dwYm6dh9Xy3uETRUEPZrin0TkQKRx1pvXxIoNFQSWapro5z2PdU5ClAC3zisqb
DjX9vdb2ILrhSNByhRV2/IS9z0/lugc/VHH74Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qwVz9qepk3J1bxUCOZC+3ZtoY3qbZiPW1Bkyyou6j0YnDBiKN5Jk/5EfBzmR7Dqzep408KKnGwkg
I8IQZRaFJRbCPYH/CX3nnRBLW9hg22xZDUESYSDyQPNfnaGdXEa/c/+VYUWHtwEjEQsjZtsNsAsa
iQzYiQoN87u2pFro4tg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J3IBWs5TG54OVxD3K6WpxUqKy5qvpCmAWVBYJUQLz+wM82DQcBxD0CAagvYWxWUkhwpAUzKKi1wO
YUxr4jRVrxo1FtXZLUP1SjdxSbP9maRFzxJ3+/buydDsNIEHOXkAuAgCrNwv+PUWW+ZIH0FWxxIy
oRAA6/AdlpE78/juksgpt/1tbxMQ/1EUHnlEY2bst/hSr+kuuOzrc/qBqnFFNlg/OTPvxFy6jd9h
MBQXulj2wJ82hPCq7ScKTJibNl1EcNHRZZptGiphEEhpcBsvQyOTNq6x5zpcFGceUXkKqiB5Rti7
2UdBYt7dyuUuPqp60TVu2mLCEdQKcryOh0M1JA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 452528)
`protect data_block
azQoGUAH6Y4js7lGt5Q8UjSNz7BAz26CH6rxZX8MRNP0xNrQm02HLZOq6C0WiXDmKrCZQZ3B1zrz
jLndjCYkYJuD7TOjFux5fq5YD2dU6hF8SF9NsL9op7xNJj3mghCNw0d8++aT4VQa/CvnE4IEI0Nm
bTNq55sp9OiZYtNOEB3N9F2A3XT+vUQnBW3wVkHLF+TIasSeIZs3XYsKzRYNJEb3f2dum7/TXFBh
GFvYvm+2AwT3xOsHVrRVQhI8PHBT/hqANOkWzvR/E32epQgVbA5gKtQwTassEG6cntrkqGYU1peO
MPQ7DN0qNnQNgOxDicDEiuXVDVkGQuJGDrEE6uiNlkLglYibcLnEIlPHLq3NbIAVjhiYxMYiEV9e
newTOilzj7aOAeuYt9WkWo12XvVr0umUrpo6QOLn+Y9CmKAPWwlO+LzPBK1k64Jnv1FS6hlHKGAx
Yx+rRB6oZ6iCe0vE9egtL7AR8FUquBEgj2Lb0MMHK3x/R1AYsYPbUyqwO8xA7YvMToLb1Y8OaXQl
khpzYCuQB7bordRzDCQLbwIVCjz3X+DoHuLe0g6k+A63AC7GpU8rjOS9EEDkFqQNVtaEmBoIL87J
S3+IMjdtD8YPtEUldRHRe1r90y+r2T4dOrOcVryC3h7bMXvcn8ixWoCLoNd8athbMLgMPrEdhiaY
uS+fLA2fs8j7/1wtnasn+j5VMfJXB28/c00n5lO6uMNfCyq4mht9DZEHxH9Ha7g67itMagZYGy1w
V1tQt47mKTy2fFnMtU0sptlkPot39QrSnA/DJqVRl01Bzep4yq4Oouc+1fGBqTOWZWMOH0O0Kmfx
n9klPkk9kRmB0MpuD8siC7DbPXOqKZTT4kfLNFRPThzdpWwuuS89ffK4MsddxdELTdGGoeilGh96
GsWJyGfEy9puCGEvoG2wjCRzmgxbCaSx99qWq4M7gn2iFOpEFv7x+Jwx/tK7X7IWaB2cMv5e/GSp
9jb+AxfO4uG77UEuIG0FK4o3Z99keW1QCmRGXTjdP++1MxO/FO5oZKIfb44yT5lQ6C2XR/jpd17M
mHf0VRkbJiLjrVytZ3aAZdBGJQwBELbILX3kZzegl9xIBnr7K1ATPpdWfr+b92x4HaXNAz1jWFeR
E6gCCtxfigCjyBnFSWsgk+ql5ZB5v7+TNf0mZORAtahg88SCVZZcVt3hKOXrnt2dxtj8Nqnqd4IV
hWcRRN4ccZfiH4y3G7i/4MXvWJpxRusqfqmyJtmwPYxbWHRY+4tI/L5bRhB1VHqtrAONUQZr/jFh
qW9HtlSA0vbKde5hzgXd/2Uz0TW+epdk3xrjc4VZDXuOQxHQT6ETAocAAiGlY22TSMWKi06ERhet
41pBmyknBlCLgJYWPbRPrjs0gZOnso9gbfl7XT+zEK+FHU32xFJKovDz/JihV7a+6FWWBcCA9gpT
QmaS+XKhF31hdsDpyR8G/wPrjCnfngFCLZH3dAtJZMxZZmIet2g1Nu6no5bNKgioBwSZ8Qz4YaXI
AJtZPD7tOP+Wz/OwsYh8C7FIBCKG7dCvZSqU8t5w+Q/8lHDh159+Adxi5/w7Ovjn19X3X4jijIuN
ksT4zPDxevjkfoS4biTHhpNnseG2+alPuZEV+kOmEP26I6FuVRY0wcSyDE4NUKNc6eJsfMEDHXqP
79WEvaC7k51HvTQ0xgSCiXrjTb9Gd6yVw/qtlrz9H+tS+RONuwSUVEy4S/LGOy/sXCaJzjy9tV+M
AyLcvpGPx3dR1toExx7y5tGvgnvJdv7aJ4sm5VjR/B9TNGPSBEksp85T5zIQ3vT0A4Kh978g14pw
SchxBZHskFP5tlPPZMqafvraEvixr2urN0vZwYBVurAR62L8AnubkOL2LOjyFcTsoIxNTP6NWWnT
p8k07k11IrGk49kqq4wet8WabkltbarqTf2E9RlQU0Ep4Nq63VHdlA/G310HioClmfmH3H/SuDnG
AdX16jxvBEmljZsKx1ZcKhBYaHTjlEAEpNzJu3KypdKljbS5hnCGxToSddZfE/HHrm7Hlm5NLdhT
XZfEPu+bXUAqyXyZ3L/i3UJfwsJdrcO2V3Y8SjRmxXrPuPkPuOhRZilwVkna/z+nQdSbB47LkVbs
QxgCj5ogZwNKhv7VvXm4vjqyNdwxaQFgdL1mwNe6DoCpQQoDgDl/z9lAHZzIfXFXND5hPJ9pcY9s
ZvMXF3lvUJRUOuBB4D92uvyeTnq8zLkiPAplahaTIdT/m64XNjVs9AIbBMY57Jzvk7f40+V0fTqb
WkldeSimND9JhYDHliYipaPikJdM1+SNHTlbcfVXs+o+MuwJcFNClE/u21xGXo94vnhJBlE4YZPp
f2xlOcRnaQT8WMRB54c2ovg/eDj/Hcw2GiVMCHQRKeE6p/M5Y7glYVXrJ5bol9QhtiTCZtP0Rvpm
omnl1CfI1m3ZVa0FatqZA22F+jRYaoCM6MFN5Of3nl1735oNW51JR5GwVjh5RopiZGhtu09nr7PB
iIDBfS91bNDtPyFeIl/l0Mp0Ieo4Dis9hl459D6XmBp8wM6J3Y+h4PZwCmBCQ0pYNxaJyka1UeES
oPt0M0+gQeo6LriQWyREB42jlRCarIrjZ4heWm7ITJuelyVmFRkePrCaAx6+8fVmUkWk0QSdUOZc
rObqWafAXeYUXR2v2Q6803x4RPYEtN2XEWiWqwV54xWRSfPpBsDjk6poyAcAgaORiSv9JzSdpcig
H7AhEZf0Ud3v2w5QZ2oJhDBmkOz54zCRIRUth+PnrBHQHOhGc3RtvgFUwHl4MrO1az685pSBurm4
RQj3FEmB3iH34M5TrCd0KOl3y2wYfk+VbxVpQtLFbFT/cOISP/eUtoqZmGsuGI0QSXb8gVwdTZ2l
l/3oaT821TyHiod2Z/BofR0BSjrMsFujoR61/243QCWNPynLYASqOyhB7KuuXnWK3zL4AAGLXhIE
mXCAsLKAw6zFjJssUnq5PK6h+3tC7YrZangiNDYy0GCfEokk0jl19+EMmyhZk3IX6dj0Ruq+VwZ0
egxBvULsTTlXmm0rnllxqIiMm9gu2IHrPPJd2/Yavlse6zz6hsvBqighMWTpTt9RuUx08AqgckWe
msP+p/XmNaAvnGk5VKI6KWnQFKJwH5Rr0xsTH2LWK4odsR1dBynw10nrV23iIe3sDAuXPWQCvzDT
tH2niSSwP7yppf3gJW+9yMwm3Hc6tyeE5j6lydPOhcOrCMo3ckHsHZOnsi+hMaoysdbOlRabC60X
7OcOGIxd+p5H4VzweA8tR+xMm4XGyOYmY4tgw5V2Vg7ibgeACq8eCZ/MBo3t22jGdIPDl83LI3nA
jiRcseGo6LUcbr44v1LpndEhEepLbh5Fs+XKsDahNsaWy8OELTEiZlL70Amb0xahhMWxFo5wPrJP
E98O5h60je7k/0yK+SovhgF+quhzjx3uyABdhGfahJ+or/9GpbwLEIW74ykFrpnmVQKI2U1IpGz6
AeHQFw228GZPpYNnTYeolcO3a6lqGy+HJh0Hu5EAf41KOk0FAQgt4Nhzk/Z+kg1gu4fsaijmEFTS
uARW8xTmBYBnSNJ2TP03dBTf21TlyiwabtRTXHkjGNJNIQp7SyH8+cOA/+aMRm/avzrNASBojrQ6
f+TmtzUB06sVKLNfPdZvELbCWp9KZI0d7aOPqhzhCu1s+L9H7W1lSKCmOUgBpHuDNM0gQEg05ILR
fDZ3K896YukJWThfUHhdK42mkAVMbJEjlsqRwJ+t0BXJUDS83rA734ylq8amoUFHcy9LFvbcKN1/
palkgN3OcTH8AaW4/pWFB4Q+1Y7sVJSaQikWjnuEXMUYru6nsdNMB5fJpX3yEOzmgjjDl7yjpT5j
ahibeGt+5j8jdyXtGyYak4XiiGLfPBusHY30MSP6J2eGXQWPTz9/Ibqw97YietIJ8djxTR7Zh0Fy
lVxaLwN6tOvO13uajpM8vPYHC0dd1yiyLzwcMuvo8pFCS9VN+6PEAlxSPE4ovWSFfGKXCWHwQZl2
FlzhBkIKPQOom9Ujvv92+6Dzzan5wnzlIUZiWDlj2MNXsVscNOnKiFN/hcGWCAwkK7Jfc4++Ifon
5+hwxjtJNPS6sDwNPIag2oFmS70gjfRGthkOF1KpvOh7U+kb0uSAbUwp/34CKKCE/RIr13PQtu2Z
/O56kWaaw3AuIs1uPZ+PREOBIJ999GQXEAjhOJF2nEp6K/rvGrpr9F8cspSvuW0j58dltlgQ0quI
o0m5hN+tLGP+TeP1VwE58ZfM2SkbqGtsmvZQuPozYXtnjCiJsWVb2q9dIe88WC/X9t3aHcJlLyrE
9+6YdJOUwbHIY5Q+SysHwXL6z9EOa2hKd6nFnVcTMpjFh2jIls5bUKs1grR/VioB25o+twwbymZd
YHVDdqs+MqO/fjEH1wBVr/7jMkil15o6vVs4UoEc/CobY8qklI36tHAt3DZcbALKcyGp8eOrQTRt
b9TxS3cbIgLGIVZDzCZfoxObaa/FWGtcsozSwgz0xjkmzCWsNhJAK0pleXpjlhQD55VIp0sbTmw2
AR6t2cOSjnhf9SaA81g3CieZwZWB9cNU2tUcHSMTCBQlxVY0QqbzDZf6GLc8W4l3PuRPkRigsBIG
nGVBTUpXLKxxK77eXm2h50yis/XCaYOiL1PHPgtdqYgJX5aSXOsoGiS8BmDgOfkzd5r0xZmjdxCF
q5MQlISbYM/ppIWOFjo8VicX4KLI5IJRL7ZMWZgfigH9YI8b2afp3zI27b7mrbm1JUvDYYRaEyrw
fSTcB8hGpoRQ3oEHj3F5EyhwzqZ7KKkJKKQ43gLy43YYb5025K2gjQhmeMOdKI2R3e6CLG5v0UDj
f3UPtAabE+oJmFfauhmq6y4ccRtZJXDsWSrL/A+Wb3AUR/8Us/N5rzoE+8R0EK/S4Fy9djFabFa6
2Em8uyIXIpaXKrHBRfsq4Bbyy5zKqie7XYB6A28TyKf1rAyqrsF82N4xOter+HkSY+RaQwvFrE1t
q9E2f1Ys3LWzyeP3F6EJVJqy27QWuuOt3xVrKi4SkAgOGCPMTIKW4tUt1SLSE9Ky4OqYmH9IZeLt
5lELL23rAj8YIV2gvddCF3WfGbMrF197i9qyjGdHnUSJCIJEOLb9/ToLK30S6CwLj7MH4huwv8wB
ztN21+rb1Y8dwcUokf27G8KkLu3wry5BVmiHbtPIL/GfCKuGOpV+fOIWl5My9hZM0Ra4vi8LqXGJ
6ja0sWTSYAjpyPi+wp65Tq1N5AWCeSDYUuj9pABvnTIsGkpNVJc73ypw0jy1qV85FWk7zOTkoPLB
9pv7B9anCGulmP8CBVQF2UNmxYXTDtqd3AKnmJ47/S84vCuEvXL1ovywIvIoOKQG3f02hV7p+Aip
U4yc6NZROTnVKvjJU695fSh8tP/Y1Zdb5Z7uA5XKz8bfh4nNlz3ZbiA2Xh3qR6j7mTdNAUJJdnx9
jA2YSjzE288mNSGMS517zC+Uoj8B5k4XHHj9rJv85ov9plg8xaPYCjImMnzRfoJCYM0djCwzI7yn
FTxqCSmE0uRvJN1CN4sLAQAbYAJNPCA23covEOFUwdhkyKElrmAI7saznYIJhcF0HldB9ILCJbHC
ms7wm+unvpBfU+CTVGIGaY6f7nc2nOxE4kKsW3jxgtdyBpeTJpusrtf5z/JWTuovb9Kjn8Y4Y6C6
jT2uZKFEHedJDoISFIjB2K14NUeB+/boEARpRX0jnEfomn19ZmoOpMB6bUm/bot3TK2tD6tXK351
O+lDpvxiz33e4CmzU0jXWPJd6Gaxbupn50N+YYxIIfGVQuoJZi/ArBU87KzDlQsLYSpGML88hqBe
dwqcTY0hyU9t5BCt1/QZQnT1U6eTRmqhjaxflfZjLNbYCV9Qx5pwLD3DInraKjsIy9QPl0nRgXxL
i9yP8pObOWL4D/kJE08OrZLeaEOXuvDkIFdYUntqZUdCV2hB/CeRXP5ev7U3qlWo+nJcwYDKU1yA
SO+7rJF6RxF5qp2V8kFMazS67kL3xppdaXZBcXXCTnBrTWKi02BiM8ryU69paQI0ZpCXh/usioN+
9QUuuuZfNQA5E4jNe5pTCykW4Xt/hF0DOIOx/MAnbU1LOdjX/Ah/r1MBdUKUHP2YdV1/2SO/1OPg
6wMdcjUNu45xzSPu6H4uHmt4bTshD+cezfBZI4Kufn8eSy36Ho11Vg2ZiknI/SeO46dsZIvgz20v
os/JvVyDxksVFxPIU6hEl0LSRE17nRUpjDQlywAnH0woEB+hukEF3zzkvkvc1nTzaEsmzSCfCYWs
h5vCCMpYdOw5OcspNKpOa2SVT+82YmlPFK9Y6GuXpnfNnRUFM+TgDVADpTLcdL4/oD28L3viWTar
stoeamuEmcTOblNUxUF46evvJSm39t00VFXdYwTEdk5ikgtFARIVbWO3AYTMOSKGzO4rIObNTaDv
ZHvpSYC/yu4ehffUIcSWnjkYKr/rtPnE5xC0gyRfHxiogF3ceXyco/AkL02oE7DcXCEW6H2SE2pi
9sSDma7J09PkcIcwGHoZVbEQq5GK9Tji28qmxlhmr8ean+8WYC8OZuobV1qMyKYh8mHnXUK2+yHx
Y14KYcMisSZ9H8ze/+88kwlrQvpMs3no4DBu/aMAL0SB5RWcNG/FlFCEbRyZigTk97+n7GFt2Qog
Uvg5v+znSvU280Ez3tGw+UlmJRJBEHd+hBlbqpSq32csOI/tLPFqXNS4uQNH4FchUwYbavYxIdNK
+UN0L5lKkkSaTxpCKmS0xtbi3bkZtEwpj7R0oAwWxMDrJPh4odcLOdfK7k7fFFW6wlNSW5gdhgvP
w6NAMZXLqKtYO6Bo7J82YkwZaRoDO5OeF7g79Krj3bHNjViClXQozZ6U/5QmXmS2aBzrk8w507j+
c6WEu7a9T53Ggd04iih8iugGUGI9oXeD0rhGamvnBHoTVbHflKFgm6cY54AyCdm3sA1wmXa4LeO9
Nk8Cymn0+saBIgDySGius1Sg9JQzXz84Ofvb7QC9NKpA4HI4wX0eyOIC2EQonnrQQt78YQNBlK4b
acOIWzl7tilZxiApFVQX+SRi/yoxUAYrEx9QLpT0M2MOsN9hRkMmnDAO/8G8vjXCpqLNwxpX/oc3
x+N+i0e/d5Qs2k1kBE1ygLMu8q9OzzMOuUN95x8X2ngV2gszkoebBZWTFj+oAbV/OAmz0BqRdrvi
6JIVwqkY5dnFdr5paehWieEsqFZQlMva80q8MEfljNCUs7+NsY1GGjzetPq1Z27Djql9fvx1bDKW
leE/VKWECjNUNGwYvEIQ5Ee6jF4xKs7mW52/c61b6mspBH/tZtmXMlWElaoRK9d10yaWXko8t4US
beiLwchhKLBurEbpldgAlfgk+LU2Umbrczfpz+Isdgkbs2USXX7f6w4UQzVMqmIAPteQId/x/C7F
QAYXRNCBeNn/toicrSDSKPfsYMHHxG4mpXQ+DXQFVmvwOLT+k+cAWTWOMNXNugIRrizPryeJUvNw
cwknKUskSwDKb6RRhJuq6MAXh0aAhVd7i15SRHAS4jJRggdGsHq2hCHVOL6Zd2MUkSfzr9JMmwQE
BP3OmVFku4eldVcxdCpacHLCE0P1SnKNer5HxF2H8qeaYycKaDcVtgaB4aZbDYw1QHPaLzYN+M2Y
hJMEQ6zcsaj2kMqjhuUAB2cHdFTAEZ1Z+TVoLi9FRvVLYGGsqxm8ZKtVOpJaW1d+gs7w26nRxUjl
9PtC0/e2qKj6KDPr9oMb3zQQqBTfhED83RhwiWK/5atxUs75I7xCWHwITHsPjGpqcytYuO7JFfOZ
M4SBHhRVqKc3FS9E5fFrazRVTdWA2x43LKcI1NS/VKbO5+V1IZdwxwjEe29aGCOaa/G7fTbP8zfc
g5O0YlD7DUBCAkka55t7qpm7X2pKIAQ6pkAK1DQK9m+OaEx8x+5dxmwp5MGWSIIkE8RXp5SFDVM+
tO231WaGkPmKjsLgQCLO8mJCqtXWrh/tL3UcKW87eI1GLQt3ArHOlGOzn5eKMRR6pyDVGakywORP
wn9KKqWlMRhmB6mB1SAz9wSkhDqjss8vxAU7c03Izl+dvfalN0eOJMRdj1l9iafosy8ahlEiUSgC
meRYAlunMZE/SBp47f7IZPu089+PBjyUjkEWElulx5JAkgGQyzNOhHy1v3H8aVAdEVgLVCDfOdEk
uSQJ9piaG+TDab2y2QLgC2HAePV28WvpoB25u8j5dCSnMlPETsL6xjzc8ljr9l4my2w7cz1Jdcxd
3HWT+W8m7V7aKPDS2olOc5h7WOC/gma/7jGcS4xRwQ1TfU7eIQUYsW1+pzet74u+0QrH2VBmpRVE
JQZ4kv3qG5r1ZnJGyGUmL5LnTU1I0RF5/pxNiPmbXdjpfefkMSBcLxmP3bJtI3bjCObmUrAk6PRo
hmGiaNOPsv+iOmpNW2LkBFprQ6tFsEKT/VZnB2ljtvOvnQzH0YcGlllDm2RVGQHjaekGG/4B6LTd
LTptDYE2HK9TguVc09oIWy+tU+ENloek6YeFtusD75TkU3td5uruwjaw+Ym0uRcB/a6464/jGE+p
qwfpXM0sZcyMOkMGNlwWYm9IZXWc9bUthvwPTT0ElkQ+25OpQWTbidCzBUS5vnrXrJ30c6YOc40A
I4PHJFvXGN3zkUJ/KZw0skHruN6091EgfplTBoedXhAcNrRZ2zxOboOoSUvzZ4Dz11JXJfMAamLA
bFOVDNeVpNtwZsxaj0Au8vd7ABfPp3dLwU09GbbfwaeldAd6VSYN30WNRA2gPdxAaaFMs0kMWvNU
y+6+r1ZlCSfM40bNAmJ+SyYqGJxjumXjPZycZgLEJkEWkIQOONh5LkIm5Oo9m5ODGtNGYr62sbNj
i/z0Or4BMUC6yg9d3rQFEr+4yqXeXcRH8TiO2o/zXT503lG76FwNmzmJY1BRqbXHjKgkUm8rgzl0
yH1gN04JEC0Cr34i3WQuCCDJwluAPRyCoKYsI2sKAXtpJ8knLiWhn5piV9USwTNwjzDB3q4hPxUC
hZxmmed7NNlon/FvwJg5spiGH/NovjCv5WeuTHtyRJ9Sa+VH7OIF/TvQocHkEzhPTgMfmpKu8I7N
x6h/wFPvzUvKBA4X15D0qHR2pTkRHI7kNm1aBOVz+/IAATYfMBSKXlaCx//fHaNfv4CBFlTm3Ve0
N6uUBb0aTH4kC+48cQOltVv67n6Mvz6xdHM/hjUW9gLgeVz3HsA/uYt1x3nSpFoxH+mkUt+14L8P
AkiyAIoFmtoOiYrgEkKg6SERN170h/F8UwXagZucPX3BB6O6JacE3p8VjrSeEYsuafPzftX42H4d
PtFCWuQI5b5HKmMbFOqLfhwYYbhv5v8U1h8KNKZdKgn21zJ3YGm70+C78nEJu9eaMs2QRSUukviT
HofrjqcsJHpIdWVhiZLD5UYSWKpSZM7E3rG6MBbIJf79dgrJoCcslKGDTWSXdfhegvySpYx0FGHO
oS7eI0QFMpPpDlCenIfg8Ta2lM7k8X0r+K5CObEoDnm5EdecHpjht13P5DfvkS7+dc1ghD6VuLUp
ocRnKnwe/cUJ6qoAwlCfH64iNd71g7y89TV+ZYMRSEwt1twbECKem+VoLhWmtv/E1q0IMuYFHOWJ
5jTGdtlzxZMlNAx1LEqGOQJOunk76UjyDMq2WDplsBrMFd4YLJ0m/ziJS4JpTafVUMj3JfXgoSee
EaT2j7NQwVlY/7nbbH6z3XHXwhbyzBxdhZ2BNOjn/JGMoCbm4qUMEoSoF+2X8MtbU7H8LSU1vWoW
+k1bqVK4FSnbBOjMaaa1nnMbZRlVkuMMyUFXSaubszHCjg55AaAWuXYW+rlgejTJ/5yxa/QTCUpP
mKO6BNlioVmTfSM1c39uc5iVHkVL55RmLPz0BN+lqNqHVtVucxB+E5mIQECnE/mCTh24Xzwg1r2R
h9J2J37F5zKbNpMyYkJHDDy3soSSi/PcL1gtvo2ZUJJSiUYxpV7qAMlh7I7dhltsqAo2LXqovaUU
tyiHNxnacKTmCDn7wdkrVHoTjja2U1KaITV38n77A9UJHTROpkuVSscLdsjAJ0D6zl+8NPnGWi0u
vJiwvJqxcy6eQEo/2N1HHpFBFyu3MsyMIn12SNG+ngMF/kAvqAi4La+KdmhoBnA8YpGt2pJ6yT38
q6lJOOKwKbaB5EH8YT6jzyI8a0Acb1p8zmU/aCV3WbzDsS981k1Kx0CrqF47Ki4QJifCtg/KMx+3
3fv8oMRgeKke4QSEZbKLdUmOUR3UJamG65oFUgoV3DRx+EBKNcWk9eUe1qDgPeF+cYWvECUTCAhr
Dj08Grms9yuV2w+ABbiMRqK9tcueSQhmPmn6FbOmBStlTXyEPw8zxkgEDwC/9nDf0dt07DTxcxu+
IPXiF2pq+u/LMZT06XtQq/n8CupZiO9hS+t7FH7qIr2AzhNY66XWtUTzKsR3uy9XUKO8yfXAsTPu
erT89QSSIfh+lsbM40JC1ic7R+xTGbACIJ2/Rq90Zw6184MPVUHhVz5oHIJm0IDscfP63Pt7lqz/
IoxvKSEo0J4PjfmVczujTL/26LpQffwgAHXduq4mqZozvCGGHa3Ib7z18F52iB8VAg1MBb7TTTDZ
DbNo7zoSQ3/Mx7m3dH8dsg5Yw/3gNqcW0WIcWeawmyXnRlBtBNYmKmpYFAE2CRGFLpXWqSr5clEN
m6pmcj1lgYUjl/maAc4m4hj5Fb7j5E2YX0iDFKc44eJi5tPBAKbvyCFaE2AjnvzM6jTS0+0ibekt
yKAdkwe6Xu5TZUSlkwwApauprfAUdCTwsNdM8obR90VDhqrU1ngtoGN9EGPbwZAPjivjXB3FOuPF
Ap+S1JXyQiPTxYl3NexpmEUDW1EmILhr+fqfV5o4k5xifZgB+oLG508IvnrsC6OWNgs8mVT4C5SF
1nelcjI2twr3gkWTKf3eypzItG5eb2bOpsLh6FD4CuC6koyznYO5h5vq6th6+e7cyodHujLbQYhq
N0nZjs2t5WIO8eEl1bRmzwI6VAl6tfhuNK0r7AMyt3daGxaBMV+cq8VY2td/spab9P4eIm/q6RLF
3QjOoDRNuY9XDkyP/SqJ6YCStwCd7s2zj5eKOCTLEq2ZxzamrDsA9ciAMtW6tRpzrngULKZcWk9S
2MOBmCbo/vzco23A7jD0+eWf8TtDn9PiVgjlu21FnTUbk1pmwQ7AsQ2wQzEKBD/4ljXXuFNDSHbr
BylcS2Q5gBpR0I2//ccMD12OX4CwuMXjZuS1H7YPLMJlFa7fc/T7yxts8XF89c1ZKoICLpZF++wE
/6/5RlWLKH0vgw7cD6emu+q5pCDr3VEYuTx2ZLRdI1r95RR7t3Z5TpUUU4C00taNs4wgq+3mnAd3
IXy/SCX5MKEWb77MtyfYurMK24sv18SCKYoAlw0DJhNH17BSGnYGY1sIJ0lEEWoWRivZ6qCbX4Ml
gfW/Q+dP9k2BVour3rbxSrp3PM0kEYs1mog9/GAnE6aEuikeVw1OApO/UAWoeD5qxYxmC7OIukRL
3E2fGY73UwPS2z7a0568flNFb2D8DO0cAqIvDfHCCulNSZxXHszu8IlRYH0mTGV5wO40wZyjDSKF
OZMyISvH1tXTHwNFbY2N8z5z5/vewWK27fFxgSodOaCW42XENO46CVfmiltZzx9sx0UNV5bEWh8q
wv7Jtut7hgsO7CuTwq5vvk1R9ZZuWm1qezu0M/smMEdU4XwWPEDsBV+oRgmYUlmfGXzbvKCLTYgQ
y87PRL+0FCJYc+MOqGN2U0bHnJOXElrvYUeaIWeZl+gCJfqkIAWbfwlBn0KYRal02aYTy6fMvRbd
q5rf1gwJBELXLE1e8SbbQVtajrJez2C7Poh2XC/1dTRMjXVPXKnvgWu99BWljJDh68zGi4Hvqy6Z
8ly3JI4BWhWKPsHHFhNHxWyPswqxHaTrRQO83EX51ZTT+TOQxU/owhrUNs2I7qDkVISpZ1QMP0st
nS/6UkSWQeyiQOuhh2lrBSVLjMbdNL/8Glx33RhNGDJdfeGalj08jDgmdXOyle19gvcScIRzkSwp
xsShMK8pw9wGYaOitzKRB+0Je309pFQqTh0PnSDoCtB2FHP7tRIzpoLVQos3ta1pTUwR6KJ8oRXp
3T0gW9oJdNkFdOc6sw9BFW8xsxamrrjHSZt9nPgu2+6MCRRMLrVAL2yCtYMF6lWiQmqDZx0fUtTL
T30F/RmKYqrdgxQ++n2Leg78giTdPlb5kBgBb8l89h/fcBauvgm03u3yDx4nHy8VUJG8iESITEsQ
iFkU1PdBr9XJCRmyTbbcxR6LNdcZwr4ILKQL/rBNzlVRC6eNzvSeSj1h+ACcrqstPpaxSj+gMxCt
iBG+hqHxbTuUGWobJC3a30szJTPDmviUj1dq2lFqYLaau7kZxGHD5er6wINpnxiUdB0SJZ7CjF0W
j5nAODyptTyi5FgAnxQnXDFp0ShqoOJluAyLe9GHPK/4rGa8X1iqIV55SGUHAd5xAxaD1oi4msy/
Z4eGsB/MpT1Y0j6UPWA8HTAsp2lbQrR+X/Ly6y27Y4IQobVpPB+vyOuqD4lkyP3MF+CN++SnN8pn
Kwq1IqZ4560ljF28EuUZ+vx/Ys/EA5+OwIlrvSc4fKamU65cf8r4kSvc1XYbH4JosEqfd8oaKl1W
DaZqHlvT0cgJ0q098woIZbKtdAsQxISYR6K8qXok2hYo/+TjQEYDGIRZOoZ677UGoE5F4Evpbk23
ttVS9zy2EmZTyjQ+xS8dUSqTlImYcLZjHZO1CPgql+7GDfpLhJO6ARMK7o8n8CAon78HxoHkLKkj
vF/cG4lqXrk/R7+psyFd3QASZ4fYacNkMVaoUQWmIHFYI1AS/v8UZnEvSVjqQLlyhEJPE4zOQU7z
Em/VbnrHvdTXOP0awlgQh5NyTHQsjKjNiwy5TPGAmkxI6lZJu54c9cbPFEX3k4YQfiFOazC3fQ+c
UohNBK91YcUqr17xD2izRX+aU8EfFQTGFgeI+WHChVrAiqLo7fx8djWyVF6cdq4q6pD5LcwAR3A+
6+Mcn3/+zVYCLmNVEcb58zdOXq7D8VbnAn0df2Aq+c5Olgg77jYyAsE2O6gbX2zX37YGPynyb8ri
/DIclsRxyH3NsMuSfz18zlmJHzunXv/9lleGPVgxvLjk8LU9LcdXF9pfkkznRR292+mVULNBXd7l
kDqdqi2sxskVzZ6rMDig/cYKBfs6gjp1qr/hvE3CrdNmPXpRm/l7mvLS04edVlboXr5adlMwSJAn
GsS9qKocYVGTtSgGl7AV/yJUEUW24P4oT6qfiWqjoxjN1tf8iZ8ePaOBmUNFbR6U82JUbtMhVDbH
16bx0rJxvGO6+tdGOhGO6tLaIFWZb+/pZf5cyyl8+UwdcSFZrEe7VODYZ7csquUDEVv5LmnFyLzL
TdvZCcwJqCJou+RVD4Se2BnyGK4+szhvXjOJVEJH6hGfn39Slgs0nkmiDMBL5jiQpQ7mfV060zLw
zqt5wOO6MweBe7GHmVc2b42JEy326bHVUJInMD498JP9eiG+Lz3rzSZoSr131BmpWTh0TcBw80VW
5JNagUfBju/xuv/44koqI+Bqa8dlLeNhWleeHdH5N51CfyeazLwM/PUTBevuTmEwbj0IdlJ6/IoR
XMG9BibHek0lC1BkW6/potT6GkXbWZBNVkWNzYQcM0o/ppNvNLiLDgVUxpbKlDG3lk0Swmdhm+sr
uMnJy5xuWXKisVTtSG0ieNgPlPy5MIBw/iXhfBeBp2mq4g9W5DV1k4+Zxa9zK+5QPJr6PhfIw5JV
EpaNElPoyL0vsApCaUzSWBfrFKjlizGMkuLOS3+BlhzfMmXO+Oh4a+lvEtlMZr4Y1eC5pITtmUnO
3F99ozHFS3s+NG4zkgIteamEj6FU4d7sgLObXXqjszKDz4kFEMuitBP1MAJSSQ2mBY6YA8/gUDC9
C0ZHsPHzMXsU4p0gPeda7Ipuv75UDLLh1Kt74ZRWyL8M28FCjCU5txy6WmlKwb+DJ+guxK1dmITQ
TpucqXVGH/e936oyGVQDDDcj6D9vJ6Io5CuwhD9v406/D/IDLOCw3++BEaV11fmVpPmruKrapydv
GMX353A2rSVTecz/aW5EWal7GSEf1sxevKv6HEYgCLiDT3FPhMevTLH/4yDHUzD/ICnsLlOvPEPa
DHOjclGuibV/jtm4dbBsSiC9M8WRDV1xCkbmWV5PnAMgGHBl71Nvbq0ySp98i8RTVrxes48Chaf3
j5ZuHscRsWL6ctIYruFdnPFsd9PmQ4ZG9XX2YIN3XTy3+k0C4pl/9oe+toYEAjxHT2ve9sLMyKt4
4KcMCkCn9sZS+mBMHLzUbnrmc2/Ah4EuUHKohRrJmXDxDluxf7z2/b7f/cAnGozTUqdNGY7b60W2
J8Z/ZgfES5VF47bEBA5xzKBqBz+opvDeV7jrCtq+lBJky+WCohtIspdXvtlbHYtKj0p/DcQ/cuqj
Exi9El5+Eb2bYT0rHtXBIQTTGrJTC48sIxBINgV+BU4SSl1hX/j1W7Y8DJl+yqGms5LObEWxOqUP
PAONvTJoM/y6sHgQiDZjDv5dAIgXHT9EAGqu06J59ywlduRX3co0B0joQao7rQiATSI89fzOM6oW
T0EcojIKyLfVRKfdqq0eNViQRCo6HdqdRLFmIzFzbqkyNPpxeZCSL+buMDboUO0oGJUhqNLyoNNs
SRG4wszLr4+WOWR2B2X23G6F5dB6zBZeOBZfXhiVJKui5o1xP2sTucbeXGqUCmaXWzYUWli0sPOk
Qy24el7T2fPsac67osbgffmrmummH+DOfBOzFZSiI0FwD60Z6Z7X/JJUBijtqs8kGO9eul9JscPI
6b9mdgcIhGyo9UEz7eAXt2Es/lUSIdSR6fG6bUCm1m+RWMoDE6/zDnK1naBuAosxmp4ERSlYGEL6
70qAEcwWMHl9QIwNdQitn8/dCFYJ8fxPqPPbUBOMCctbx6vut9vtaovFGYF5DkzjoJthqcMApplR
EPUk4rbwilD3GEKu/451sAPkbZcKvTlA6hGfXH447frJPCs7edJmAT/0AdiT7abTl5XGFKMQBdRH
o2KUHJ0gJRNAkQjVL3IsuKtU6yPUMVKGqf6hiEkC0QZ61oA1Da3WkkBjxOpequ9lzxa5ZRRDNOG3
vuFkFWq4RIcLoYq0vJrqebWaChq0b2/5cPf9KJfvUmyWVmNQCl194SoZyCgt/lr1vEPFszuhKP6n
/l1dvvWorKogpjNWw/NLzVGT79ZFBRdclY9InTDUezqt8iovz5UxqXgTKfvr+tSHNUgsmb1/e6Mf
GUGzjq7zLg0fTuhFjXCk1/Sizgx9Gz112xMCUGBJ2wfmpdC7khgrAQa4/gRSkUYyT2LBsU3oF48p
cYDNqqfQB3l7wz+TlSp9HzQPi7zwqF+lkX+C+uQ8evTJQq8K9Wgm9sSaa0rI+1utbWSv+mNETERZ
fnOVBbRVLxAHKKDmNuv8SEIvDCeQLTd89XaOuATn6Qw5y/JnMJeDkQanUpu2xTx6C2vFYlgQD4Cf
RTgdOjnVBQvtfhXa67czCuDxCqCS4rgT+OkK/0TKqDP5xovGvU1NqfJPGG9KopHE1UYCqZPNHu+1
IozGrSXFc0hxPEHRrCNf7OVTjGiQpfAJSvf8JQEhbQHefJRCOLGvVgRbVzj0R2UuB2suME9GMEr5
hw+bIvgC6RecjscFWRK3tHJka0X/7lE+4tHMCIIEfA7qnv4rSgfaxDGRlXEgEQCIjquqAIkrN8by
//lFynt1Br43T+yK4651ajL/D2MTLzbI7wjymtRqG2neEYk3GUsd1ef6+toUUNfGPtvmS+y+6Ifk
uEswixVKkdKposySDY3E+rkuFX2riXVHBrDRxaXyNbIjRUpT7+x9y5+aeS3vRLCCxRDUzzna/2DQ
SJzN5ESOfGUtT0IwwKZhCJCy5Xcx3nNr4N3Uq6jrSDP3FDDpnDWrpJXV/NgUl5StuxC4F1QLdfk7
AqpAUkxwK9NOM0ENtEBAUPviaECGOnpTfaNRffmU/UKCfV+1xPHNVk3T5HL0PwY+AzakdnUWAklH
HKWuqQjZL0yfNcEDXw2CZAb384IIAMmGIZqng4GGaqv8eiv9L6VcRY8TMwH8UK21xaDbcqtvkHZ1
yCdNFnan5zr+G5a3tiY4bNQczfoA8gsNn2IIftUwtlpNZ5N5hRebTY7Pz8qrnO8gBCAvT1ABF35l
mSA+UgGytXoTofveTD8lOn7JC78eZBfXxXto15glDV7wHwDxjT0INjqbVqPELdvFuQmS1ukScM9T
fDVoumIruyYyvHHcZOhKiNe5N2s64pbrta0E+/2MJFLsw1R76rFkov+f0QryVHuA8DOn+nhObRjt
jJmBQ5r/EWkkorW9LkbP3doMaox5DsbrSjLB4Aer2gn3tGsH7V0uF+WZSu58elvDygmBEsamedDm
qXcDZk3X6F2FKAOtF/bBXd0ea+6zFZe2t9RljSIYAaQk2Cbumz6zKKZure0DAnKkwFYKSbNMo00U
JaA6aQpBtI+vqfjsxAWWqXSMPqUVU9kj1r9WClhyv0LL3H6HSq33E4TlpltlMs2FsOQWdjaeN8Vv
dZ4mAYFIbLSPO6CS5zQ31tHfTMzC6NmFt3IiwX+Va5byiMWOGQBW2kMThGQcvNBXtJUMRRDlwgQY
PjRb81pQeep/0Jipq1wyfi7le5GMWCw8ZEr2h/I3iezB+TrtHya4JDPx1sKTNvrJxdV7brC1emb3
GwvTeFq/kAowkSrLNb31uzRmU0XZHejkgqhPodz1XeMI1hETcaXrqja7CJt8wFqeupGXvPACEZqy
dzgEmvtYnjo0K/+XzUqmdKa6fFNdwrgZi3isMkJFNr1NUylMmaCKtB4dltEk60kOjLLUHo7uAJJ9
uNhLjIRYQfhrJaVta+BpdXkU3Wm2FYkGAJNTr56GdPDYwfciHjsiqZZX+MduxXfaBnm1KaLJcByZ
IWopNwi/DdAdsI+pazovVo0V6ioDMy5B/NKRZMQQuINy6NW6BnZAcqARcBawqrts+MejAJNdxnyh
c8ukA2Eokoo6M8PYkW2IEmo9a+gtTXbbNC6wVt855NZqHGPI6sQRNGskDIPU0T84qtNiVt7m7t4G
bRkY+HhVm8sBfojiOzc1r3zQw1N9y6JB12RV4XHiWPlVW5ilMzdCB7/FjpUZXleTTiLOI2nPzGAh
+eEYiZGsTtPozR4rZ2xbriWDS2otxsd2FThgXGcK2XmyeWh10rxpHDKt/opg4mUyeDJmXpqXUBvR
trgfDhW7+r/i2Qqe69PZ6GCWLEKzgpCRL2tu/mfE0UkGApVvT2WhEyG4LZX+2OS4/A+L6Av5Xr7i
vCcpwidnpAk6ogNkXKjxeSHSVkPfMZ7M/oDygLeP2XDV27xQirGDRq4G+9CiQqfr/Jo4og7jsXTH
hdn9YREtVjyfdcDukKYSHp9LcrcWQC3eJ+4NM0KAz/QOVpu9vTWMISVlzDDVCrQz/S5uYMP3Q5pW
lWmDSO8NDYOfMjQSuL+fMyWSVEPZipJvAZ74htnZT2d9W+X4OiS0U3QL4K4nbN9SjpESRhWKQyH/
3CCkF/fAONFwh8ALZf1alEiiAq9jdOZA1J2pCaQoSAX08bKuldslyT6cXitXf2MzLyFacCw+IZsB
uCA12uImiOhanSd6xiHM2sSUMDP2DedLWK8ExDmF+gY87m5Vaxg03LqbqgIGShBHKPDxqOlTsKRj
86w+4m/uaCXZTOFI4piKMWQLUJOyxpFalbX2m+mmhXSmsnJPlOS2D4zX9xpIoSX0R4jWgA1PqI/9
pfN0ODoyrd00QudnkLjfjenVD/eOtzoIDZ21qPLagCYvhhgWb5aHsl7lt8jWv/RYNgHeJfwSZg8y
qtpmUnwTDn7kp7EeoYaluDrl7iq6OZLbstsNJ0yYZasDWo5TPZg5q+n9LFWFCn8CUnRKXkncctLA
VdukRU1D0IBJUYpdd/OIV+TUfdoPce4QV9GOsRM4OjY8PxYgsY9MspzlFsqDG6wJ82MXKnjvlCSm
PM8pERIF4WIy09PxHjoAo3EC5Lz2Dm+cu8DT1X3i4xwt3RAmddJZHkg67M3dDiDnEHQ3MSJ9Phst
zFGOMR8fQ2+RMrJrdgYlgXF7Sm7uT87WLPNMxaWJVvIAMf3qApSd2PBN9moXWrAeVNRHhidNPF/7
ck7p4SPGS/sY7rS7CXvYAju2Lc1bnqmu7maC79c/J3jEu/0741Q60mlNKeng2B/kTujW8gZc6yV4
GEztSlD5nz/nXHlJB4YPyYwc2LXdB/Z3CT3egR8WNB6VYhFcBhVP0bbZ4W470iwkgu7lLdaesQMU
4HSwwylq1imhrDf1c6lcoE7GdPXfP7mPMXJUM99uV/n6A2UajBP2lvVencgssjaHPnKlyPKbShn4
/3tTWLo+XVSwwXoGfiNGjLx+8HCPapMxPnWlDYvWY3Np36vADRqboBBXr62KWjLD+FtKwCNAuu7v
NtJj2mUYgiGU//FpPMYWQo7S2a4YLa/EmN53NN9eGF5pDthJ+zv8Qul65nr/39t7b7VLDr9oOvjc
AX6GGUVn8rUP4Rt07oro7tRG7e3M0ElK/TxHQBP3zLeNnZnWGK8P//WnEBJkf/GoVa4FHd+tzeeP
eTErJUt7mYlTFDPLk09UVQsfBHCkNigbWN+X0e8FP4q9Ns52QrzddkP1qt/7qOu/JZN4XH3GRT7a
tkWhY+2k8niKzn5FQF8bWSu/weTH+l8zq7RxW+/NnE6JChH4tRGo50ldfhT642Rer/ThUlJIBeTH
6UOI8gJ9CbvrLRPywdcop8PAfDqETNxGUe8EDxY7HTV+hFnLb4Vsn8/TMvRhfUb8LCZe61mp9FD5
zi1rHmJ+EO0YUbJ3mBOyWhH8VR/OIvTA1n5TvapVOFH1gs0t8gluxlKxIUdX6wHIm0MDiNVf0p4p
V04vP+IJTb0/BX6EFAAyjHVYYUork6OOHub3yiiZIhyEYR+DIG/gaaaBue7/tmrtbs2eWXEQxVWL
pcqqiNtJ5UFvGdndGc++NMlLTQkGmqCPS9Gu2wI+p4MfuriX83lNrAQYwk/TS75oCvBBNdh9aevy
HidFt0rWrm0/bia1DQ/KXEMMWlCUfHzJPCbZ4sP95PvtEfxyL4Gs5YkEcHb7ZS1TOBItPjxbFbex
S85emrnwV6KHw+tkNroohfvL0bY4O2u+/9gEOmEcDYNx+kdVBFC1Jv+cFCSolipiytcCkdZYnqQY
h39NA/2yVqwBZINRTLPsGJbIAyk4R1QDpPJR6phgB2gVje7+ix9XYYlEPOpE3qx3smdC41OwyfFu
o4JDuH6oOOs6/SrlKjXRBBhzawLPUZmE9+DpqO39n/hd5hKg6OqnoZHFZnb2JV6/Iqi66O7XKKda
zZ0wS29G+8Ktm9zsnfyrVXsaWZlpYDG1pKwOVZJx0MIOH/p+31Mkm/QJRu/is6zCT1us+R0z1eWK
PqO1RNojKjib6YRKyup20KdfmncQBqntaLhdYcj978Pm+k5xgjIpmAX089j7VKPQlcrlGtY58rJI
KJHwTESdXJZBWboFDrIpPlC8fLNtfINHmLzU3YVPKvsEy50ScBC/0KfLyFIv/03L71pZ3jhsEH7f
Egxf7SrXWM59j5XPjF8Mw6Lmp4vmuSpTwpy7J1pNK4SIpWz3GKWXgLim4+6qflZBh4RcGnM1wbek
JJomi5kHdUp4ULkGyWjv32imI1cd3+dgmVlvlrhpEarR0phj33RCW2O4hU86DEzLfofcQpKgcVuh
MhaUCh9SZQ5U8tpk2kOH7lPp4nj1ojRfYn4X3JOpNBA1p5y56ob97wvOBGkJPeHaIF6MF0JjNCl2
qdamHf8eOaI88DZH13rKYvfZ0wBCr6TW4bsLGOaR3pvWFctMA6PA8BmyHaSPtITy0vI7k0MX2rE6
nEYQ+lI62b4mmt7TYyzPL8RH5cYcnyZkEYdhYqP/rOgn7DrXV46MJqcO9SED2+BrDuIIHI6S1gCi
6tPGsPudm86UIsH0pv4D6FLTk/Dr/1fQ2Dv+2qrgDRDnYYmLk8yMUO3xKqaqW4b2tYV3ZDVLMlpE
DZMwH6NRNh+YcKgmIijCIfWJ9L23BsgsIoqdy/3tpDHbEKNg8P8+cLlfoOTD4PQigUNTN1dXiUQd
4SBhJgqGaFOC+bdQOpA+ogyk/ZfHIvUjBuvKDej8dJu6W1YCmKwYCOjjaKKA9Zl1idc9c5+7lBK2
DcjMt13LlCZiEjDZlNe6oycn0heM7ORwP4RfZ8GUbYanpJt5i4lAc8w6M627hVGBA1kxErai1KCu
RRvE7ihw7+4yAPI3+it3wZkbci22rvaG9eg1vPdBwKJCoToRrvsS0UI8BiOVa/bquoEn1OkVrRMm
BYe44yAvbQmJ665SCvxFxNdMiuCIO+AroL4SgKVw/alvsfnKYwAf4DW+lsFQ29eVazGO1Aa1K73c
mVDxEjtOeFSBPCNldEu2U9XrfXIb3FDJ4ysJQa9NVTnLadKYVbRkgQyjCoGg6jabdgOSRGn1Ulhq
7cn/1D/WdBRllV18foXdRCcV7sMT6TIKkg/VBmvarwfzZxeIly6l8PuG6lOEIExpxBleSxey0EPe
AupHaWGKUiRvPhEJeN/ZnK8+1ze1q8ggieTPAe83ZD+gy5Ksjf+zQQ4SWb7Y6Nv4h2B5vZlHuKi5
jwAW1SvlyQezAl5nBtFseGi9+u3R1K9oqL1pMRo8tm+5faM5LNXS8IJhKbFZa4f2riU9hcBsUWlT
4UdNjaDZOdyDD2ScQ7Rpm+BwOuk0UW0P0ItDrOju3zeqjm+TSG0RfQp4xJAq5fSMwy2YWGI6Nn1q
D1Hlq7aogjSRTX7WUBv/GACCEphNN9gc7L5J7u8FXvTabu/EjGA0ifA7gfJbepUiXudnS++wHkRL
fB9dFZDAPpW2Vu+YB7FJyeMym1+aXt285jgrHSUUQsCTR3WAl5BbrU6/txRfZo2x5Zop03daIASG
auErAu0QF+Swk8PHYMceE4M5Ahx57K6dRO/ifvGvaX5VU20gmDj5tVTotLHsxFyoJ/8HOwrxbrDs
/M/4VUBKnUUan8ZUat/p8RR6wb7oJr6Yu1T21nwJtRB873LRlBgsGjb3D8OZ4WN3zqNbveSd3N7q
1WVgbQUIYiU2ka4bpSZtaWcZavcqs6ClEiXuNWhVuc9D7KQlnJGRuAolgSPrFMDRc72oJFyZMveW
3AgN447t7EEDv380075kXcTYSTYiVMYsZtEMjPwY0xiNzLYCy7+spNPmi0GDdaltWK2v+jImLND1
+OOAopTdHCydSF7lkU+TJxvjr8zEJQM6BbSFC3kLM51ecKSRGSMbmEx9u5ESs2NTSLSgn9hxRlQS
elJabmTp0OwEQzlVhf9RQ0ZptGimsl3BIeknQHjWo+jVSIYeEIvDsiFj7ncKgdb0z6zzKeuBWmIk
0LB3wu5U4FgUxBt3PL3khOWvRT+eYHuaARSJaBaTFoCgD9t3llrD64QLOAx/MigGHSk7CLZorIEP
8BhVq8lXmHNBQB66YGxnuNpS7NdBYkaVoqY8okp7Nx4NYEiywxBsZ+iUuSQbhbhR73DVC3IBsyZW
4yp38oSfHUV9UiZQW0KQCLM8PebcjW34+5J8AwNKwTsbVyoTzuDjQS8xXYaqbZvLhjIHEn6rwKwV
1nDTZ/qgvI994waeYcTGKV0Jxe42f8K99vGuzaHcuwtUicxzlij/uwZfEzw1i7QeeRb+28tu65JH
thuiM3Y2SZ4JdCfwPY+ayDjjdAH4bXA/WWTieP2FHZPICh0S/F0ffWZioSwjSN3hrFs+hb6ZmZxt
5m3buzj0AG89df7M5ZyacZauiqg6vTcWo9Rl6Ko8ClbyS0KokxO/fGYAEonvqaqOUOXirM7D1ny9
Gn8IlGuir7arQlP8NLtvizR9xuPaqvzzlHiVczW6g8cmW9eEnColl64wv0U9SFC0ZE+gqquRpsck
4OUnRgWMP3FUMx7Fh/Nc/b/5qaFbrmKpn9hL5OuytjeQHBbVNfRkn2m9FxOpZMp1rK928kVS/NvE
h2m7NVPnomSJUOhDmdIg7TiybAJVn6LCgB5XbNGij01C1ci5Jcl75zSAlEMA8p5ctFZkZI41mT4K
ZlfDnqQieSJtqGQTLLqRhEFkqYElNv74hctR/fPfo/90jfxaq9oA1H5CPE2IBFnRds8IETRWnKO2
6/iojR5lKdL6XpX/yYUYN7IXUIyP80I69eqepcregnP6SPTrChS6lHpSixyYZ5mBjDGIAakNyYc2
V9Q1mZxpmHwr5hIKqL26fmeBGzuEgTEPZ8J2wT0ymAxLuJYRBnqPTDP12b28wGfmwrSh6Ozm5EoN
CoBIVNg0i92pAlhGAeobLFD/3pQlZipUglA7njildFJiNurGCrnkzRISoLQirZu/paQs7kYUZcjX
EV1FGn+FOe0/eCpMnH8zfBspEQzJ48ZLH7lsTBg14Hgu4IPvtell020fcMk5KWv0aD+GBEuwt+gv
AsDE0F7YRu9y9+qa6mq710LxHRCos4blGgH6qeEziM3z19xxe7wYwyB+tyl/DlOojHwsBBrIIEJ3
ZzBmok1bnqN7AFSC28SgtTc+rGmIX4IVabl2Zq0/Bou2gYOiTnRbgcuEjmrxgYdJWnPro6ewpFmm
WVwvFeDGC6AcJ9HWGID/wiWwqkdMbPB+L6eGqeu2fES7Z5biEVtWfF4yiY4OnP+TwKUbc4lZq12y
g0VcpaHG1ieKoDv2eiuTAQz81X7o3A5Avm1riI1WtXfNbLNmTEZhgS8JrjRsdNHE3aGbLuZjJNqj
lYTwraxl1sSXP+iStBWDHzbenxadeM3mIb6cel/86GUN3K5JBXH2DyfJwzJSe8n8IP71lI2oLZMw
U77yl8vYM1LQkEjbTMkgHZE9yqbhWs5PIYdkqccRTuseh8i33sIjyYu+/hYJIiLgzQtIU+HgdiuN
3x7yxwQ/CZzrVvg5XHct3+kx4Mcd3rXY86yPKUGqVEtZNT2ytg5j1+TMxFrR98m1afiEVcylplgn
XOBt5ICRqZbW1oVMOyH+DFKcpHcDOWqATXVs7QN1jZZ7sDFuCYqHt7+vf5hGWy1/S7Zylv8YY7wY
Yszc9k1EmGgLkd2AyNabDnOHjHAX90bNecBpr79OrxdYTv7CEKsfLdrBk9btEVegK/uY0ofAMbfM
YJxsAFH+KlQuhOJS4yvLTcMXN52I70pOuMzVFAdEVRCwk8YaxqpjBho7sQx5pFw44GdDNycd4uzV
7Km3eEVDpOxwzCUEJC/eXsTyelBE8N2E7L6wUxAFmEF9pQ3M2lt9EdWxhMu9t127rFm1ZFc74zoc
/KB/0Yqs5IiMZ450K/t4OHN9S1SJBAHFh0/le0xeaJO8iM/IZxu+nUUTJhEsj0eG/Bp9ffsB6QXx
QassVMnUKSQn3P/5CFFCa66caWhNuLrl1qKsbW/8rDtPztWS4/zm/T17qmKHFY0xi6ubyXSpo/6B
9bktNHSQamv1wn7zz7Qas/zU1Ms61JGSlhHZOb2r5LeqpEyeW18+p0Y0Nsf38Zr6/mXlYFe+DKYA
HUYxaR7CTpCa2ChclgjXcqLdHwKvjuX1AStBqVsOdt8PSLSO15cOIGpnMsr6SMLqbujq6kJLtEaU
K0mSfv8AV2ivI79flwX+WcJ0J465hR8rKjjF/4KPIftgMps+KWa/911WRoakgc+JIt/98vDEfR6+
LS5bp3hlQhuWQUeriYCemNQ2ViEEM0Bx2fOxIM/IH/zrMrcrHdVO0AQPIW3skzBrs+rlicIclpkt
948crOw9RInAtf4w7NsKNrPyIZhcck1ZyFVLpNDTsF+uaAOv3AFAbxXXbEi7S5Iu9cXOZgHTcFjf
wWoohcAEVNoWAh1l9wkLiPN1dGdvdJqmcdP/P+EU+LtQ2f+x2LmYcztN6LTUDLgILa5g88TmKctH
wSsf1ep0hqw1RKDzVBGBJZRCyJDPbc6G7Vz6XvhZ6c0dS/j2RF3VhMMRkyZX8c+4dMxRDaOMMLLJ
NQ67lXxiPqlBE0t+hQsGT/gKNLemq8tAP5Cbm1xZ0doEQORnRTvGWHnW7lYw02oJ50BspHyTtFY3
/ENnTubrr5mB157HOELiR6sBaKwzEcyMfk0hLjX5eEKEz043Sn1/1rRig/eaqqOyas7+jFRlU5pH
uSrB/Layt4ve3RT+x0ECQHJBQuLNnJuGIgeBKPIXnK6ngQ0ifSQiVr4sEcy2S8AJ3BWEHyH6IbwC
k98Tq+G4dW92Mu016O2Ll9JWdRtgA4jZIX87Y/TO9qh8++T5L6B17iKHpPvl0IqU//ROfKyJ5MWJ
4yoZXi6ZzEtag1xLbKdeENoqu+sMUdfqS+kHiivv3+btElpEilUHAlAytP7HnJzkiufqDkGYHpnX
TP0zJT1JxVVF7EDI89vzvJp88f3usv8RxlLp0c2jCviDIJjq7mMlPt/2BdBO8qynfglMupUH/phu
YiToC2+Yha0VNMklQbohGCZOP5pCseHRoO1mZzRcT1MW9fUzg0X+dRtc6aA3fcdykWxsdQZPXI22
UrJp7kkh+qPIia79JRIjrmQfA8w8P886yy6ve7qnqvZ44Luwwcigy8WL7yUT5zaeN/3jbwrdK8Ko
shpuIqKTiimWm/HS97YVXy35a8EMi8aZUmGnlsqYbYcgj2kpJf2Q1+dFgxX2KMOe/raOAsfD1NnD
nFl/IFV5RlotRYC3ftK7Vv90ZOaQyRD8soxZt2z6cPtjNSf7ZEfbDthk8f/4M1eh+oQ1F2hQ5diy
Sv/iFJg3jlNXVCMBJMI9xz7VU7aJXSdOs4FnoDeq7aC4HRd27Ag4xR8rWB5ALj+e+aggw9Crdmh6
vvHKx1SzgUQGhb15AQcd365DSxbgemg9z2ewO1Joeldi0LJ19dzDdpTx8ud3SeBndIarX0MbfCsM
7BC6xtCOyOJWenrcvO6AhZRI0j2sGnc2KiXrVAAImslMtZc+tz7JDsD2jlNQFRWFK+081f6+CXTX
4lP9K/g/yDbsnYtDfFwbowKzf5B5smq0dovPc/yykgzGK8377u1b47Xmvt+LhFOcy5EYggpv5VOL
RNDCl1b30kNtiWKruTiIQDGPB4IUso5hIE2M5OaYAlHL2kE4kN8tWM1r3TSfHCORYd4zKeJ1VmHj
Gno81XezzeMyUCZ8eM/gPCHdUadVXEWr+IajCMfthLqhfP70T5Oi72BddtMAkK8aZLDDPnjnpRHg
aO5Un/N0fZ/qMZDHXvawSKOGNQqjSUyoHmQlE9UGhhygKVTs7kl1Jg+Y6QhICTZY5BAs2y42xrHN
pl3VLVyuUstAxS6T3GbOsgt7tJSYQvCXGbMK/ryWDscj67nk6NkIEb+8Pp6Tj1GNzebAbsZUskKi
342mXsDHUF5LfmwcWG6xghPmg424pZjCG6JfpyGyE9azDsk4+lvZuIeq1mQJwbhNspdS5nxTzGBd
fgGXSBIrWOnC3FWV29g1iXzF5TlGX/ElDEUPOXR9yvtyx3wp3NWjtT+3fUFoM2YWByzuXL8bneRi
3L84ScSUf8YrXELUwlno5RDuFxqE6GJpNC5drP1L07vGVEXtMI2zfD/opc5o+q+zyO6xbGk5SBlg
QoXkcRugW/rBqc7QaNwrpsxa+6XGTMBzNn/7T8/rRzJlEBrGuunBnBgR2VHc0uojTsrMia4vlpkm
E8PzvGsKHa3txPuwHdXQgXeYmMpy0xvJVPfqf6GmG5SHHFoBTqm/0TZQ8uL+CdM5uxZfbkaDtuF5
OY1C7ZS+9af+pabUqomdeP0wzi48Sh0zO+x1S53jRzwn9OG9FiEPzC9Em9rax1h+7mbB9H1AnvJl
V3J48CApofB4TudLPbA/6LUzHs7VcKpgGupy9ZTPuOvp/W7ivt++R5uJvhcnnaGrtH55VjauHYqi
+e6zvLYFwcQvFJipqSc4CLQgyzzEVMr2euLRbVle3RfXYaJuOgHB4z18ZZzoTaT1A1xk6fgizFtd
EIbPgfzpMtHUbztPkXIXBKszUCAQQcZMxvoki+iXt9NRBDVABA0xsoX83FFsr+A43lrVr5HrnJ0A
kwd8d9tsr7YpOnYue7df4kfch802MbSwXNIFZ1/X04V/bSyKwPppCD4oUqgoA0cXHnCGgP8N5n8b
hfqmrT7GJZh0NoQb6JcXa9AE8wTj+y3fAxLd6fUQBADckY51gwfsQFTrMV9mSQZQWQxwMFz+B9e9
2u0Abg7Ge9vlRbqZPjX/YT/6GOrR3Z7g/Z1L4dJ2gMgUdLwzprgezPUZSGHP9ZGVg8m0gDaJUkoY
95Rg/ArBlM4aTmwXbKjR+ym3q2RXcUiIl2/3evpoZ+GWtcx3wh6EeVs+yfJgEYoBxvv1Mp2MCXs4
tzvUOqh3ABpNerHXuvIpKKMobz/360uZahWajEvQWBuozYDtwa9sglWuXLCXoVqc1AvhBoQtjSsv
U/o4GdnVo39AkQSAf0SM9BPk3PgLbsKcdEHDvEnii7dHXfXPsDVI6+Ok2tpeMYbxMBZ86wwcxRkt
YYXl935hZVVzyHH96K3cuGikDFRenrbGYNGkc2RLFCxnOFQu3wVT1Xhj+ieGr/gVFHz+mVcJW9L4
9NpKVX1zVe2ZuSRAfDwwYyQHceW6lIYqo1vGtdcjZmSkbHpJXaZ5Wc9n+Dwr5wRTfrv5wlJdNjya
3OrDBLlboP3eLzV/O+Z0bcIesB/9xbIGPSvZ7b2cfoGgulnI1wfbUakIAXo0S7Qlswnm776w2aGY
HPN6XzPLTkPEnmrzBnexL9tJJ6VrNUqiqxArHVPdTfjoEkz0Jw/MNykF3720vu64ten5SKzYkZpi
t8s2AkkNyLVA8ixVst5dqFTA3e2K3MzKd+Sk326TFd+Ax5axOx2CmZ4kUCIhU6J4YQL5EVs7MDZP
ZzHV+ybrCqwzjkZZP/A0oenparMkxd5Vgo7ilxa50M8+kcXuW2dv4BNQMYVbLrakWx87qx9fqVS6
2jRYhCvCCA8KmMQm/E93N3QkdNgUptA5pmtQBZY87n+FpdDJepuCoNaDuqfJ34ryARNOYiIhprNh
Hib9Q5eL8WlihOKnz2DTRDOrpb3jWa4PMcdbAhYDpKR1Tk1ss8Su+AJIRoher+SI+xTXKCUyQIwd
hXck3LgGcUdmrA3Es19HWCYJOuijxNfQRvkNI1HQv1xNXMc5Cmg0fZhxy1TVxhwZ/1aeXe/8NoJB
TfN51PxoeBT9In3Egx+UohWdQT9tN8RdEkSrF1cnPujLOlSmh0LWyLhadU8XYVJTNagcRHmSBv/Q
kYGlI1XUcoV38+8+r23GT93oQuv+JIOsfdyUitg5krYsT1KdVFsUa6ozCCFAHGgQqkvCAKuZySfJ
LFhTNdJMzMCn86IomMlMDcwkOLypMyvFeLeGY3SIEdEyqhQ8owAIxLSXXuljFXlXWqDuM7KQnc8H
8PM6Cem/wdSpGXseld8p0QUJak8Y0k1h3/EcKKhV2Q32wIM8MnNMv1P9krznQ5VWL7pzCCoW3hSV
Vkp/P2v3DK4B9+1b3Xe9CUmipFj6DuGctHKUc/QU2KRyrOvb2MmZPE58u6q9hVQ8BKZ37uDLnATT
4nIJ2QFOBKf1NadSyUg0UM68zfeIpE3hvDbsiNrYSt5RlPxwnlcrZUKUpUVwT4Ij2qBF9ng5gqE3
8lcF/yJtXdKhnOjFrXcmH0tcsKrQ/unRtf9HGcXsfumC2upNWdzUVztehbQDYf46L63CXdF0Y+rE
trH64CZlratJ7dzUUVmw0ugtungTXfJSI84q48pzi4iGZBeDVHo3D+Z/S9kB2MjiboMdGxZ2Kre6
uWmjgD4j3O2gxqmX6qrlIKx5hj4Bg+7RoKhAfpz4lASPJPwOxmkd/jYMyJWF4lhuUrsnQzOf0B+H
qaYSXjZRaLDkkrLnAONzuEGWjyXLPBQ76ZXOW0G9T9mXIFUil0Z8v+3rl7qIKOpERuzKprjhMvO1
2WhhqNxrh2FkvhaAvxkfsoEBKWyo7yncnuhC/xvYgTu4QHnpIZ1W1Rj6WkeywoQhGICg1/0CkOk6
H93JSmIpt0rxn/IyrZb9eHvzzOpkKa0FPNG5mRVCb0PTES4YrnZgD9rAc9SkRkTZi7e3Lg1DoYh/
GBYmjbGUv4zcTW3BsLoG1CnFvpaCLH7MtkbbVl8Po+O3q/rKNnF7qK3FGr/dkxFzST3ePhei0ecl
vy4Pdui1xsieYk2CLxSPkj6qqkt/Fc5jrHH/i7iZXAFCcoiufWZbmBPj+r7g/S+D4lli2BMTmJAg
fGlKb3ZZqeIRXWnfezP5+a2YUmHEZM9OsinZpqr2RXHJ/BWJ3w+A7QiFYoJ6WR2ojpSgB4RmcXmx
RrUfqNG68oS+1D7+/wWRcWSjEzAAdXFOB1HKS4GmrNQF5F/jHGAgjMjXdG5YXS+418RHho6qoPs1
PFXwIfu99cFINwFfO34YhagfwGhbdZ3kCorciertuWQDcgZor7Ba1OQ8ydrH5D/hR1Kwh6PsLcpF
iynCgm4KLnPmswVT1GSHng6IBnqZUDQoLHXeAX+c5PslccjgZLM+iXmgZkyrGKUdeu6MPMST3xaY
zC2YKseL9MUnlzAoNIPsy6ULBLzbp3jMXqxkEBMhuDrzvTFQosd5a/cQ+EbXuBqUj8OvXbx7Zk2b
yzPnGCczl7bKY2Vf4UbRMM7AJMrT/9c4MJOOM3iqxU0jnQZcOwb4OrP+LlNxnpueMMV2uH1qlNTO
EDOnY58YSZAGqAqV2aVK86XhMXLEc+OyyAwatWuGY5XDECiXsHpTJ12SKPO9VJUIa6z4iNBByq+d
eXKgPJ0qTuKlPS8R8rcE+6+1fP8H/w6K9m4zH4wSq1GxtPuniEbnXkAc+zg1MfZ0rE4yYAt1VbTw
QD0hHqJqIRSTddPA6ph2ilEMr5lHBzhrn1PnzXZIPC8quEB7e3lQmQzo6+Ifu+M7RRDP3aI/tFiG
/JEntXBZdhnkuyK3fXGSFGmjONKQKUcRQLHUJGjg/jR4Y7EamASB5+4EukPFsEgWOMY3k9IqxrlY
vvBvWe9NkIOGQtf/0hXwmKGrgKxIIWb8kqpUBba3hnUzrF4QlvYqGFfxnIw9KVXLB2Rm+7Euxo+b
FZQz+8yRLJy32oscTT0FmePbfGWnotjEJzucFjEn7kHDRVKmLV2Ns7LBYFfj8+ehkC4ZY7+SJJ23
sYBmnpzE5qBeiK50aQ6RFPiIjSg1JBHCk9RCmh1xuKkZeByi19YgtJQZ8HH8PO5Dr2soXkBqo8AF
4VzvWUQn3DpUksKHFyWvKGGCFaiW58QJcElZD3CvLgyOO4yyGARZ/sZzo/3CkQb3JKrpiYlyEF/g
ZqmFySZLOIKRumAPtdWp8YqSGI1f69k8AwGRpqHMsgEcrVThVNde8BpvAYwYDlvROPBnJ2DfDTbg
5JRD3V80E15/Ha4CJQOhCgG++zY6VcqMZKEwdVkQyFgVBk/0HB1j+FhKgM6jTUILB3+LkKRe4uFw
Fsc+zbQvb5OliSPhhpyae8vNG/Fh9kInulTXDW+dAJpLkoi7ECRnWgAfcUClRCymmJOBEV4EQ//z
EkD+lvOvlSCMr2QYhRCt/ywZZHY1HcYvBabPyXV7v9OrXrRtQZ+qhx2EHHTqaAH9A/UmMttDcLT0
RD3MTbgTrH4+Z37zbJG48bqL3CBMB85oag5hRyuGyvS2gwaC2awjU2b/Uq4i3cOWfU7Jp+T/tWoA
0vuNiFKQm8Eq14kbnkfDeVvMl3p4wlcmNOem8hYhBPT0CvVtEs0Y+hd4Hc2U1EB0DqK8Y7bZrK00
Vw4FVtvWyS26REI0BfSdMqg3onN++RX76cRJr49THJ+1SuOpVlLD5Ugj2VDYHSl2oPHhCkQb6kuE
Q4GsupoIi3lwqH/7BcBrQP0fXLAuuBCCawOe8H5IgBDkTqjbzyPBP1SZ1TbiKWrL8QW9jYHHTXvD
sWJ63yi6RGkpD6R+rVbotvBed2PCQs35FUPjSi063/PCe/cDuE0+td7Xk8lsqMPUsXMFyW+zSaeS
z1k15P3iksF+T39s3OtFWNzY1syLGQ1d/c54yEz0ClUJtbv4gEh4Ct8CF3RTc9hSl4f4jxPw4Y2T
O1064cx1Y3Q3j9ywmmtDzPa7SLHEMbyypJU2KWDaHLXuykth5NAsmu3PVohgEsnsrfQ88udH4P5q
wC6X9tJlREqEZEgrWzn8jfA7cpUBOKZo6sTlNB9ZpkVruGN57U+4Q2/B09DGWZWXpnWyHRPeTD5R
JuVE8EUwXAinhIfggg4B0IxoTa0GNxkXH1B5A14dSWan+qVPkHk0gRx+oegYFmjlD6roAoA91eRB
hXZyoW+4dxjJ0/aVFXZXT8aGnqHugNRCA1B0A46WZAjIVlaKhx5qAF3fh4UkeILthZBKgybsoO0k
BquyDyHJgbnsrFaOBmOUl/6zp4j1qPXoFcPtmv9ljBhW34eezQm4Nm8KXBrL4Zb4ZPgyREgFeO3p
fis7C8DAUzvSBBuJsat9/lxFH7mrJZPvXSHJJJV4dNF8j0LE7FclA/f+48lkXKRhuGPhS/D6SX7s
T/rsvZR6Gb7ZxXQ2pLWxili2P/jonZX5vPdTPWJI7T0xxL/s4qp7ZrrYBv//1obK5sOahZ8320PX
pVN9j6HcNQ52cg9PBHenhvKjB3IJPQx/wkvaGwn+8aDsufnvQoh8of0M6dMzTQChTgieaEU4aBVY
jOyc+iAtmZNirUQuc8qvjNbTI48Lr+/khSrxU4ywM0/WIR31fMj72+aQz66hC9gsW+NjaXbb9G2F
px5qp7oSBY82APi3PIcAGL7+8ywZf4ujy2s0HTbBNn6UvdRRhmePbBOg1SawJdCYhGCn/ZceSfnv
WYmQq1rELas1hSyW2vlAc5kLMs8cI8X3bgDIFJxjCxgEYwrdT38oSplOnuWP8QkWFHbFYRcsfb1E
+Cnz6nufb+ghtGh2CxKi+dSnucIKyUXk7/2H+k0DMuYzSUuscbOn3z1veI/Q6qKe6MmALSelLlRu
LE/oiqPaO+Yv7fGZtZda8WEdf8DaoxvHwmBqP7GxYI/xdpLH6ZxJX0TCnZTZATGWRTGNEc5qhjkT
tLN25dXLchZjszKQkDp+gX30gE6W+XHBvlDFcX+b2pxC3nx6x3Caf/+b1PVgzeBA1Trgq0KzTCvr
6kgwvaLYwtTsecnVr3NYwjlbpGmiM6VktkqWX0K76F33qOVwqZxWOW3fgchU4x5I71DMRjm31xuD
nXTsrjqHKtss63OeQaJ0+Egi7RT3Oe625rb2acS7+nEPqRb4KA170QNBqe0oFNcBtH777pduJdM3
Xn2sXFH4IjtdJxTzorQRIprh0bXv6I9f6iMfKfgZ+Vgc6w/vTYYDJj00W5wmCxztPDhJEPJe1s+5
xCWTajNb2mSClTFl9Sr+ao4uigALYHqFL4v4Bouqe/cogIX6k++TAYvTsd/8blk8Ha/PCggDzjE2
mKLw92Vg6XexeQn4waM4uPM4Wktqfo139r5VQnZMC4JJT0gF1w1BZefxWJeTLAc4O9D0cmWb0HxD
Ku0mznT4XxFCrwOGdOZREgqFg5rK/oWbVk47KqU+EOT2OK3J5M8FFplFA1b/MsGgwlDy2NFST/9Z
Lqv/mIFucaUT1erGjm26x1X6/nfjlLwK/0dEiIxl2UMdywqxNUblyDEcPMNXgVWq7/nxRuQBTISY
0bDor0wlzNA4OoPjNiNMtQCwOrwHM6hjmodv0DdMy69wJanv10VAlB+LIYmGS2PeUtQFP/jTFi8Y
jB2JLAIaVVTwMh1xUTV0UnE6RoIttVkHeaGr75wFaeMNJGgFBicX75G0I5TnHUUvRJvpmZHJPvsg
CX/7/2GnhxErmFjz+KuLiBQulV+JT+h+MB1HAf6dmHDr2vxRRrn8hIU0sRDBwkbqKflDj4FF8/uz
1SJY3yNxK8VzAcDyJS8HoWaA7pSAJPYZwV40WwypZENeSTWbJ7eThdXn8XtxWzs+Phkw9IMVl15p
wVPLwaKKbwdoTDpQdm1dMcQlC/n/Clys509LIirLvGsdBFmY2MRLCYKx/NIvDiMcTFcuZIDOm6JM
FEXU2jijV1qShozVjBSOkfNmRTQewck+DsslltNhLOyakS7JhD691WsOzelU0wjtQWgrHhPZoHcn
PRjFu7YlyCWklE4CcfVDV2W/t5ManAwRpQEIWO9I5loeT2sYdvTpxCqq49Uiy8hJ34/28AKBUTMk
YQM3KW7sN1s26VsQPNeLBOk95mNLSdP6ZRScaClEWF0vu9EvRqkZuvMqsksuDqi0PGxZh8Yp0RD4
8CjYuRDSFyrFnQR8YG/TtUZc0qZa4s1309PkrgWW+xqi+yhzN/TUI0D3k/HPMRSLK1PPAn3biNcf
cqPPclBDYjbpWq7q76cgCiq5pfFFnmDRB10BRr0xiGeUFoE2okL/wuPzO4f3HDxkVCf6pwYI6k3E
EXjCZGxwkTqZ2M7Qz0wu0NMmMvYAVNXNmgKN0JPyz8pTrvScmEJbCZmF2dQc8HsnZSgLHxYuJENT
W9V/uq5Rp/0KLBbjYk68jRqIkBexqsb32XBixm4g4JF3kK3b84QEIeqyqJFNmSlhvxVboNxHNBbT
1RsYScYeDfJBeWdy3Op9eUqkvbmulv6Ry+SbpdE2XRqsaROfOvJ3x3cOoXy5iW/oKiJdlJUDqcta
tMqWBuB8yAYvz6NoQoYO9+8+a3eKbMUbG1MP3F0GEuHxVDm42WSqVQaFVOHdYvqnNA+V/f+DL+kE
5l2j9+Lb8EeWjvrVVe3sE3pBik+/AikpwO+OJ8dsXqHrWcg9m6PBkGAktu0FtNoHi7m5CczY3VyJ
TlgWPDZDUfRD5tFysSNHdd5UNXevW0WyjjgdlgXIPCWRyZr2KyIEzNHqPnpr23QcdyjQiqS4UZph
JKmU1fzg33BLwvIUoy59QBHX7Ga67AH3LZrYv+8TAiCpOpR1NLTvndgt/2dp7j0pHkcoG5d7NqLh
imOfw3NQQGVZpvNPuCfx2K1WAgvUlz60i46T8z5KXp//E8/3AbMx2oCcGhlfRwI44wyJVYMwxtZ7
5X6Oj9ubJfIqO0bPBbmlP30WccajbvQQKnuyhp+X7FVi03uB4F8b8g8RVqa/0d1J9cDa8tHuelVE
KpG20G2ldBHEGgklyzlPQdnfSW5q6Wi/xXfiuFqocF7pWINttJB6BhF/xdaukhmxfZrARKKtPnwZ
ur4cPURNI18wlZBuHVSsjA7ntEucbLzDMOX1FGLp7RlZF8opxpXK2DeAPDqU+snixW1TLd/ufY+O
No6dBFhb9V3KV269+FF3j/DeYr0dfB9y7DoajCUEsAMgcDheqRk02q5a7OKofPl/9BrNWg8fAhJ2
Csa/DdJyksp7ZSrOft3zY3gLOoOP7BEcG8FgnU2/dZBB+5X2ecIlHDPz5KrCGT36O9J8lIJ9UFE5
2kQjjLLIPIjfxY0Okr/JUNtSsiVtzIMIzvcx2lSRi0CIVYz401NvmT6hEatBsO0ttOEaTRDCj10N
erO/8FDo7oxQJoWnCgTx83cZIDeo4R02NyLJCn6+olT9wAnJwrVjatLr+/3f6sSFtm4mH8yl4Uti
u7Pv/+bx35C3KaGmZH/EhegJoJ2E3HUp+3o/h92fxtXQjGUSKKI4kAcl3tjCH1XFgsf65ycB0gdV
1D26cdRwiOkfNQF4nHdxpC0fb90wRohJX2mBpuy0e3Vh8uRoLYZN9PfuErv+eJuB3REG55WefVH4
5EAxpr+F/UANamr1YaPlUnGKbXOgFhfDe5ApdYUYUE/FcMkLpcHmX83D2FjWP44d+lB0wM2JNpHa
Vr7lJCTnSdviEtpz8ZtZgwrCsjd7411qKgPwxbn0jW/0xbMMve8tZvgA4GrPmp6bqeGilos5SdpG
VzFRx4EyHozgGzzRv72zn7qht/bf3UO2uzu0NRxENRtaETlJ8pPMhkrEpkr9Tt0T541yHsXr+zbU
AiFvx7vP/aD0Y/wV+qc+/QzXoHJm4jR99ck1Y8E2SFDLKeNieH6dMRHNG+J1MFKqzd46T8RXe10e
+sXB1JGA+7brhBwmyrtPaSCriw+B0LfFuIlG1B048x8E3ISnYuvXIyQ2Qx7rH9uBGrAqeHosth8p
26ovRhItNbOH4hdgh72GGds7O/MiuX0yDEp+kpVVgvUisUAd+MghtZ7xqkqe2fcE+lbK/WhDuCDQ
TZHXsBNjHQqgMxOCwQZ/bh/lfwj8DhwbO3JiUPgmeOa+AgfmOEYN7qTs3iplrWYc5hvmvKLRFZYi
VkZW7rUkK5OZ/3cOaIuABsh7egD+37xMdjNkDh8wmBLWejL/23zVnqCKuYT6fL+OqDDh/hZHw3vF
7AY6QqktBtnnrFd8Y4DzRAqI1Lhj+UrYIm8R/FvGVgrqMEHTkO7EKXkZfkmesA13RXaxl2Uk/ZOc
5LFwywKlWCtAbcxJI8qP0AzdlUeI4RkPPQKNdknKplYp7FGmK/e8T+UxMkSR/ceaoTW60GYnaL+C
B+FY2efESr6M1OKtpvm+Vyq2aNDNna6g/w/dZl85fLvezH4cmIgxEzukz6AOq0ydLk5tDQGCCZ+J
YV7cA9Dcc7AuhKzy4JYo1mKsvp7eZeGvcgpSnLjwErMUf4i7pQuVBae0CFS5a+A8Gbe0/ir9Gvpp
/0/1jm2sRalqgxGo7kNM5dKOWM6T3IIcdMnc0f/q/g+5c4bCuSwgGTC0Owv8O+kpEwmWG/X2pVwW
NQhpWPL7AGZ8EwhLgznNneqwqPAuKnbYgIBELKMhyvVK02TK57LKOfS/K+KD6f5AIlf/LsGKJTp8
sYNIV74IN6VpA4LxLEKGUpnqwJF1pPkncLlXU7Xgt8f1FdFARNVzOao+5czwfmF81RD62m5Mequ0
UHT+RXUvydb20bAHhv/sjotpt6iB9SOTzpkK46UWUfzwk3DgHDM8FobYOE8nz1n1C7LpXGNap3nr
ZGhA9FafWB003EceAf/Do/gJtYQQ0emCealnwSwFIyzKCg5aSEyWoLI/c0Rk8B+VHQDppVtRp5wT
zVAokO+KU6XsdNdwCEGlL0Y+hrF/8Gv01zQm5cDfVXNduyIaDxmEYGRfPjY86g3tzOipvL7tME2Z
pzjWuWFrbJbl53DVnegtjt2pj4ZceAAJJdriCARmEdguLTbX8FyDWnnm/Z73aBiF85tbb1IzZf/g
Mlt0infJpmEC6wCPsIkZZJrGjY6pMkZRH5AUy8U36ySz9nW8vl06LKo+CG2VhWnJNIZaR6sn67JG
JvAueNTP4ZBWGIoT0nxSpYx62mRbt4Q1xpOd4P7JWkDPFsMkr0fQ/B6+wRTgf2+UcT0iHrdvq4aG
G6R3UaLcA3lfbX6TeVx/NgSs0rxxt4mcbifxSl/lOXRXjaxGw3PAmThjLoos1sd/ZoEJ7v2IGAKS
TN9b0nMx66cfA35vtLzMz4mLEMMfbkOVj977/fStHd3afFnsB+IFYzO08ke4gEJ1EcIc+rhRSFqy
8QA6BCc75oddHd/2yWpyWMUP+x7Xw3FMQyr6nxQ0Dp3rA4WkLOs4rKYPOQieLffhWtZC90dkB7i6
rBCyy2Qc223iE6ISYwtAmATtb3u2xTcrkpwcwnsD4SfKPI/JS4e6UCdGfr4d5jRLl+akQGLcbl7W
BdMXSyuC1J94ESBU0V2aVpu8KYMYGUDVobmxvE56UA1JlPgqCGCRU/TWoYFUa7Yv89+YjVgMPMYG
H8vjvHJdalekXXmq0XO0uhDlqZH+dMiwMHY9uhRurph8s8dmpQgFLTOOQBkKaFnw3JOHs9CzLAlC
J8FR+K2etnVAWl5I5Y36mLqHLHr0zKlR6zbiejI6gpYRXfSJQ+e8AvUGEn2Y/eg9DbpOFs/iabDa
f0G2HFppkBtRZMSpaFQAdA7La0YLXdai20YHp5h7vk8cYFBXauW5CxUJxMYuVXxxLT0QU5LXKBGd
gWbJoPVrGFH47gHClsLHx2F5EhUfEkSlNSmbFvu5p01AmftOG8jf5DqveTRNS0C+UIlCUob1BVEo
snm6CXyODth06iaPymUT1YUYAIx2C/k5/Ezcjp8Mzz8HYcuhdsd8zJSyAPi0lQkywQKgSUxO7UGk
gXRe7LNEHcJYkDKcMcY9kppIDczMHN1FGjXMLBK7xM/6vSu91sgsJd/mO+tM1igzyN/uo4drGuMA
lBO5mOobmuRp1UGt5lSRFF2QOtSIIJTS3l6pwC7c7EV2+csSEuQg9uAAy4Fhr9CcL1LLfXz/b8mK
Cy+za1E1vkNU8HVN/ixY4vCW7UJ4J0FDYBjuWLDmoN8ejp1z9f6zretuRFE9CaVFC+J1I/AE74nN
rGPuBiD8oxJEZAdgVqLmBumKytXHS+8jKj2D5PdggKG2YJSpoM0KiA9YLnULoMjkY/kxEwgwTeOT
eC0jiIT7EGl8CpAsbD5P2mws/kK+DeKZ73R7TxRX0uj68pvhI/1u7U/pzn9oQhGh0UGNtzO+ENeF
/xuzb54h4b8NCBwbB9zh4NQDe8/nl7wz0zxBOPOz0I8Q1ncLdJ9+KXb/m/ViX4At/enBkQPmHgXm
p4kIaFVq6+vEqjHz6QrYyv29WZVqEUVb0A3MPwBxORPOQUhF3cGEXdTnxjLGzoPPT2BAaDn8udtV
KeWBMVxbNcCndfRDu5d4G96WWdHC/FoXiIQBRDg3U3Bq+kI5ee5dv9eU+2W/BKo26Vzyzpsj1XHH
PD9W1RXMCoTIo8khqmEvbf/pSOiqeRudTBZUzszv+f3YaQx9r/GSQb6Vzrz8BACctmIqX5r0l120
dxhkGlKegWh9++4rylnGp1MgiiJdf5FQVL+caF4+hoOvdUANhuk7Kv9g0HQ6z5pkTc3fxfjF4yTQ
BcPqbTdEQIZehF6EphjAIaZ4rzfz5NtcUEF0FZHzAjJHXmGtBG1gurKNFehxMUGm/TArPThnO8YV
XAvUOschnmzSsTB5FILRhW6dwUvf7DaJzZwHhIqU34VJq938YE62DN4vD25F++PzdNbv2mr7RiTz
GUskn5rdgp/2tu9wbM6VKNKDeASqgtGwgxPFlQCZU/DWa1JFTfDPMqhPD9iT0vufW7/0dcf/FXY/
SxLrvb4wFhHnXwdMhFj9Wek+Fzi3yEqSa//o92qo4tHfFdr2M8Yd4XCHSeE21ZGcx3j6eD4azcCt
mwKnWMFzde2urKeoHAELkV0qcZ90Vg+5t2CfLgNR3Tae91d+3m9FMDOXLBZluRK2Q+Mlx4vugfvt
6/P7sk3/nErB04sa3sdhOzJOA3cvtOFSjntfgKH9XTci5ZMtG5L7Z7yNI2taK8gskXBmnaRb6Hvl
gQ4AKd2cKzFDk3+nlfgM6qEaNMYjB0ANCjgpDzSt9MGQHlHcI1UOgrUHrQt8UIYhAl+ePfdA0F/v
5qRDdOVYSt/VNSouQD3Bqo8scq53d07gxM7UeDDrrIBe+7MIHOEsTalkCyhLAotcIwkxb/i/G18d
OAEc0KBpjSeJ++dbp/T/w4s7xuDhe26iucfgcfCUUEwqhdkAish9AZbApR2SzlZW0/xZU9WWk2vD
Ad/Q56lhoAxh4KZTxS92t/i8ypNn1XgSoQM8wIesZZ6hODSHarfrE9yyAQ5Lcnqze61bJxoACK3P
M4iP0lkzv35cfx+56ti2t8ZIeiqa4v9FwPAQZRgFBAoYyZRfDRK8shAoNT793+XiWW7VCytyfwEg
JTEXYCfUgSkw0uz3/9MryZz4XYxACdSR7whyZWAa7P+sJawgFBQWoAr5RMo8IYpaYQU1ycmK0XPH
PETsIKNYCDNvhjDZxX+XG5loIg7SQD1n/65uPjKxr7iO/hILtlb/2WgMcyG8ejaNrtJWtBS8POc9
WQBdBSAaTPT350BsiW1LLwWoPx3n/yG7DWeimop4+KIPN6nUdaGiPbL5vn5pvuPEHOu8Ca1ysDr5
Dgd69rBcQ3UJRXTuVHmvQ176wFsPG6fgTD+Z87b+BSc3OpeaAZyaY/KhvlVFxOnWmowuV6SxbcdV
S7WPIp1pYaGuMHIwDyTbhkmMIm2hGCN3gDBNdUiuj4FMLNu2coLK3Ul5V6xzKYxDJ0i3u9mEkFNQ
GU2aim0moBGwhYgm/BFCUoLw8DAv3DuP/gg2DyaxDHfMPcvqIl4dblyjyRq5DzjTK5B3R8ISsbou
1oEvLLPA8IbYzldwY9yW1kUuPBr4YPg20YxG61U9aZIkiqPmMBTs/BQXXp8zbQ4AdZq8gcTg8QU0
dfwWsTrzJD/ceXE+z+MOKldfLevm5oRmtvV9T8xxwt1O/5ZM7bXUeseishy03FMvo/QLdxscEXqR
Kst5fBqtQV7BktampEtRZWcE/dK7FYG0U1FgaxfnLr1jAVDOgZuqrRdyHuNpbw2OYGKPoRLRSK+T
QZ1Thmb9WJbrgTf2vZ//oKpJZeX+wFBxEPdfClRKuXg/aE6Ks65Io2N3rjqrl7NOlnNr3fOdjKI6
M1m3/Agr9NdjmuLVP/LhfaJcCKK50nA2+wNbVbxQFsTV4VROra3WzzC30M3GKzePFPZpWrcG1AS+
+GrnR8v+heZGryk+EF2Ea6X+cMNVqlSzvGHpEcUykYDhBG52bUuEms65gEmr6UfWZG2Y0NCTCyEW
2mwsFgR72KDS7pTbEZc8lmW9cJ0xr5DnHZ6D6wn09t++vQCBg6P3And0vv/tCUBg/prDZ0Ou20FD
rokQkIQAxU6aP7AJZKEGcir8l+Y7naV9AV14Cc3xljyB3YjZMQnQ8Z7OpCT09W14A4woO871HYmX
P5B2E1wZUzWCEnyo5eTIkTMz9taYWyA7xTaSf4gHT+O954Gr8YtGpvz8BkSPzOtuMSx4YsIjyHPe
i+osD6oVzNYbrv9a7G2OGvgEhn1cn/NKRaWt9SutLPU9VM0MpYgX9JexEVIi5OVbRcFNpQKSdiok
XYUj+woA2Sv6dsd/B+guxtrimhzsteVV546X5jQUOlcxOxZpM3BLow0w+RFYl2Z/j6GGkPD3vmS+
8AyNGxueZRTDDhqngpZvkeoq1RrUimqtEUVtYkkw9ZwS5knciX0d6/M//LPQplvFKxTzXohy3ZT6
ecWOfHMHf9aaAkcba/KkL+EX+oAKdKbEjroLuozVH7toF9QrKpdM/Rc1qdMbsEMANRaF3lgkNrm0
LhKmYmTo5E7skNJJ/zRL6hdklAPu66WS621kTDe6k7U7VFzgvJgLhtfiJ1RLNiVM0LHOATjl+P+T
Sap/dke1P467nbiiY0Q3GJxm5Iwnr+5reQvv2It9mAMuOoWo72jEDdiJJs4ZHbbnT4YQukF8RnKK
sCiMMksgi54ZwkigKikc5ujl894Zxsf/qNpJryRekeKWorl0NHs8lWGUyFbpfu6TOBKiW/cSUhm3
j3tOLFZKTgCIO+NdjEnAJibt4LD6lhWbOG5W3gRWbkqB2HOv/zlnKrfEEo+kDPgYJPocvJ3QI4cm
YWjlwS02ExYGBLi49Sp9C1Dxgma8zBZrDmMTJLd9laPmZxa/xQNsulLKV37cPBGVGqJXoPWwUXKU
lbfhuiY88dxSD0x+u3zgPJ5+xXyALSxayIAtNjFCBh2n3qsg5hgINDHO/73qvy4cFrDNVKlfeTRA
61OUqoLLrwmW5ItI2VU8g1rwggxSGwMCoo+g8QTOFTVaBFPdLCjFb/1RF8QOHPBTAGFXEW9UAtuK
kLZdUPxy4OQnjkNYZY1efaU4q6E86hxYKywTh2t5a4O11Hcf1KF/I8gNxz5C0WKeqL8oOGn7qsp6
HHAuSH2jAlFzuz/hpNn47f3p3EnFRHnFiXPjHyoO8BkRu4zSrEjNRf9ofprugLD1aast0/yEZekr
5+M1Q4sWWHwcqKZNxCmhIETE+G0kcdvN9edOd16qdVISMzht6O1aHSGKeZnf5sbw7kPk/g4hnScc
+w/b6YgDncDoEgD0GYOc59KtmR5eHnNkn2XKtHKThuFoj5KZodzsKKu6YOppr5NGdK2VcfVLTuco
F12hoM9gsDH7IlrBpl5kRpVk3QLPteaeaENoMtf7u+eGKLeQhahHuG9nWJ4wp+PYEBxoPM53I8gN
PKKhM15rCZo6ZS75OUwICCAmkjNa2U/8ELEM+zGORG1L577G4wOABAWVFha78qHmoy2j0j03twoC
zMUy2L+bgSBmiEfpX1HLLQqt0TtgClPab+iJqLzuzQrYcBFnoxmYnoLmZ9brrfi0xn1WubXUtj17
yBVq2WnKG6AVfBmfxC6oFrqm6l3/DxaBju8gHqv4cj4R8USqVNOQaWlGOjF3i584YpvYZ//CGNtL
C9jvEzgL5J7Ef/75PDFoHRw/+zlPwRjJEUBa4ZFgpo1whn7UtforYAfJsYJbqraPr0brtwfSWjjU
ttXfo31VnyJCBwpaAX+nknBzqBgABFouHMZ4W8am2Tm+SUNdEkQ6Fa66FLUiAsK2sA27dhM04jsS
o8KUMqJri8wVNBoIaQtOxaKdSZsCisUJHTcUrZkPJysx8km3SQq/jvdEdfxw9Sr2Ijfubsaufgp7
ls/Bs4b6RQvPrDxePxNlsVklM490ijOUqs7XVya7oZb1hL2iBUNcgqDo64mqgJHY3FhhOZNKN2OL
DiYzyO0L+iaTdJSAK5pY3tJHEbihxH0OfJpElOtYc1dGvk0l83niTPgm8/DN0wGOD0lney6Q9SA6
lW10+r3tZeE3A8qmRtoMQmhqt4kBFKvWa/adFu01r4gP/f345k1q6TTIySXNCr/KkvaSUW1YIU1u
8dxmbGxJkubQsviSJQB3odSYyyxm1exLjpAnRukpdVr2kgqITz12HtUc8fvMk4DPvDb+VMVU2uQU
9Wx/r9dnz21TvdN7KImIeDbb7THozza+2ODWOvRNtR28ZoCP3R/+k6X3+ylHsorXhAKukuWnRrHG
FL6LFWFA7dnJ6/nPUl4v+BndoufRNsFUk0l6fr0oPCib5wGlnH/s1phQf+05fJspm1A67XLM4sW6
F2zawIXWSeAOy96EH3d4EX3OlFx5OXkXPgHmie8keCgTedqCKrwGmsmS6pX2op34tybbO/ryIbZY
6iXmlfEt3pbknvq11DMwF5khlDIzUg8ojwqxy3PvG0uJ8kC+PSvGJ4WA9o4qHgT3DLnm4O1qKX8i
KpgLdA9IQvvT8qeEDwvtvC9TaZ3MFC0aDKzRfpRHULyj81zoR/1+tT7In3F+lPKnTeu/tfKtni/a
QW7BSxUVa1VovNeArGttjB+wwrGDk5NOB/t7SBW4OkZaKCsT3yrae9ZVLX6QP3uN2qAZM7H1OCpi
Ieob6rnJ6FTx1X7t60rsOZtVYGZv1YWQlqQ9BZg8X2M1eNwaBh/v1XiqV4PcDDUqo6yGMVOdXMGi
7HZqli0TAK30e+w99Jbt8PE4V9lySCjMLXXrfixqKctBR95p5grYLDZhU1RrLYv7nnHhsktNcZGV
ybNrh7yuGbdTLtY9OzR6jMyfDLqMwdBBsmWMF/disFXfWK7s0RRIvTD3CB2Gh7rHZD8T96s1Ib1d
cF2Njd92ZhjyOSJKVll6uZP2l3Az4Ir9wSzrTbiCnUG/uZBQ1vYHJovaaeJom1QOWUMNG8QQLhqW
+UPpDgxtaYKAAWY3Gx169UDyUwiy5fxJqk6nL7FBKyPFwfGfd/h23cegeqtiDmknO7/IhoGXqCPM
a9vhkL2bMgDOgaPkWDrV4AlH+KNoE3JNM+nO2ArwEs8nUW3y1Ojc/mJilNCdoXIWefgru7cJ6qLy
0w9UP4e4tqKgfHDDlCD4MuvZvqnJrnJTJ2WysU6ll8hWBs4HoBTHpL8FISbsLjeQjHA8q/eXOreC
3Xj46hf365MNPWKi3tIBTflMOOZn/R2aiFghChxb4Zfum/whxkIm4nIbZXik4uVB+5ob57pviVQ2
MDcEu9F4aVcUpE2VdUVIHsgnKqwMocPmyYV86KT4290tEHVy9VDPVBLMjLVtvWjTu0z7VCJee5OQ
v23l7u4FO94X4YYcepUSEPfm5WM/31PyPYjzLltvgNBIvZ+YhLfIfqMnblAflQXBOOkdhhIrzok1
etG1TNvU8dURre9bWFIv92Iob1w5/RLvqwtJtvcpzazN0CF61JkX2YaXpefa+8mUUz4waYn4737s
G7A1skX6FAcmsl1bf/xDdvxIXCytq5gPHDpF1264Ouw0FyjQbEl0/Or9xfyAEfu1IrkkS2HVLwG7
mCye1EM/y7vQY0M3snFKPVV6mIWI6tXAt66ySxRLfAd/poAqSNC2vuTMkhI17xPr4BsXw6IlpRCB
owMeFfy8Dh/xr3TKra4QQk1WjXI8CVbWxzwKPopAo//i9Xtmkfc7rm+WoLXIh5VliseD6JyZkpI6
VwUrUcMmb+ln77hFeq/gflztxsoRE1C9bAt2DXUU4gRZlw66FmNTR/pmrALlTmbhikkzN6fl9YKS
SKy4MejOzRhVha9iRWBBEhptYDedVqrmNbCmAQyhXJWEqIrApZPCSQSdXaKf9d5kiwwJO0SHbngz
FXMf9qrM3PEnMRCq6bZYe7z0mXqcsKlGxG01V/K6Iawf5EG8BOY85OL9dn/gf163ZJgipLwq2hqN
QefEm+YgqpSmiOG6ZIE2PhBUKGh96EYzpqOX8pozdDI+oewCl5LUHmo+BzE+35DkDw8VQM4Pl/v8
7u36dRBlkgHrJ3sPFW4zU3CLfiFQF8OIu+hoFuAddbZSSJ75daipa7UCnezxzsxu6jLxXKooesca
lcF2nykkr0Uynh4FDZ+LnTEjIfSDwK/Nawupq/oms4kY4eAFQPmlFe+tSl0XgfNM4yvdoSGOSkNL
lcrFhBGTBy5ciralC488G2Pk3VI9pxVkSjME9eiYfXku4Ji+P3FpP7ngayx1OJCqBtT4twQnvVdR
dC9GDdCuw6CkDd7Nk0AT4RUkNVVrDRsPu5o6WDwBBIolioTX7nLO8V1bYSEDXqVHQnTj800zqRd6
YmGzWYIpefI2K0WkNSIahME5kLvYZcdXF6jvfII20R39EMuL5vTVWIzoMCrkrPY9QN1csZZHumNh
3Fnt4F0yD2Y5bRrHiK+8wwLepn/Y6Fpq6A1YFBB8SnR6LfoF8CRvGh1IuckX/eiyhWlASSWw14pJ
wSysLF5989M+zQmWQHpwKEplPk6jpdhQj9ARYfvh+Hap0exhwDcFhnbNA31p1ZDNpd4ZbwGI21KI
5BnkCIiJv8uwuJxpFL+tEWBYJe2s2INm+f2hoQwIwN0HRgf7ioD+G0o60wq3vCf4qE5g953wATZi
DVVS1KZG08NRdclOM4B5Mdjg4frfgJeJM7+2r+0OE1E1NS0vAqjdEavDB8Q5tjwY+PoIk5axBa82
E898rHVhCHXaqNQzFb2TjOXU48LPGe3BMGUysH5GNVG4xUxAZfzkAwnxYuPkTMnzpV0pTe7UuLqH
h3nunGns60yhyjlAQfbgeYQclAuOBont0ds7guf5HlSFtvXd2MvgOwD1vYOxvo+oWO/L1/nlN7G8
X0whCjvW8hmAM7+FIopnGtTuibfmn9IrhHFvaijy/1dXeyssxP/k0yOvOeqdPgkIpg0p6iA8g5Pg
rEa/gpb83bYq0Q6kFbqs3Z5Wbw94WJILavxTdhjdiWgmFZh3lMeuduRTxISjHr+hiQMedT6wIdys
5e1r3w8bV2jaewM610GlVV7k4827SiqXGr99fT6rBb2B5LswocpaCAOvK12yLXKjktk2NaHrymXC
BIl8Td4FExoUXc2h5gdVUFZwiR+Vkc0OKJdDmGRGOMGXjcMwXHGdIEwt2JzXfCGkyg4UnQLPcTo/
LicSLOgvDzpGHFAmN6XS/ghPsJqWvIZxSSkNbQPR+9pfARGso9AIFtqsEIhc7KbT3/fLIUMOECri
o3YpAnR2fJXtPoyFA9NirQ3jsLu/uMDChSJ/fu0kbYhFysjHoMGeaz5eFZsy27qr6C0UVmMbQhx5
VQg+udEPekJ6W+8aRWaiRf49ilakgEEThzXHGsbOFrvG3fE+S32hXcomKegwiOV58i5XXmius1Nz
PcRZn4LQ+x6rCZ8greTzekvrro3avPr4cOs6V+O8C9B0CJHVTRztJda9HzVPT6VHERKP2S86Wlrh
kNfNMA2BfVcyIC2i+bBNU1cQV+x6YfqPnCPvDlsfs+KCX6JGgDX/cljynX1RVn2ZAFO7wrwyVbuc
oLqtNkKcXQWJHECdNzX34KsmRXL2nkfUBJikJ1rs1VHQM/oPZLb31mw1AP1kwnW1MAO8rqOglMgM
N8IFY3nvtTiv3wkuhRzF12LRqwM5lEI73z2V8LzT7loPkVs/Ww5fJOrEj9e6ib68IRL4RymX0183
cD3p0EGLHpNXq39WU7TUpHcsGD07GMXwqMJZhGHtBDY8zYruJBJn0X8dtj8jav2OSzI8NbPZD+jt
FB14N6WCr3F9+FtzXuknyZ0SDUPHVsa2aU/r7qeG+Lzd4Nx+yuBwS4SFMF1Rxkn0PsCps4P37+ko
8TLQlTx7qvQ4Yj54iGnnfQADcLeWgT+ikrvTlmEeXSH2y72Yjof4CvDtKWDU8xGntThTsYVFaFyB
3VbwoKbO0JGBRt+Ff9SpX2cP1wLn4v11sxnPGIKGKySyUJPRZhDJExPfhRgjnVsonvUE0E0lIC9U
lqpMxs3eHXD5t328F/KFMKxVb4ync84VmO/1mCfxGNdvzuuAWb6kGaprPamEvFlDe6ckrWg8COVP
rbY/QzCiyHK5/rKAsdcEGveuBfu+6Q/F/1+91TvD3q/EPvr2yHNRCu7a7eSJlbABy3CBAcmTSmdW
vwV/44KgSxwZTRpKi0s9JiQ9IWqMAk4YYQ656bKNOjCu49D9BsgnUo67UXNv0ebCbVThwmcWhF6f
T5OKI9NdgCwu07mcOUr1ErZ9RTNLVI/cu1yvqCrga0madQq869j5rFBS8vDn8TN66HAAYnAZiwPU
UqQpG6+WbquKy9sH9dA+ZwwHoWxHgKsNo2xlnpzL0weCy/PXMJXqBjqGy450WFu6c3BYtyUJXXt1
cnL+RMuwabqsZAuHppcvAwhqqhqHFU/b4UwgmbEQb/7FZUuAoCluMGu0FHpdXJR/2oSoaZpwkkvq
aC5sjkcu8dYNXggr73/HyuTC2WLAHsuGiGpXNTJdOAYS5OdD9E1x/U9XUIIJmR4Y8PmhEDN/pjkt
glK1V3L52bGBCyfpQ7h8+xm0ts/7vOFSJdzsE0bcl3tJVXCupjpwnkPJuYiNrNvRs7z2/EH1FT2J
MhkNYILwrG5PY6p3dgjVSP8HHfIhVEXdMHqJi1tgb9MwEBSgVoZKoBzzNe49OTMBgwKKcXsNmMKM
tw2Izmfwu0AOS5X+Kn/pC5emrD1enQSMJo/Rzy6Zertkwq3P+cbvLzsc/pOJPU3w+aOWJnnC8ZN7
0LngGLqujqi+f2GCqUQUI4ZI441WuvEgJs/6FNxlLxraqw8g41F+kmZhezQNT5Jt7fdJfm1Sdoyi
r6lIA2erl7O7IpqSAo5cefGl+CKWpB5Mo9LtsrXvJ7+XQaibBaB8kX5Y9ttelepBnK2mB88Hgn1O
9sEDlUvquOMaDy6YK/dY1w59yGmPj+VDV0W5h6l0y3xsE28TNsKxVpERYGLloiDeIBujXg0YrZzC
IsemttfsXiwU3fb1CaZUTDfY4xKq/c6POLXlkMjfK5NfaL4A/NlQfhk3oib1D62T2mPi6RaijBUK
QeCNzU3NNB5zNUdzlgzkOTRnXr1imGRIR6g0LUvP3ibCHbUUZvNvzDnfDKsqCn+WILbYbmvJ1VT9
KCTJEzoNdxpjl5/PxsEIVHfnfWCiumjwCwJDJDtgDrpIjgin2mbBF2tO0zJHcUXisrpL76pNgV4j
EXvKHZaCu0T7UJW/cqhNaM2THPbNDs+EhNgLlu3YTcqIHEWYJs6V2eitl+23KqCEkCxjENCwNU9M
EOj1QiXJcJcIb6P7onAk0MWnK6TPQiHmHp60byMNGGcGijPZDn+GBnO5Yrd+53eAA0c+K13azJ6d
ZxFxOepM0T8wMdm/guqYeBKm4H58eucQhQI16Dhn3TU32K1kbR67PzUYdRf9CTkztxJRX0rl+tAt
c1OVOFKI+qmWm1ajlCg3ZXn4OPwXhmIApFa3ROlBTJqwasNxOsmRTlY0xeV4szz/jWqKNct6bJ8Z
wLhY9wpkvL+yjxbcHayBTAXzW47jqV2s+UNsispMTF/H3qISQyV8jx9iY2r2GXuHG7jHXObkf1ap
3TXStgNrgvHAFCIONLH6V/mJ6OGGCtqip4H5OlbJa/Tnrg41l1GzZN4/zX1H9WogDURARwkPoKEj
6oHBqP8ZTEbFe1ILZMHe2MUxubf+7yf9WEQzi3RkImLIGUC/TQ+fw6/c6QAOgJazcfd0x6CUIUko
fPu47xlbx0/lRDZjMlA5Z/S2lNgld3uU8Ji7KSa9ufC+53zxQ5yn0fTeeyN0UiIm0Qb5NmliXxPu
x6q0RnC6BES6m79DTdqVIXtxs/eRXfuRlxFo23HRcWScXyS81gWoYumxk6XgzDfy8DlpYwxfyEIo
XNC8fJ/gXFAdgBkQ3/3wEOCLSAFtKRpE3uv1LANb7hgtWL1xRFzr1FRL01PdeLDyLVoUyUNpKomw
O7aHglGYGkhLzqdEYAZ1TdJt9Mgy5v0MFan3cxSIhXs6THcjiMLAzVM3q3YsPh6iEX76xxzgz/o4
Q1x0mcXuzVsCMgCcI0RQE3z7YJrp+C3uWeFBqJ4QF0rwnrgS/3XAvFVxPk9S+SKTutz9m66Sy/1i
hKFLlVgAI+T9GDoV70sJ7loog/451zIp6KK/6rIWJ6wpuUHSgU/XexWa7sV+uIDbUt+rZKPCkXjg
hIE4aq5rdkjY0aqi6vDY06M/4sh6KaqAy/iCgwJOfZvO2mknvgOwyBzIgcv5FgcLycHkndAl+wwp
LGJvboi98HAdXHXUZVkeYHmfctnSa6I3Y27GQRj0gV7er5sFY1X69Z+QxibSKRRcoVDpus2jjd0r
e6oxEKQpIjCDhjiaWPJc4AAp8I3JOXbUUvUe4EYBrQP84fLuI8LuvAHoL67x/mpI8v7Q8dRFYtaV
4TC8iOEhVq22c+1vwrNKCcBDjSDPD862rJ6NGSFZJnakTPGVJEpRZbQZAxhum4jOJ6SBJ1Pp8xPS
mbAOeSCkhft10vUpGfQKmKtn6xp8Ugu2gsqHGyHenOBBV+s841XCunPMm17Qeotfk0SSvSZhFp8K
ps5XAZU6oSTcpOPMag+8hKUfzw30XyGXgniH1vMMyCyJv7wfOmRI87OKZt/3FYpJcfHm0u2a5xFd
vLQBDsi10OHgMshm8lKG71uMUDV+aopDQsMElqBFYR1LTj7FIOX526N7FUtXKoRZWdLbwDWRfwZR
S8QpMpE/aKkBfvDH8jUU9LSntDBfeuQRrmkw6pLxbSEFWNvlK96i7q5ob6uTzuf3vLgIyHmINBmJ
WDv8VqWYamzoIXqx0dJiG0NUl/tdpYnkgIT1G/p42AXEfxubuMutyRP24O78DEHpPCrDTEGLUNap
rqMv/A6c0yw8DMznRmjQukO3BS+lATt2MspkiKAuW2yXdCAfq4Sq0y23jxk/BkCGod88YMl4BJM/
zEHlrG+yqOpZeE5bbdHyAV+DFa1/SMcqNlhXuLODVma0kokB8jmJTBLFbMvXsi+dGRMZyYC9F6an
1aixQDoKOEMT37IZDrewdCOmULczXMfTgJyWLgPEO2GZ7pLfudaUedJ7cBb74IDeFRoaowqFLaze
8/Vlvb3accVSRQbsrfZJgz86gSP+TukuD1FDNGFbu7BhrMF8+Ih6rjdA32SN1jnhfWRc+RV5Tml3
UKn5yM1O+3fVj+j+MLmeXfWqvluuPHGDq7MdwQ6Rh0hbD5KhpZZstu6sXaOqr21MNEZBIcG8iFof
zpw3keAC47fFLz8YyhcExBYXhGsB3kT0JEDUEzHtJzQTg3TPVXKIynIzLBiCKminWrWOynP6tY7u
A4voi6I2oBmeZGAOg6LWZhB92c4sWyC+LnVMvcwceiRodNl6Xvv3fSMTUHRhZl/KLKtQcT2YAOVm
T4082o1fcBdfRaUbh8TUsmRHhnsn0LIGyR63kR6Uz/WkkxAz+K/Ofe+i8OIU8VJgRKrh5CKBFU9R
AXgN1XFBozaxubMIWbqfmvcuJC5Ft2xTa+g+VCK5yvdQw/kOJIrjHxilZi+02GnODfdvQdqLq9Va
u87JpSChiIzXzCm0mXkaHZr8WJVl7gfF7zDXg8k2URaQGfgeTNKDhtbquFjr2qRcyo80nOjBC4Og
b3UuamfzbnqECXDQ1Io1vYJkNFbkbsk6yKXNQbY66zFI+WIfdS0E2iPvvI1PgKT8HAVcmzyesqBX
chPQtSAf8UnS5lhgdrVToUn7dWAFDqtyhkzithY9/rOD4BDcxPaZTj1qA6tWq6JVvJjyOLrC5bpz
pd4IMSvc21L+PLL1UV7aYxtZ6oT4yfdOthuqnxJt798k3d795KGkHsVJ+Yx6B8jwkOiGriLT5Le6
AzH8fD4Gp5bOhKZIG4+A//FEPj2ZBW6iPiUmxJ8UHncrQRfp1a0ZaBLUXV/7U7QbkbsR1lufE47d
72hPOkuqf9E9vsoD0p0D26X/5I2qeCOk0Z/gvN6yRF83Ni4bnOZvwjeY727I5Mzis+x/CJQPBMJj
4v+AT6R/f/mDY8Dy10w9eN1XLeqxeuU2SOt3VgsswkLCQQzqF6anjlVDSG7A5lOy/etsi7P88His
0iG+12a0VyH6D9znsa6GFobwEpRtljdev7eyfvCJdkwKAqI6YAAlfd6cbgBbR1mvMnHKImRPToD7
7l+kZCwkU4Dy5MBtH0Zh6Jj9K/o6mv6Q0HR8dLz7nSqzz2aS7vnutEZFuKJukQh0xMb9/gjYeN8L
fSkoo+KVOF7iPWSgAJ0a4kBMAipfwMEJNBOnan/GHQadSnsYz9p95Oq9hwa9+DGC//H2iYS4FHQb
fNiGVSDKjU/C42p/e+De99IERvZiYkfbjNUNMbEH1huHUQ3FcEx13dH1Dov2K1Z4qXt5rj3wrNZw
TAY7/0ScQXaHhEN+/ZknV4osry+oUVbtFFGjg9+XAGolaV+NrkFjTE1wby9X3JJQpQq0B2iRSVJD
k8Aot4zDxGRWhwRGTsjLuumzCpPLpVWt1DV0jqRR3eq0ioek9yC23Hj7w8d7KsTQDyzZ3H6jA2s4
juiyhuVMvUE66WHKSNrMemJ2grXUt5PtEx1hZE3kRn9zVtmnz59KwkGcIqQ+xwD16vKoH1wWWZTI
3zSlrv7k92RjuB7irUow4OkeyyVoj5W1AuerW1uH4TfJ90k/8Gz10oSoeOvUPAszsesbepvuz4Q0
lN6/xTDHdU2WORHjyannxfKBThWOOXIKJpj+eoZwcBnzJahvy0oYHq275Ur06jo2Jsvx2ofevMqG
72vthb6irOzaiwpzDCZJ3eBAkMZN2RqbBgEYmHKRM7P8z5YIZKFMDC9isLpjjjMtkn/HCHH8V2oV
oXjT1ppr8O19p4c6D+5ic2QgEe9K5T2x20axDjlNJaQIPdKpk/G4BVPnqH0zX8RG4UkCAbyuaDGi
BYj9pfZQcvWgnC+wXG3T2BjZgpxl1f8qULlvbz+32O/TM1NGqlNQMJyWO9vffWHwEhZkuqWOGFhy
hjdjnKbHRIUAJ2KpQvUrKMXv6tISVPnMSMn1DCc3Vlau9gpIZJ4gsYHUzgKiNkbi2HC/jw5hXqnD
x3PeuDiw03eGr2zQCHpCnNIG1MsAhD9DEio8fQqZ0dP11V+OY3x73kPyiOeRfZ/RuzPEtzr/OydD
3vPVpUzrXj1dSvHbGHQcex4hhOISwV0o7LNqdlh16ZSmvyRIPrfeYD3bKann1rRCroAol9TZ721L
zwLn3gtpupOxuFLvOf+Ux4jsDglmKDfNMpNI/Ig89iG7obg4L7tbmPyUJGyUKpegdbvkM3Rvk+8p
GXQpjyZGWnVmUu6uECsMLZPHjU3IMHo7cXGrdGdqa1ThTFpG35cBIpQlHXSBkT+UHzWj+E/24oE/
oXsyHKlK9vl3vYp3PpT+FP2zPrqOCEIhJZV/gy6R3hEnUKLxIQK23OAjRWEwj7KjVyc/gxBtn4bc
It3hq+ygOPQeDVszCLUvbNI4J9++T/ePKpyut2lVNtKowJXQkrpWIMTZ+43nSt3aInf4EqlnIIRG
vg7Fo8W/3OqGzG28k2nPF4nwYEceEX2YISwRKFvn8rCgzbV1YiOUwh8Ak97XmJ8yunVfSBTR/Y6Z
BKkinZzNqGNxHrwWs+GRK6f5maxNBuvpIGZCnmJsLJ4g/0ND8/l2OAv/O+duHc2J3Qk+IGexUZ1g
dt41yV/8OrWXY2/vtx68Xk0X7TFkLYl6Tj2v/Z6yGExg2FvONsVBvXSEk4KEIb2daE7/iw0UqOWG
eB+z7mMhiaPoI/9i4EZBrnITCm2g02L8rppJ2O0lf9ZUs2nUxCZ2A+pnXecYFfubEHUO/D6601Z4
3lj2GfKvVn0CTY56xckjcI9duyRFU5Ox0a2edujri9eF3vtNGfALCcdnCgZ4raRy1n2LvXvBQjJy
CCiZwQ781FNOPchFpa3mNMnGU5Mj2bzXNwlMu0QlHsD0ghO6E9/S74OAJ/eMUC7vT8jscySLup9U
ayQ2mcahRvc8XF2GsHtEAUsokh1M0KAtCWm/7YjtMet9zB8RpLm2BQBidYCrJwisQkB6BLYP+gtK
ez3dZQQ6OhmyLkxE7/+xnULXbtUuSwVEeb5NWEUhXWFYo4hoZgcKXqZl1VAFooWStQ+3wtFIQ6UF
8eoE4MocAo7WTnyV3TSDuv6iczgMpY/z8UY/7m2+C5NcU2Ah9jrr/BTrXu72frKoMQcKrevNjDe3
Dih/oHE+5repqJnskjjc4keNFtuCze2Ig7x3RHtTethxr+5+1FRPJF0+avf/MynO+wc1lR3C0ZSX
VNTcQyg7gEacFlX/MJPVj1xCQCyyHtLJBGpKakkKaWBS6wc+VoA37sEgPcGcnwLtAGSq1NkvIYZN
HqFIjE3sLxmdJlrZWcNQnwO+O2k1YrkV9pjQAqYwa+rpSd98XRxBs0Dz3nW0g1/xFjh5hM9E5IdO
lAEll0sEEvGjBLozBkWwWqbEcARMpe+i/uNw4six8rU50s1gjdBksQHz00SBEuu0aF+WqsQYY0ZX
72rjawrK3uEFRnlMB7lX0V/J5PvAngMY13GZegEUCcCc/g49b7nqbQH8/a5SIua892rkHmW1Cxhi
CnWsf5dAuuJppMoLFxLDQmnD5OVqLomvsU0E68SFBaGclMFxgVLpWJC6up7tpEWvXOADmTeBtDDV
sQEW8xr/Yj7SyI22jBPx2rGV6yxHSfLi3pk1ImgURyG1zNfudfTglf+xfzUIR37d4+E2IYlxUzWt
Ceg6aStbr7myN7oSgbbn7To27gMVDdV1IYHX2vgM4rVYU9K9HQZ4XyPsoAUDk5yFwnjnKJfRJ6sj
RgIhTXSNjUzr78M+MDvVeRRyi64MlFGreiW62NEicwRxLnwj9enIjpH4T+WD+LgPzQzXMWN7gHUY
Ga1Cow13W8PZsYwty6cTJaKstMhya3u4rJIc3tAmydlF8TNEk383tmqkTp9A62Ehw7UNvdJiOxfL
1hw1GYzrSoBQ9OuSLy1jWr7cW2mLdw0v1WZ7IpIS4IV3OCuODNPKzb+d4xnp38y/7isTDS/Wg8/s
0r0+PDM9Wkzk9IJ+RcyGs9+E6uU9gT3zPxiYdgNv9tbcmIa+HQOnKe69GT1OSKqIa/K+ti0tYn9G
DUQRlFgt6Kg420Frc4iK1DTjHlrcn4CoGl7+wduLZNiY7pMIyybTlAiEovNSPEFYK2Peb8EZrM76
I21kxWSGsMl0uw+5k3fdWBUoMeh/cbpTWg32Yv4BTYZHICBiAXqpoVEcghO/G7qwgBhFJzSLDjeI
qjQ7SZC4e1AWjE8BPLJjuw94Dc6D0oGmfsYez4Zt3WWYhBy2iEG8boZjhhfKgS14/j4RImShjmMm
hC3YfAKIawRzmD2M26fsIKd75yMpD+HOLwoQf9MBUnf4fVazygSPy7QvNmPhbCueKCOMPYxO15Ba
OZo6u842gbzKHXMDi3DBSUmryw13tINpx6GvvPik1gczpEA1/H/2KZp7xmM5JpdKHAxQdWtka5B0
pjXYdp6g0CgtoD34S6veHGrLilHuCIE2wib+CN7qRPym54FcHv44vUDQAoW5hSfCyWdYzgXfNmwK
blPm4lv2AuL88yDbyRXJONPX0mimiMkRsTBMHuZRFDtq9rNjMSosBKYCB7ELI9gyTiPsEY5QoWnJ
ufDIgvwz88ahLFGiQruHMRq7D2ERL5cZTTYnNWL9TGJfBsKZfSrKDdN9/xUF9u/rdPKc2DNiT1TY
69qr6GFw53TK47zPNuCF0VvtgtPf1j1AoUGfPJZjGdoiX+DKC5gMhXXWokzcnzcdKdeuE5Ssm2X4
68uq2MdC41wHHLmL2/7fnCwmx1+zq06Ij/XUDoUWI8mH9yHIHdCEM5uMpGMCFaWpWEi1uataO4jK
YuE0MyQhoFiEjCiM7Wh/Cm76Ek6FvMm9cUkMVgMM1dnwIiu8MUk5n3OC2q+AGvN7pPObxHyiP/mX
SE+hfUyHid+/XxpKgk+u9DoRTFPJxIzP28VPMNtgNo86o1MLiOzndHdLYHLYQmxgElAOVGalyIJR
TtJ+btEbj0NNh9IBeiRThkOg9inhNr+7y3Wb4krTYiUPgIXkDLlilHd3yOQm1Ro5UC6jhdzzE6FB
FEmYgagNkSpqk9wvxbNM9l3YpztDEfxRLw7EbxAdUN6cC7sZpC004da/Yp8xrDtgjRtQXHW8TLa9
yPMsw7VaXYQpPFY1A5lvT1GKej0VuPojiqja8f3BiIygkyVoZe93/5ZHgR4FtjZt6aT8HIv7I2G4
vfZs25rRH4tO0iiBCMdI2MiQiBkwsohuKyA5Tbowd66F6V7ptt4b0Z6gIaWfdFeXAtizQ7L9rw9Y
gYssQJuRvrOwnKYINZEYFlpsrprb+izzJA7+NPAF62AKo881BaWJiERsj2m7hYq0wlawXdq9E91n
Q0e5uz1vBkteBKZ1SERvy549a31ehcXPCGbcGo90d3XYAEJbdJvUV6I/RFLrOmewI/bWIqWJezNz
C434aRPJgDC6wSQuDOSMXV1Ns7hefjnw+VcprhX35Zww1r9OmlXswE0FQlt9Xc5Lp5KDeKC8zbVc
1XZY0nqdMOeQOmAw2v1nKiDsBqYp7e2I3JH7KERd6za3dBcKdRk69pGb5cm5HjQK3E+48NBA0RTo
jPHNJtPxMd6jSt5aWpWcVkNCPRsF+jUb8kvlZsb+gs+m0zD2dr3zljj68VIKcU9gZeA/Id1nnIqB
ba+4N+KE+DkuAeKS7rCasGljy6MvOkAsxL3Kodxj3pGKR6X6rwy2acyBXEW9MdHZmLDIaqq+hg+H
lhug2hrVjX9LxU4F1OJR+3IbwRCfIWudu0+ghSkRs4dXOJXqutGEHkZ78Rc+xxGPS1rIw4tFFb0q
tpqFTM6gk56swRNfjwT6lTfXco2zBafv+DIFVTwkHWgD9/+nT/FGtwWrVw97beEE/6FAuvYzDvEl
7XsvjzVmvcZZcrEzfVv7U0vZEsa1OiD2YBudwwcRS96JOKx8n917su6vE4OBZS+XadWGGES475vw
W/m0iKEE+yVOinG4I9UCwkl+hWjAYYYfS8jQrD8Xla9CSiY3hM75d4rf+/7Xe9E06JuswyY6Jg2A
0QUUHo0E1a/pK/soYTEFCGcgYXRWZ8p5toM7o3rDlL6pgWxwxID52O4JaSEP4ZUY7d1B/yOy+pGH
V9VJ4S8UcoruwL+1ZwY5s13Qk7sbptdh4/twZpLCJ6IRBA2MBIDzJsmhSlz03Vr8IN8u12ZZSYOF
GRsvJaeCo1YFjcNDZt2pxKADxBMCLj59S3P+BreApgrxOltrQ8BFWoHuObYczj2KiIF4nGJlE7yE
Qp5579gztbBVSe9MmPi1d+D4R67mv2FtI/QIufNGm8WUJSIhiN683rPxhjcDbhr0l/3WSMDHON+W
BtjEMXwezELYZUMXGnYJpPSy+O8miI/lNckvK6dfBRMDS1gXivb3Z5bnm78Y6sIWqEhqcntRrjGI
c1nUYr8ajiLFxOfBxI8snMxL7/qON9udEaCPnhn1JjceT6uLl/hOhcqK4tIS+GbLvrUi8WQEN+/S
NHfuTiaJrbb3XzcdtTQCp/Af0JdHRF/Hgk3kPZPxX9X5/HIk3t7fNPJas6BXSWLol6GYVEzXZQvr
mstF7fP+H0wBQI3EpkSPLUQswGzaUddX6EnvqU3DoWxl2FxvE50H4/T2+KmZ7dsLc7hUq1+7w6ya
JR3SHWOBqh3oSAV2I7YITmC0B3eYKSVoJnxCFiAFkshmaXOIT/QpNkEH9esQ9tg8FXO91a9VOQLU
hROdA+SgC9bCzwPXPo5aBbHyPwMIYmpKKKmWy6qYCR2VC3DbEoBILuDVTa4A2qIn9A2MgtQAMeqE
hz/OR0moDEMGi9FmhCdLkblkwd+i2xQoijlgi/QrrKPLXXozpXyjE/77nkGq9M/pdTsWLkFyiHkr
OI1QShTSBH4bNt5if/d5DD33kTFSj3lm8EDCowTheBN8ZSlqTf8E9MYIWgw9gO1SPKho6Bog1Ku3
l1GHhh/ypn4BuYCujRdySNK4a0Dvf0aC83vd9Nospk5fGUj6lvL2l/OT8o6DXXm/xHwjeLL7cH+7
6NK7ajk1urh4XiVKNNf2rMDCTM9mu6gXwSdYVs+C/1ZrGHPFDBlUQdH4wfwp6CewImccuYOtALhZ
0y79kUBhq613qo9IA7+SZrmKUgvuUt1fOtOosrd+G6w9r00qlNdEiD3WlB+Wglaa382QX+gz8j+a
To6ogjdtOftqX0R4Yw4c2E7efM+L9RBjnOGtuI4tPUkw1rS++8u2DNXXX+wKmVqbNhrVb+vKD9iV
+AUrq00PgK/VhYmsfwmxL1JRXFgxiWVT1XTadudku6Gd4WWuQJSUi7q/VtdAvFx5O6/u8e8LB57n
Yqen0haxsICZIgF9TId0Y4Qosa//cggoJQUSYPkl1L5pr2uupqjnjbZJmz1Dcvt0yX+J2hr4nMBu
Wur0KNnG/HSpU6mSg/wB+pye+z2ph5Nqftl3XvjjK6Z1t69fDgMkhAlVo8EzL5eNP8HK4XCzvsKs
nQgHcioqLRRvRnbIEe7tMmB2I2C7dJZzrgk2oR8P5JHuCXtg+Spfq3d96cT0U/9CZR4Hl3KJGp2V
vMyeLqXFauOK7eUiddoZddekU1AEy/MTRsNs+2PzKLVjLBgoOnko6AOJw6BMridt6OsjYCzhWjPW
YleCe2AzHcX8LOz+mMXFnN6eqD+WOxws8PSvP9ekJZ0nYsV7sxwS9pXn/Ci8a89eWdBH4Qc53JRX
BivwaIrbWhE5HWqwzR480E1lilHfDddUEJEJLcfF6AfCEowqKp5q2m8OxZYLqc0tZRtHtAG0hEKZ
UURqLDvS17LQi2t7xtWuRE0oA0oIWYZtULs3t319SIGuH/0EdR/jOg6vV13wNbvQv4QD7EFatRGI
iL8c6aMPTCfNQyyML2oWqx8k785Ve2ZcFAeHyXK6StRbQsfAgWMZoq9vH8z6bdYuuIFGLKM3/tD+
SdvcogXz+G+V/YorqI752cQNIXWEB+sBq12GbNtG1Pk4J9uQqpUV0knfgAmnRwLm+1XLHUsq/e4J
oWPoJD3u30W6fQYiWXCbE+AkIOCtQR0mEjWhp1sNkSxuzlgVR6hei0cEP+h0f3OePJ5KyY/A5BLx
HpbVfTe9WTXj9bybKH/d+d19tHn9N72MRfW+D3V5p66XuVjvKQe1VTbJuu/9GHt4AtaOwEAxRysY
ZdYnpblbO3D7u/F+JQHlWNYaYJ8io760yLJWtN6q1OxxrN6bR0OwGcr1k8C91OBN5FuNjJqw8F5d
ETf9wxekSo98YZnVuZawwiekKXM0dY0TOaoE/e1mUO4ZyIAyTnblINaISc7p14Ah0KO5yP9C1Syg
h0NbK7C3WwEDW7154RcuikV5XEVpNuMVM+JWlnBnycJlRQMPfrFzHaotzP+q40bnrldOp72SF0wP
2hOo6ub6eAFq2/X6InEdNaNIpM5CfNDxwP4yJpzhjJ5U+Xkptc/rmP0Od620dXvFNr+t08Yht/RI
ooj4kpa20ZUXq3P/1RenFmJyiElZOHbfJ0uu981h/ccuO9OzPE2stDhSNI9qtR621NMYs88TVxm3
ue8YVy1PqQGZmJfZ2TL2jUvutND+/AXbbChDl4aNFrEF1lrXZ+gqDFsAjwJSWmlLqwjXkO1Beark
vMRmWOshwOrtELW99Sq3g/I/o2KiKl746tqB22S8z4sewXOEt3wHH2eVZi1bUski6hgoqfbfXZC9
p7OTPm59t2aL04UddBKkc0u3Rgja2eclcvKJMUIJ54ZEs1Bo3PLXGsT3ccZsmgAImH8G9u+9lmeW
gYBfSrflP/5NgdNAn0y8vxHRTjENV+ZEwxH7OE4cYhXSAyVIHhBnJMR3dQOSQFrbHOBy881a2u0G
MeodDJafEXYZqxnBY0iCYYzz07jCDwp3UEE2zmOtHFEowzzxaKNWM0qHBFuMm5WPuxqhNUb5fQHR
oNrIoEZLkWfj16iw3GrNvmwvVLsnOr9UtTu3AP6L91Mz/0saS3lIJCnMiNqWlXBJqslaOtxPOY0u
oOpSK6vOGTXnir5JMD5BThtJUVzT/yUlIuSCsbX/SxEVQqXUmifBPLOOw2dnRI8Ek2QFR/mwdJiu
CVaI66r8HuvSpQrbySCMtVHRPOx+gAy9l7ZL9JPShWFj2uyKLeOJzEcxZcHTuGxEYJxvQhvp4WeJ
E818O7A2xAzXiI2qTUVzXsPOSJ/JteYTj2DAWmE6XNtgen9U7rm2uCVr9J/oMu7jJ+hS9DfHmEra
j+VubgrUZy1zkoPwRX8MBdhBT4+KCW6aLhuzdS7CVII8jo3OMTdg0YHa+QAdIiyDvKoev+O+ekmp
U0RPDXugYzPOnhcbnJLI7kQ9wr4VpKHV9NL1bSrijtuPJeTvKex0umxdX1eQaCele2cJ70/QF73Y
xLDDjosAcn4kQIGzwrKhfD9Ec4RH6UpohTr1Dj9XtCcHK+hpn8QJeWKW48txflk6+FQOVrXSI4Du
+9UX5/zMKsPNhb9q4LygIIZnA/qvDgncZAitHoyPH8LS2oNBXBmJd1WLi1xp13C2X9lCEDqhJT3R
wwsMtD+B22LDmzTtne2d8e8SebDxryGRmAPNn8oMyuwwUU2Dq5cEpV2rF3VyvlcNMMpcXtT/qAA7
gtaM8kNTLKN6xPM7RyVJE5NqCecD6hvxU6ZKycpfTWXs94SxJmd/Md8dZpbqvxgwJF/GNivp2/lw
bJtoXdNEub54ikHh2BT3k/p7Ze0x/SMAsA9zEaCrbddnaM1T3oywFP/3BtnreRb8GF1s/qKPRj/A
GdAR5HSyttGAU3tBJ/44KLWWB8d9JCsZDGgQUeW1ZKBSWesPvgDrMkoGwuhFy00pwTGTcOGWgnw9
SMuz4G64FrSX6GqW1Y4el6RGbiFyRu7t+Gd5GWeaNNvByyHMGk9dfi7TXwZI6iNfZCjU0dA6RGC3
kk6Ie2j/VrBy8gRTWw0VPns1IyH/tH37+eTO10iP99c6okMzZon8pAwIdFRTwNz5XFJaunmogyJn
la6p8L31VvbsbQ1HSLORnzy9Ub+wNu4oS4moeY0ee+jjf28HPTiQ8hu/VBZUIVWZ8F/Cyt9M7MUs
yKtObTV8opWKq3P0CBu4iL7xyGppvEppbk/7OCFp6I3P67CnxseZxoN8vNVCYJWe9XMK+AA+Q6K8
ft0sX7xYl3uTqNg6NO2VEcpfBajqoiIFSxNWZSE2PKUxsv1ZUyyOIIG8OdXHSLpc0miD1K5HyLAn
rThTJGU5UqYiIQvxHJiOLuDox/f3KTe18/J1NDA1ccuHw945nl9VP9wg176JDgoV2vxwj1pJYkat
a7yCcG6xloVNsRBHP9bTUQHYMjWbOTJXK8zAkzIfK+8c9GQl42k9L46LrrEy+Yjswdowx/bnuDsi
iILlehwIj+duZ4j1F6BAmJ1npRpxakEgUNu6qZ9TOqh+OmJHh1bSTnfYBg5IMIVMmQ7uXCylvOhM
nt/elQQY93ecUlxvQY4XvuQCpqSRRRrv3tpXtlDYX0GscSTgjIXIlO7DDzpgIRxy9cXwh+PVxl7F
0hwtqsYgVo9Z9jcQOBwvfuhWzvPc4JU3gOFX8OdHJZqL7RXUDOm+rsBKyjGOh5pBgrxTPa270RLO
SqN8zROrFoiX7fIdXjv9WMVjVCyJN7pM7AUc+nu3ZTx+6K9D1a6su1z8EH2S+9gmFQS3E51uPigL
WVE0iTULD+S409w0VbVYhq9Gp/j3cCPBCat5xcNgdvUfoHDPsQHEsDJRqOVK0gaq7ksxdLzVRMrn
bGAUscmUQacJpADaIfVu3s8GrhF0dRwAmHgU0ehaioVrL7jhcG9da9ABt1nRZEP/Hp+QZ/1n3RQo
BrCNrKbozBcIPX9DV7sgPtuYDlgqHQoA7V+6cUFB3T8Iyg9Vaw8pnaq9c+FWnK8tdKtOZ4msd1ts
TPpcRWi85AZZRuOOUtGxUvGo7Lz2YPfX90w1Q4DijXNjhJnx5oC29cFmh9robvd2rmcO6LJ5dpRF
hObdz/2/LJnFr1OdfhfEEOQzOZ44U4lrkJjnUzw2uT2szaxcSRzAqeQMS4s0osF7yerMeXMJzP9q
y8472tUDiwhylurNnGmY45YyM1DXdq+oJxF08VOesg9TUDF4J3lNZ1GOdMNZtvF5tpIueWRL6Dgz
WSU3UKRhZYtTkFeLS6ZehUt24Q7aSn2GSj2HavZaXOE6r02sUJ7hLK66v9E+3mhaG6mmEt3ZA5uC
znCpQVpjgx4QiIxkG/ZN6xeIBBAwtwcsJmg3u9awBnLKoUkW1fPSzmv4LlcB2KXBfyOP0v13f+AJ
b6o6Lm7Gzc+r4UlyAckNxihROrv6RlZ14JWcfVhGJdFcmitR9+vwf9YRqylxKsjVNuHdR0WrGlJt
z+kiYbI/Qm0HTAw6AL3Neu6yEGcmsT3R58lmZGdaPw/H3lSu++CxEIvnJFoYnrgGkRLa3/iUfO+1
iq0phaoloIrK66DUTS/cq1Eb9BJ+SQyonXiafbtT/mACxKu3/etNn3cZ2AWp1s5XImaTDBHky9un
q0hya/ZTuuieq4HvuOE751ZOjhSZoY1CiaoZQmyREkdBsVno0qpaM/O8hwC+vfhDgwig85n385Ld
/28nAi59Pm758z3RRrDoU/RY5NsnznlrryTrfCjcsxHZOmrzrwgnnTyKCNEiLcVGWXdpDTV4dHhW
slzERMfSZw/fMudtrTeNlhVSTWLEJ9N9BCHc4erUgwIdnz1Il8TCrr4lqU4zCf8d7FBIV8GKFwOs
Br0VoVropMhBFzmvY7TN1YjO/6Wj0hpr5MKSAlTLoNtseIvmmW6t+Qlp+nIHY5KpoDyd5stuYlpo
lDAcjOFybVlP0tK1PFj0lGtwdSqAo+gP0ULtqD+Z89XqjFiCgUkJaxWsTY116OZkeCV3mZwMBKSx
N07yltLgruJJAHIn5rxwgW4vh9giMKw5KGF63Zj1dIcq3938Sjg7uwnDxBR84Hlm4VouE27TdAhO
WBPyu1cTr6Cybb+J9O27g3F9+zNyNJCsoShA1+gtamid0CnLQhxm22Vc1coMXCruWhZxVPYAS3V5
D0gyOghDp6HBcxv8dF7H/G8gUxXSkyjKJrIPxB1m9UEJyPYMa+z+8+7j0xPdSWHIumGDKU2eSQZj
HknJV4DLB31SAucdSHGKFbALzcP5MHR1AcNJ+igiucP5KpXA+0YNTqL25xmFTguINYUCPSBzZ8Ke
XEowNaIm1DJB/Su8gS3vbthXoyRI8K0I25fRlfSVysdwgvGVS4/BP6OoI3eN5+NkIeOJLTYL9byy
X8P2fjwPGmqTcwbyeBbWGgG8GpY5X6CsGlglSb9iosJPyNxBUPe79YRC6ricqZr++1KFXaRLwSt1
PoOzvh8NBIwtH9AzrJwzEUYh93t5dakXzNsPhVXze1yG9rB3+XeRT+ZOLKouvQxWjCYcD7F0dqc7
+DHpZAZKEdPFXM8uZOBD05Etb+hLHmWRB7f0R/ztJMtG3LaOcZjtt5RZTG5MNkl2XguOFX4iCvEZ
eoOrDBMAUfABOTX/LZkQd3ay2zNxkd2QHP07VesKBsJveBHfYNTcDpt/l6NkQNV+cECDF9mr0viI
C5uHE1l62sBq32RXZNwYFr5Fybk6hfl6PguFj67KYnd9Ab7cGH49oiP2Lo7QHPVQ61n/07EO4ipG
f9u467SxrzSN5X4vuv7pvTK2Wx68+GS4GHZBIicehyYeuMrXhjNDflklF3aDtEYOLCqPSCVWW1nj
LoI/HPjC7TrLgynDNjB3piuaTUC55pNkNRxePCxlaUC1Oz+7Pxw6eVW+H8uqQe/Wskg8YUuB+hPU
PI3ljfCtIC6tkb1tumMdNnHPKlUaXLwNXbTWmVwDheqh6y8UnNTEgWj1wE0qt5kR+D4Lw6y4nL7j
AeVxsqjOh3PJTX9VMw9uiUCBEQnI/v+2zXPOSJ/ECdp3e81JvzqG9T94r79Xh/Qqt0RMbf2W9NlR
h+xyJ9tsxKnsCcHVsj2Ww70dsd+D26Q2VNBCp0QFdnCOTe6bGpQ0QsQD6o1aL5Mg343NV1MUBGQD
xCZuTNrjVFa7OMM5CwCIDM7oLGGS40XZyxxTfdIi80oYawvspHtLW3HnqVAiFsC7nm72CCk6jUr9
wR8bgg1lsQZ4Wo/Ockz5FzePhcaBMmQL54PEQkrS0SoF6N2w3hymfJo+2KuSrRiaa9MJwVlB1xrr
5AYoSSsc7TIOBBkzXrEhbxPEiY0d+qggt4FeSPnuJvvA6cOAollRCY4GqlmMbvuJabrBevXIrLTc
qdp7oo24Txd3andEI5JlOCToiObVdNzOU7bCvKb2XHNG5tqSCVHh0/HTQt+A1PVHi/H1YOAbCQPP
7Pg9wKvcMZqEspKAOeS/xOHBbSz7AJiXgw3j6LkVgJFSgOzH0EBkFSoDPu2FAl3AGLbpgUeGCmWB
aHvWbF7GOqqZBLh342T9c5J8O5kYcylrezLTqViw//AEkpdqWJf1EQf2BXNSmBSvLB5vvI652xDt
q4vazd65kXwvQOUv9HaMYDcfvCapwtJVQt/Sbnaq76bgkQ2jXi0yPvKp5twA/qegUkW9MqE225zC
/ivvIEXrLF9woodYGc8hb814MZZ9rzo6CXFG/BXSnx9FgIkR1OFirlkq0ABWcR/CnTioScrAgHAh
90XfTYz0fBCXTG5gsX1r6Zwn00vl5XMGJcfP5ZAnTBpD0zR+UhhdVI85d+P9Eh2ufVadvDH//iK8
QrHba6zjbl99vdWpAKTr7vC+T9MtNZqFUHxK85MppTNZcZKBysrlmJwOLAuTNKwKlEpcaSfteRaM
gveaxps4HZdwDP31RZkFVy1CKVmTICftVgQFtMLske3ZyGmnZDznQNQc/Vf2KITU7Ot5+8rLtHBN
qEK+/4lHasQbFofcHLKykmZi8VMbL0FbMnZDGGJn/Pmk4KTQAzqCE+JgaajiDzN3FhmNvhB4wwzi
hrsXyv0nrgadQxV0g8U/SwZaOgSmomtDakf8ERY2KM+V62VsmZjvx8Z8x7SRsewjlPpe4LkWLjI4
0tIYh7vVusOW7y7F8DVtCmEX1UxvNxe40/LggQC2kkYUDa1GUEWkcuwvblo4kmIbNxTPzpIvtIbT
XKU9YR4lEB0g/5AmHqs7EThix3iLatMB6PDrTKHKmdy1uTvX1M0G+xbhjK4ROj8x4CgS315/quuM
gDVqlAsGwadqZWb/c4DKxPm+VQQXkUr7dbmquw9iFBg0LE1qLbKc4vMBCoYf75XpRsLAiof6ZvU6
gn+00+QEVApDPheDwGQ/o7MKSZd5dbRulLe0oH2IUuMEaQBzvUNE3a+/IK3mSPI2LSjYMWZAyy7J
rXBMdTI0YJkWZR/hkMDMmnDBNQarH9dmigxItNyb8kVfTJQzwnvH1JshCNScDYdzn18cHer7QKJ1
zbjfn3Hffy9boRfDaKOArqRD8g3tvrAVEDJBYqypZKLXEHNGXV70DsWd6pz+SpWbTC/DRHFQ3K/8
K1wIA2MJjjaoDaNvGfe2p27C638u82SoWHG0nYbi0391XTfVjAfARHjhlNlAwE5+lQmcH58XGq8/
LnglQnhNwC7pcfOkPn6mjWfoPZGKuCYGPjWYjZ4cDAfByIDnq2OR1YhQumPOYbSALHv8RojD7pEr
m7SLmDVFj2/+wndbbOnEiKUmCYCui5lJ6wVPoVtInG/JfetPGSAaS/XOgUevJ/NIGN58avlLJgOb
WTK7+hjedPEfHY/sT9uZmw+ovRaLJlKwKMVCPiTUpVMSu7aLOqkMsueaA32tvPalhxqcUUe5cKi9
v5MX8JY9Cc9Q3vQSfFjHVDK87coSUgAtIpcbDUPxKdID3kNFMYYwQX5bNP8IM5zqjlR+ZFe6hDaX
1Wpm1XX6PahHn8pL0uSMNDeFs/8t5TbXzFLgWv/tD0UB4lZgT4aypuyY3g8s6DkqIJix7CEvJyCG
s9SSN6tQjf2fKlfYf4k6mmjajalmjx2j3bkGnPgdFzw7rnWAvLC1p0MEi7juqOLhTKObGMhIqkSf
ojTxbNL8V6P9AW8PC4pKUCmKoHz8gr/TEpnTPkB//eTHWisO49JvzfL1rP8R4C5aV0eMx+SHELd+
K59droWUahylt/gIi2THgxF1X/dc0l+MIiRU9sotoCxumjLmHY2GPV+F4Covf1l88v26IdX0YFwB
MzL3fm/z0xyrdp5klpdsCa990F5ODdKGUF9qB4fo/Dn6CFiXjOlZI6wf/FdEUVDAVHL3lteKCeLM
aV0Vux7+ihwJfW5cOua4hNN2+V+v4tUBIdTCshj1yBMd6Q29C5rsaNVzkcRyCnJtPlCKOdzzKRfH
GPjIOZNWiex3+olruB6k4ufdXqaDwN0VM+y/DocgWYLwJp9BZXxfekA2chooeVPrVX0KHWa1uGcX
vz5Lk1Vnleu6yP4P76oSwxjdfLlc0cn72GJgPEPXjS2H8tPHNaobG5FFNv2nDIrPjDhCDxD6sZD3
KeOfsFWB9GX7hQ53X8g/EwzB4cLPCuktx1/BWT5Rg05dm/O48TSQOaSaUE+qF6nLQDdLUNWJ5Hih
nn9zAJc2JMzTvjN2lbL5AuZRr/w7jjmeSMT7N/Y6pC10b7KpIxdoPierf6T5nsdbzDwVECw4WuYd
7lfUSuqtKrkFk/OQu+S9Xp2G1BEa1KGwfDQtmfFVDUwzk+k5hFJqkSrNsDWezoEf/R3NoVp+VIf8
7RyZPEUNmXwS6qEoUvW5iu5QhMBn5vMC818lVv+tZuNLDXWcrAxon5xU+3IptA7AQ34DXwRPZCt9
4FIE7oMKRoWuLoxXPu90lXobQwiZFCvSgZP7JbvcR3HcalDc2ztHVKdQFhRseXMhrhaae26WNpf0
YZlIeaUlBGqOvO50eZYkVEkvgoSNdpQlNLCylT/q+iD/hUCVDQJb3HPA+i5nYY9iw0sFQqdHT94O
qG52YW9U4DwPCtXoKkbubue98/MEO92D76lZSSDVsVF1VUFLZ6KVblli0yqX4GKAf2mKVfk7nsAQ
Ki1HQMmOYDHt4nc0oVgXGTo10qJ+g+hNtTQeDq6DtUVSJThsXOhLLWKCXhMheF02ncBbT8rqhOxY
UxtfeDqGsCpLTPryH5WrWXeNOzb3E3jbq3FVsUsEyQZC/Ho37tQtUgk9BLESbpLuthT62yL0gJNH
eEMKTHXJTXawfekEBYpZf4UPnSPkRTu6nDQrlYUiBhX7GM/fqRh2YQz5f5f3OP1ZuNgQN86972RP
vv1q2Db+HtEh9IJ6LN7jbARTlpHz9iG5HfmZH8lV05Fswp4XXdsrMIeoVwox1D0um1Tg5wRdUTum
dSyT+03qBMCh5Spj0GnoEshPwB5u9U5iDkmPIvNSM1QnzvluW024JLrEJswGvaHpzmFGowFRK1o3
/Q5RQ5QLRw4Kd0O/RpLDnS0xZ4kzn7VObT86h1HAp8fBVCFuA1tNcQj5QE4FwRi0rs5SWZfs0zte
FZ1O3WJFDmf4zOV+6Wis4zcGr2SOeQZDl/OVWl1G5VE9DmCWsNSuY35DdX3LCHGlHHPIyw3oTBmH
ZR4O2LFfce/gKaQ8JCJzakBVaK/o0wmPW5tHTqrWPWv8VJWmBwsl7woJw7unlUel0Zd7K2Ocy3dL
Osh7zi93+olTKjvd97cSuQ7r5n14zhTZf0Tg56EqhoUHl55UUG5OUZMvfep4Yb2ev+K0ybd66Skc
9exIOpW4CFa8pVL7Neu3SkM0RpnqmUjsjoyCoAfCZjffI1r31Z5V6uMcHBcSBL9SQ4MpYMCfgOL3
tAMhKsNDludoSMJfTdaruOc8O282f/1bL9qivVOa9XRJYcO4Cum921WPzP4uoN6PsdcbxvjkYnjD
FCVS0JoDIwu9x1P69s5ttbW/sV7QtyhVHGm73TAHgQHkGwYZtEwJBd3EKuopBS6670nVV4YkVlu2
LpkGMa7aNo5hWEclB5702CS3rh17ddjn0Oob5FwCrErIgCzLgwF3IO5pYIfCApQNXsfNGvA5w1I0
kUV7aeM2aWtq8T04HmFu0AI+qmoflS2ACpoRI9ZtkAXJg+cb4KW5eo5EV3TDaDFX/LywwCafh48X
KuRo/c9M6q3UMGSkGWX/sB4QIUMColyGm6QIMmXLAi4JpNnH/6yoVojD1ZtaM3vWNMhM24PXNPNS
eTfvZmMHeX22je+lfvEE5BOGGDrKhwWlauXko7I20Vyh9+BakXJf/Te9M38VoeVexESXuObHw4qF
w5EE8dvUcnokqDD+tajDvOv4dOL/yb0E+ifqHPXf1hynCeV7asrX8Za8hOHbI4/e7YDZtJ8IQ65V
Czlt47IBoQhAPiQgQ7Ii2I3O3DO3/ESg16ovSPCr2G3ni5twvPTtRmrNE3wAy2Jne2k+eWOsG4S3
bWFjTAJrdOy/c7qtXX30ZMse5Wj84DY1Zl2O/AxmKKo5EDeOGsGquYuTjx1wUeY1DAVy+PXWMSZA
vp5nqPXdMhxlN8w68mHNifIxtMOTeSYrED5/E85uU2OhCGxaP8w1rDE1a4NzH0GHYgXSI0xEBphn
5o/YpUHE8il3OGk6UfMVfMKcqrVN5sCf6PDt26QbmqbYd/QVYfZfcTQEdJXOSiGQCg+kwZH0f2J4
XntRpKODza5BU5LCz3dWYFLbIA5pTbeUZGgD+gzZn1CZXL0AZW6bFCTZkK3r+bsWuYvOh6W1cDPE
E8NiM2tY71RSuHhsyMGKyoQeIwV9f24uR8AekrHCrgIsCMZVufCDpdeUrLuxWmaWUBMPbGBXFjvo
lGFlABTziv25C/O69kTTZI4vfM+5q1pJSR866hdhrAecKK87RKJAnDvNWds7xRXtXupp+pjgqmJu
pl6QTgWLxEgrKN0KBTItIxfu1HvH34QKVGVQCKN4a+uHvpx15/AQ2Bslouay6Z/Wnh/muwcSvorw
GwfVB3DqzovTLnfqZtFsMZYEKgr4qtElRXZIExpFFxcfXqvcMIDmuO3T/H4lkL3BEI9IHXMYnXbx
z0oPP765+6fNRaJtBxUY9Fpk6QjI+fcVkHH/mUAuYSnw+VK2VxW7wiQZqZpL1mvmA5Ap923leWwf
tDz4Dqn+yzE5b8DaGfcN9OdpaUKj9KIhAvniIr6cUHzM8ypEYmpMziGvD5XVhJGeFb0b8jF9GXcy
I0EYG+N5WIOX87sF9bn38glnSi4ifxw2+4h6krOvXLENa4IzdjE4L+KvkwqzGLw8eK2MApjsn1td
1T81HBGFvAIZM30pCsP2Kvxy0QfTKx6lJiY7ZFcYOPb2HbDJ6lMw+z27bZ1rO6/1CKiUo2ZpOobP
Rascr9yLotFnQRgHTfTtZREbq3yzXtope7Pn9nFm/u556MEgpcK9eXslyz7+sc83tO6tRpqIzLOo
6RB5N+khQylS2tovYNOnlc+Ig1jsXpXPIrD1HjluK1kcJhqwky4K5YBj+ZyNcYGJxPT5myLzVLYL
jEkHdMzJRxLuzAR0xwIkB2kYbL/m8lzUykkhE9i36UTKRJKXgSteUliUxquKvTP4Gb5DlQLgQuJV
J9goWOzeTZGrsLiRau0oSep5E0YPhUND+pf9sMKDvJOC39G6psTHf2gMZIe/92Y0xrY6QBM4B1EP
RV8r4S5gOMxg+r68wHjgzn4CKggurZR7Obnxvnf7MlSjSUj+A8ouLeWNgNbdn8asrCANt/mBwfwC
Qcm2wpsjE+gGS/+5bGhriYJ+97IGiblSDTvOd3IFJin8huAVCYs8fsq7nt0NqhgBtF+IY3iA2U5S
SCCW5FfHGwL4HbApm0LSU6feJnTUl3f63iO0BUTr5ywBdPEFnpDwMzBMT0kCyHMOn7eViqzJslYO
dBZ8b8YUO/65BnIrZyOQhAI2CB4FSYAyi45z1Zxv2rzxGIaJ+NiKkW/PdF1vQXYE8CAQTezpfJhO
3jClU4pz6PZNcG5JiEr7tTEriKhAw2KcL6RcTDRA8pyC6ZVTwfTFxqfgEIgF+gMrfhswoE3cuM/9
7o7PuMdSBw69bVU8nSC2fORhdrFuCKEHeOyJrM6XJTZafvYSn07UVfr26CI49UbcCkbw4vnheLnp
PIO4z8l+HNVzoH73vNBVwQa+Lv66QugTx+Em5LjyZQg2WynnrBpnHuKixJlKqIKhtmgHWKvlLKyF
fvTe22Bf72yvjC7egfsAX7T623DH42y4Rum1OFAEO7gg6OQVtzH96y6EUdEV4tlj1bVHDuD6/z/j
DT08JRntQPK5Q0rTuAifMAN/a8s/fIxrhvbvkJJRvdL1aDerwgIUSAdYQDQrl+1IDobR1f2E+9Kq
EJol3VbuT/7I8En8YSQ5aePqJ4FewC/ugF/43jTzuLY+fS0iQtmspxoqS1QaxqgP5S1np6UohiYj
lviD8wqfXWrdsQPS1738T8d2fsF5F31N8N9SzyINxTvfecCYa2BfUXY7+LMSzU0LkdT/pghOudT4
59OCj80nJXCJWO8nqSxQ48ctRV6UJk3f4r30ICP75PdogLvQYymJZ4HdT1tCihYJIQ3WTFJL89f6
omisyY35pdoaeLgYihzwZdsWufxoLHsBp/gL9uzPCb3F7W/UkLJ0fsSEJ0tKKqLbMn6+Zf/ZjVwT
eLqTJ8wCcez2QzXC37pm1TrnnqiROUZQfJsfCEeqQkgE7CKBa8VaAG9ttUjOt1RALYTyezuhuc1g
aJJR5oGEhuK54Q5UZxbg0ZrrlX1cKusy3csfpkOaEtzTC76m8WGZu07ILNQ4ePRShWTj+MI0G2lr
rRh3XTatpNnaRGGIpz21nIwD9k3Vjic2OVHl+0iUpLvzWIPh9DYQ9LuPMZHhhnHQXR75OCSccW3Z
osthe4sES2/s40vSfWn98aA78qVSEZPpsMNMmzJ4WqXH16OJqwEeY39OQ7EMkPNrO7CDRSnQscxL
OSUgrlx5sYuk2kLrOQn939yo0RYeM5NW2c/UOc98f63aCT7E36adppYvcwaIcBXDmNi63KLCHUgi
z82oJi/bBjKuEO3cczdu0Fg/3l6BAHIxOgeCyg4I6x0j/h419WOISS424fjgiLsfYwou6DhM98z/
0jijxl12LDvwZPcR3PGKFdYoTs6C1Dc81V1+Q2ZWor6YT6p35JNkPSBJu1VSIXqWJxvV9gErQOYX
pdIWv+2Nskqqah7JVLzxBkqkc0a8G2uNhuV5cftACGOok1psFkwDcQitp7hVx45bcimu9xhVhNAc
y51grUVwwscZ9kfFyb7t9clIj9ZBKhq5n/RcFb7XCVVYWG/nW6iqaF/xXlnvkiDOCLMco9hUiVzD
/NLefyOdmBzTEAa4/c9zMz5c/JeOJC9fN8T9j2xK50QUii8D0nwUO+XoercrgeHG5gi+dGcwERTy
e6iz1pytdrXeYfd8EoOcYdSUgOCg++uknozuUhLVbxaq6rjSz3PNv53+TfLvMCGySLkOy+3Z7Xso
yTma1X94IChjSXoV8dIrkt8WzrNCMXaSDw86Koc4EHhjm1RygscUpGNMCLGvlykdhrwT0VuVR8km
Q8E1GgI0ZIoCo0SztcZecD+mF9IEBPSAzeIPfGC+KvIGxm1U6ZYRyLKYTphIljbJLl6LywloSfgj
7ASkUeyXUzLflif9pqOItrNFLUz6FcDkkGnNH9aHH1pZaHwIXqcN/cCASmJ2ZeR2cJZLtt4W4xWY
mzs3aET7m3YrDajDFEif3+sU6IZ4SYQ5cNVkx3HRPsO5mydzgsXXjL0I04p/r4mIKB9sW/Lu96Ja
TKpAdCsmHfhnKc9rcp1/IAtiNMBs+MOKyDhEBJooWgGRQ87lWZwCkZrjnWmYUjZ2neuCaJYhabyl
R8UdB7/uPLORkannm9iy0XvhlHoX+NfAlXWEvjBIB+JBfuZeF5nTQTur/pURPso1POGFcrbUY/K4
b3H1wFFcimaae5VijVbS3WqBFM6ylWiU1/SOKkxWGhjMIQ0hEk4uJqSTrjPlQo/1ESVgxzvJRCbX
a1NG6psOWwwNaKu7m+92e5803MhL2w7ihQIOSYV1Sh7JavD6jt5a6JgwusAt65WHfXcYvsbDZZJZ
o7otWJ+f6xAk6gGrUiureQAWw/NSWZgovvyCT9kNlbssYpzNoQQIiueI27RVKeOrEWnpwaI9az1j
I0o4hhsYvzOquXSQ5KlHEz25VfV12528PhaJIN8wPvKh9b+vNs85DYp7hch4u2cJERgU66sel6UE
9pzKQ++3D9HI/wb12Udq5/K0DPy2RcxDZtM4B8eKRjb89x0F3fYgruK1SQAdJfddoIUqfHQkVp83
rrBNTnK54Rr4GpF2TOda9YbeKMonUidq6dfdVHG/uH3E9yZvLHCSvqPzzEWxYwchNMqrvocEIhuR
AyukG+XWleO+uBxYm3XajQ5mQSxdevNfUvvmmOA3/VPpJaVoOLuVniNZZTtyyIWZC689L+/bGIvh
fSxlKplmEvz8Z3cQS3cmJYx/R19MSuOFBFw+XunnbCHfntw2MoQRTX5GZkzy0AT0XlDOrljq75Jl
hXIEXZN2h20s0llMoeWMYycbeVeq+twTjosOU/dUnZULDQ/GZ7IFt/xUAnT94+UINVM2Xs/lzhda
77lyQPygwmSjkLoMfBQxmZdc/m94Tg8qn+QOYDfagEEsmVjyrOhH97885pRtXT521Oiwmyyi1cnv
vooe3hkCyv26ruGn0pfHn7cWWrOI/TQNO2nd6YyShi0OC6GTbjp1S2c26SQD33Kz/0x5Mu6zGoHJ
aRJSBn5HS6x/qsXpa8ITA1GCs49UsHdBe62JyvEEha61maWGS9KUPxv/7IV88QqQ+Xk1eblyN7d7
LpRyKZlYnw72Sh00VrMOAauDNEd4AHumEpq9QKatylbHpeeJvoQDzq/UJZ07B3vkqNPH+YGnz68c
tZB//1tj931OlbBBHkz1TS3/BxooP5+7H95f8lfU70JSBVwA+tZ8/Kr+bi+lhHkpAjL0ttyF5L1c
wqk9BwqxpVryCisAlFO0Zl3qTgByyYBVVU1/Pkm5XUpWwR8JrZH1Mus20oqdJfUV2q+r1/I8JRKJ
/k/SMNthaYHlOxckIiYaSjYUdqffJgDv4yQ+6GDTqP01E7gmGwDlBbBTuxn2k5JDc8kyP3Qh46Dv
8/jfATCC3ounILY3RIC6PANHCzKzTYOehGzGLgN16DtJvXYNyyyyuYFgnNKrWljkbOGN5IpceNcA
9FvfE/1BhFKUjWIRePPHfFU3o8gQCpCpuMOsn5rxW8oaAi17qxHOam5IWG4DutHX0zJP3euujW3g
sOjsBXkwtBuc2B9uA4IO/c0o51AFUeKgeAAUMwebIQY1tn2fVy+1iVGqg61MEUjZ9ZQ/h1bdfss4
1dJT51+JKsDCJLqOSGn8uHoJpRofzudzi7EqICjTrlQuhQDGERqTuTXZ0LnvJWvlHS2QYrXa7nnV
S+ERGnNmHgd3JqhC+Aaf+b5h/xwi6TTYl6qARCPo/KHZrLaBhy54QWgtv9LD57xwm7G/CTPQjlPU
5clhnKwRjEpQJMMeDhzGOdwfLv48J83S10LZr7OAbjlE7l3bEzwQMhI2jtWb98d2ZcPNcEClyZkZ
3imtbbAm0i2tWJN76Pe3LeV/1WrMV3dtLzIqMYbuS8acFWVJfwdluuyMAwJ1uxcuHuyw/LTCxAfY
mVtVv1EQCIT/SuDa9Yyfn3qtao36yczrAqur94qkdqD1fhntw6vPjtvoDS/Zk0tFoL3XAZAzGm9i
FhD2ZQjinuZFJo5ue+ef2KHaOCca4u7incfnnBCvhc25IxlxgHjaRWiVVpMCBto8p/AOo/BhJUWo
6Af/11eThESxpR8g5bjvC8Nju+kVIwxNtQzL3ZPEWEhod2tMLSGthcy4jpKGRu9+ztSwxMNhLVv8
O6QFBwTGjbepT4tG8qlD9HRnViIEz53V70l21BGZCHj4zslfDxoA2qL/EeAJF46tibAj4MM2y/Xs
X1XS93VoovxiS6sObjT8ENdcanUvQ5BCRojdLHfZZ+tV6Izl5Je0gpWvW39aA3CCqOzekZkWddS+
EYubYE86be4jM15ddd+o/c1cf48zfWsL+KK+1rVeELw4rMS7GAZk7tMrIs7RGEvvzQtdeuk5NzH6
r2Xb+rrmE6iAvHUOpDjiM53WTTmQynoWgIccbq69J3zoG2dp5pHdJiGxGcHE1DvH4EvWI2VquWZl
TXhx9BYNM9A5HVnLjpnWHhf+841SOqGIJZiXCB7oTG9Q0TnKZSO7zoX0Aqd3wSZJD+6Chj5BXUuK
/1EUuCiKx7EcuIveP+zWQrDgNi56ztH3Z6iSUKO5BOSF5kqDSpyUPiwr9JBDSL4KvV/Ui3bOmmuI
nXJk9IGg/CHrVwKMfM6IyLSnd636dHfe9X7nLzvWExIca5l03JjIolFN/OMKHWKxuyzMOjh4smHj
sT7Xx45FqFS/rsvtzNe1HUf2nfDuBTHUpcifXj4uXDnC9aQXpMjchd3Xkz6Zxt6UVLsudYpZvBKQ
rlD7Yo01BwOti6GZFDSTAjopNhlxZ1oHr97h5cTV2Vp5t/aR37rUKCTNl2rbYB+0NEX37GYiXoJQ
bq5Fs+7AmYvUiVTzdj/Y1AYL8keSjYYXJ+ihhehDm1diKfKddw/o3Evo8CI2+bkjVWijmCBG3dKR
C+m54st2/o2fDQIc7TYZ9GbHH/I1rN052dTtSLMlfiCC4jN75YtWO/J2J3siK8TC4Lx9GXa9Nxhd
x0L5ufa9/HNzJohSnaeaYjwAdw8SX0RL0HUnni6n//zDMjS8s9cV5fPy1koQjynyZodUm2ZQpH3i
MzG824GfrlVF8vhwUn8WK0I/HgkylvaB3a47tRAsj2W9y1/qs5mUO3OyntPtJEJLYhQhAEdhBTdn
/KoAvyW6waMhaiuVmR0Ochtqm1Yu9nvPwK6mLREZaK3PZ1DhwZjkrS4xGNNUnV1RXxO3FLbRSI6c
r/q2hA2ArKv9ZnCTxdf5nnou+UbUTCya9EqMQ/OyTD0rVfccbjNZgFmJWnFF/Quyu+88hQcyPRee
C5oj1N9QNgbG2N3S/qikfDz3wZUYrwfHejfj2w861phEMmPkFb8SNdWiSKt+XC5yjG6abl8FnFsu
2UdRnOWb7qw1PSVEq6Vp4GjfK2bnj1ZmE7F/2Qhxkv9y1ZymSuX1WUHhsqbRkRqfGhixJjf0h14u
DDowT/UZbsZuxPPuj6ZHYt2WohFfievMx3Qw+TI8winLqhEnbO1VlniLUU4PFbo5PLTEcYXVtCTd
70iH87EZainGU6ciqH8AlG4bRdl5NPkWJFyosQeks6RWboQPWUhYKqFKDLGDkN95pXxxKnZ+vlPD
4/0KoQFmwOJI4I0TNv/++NaXX/WKkRCe1b2ml9BDo2pqfDEmKTss96lLduvH35GehYId/PSevBNk
qAs6cXx53g+olqnAIr20H/QgqcWfJhJBnutogXnBKU7/q8R613T6WeUa7al/TpA2tW7AQvrsEO7X
DzWc431S+8hWDKKjXtBzwjbe+8tiFDrTCcbiUTkqXIs9Kqiw527HwNDS6Bwwh4jHle8yAyAU8Ec2
UunqZL+nk7Q5SrGufEVkvgUH2Nx4ED+6ikIDF3Nk1M6tpkafgNfCEi+cSLdcuIw3zbKOR2rWYylZ
hKlN2zocnJGviUCT4feAwiazVcCmh5icY3cvmJeQ8bNI8Gn+BFbZkydFRI4MJpSnkGBaGRNeDrym
EDynb+VXKHV464cS7kJ37NQeeBcWSUga73yZV86zR8gt8fETzxoyPperpBiYhq3k4s4budZjyAki
5ciACjxw067LCnTW1t+5w7598f+Psu37PXI/0JSQhX3k58NF/my5wBbsEw5nuGcy4xbMkxNZPnQ6
MN1FVbBK9Zeazz3DTiEULn1ofnPB0Vq/9h4FGzlTRep9+5p2Hz+sINOwmWFcg26bKDE7LVR4s24d
iHQTWrvMHLUB84L6x7ijaZtamb8tWGcmDzVbhFFkYG+DO6Xl31g/m28bThkiPXuFaQZ9nPuRTAmU
29gd7qqfILOMhasBkT1XYYIuv0/hrgpg0aCIXbCtWDNgJZ3ZRYNOY4T09JWtcr7ZsdAWUPmCVd3P
3ju9xBij4E1fi35Oacug8ZobIC+Opi38Axfxr5X/En5v1tBc/GpypgGR5AqdBclXWzj26eQnqAfK
rWCPjnzBo7znvHtwrQyFnQ3bt7JS30gFkg+NCEj067jQv8nPs75Ai05a1X19veUa8KLGYfkNZ6xE
sYqPo7kVP+K4JGpTiXDBk1SBdqVgVX0eCtxNKxKZ5ecgxpOc86ZdiaIWtKhYoP0N53Sk+WNcFKvf
mBHlLuFY420KDT93zqUbepZK6vmHGnIg0MLjT+NhI8PXX3Ay5e0otSIyqreOxfm+qHD0neCQXRwc
OAwwSe/LVWqgdJ6YAY0CbuCLW1H+IfHQ5H1PdvBZdCbBhxN/Z2RAMKL7D8Z8EhwGM3ADSIIrscQE
EUjRf6fxG4QDgADiYcs8+hpyQtjRhUf1Sy6yIvISZVcrIIZ4r1UyRnhZlnIo6AdC1iWX1EcYm9pm
yocR04kyUuJdXM1+34cVMhxKGmX3CUlJ7dftj08Gpu633o0hZMiVcgXafrxN/6QBLmZjUaSqh8VJ
VQoQsGTe0DBwT+F6iyzrxQdC2iZ+OQCgXS9NiG9VMsGy4qtLQ/KsZr4F279V3GFMpevvwhcGboVM
njOez7EyqUoRbIBwwynbZgaTYFaDmICF5DJjy7hKw6m/usCJ0L/w+e/O7aywZcDaPqZNOPlMdbI2
C3W0SMuTQ0EAlAZ3L4ut5QqI1fhlPJ98Ts+3J/hTIIVN3tSvNKzzeWomPtVnOWDDX19N29oZE27t
yfRzyqsn1kZgUgatxICdN/cc267s521jsK/HKqu/EQ25yBWyqGyTCX9H7ial+dkacQE5lYB4xAkT
NgB/EXdQxpgSMfLsOaaYFEsvmfTy3s2c72T+SlLXmCCJfm3+QAltd7X4l+eJHIEsnZ2Z5eRTUIlR
IKjnmhjBpIlGu0ZfVSIY5Mi8xAYzN3qhc73zfg/1KpIyyuPnShppMLEt0Lz8ukQn4xBTvG1z27xv
h7QoYgvuH2vMBfRQWXIUqq26mdRp0Hp2Kpj/1HNvCmoS4x2F1Po/vRIkSeQrUHsYXCMRPD93qTyS
h0Uj3hDATMovmwcJFtF22v1ULjN+5mJ0u7Cvdk1f8c+BmyEcLDmetNmgT2Uh9yswPvFwePB9pzHY
925aWjdlj35G99uSjDyHWyjuWTnrWzv7Dskkbw0YvUBtzB9uPU1Px0Zvj97PD4RgMr5SMCD7OI+2
mI+vSFaDDuhrDWY74MZwzPD90BOgkl9Q83zWHhWOrswoxSyR39Uumu0SBBvUvSFrsaqd909iyVam
bzoDLptTdv1hFAYnD8zdnjzQ3hW0hsxPYPXF/LWGMHySj9xL2PzOPWh1kHvRVU5EXTthZvqjXO/P
yfQ+qpIzcacPJUROq6mMNnkN7REyZKA40d6rFs3ppmubqlpS/S1FgPI1XmSqUeJMVREKCTnk81Hu
a8dtc+aL2NC5ivbTNpQgxR0H0pnwlzDA7V44/Q4LWe9bNayL76yH3Jd7lVMFG/9cJasQghI0OJn3
syO8cTmeEuDR/TLUfec6aNfab6dvcynLlj7znRdQ8FaYNNo5bbQ4Hd2eZ4gXhMNzrxJsZ+nBmKcx
PQYdZEW526ailqJS5tSpaNd9yYmJCnyAm0ywvbwp81G3Q0B9qIWPYr9qIcX7jhZ1Kw+HrDw9anV5
ojWTEITGypwfwlxHiedFi1UiWN2IEGmHqTTiecfC3hsZdFleICACXyAwv8iJbKZK8GOXxy/3f4B/
p08kbu/yG32Taw+WfhO6IVz14ogYtjCjIhF2UirYn5VW74OZ5m85cYB+2sF3rCg0fcC4MjINf7aM
kPZCteF1VleQIpfTQdTxOHW6MAFzYa+yWGk5GyIEqynM+QI+aBwz6KIIU7YQ3ikVnRYurdjAKtIs
RVdThqVzshZgxRuA6l3GgC1Qa6DYU8w6RrUuAka1Ukt4VN9/eMmAAuBMpQOKpJiYobt6dxkqqGAk
/TINQYJdAyAAl9O6bqCiZPN+4WKC1OsO+drHoWw0tj1vMwEbZepBbzkfv4OWEEby+yJfN/axOdBE
s161uoasGLGjNz6ToZHDhfaDkLTlFF3PCI5XND2BH+8i1Mus/Ed0gOUZzpJGqrnK1fSMEQYoExxS
oe9+4WIkXpVGZL+3UOe1Y78wXxWVyWRznQdUdlK9vBeRh7NlEnU34xWltMnWWg4wuMNetjVCZMSI
RKSiw4q/IePQ4FD3HbFJjkAIUTy7nGlaDhk1PJWTrNL17eausTzR8Qeqp3Z4QC80mPqlrMBPyv5h
Z11NVKA5EE7WgmGmWfF0WMQbuaKYjQ2eQvyaG1fvJUoDUASBx+TewxCnaeQUndoR0+O00FWQ7R/u
+gMGIzHMdfX8h4oS2xtr2iCr1ZoHL8shPuofPV607JBeYRXuUdpE1DCDMxfHIAu9Gow9SD1irHjj
xiZS144dbopr+zyo2DLyjtS+suOfe5JbtXJ1xgAckk66RAxO+fiYWfanPrCwWVJTXMrIHpmBacQg
R4ChyW4BG61nZZ+MIbQrKfeEDCj0ZCaX0lTWHKBC9Q2pkwY6hKK9uvVB+s0xFn0nPK3r8LECNdJp
jsEhcc/fWBPwYPlBC0uZt4LOZHS19M+uMJtii8ZIw6sE+ZSzDalRn9Ai9ZVxeq6C+L4dG5ysqP4k
Tve74HVvBWcSxPd7r8hd57DwVfekw1kuNNxNEr68m1HIDLZekiIlP7myMEkxbI9bqkQB6Lhr1eCU
OyhnooMJ5ITkEMwPupirXW827Y8mlS/NAbCRIROrsloeZzLYkOQFxLtRQvfMTliavv3pr1s980G5
ahijubnHsXiqgulpRD0zYOZSAooVr8mI+WbP9CfpG+2RIjt7e0rBnDInTOWxYtxsVZMqklzbjdO7
rWkgHNiZenOjebG2ESL3GNoqVtfhMgo7IZBMhaa+k05W6pXWrz0hjdD4UAYx/h6kvdeRIyTxBiJz
gt+nfYuAI18Xw6MEWzoGnk0lSjTlQ4zowySxqEVYLVX27lIbTdcDsv7Nzk2PI0bPUTW7KfdbZlDc
1LosACmaBd+AdaBORzRFIpMmUw5uUImoidSXQzZNPiR8CFr7SYJa821gt5UC6VW9Yn+Whwj4sYV/
/EGGHR94eAf01UE+3xPxcxdOfECKomvyHK5SOEINdLnbBtKrH4SMoZdS/W1me0M4anhNLo0s4HEA
PG16K5HK+Rd4qM1nXajckDJJFtP9j9px8tSgTMQsQxMq2NC11BMLJypUrOf01q6ON9mXYLAcb7w4
FQ1thhNbyF1Wz0HYeY1thh0Pyq8mwpcrBr7aHMPEmAnAW64rFqDuRqjagjQ8c1zZFoak4EYLwmN6
98oFGte6hE/x0zojrw4LoIniGDMjqXknf8I/BcALGmNPWpkEa8r510B+2AHgavLewAoXoha45H7H
ubnzq2H/4AJQKY2whuysJzl2dZ8dU/6HRHrXL2bvAyCID+W1F8DlzoojW/x74apF7LXcTVa4Mdfy
yQ2GJl5ss81bcf451U7V1HSVFbMRTif8mhK8uOGiSeU4B4n+JU+AzzG0qPUNsnE7XMlB9BfHwS83
QwicxpeeuqEBQtY0PMDpxqJzM5xDXnePhoWCWdMajNu7pNHhN15oNvgQT+XX/4H4/hmhGPvN/sfz
fd1PYA4oD2WcjwxnDb06vVo9L8+wagrY3c1EbnBGZ+kywrO1jGzFOLpQSMI4AS9QNgcI/pABrcey
8B62rLsXQ6/STYsUTKMdsqL5sMlYyCKlcMrttCpzFZWiWtqIhOMc2E4N3fIVyrc/iA3czpEzM/d6
bdZV8qm8EskfQ7NXRmAhCkjJsdMmpeT0sq1gkGsCmx57EembHuzabHSDZ24fRPLIKrf03aGEpYO4
yGsiFddAWY6EcqVpTep66Jykt0JF3a4hiji/zLuzgS9HZf179fmy3BybYymQTveMo3AoGioX68wv
2SlqV0Oo+Cu5tI8vIdomOACLVkjAu6BSozWPrzxMNeMpda99CThvFk7UHPKm/dLYtNZU4/ZB0cmv
6qDbHaKMO2cRgPAk62ujbx+3cjpPcYbW7WAQZC+3dM1/h/1/brMm2BGiv3NjIzdRbv3ISoiBDQUZ
JdalSKTEJAul2V9fEGe+mKbCYUA2Q3S2gZyXAXBsVkyBgNZ1rT3NGjy/f6JGT76Oa1S1A/Sd/MUn
KV25TclmD0roLeVqQ6hg/DE1PpY2eyjKFlzPEg4t7tvztl50Ixj7bwzKMYH/9mOEGsR/wc0Ng6jM
VAqYDdioWevwdc1sPhRkzIeR1iX8C6PDvyqIARnpV/MdCZ5lHr461S85oQBktqttnSWzMjZmYWlG
UOEw1o/hVlK5VN1XYeCFnm0T/zbzke2fpsH5JnrRcrfg3IqAsXG1S+PfMo5068UG0DSMtCrx1vm2
nHKfoOmwJehfaLxcFAA+DeoInfTW2fPV4N1K6Yk1KaL+bnBIYvvKQ0Xl4fQY4mAajF7IZNvq3gLl
Y+Hs2B5xUx1qarOX6uWPqH0+SwisILYmr/wHanqlfXh3j09wCWF0y3f0h6q5GBUI/nA6q9ypBzKv
AsBg2E2/ESZMrsiZJJya3Lf2ag55owSE4byhGDT2QOWtOoMKQ1a4N5SMqes/6R/3xlGihu2mYZR1
qR/EaUUo0VItKVL3mzMfDy0DICjvh03rBjHighALE4RXSUiRF7IqzijQH0RSP3V7o8NIii4riXwT
5HiuGKyadRKE92HqH1sozgUVNJR/APaH2kZ4tpEgcqIi6kntA33TJW8ylX6y1EP3NpKuBngGMMmz
A1qt7iIfj7tPOFTusKehze4Edka0wq62UizvZYEV9rjJQzfWmKMFIf9ecERjkZCkuB7RJcFkmAIi
K9DbXXQmfQVkhFM2b+q+zXUVxQFG5kgaUKbOOZLTdw5Ebb2A0lQ6rrz/W+EJU77q3yxAyKhe+1xo
x4c+pw5ArMP9vFmVTvuEaICZIFqjq4N1ZOfwvMSkBS2glAA9+2+NjtDNwhEMPo5SUlLd9aX/7pkN
Og5uAqcBR7OhSVsYcDHRRm1AXWP/43GiMzj+/XeKJypJofQuuwDAVAmqq0HAhq1jkjL8VQWLrTxz
M9+SexrnriNiRrkAz6G/UKwI/ikLUnqNM7lpScqwRgOmCXbtdROE6YXtW7jKTsGhH8Ilghuiu/Kc
qVIthdOQGty9zUeS6H85xoYOTskTCROsA6Zu/6SBspy8/OqNjTghL08vphUQLE1HxIMToShWUqp2
EoPfJs7Ml3/n1xLKxQR+MiS8SfAPThOAKQH4+D2tFXpwproSeAgbZ3AbcTazo9uqQi3AW4VuQFXt
s/gKZYaV/BvG67MRIsy1ML2svSjeaTP3V7NwFCKBWgCuCpo6OjU28Q/N0sEOpKuci/ehgQAMmEyO
nf63A7yiyQ7zfi3rdgOxjpNi1BGa07qT1EsTi5HIeHs07oAZUN43zzOrWqZLADifjCyv2jvxiSPS
3G3HVsWTDEGbyOPTO5z5dWbdoLDHmQFE3+Brf33MXeJ3cA6uIRsMtaV2/pVYmdRnZGejIFPlEKm/
tNysoqxgkojHQIYPfTv9dXWyLPKjFaDlGxECN3UWcA9cvCh0k7J79ABK+jd7bSWiy6VI7gLvrpgt
zHUr8AmWpNOGSu7HkJXrrYljtf4Meb2nPPwSuzVeyqupHhtTOW1H2SARRZ8Y3ZJHZu2Uptq854GJ
eJGIQ07kCSoovS7W0hi7iIWesmTkoVMcLTwcWiDEnRXo/D5D7K45XJMfSNYiXxApvHMaz5WIjxhK
Rv3ia82etrzAraKqlOHW9gRXq9+4eGBA/t9SSN7+2UE2yPH3hhqZFLgYTW0KkCliDpVPcyV8u2u3
jUTJkfWlv57nChfnXHxDUrEoj6ps4tNvcbDxHf/2E/sFz8H6O/hGPjg0CVMSk9ZaUcw1w25K6MDf
kf9B5hZsRiquQTnol3IZfli0ZprVKFKnffwBCG5/g5o3Dm6YchORtkOJCqyp3zzTYoV0OZriDCKP
8M0smDAbMgP+m0x0T1oh5Mz59AMdVdqtwmzednu9jpMcMFHdWLPmSCmkxNunbls3FbKWRwcoGwkq
dcrPx1zrxwtkQGzOA/1QD0RFXJ62Ra8U9xfUbi/TakkLosuy61b/8OUfgIcmgjcRuTntI0yqc96N
cLmfK8Kg7e9ktgDOX3yJ1wMTThFLOFObaiEWtPysZkMlkbvanLqYNym0fPd7D+0NGpIMaXAEZi5z
H0XjMhMmXOrCmQZ+ImX9Wimj3ctaF887RkC0cNYsGIyyzUqZC3fe2PvgvA9AOW+XhR5gKnFrL6Gj
t6K1bcBJzWNsJGtpZOS3sCuCUDbSBvSCRkKJAlmzt0vHxe4O05PgT6XYdoYqmoGPuJWWybYoPDdj
+6EDaRx9JrGdz6Wygb98YEGhgChcDtQkanumx2zbi5Lgdqoiw4h/KyYBB7z3K1hLUDmSWVgQwyHD
/gjSp7ebWN5W0lcIvdv8ToOl7Apx7M/jBbg00wjZpQpjMUdra1ygKVdX2Lvcjp8St54GVDqw4IUn
Qtag6NHvAiBhN1mGxva0ri+SlLG2aWkANd/FZ02oVHl3WG/NCMOcFX3qVW6Zo0+CdGSmQQ2rOu2v
YAPNEgCmggbjemal6VUj7Lp+vUDP45jBzM67DKmGm9I5Tq8YAF4TOwx+42ngqf0uFaNGpLpPKe2J
psprQodS1g8WCEGWh6ZjfNFeyUxVKcGCJfTV/OWjA4s/z0in7L0SdeJ2HHok2PoPLan6URRQ5FXH
gs3EKcfWMSYjkM/8XnBlLpL/Gtm/BCL2qteuJ9lyebciIfUi+HSfpD1h1vEBCKBWlOiw7Obr+CdS
HCTjjs0IoRsU4fqASTAFFBBfDyjYnvFZSuEXjj/oR6NjvUw5iZWmSeaMNRVAtnSKyVNDN6iFI0kZ
TvWXSWFA4cNr2Z3UtnkHOJDNlE01lzBg1PZR/FkViI2ylNyuCFCgwa84uISbzOibGFCNhrQ5vL2w
7XgALjVteM/yJt8ul0mYaT4mQaUOdjgKCMWfKLsCudsvMCHLdg/vIyvEI7KqW8hT6F+iPrOTVH7j
vEa64hr/yreDKDFaGF/O+gZtXYkFcOb3nh8JOBGnJ1ZJFsub1twhRHr3NxfI9TrdNaQn/netTBGt
B9V9RpYCErB1m3HOSUpOyvzV/Rsm3f7rykDFrR+umuZJA5WhltTjGMn4TJG+7e7szVrlqyhiyrh9
w3WXMre3w2cP2zLlA7KbT2R/oiVY84xh008zaWL0B2tZretvT+lnTYOio0GuIZPd69I0EvDexHic
hGxHuy3VfGARLC0w01aRUXKE2LiCxruPJoBPj2qD86WmSXL/qGM/B8qJlfu9AruDeqy3MIWUSQxH
Q10+SFhkk1vOaL4hvcpEPDd3dfcoZgFD78arDPR8FyrnXl1FxB/JfzvkTMxvxazeQvKos80WPWbO
vHA1CpW9A9ytrtr2v6p9qfEzQeaqWqzT6wBi6izMBhd0ua/t+YBCU4CFWEO3+Hx1MSxkdKlR1kLO
BCWkq8usyJ15R31Zyq0PPKwhbfZSZMN+M8ohx05tolX0R+6Q0mlwQ9Lj45np2BD7svq3hdbcCETb
QGR3qPB5hfZctq4Ez2usbtTSe2D0+mtD11Daeyc8cI0ZJVsW1o4qRitCVCeBVRKU9aDFWU9fy77f
QHdoIaWENg+fbciz0yS1XYoYxac4pBzrfQDOjyoz7MD65fFjdcSYfwhysFa8q8bxwkXN1S8XJYJt
HmgozNsXtZ/VH6UBG0qKTdsfZPAQVGHvAB8dv2KkrfwaJv5GGjZruXuizGXTDNMuOpM492HhSXGY
llyX/62eNWNnnM0Cxy3beFRK8o86D6ZrT+j/WEpN6RtNnVt703cQVvMu4wjerI5tTxNad2f7ai2y
FPYcv05ogm9TuVqPAp7ty9kDeHtQisa/u7uF8+WqMNaUU/72jSXAGaYxaSr2m7rL3VU1nNWN5bUO
aM/rOYvVtRKL7Q9VS2ekb81eYLunvi00fKmi5qwWU8GcV8aWud5JhWo9bo2e9GhB9AphT5dV/abi
t5eiKtfWW86kkEnvZdLi4am2P5xu3qNDvPguCtziF+U2MEJutOGFOpoFkFIoUTONojM6JzlEVnGH
EUbemBtpwHlX6M3nUWDP0FZUD7D2KCOtp/OpFG2fqFFlErmf2CNiKgDa5MKittbsrYNez8n9kw4I
7FJTuh4+0WPbK22pMpqlHxzAz0gT6PDymiNMp+7KPD4eFNq5g0ZG7kalqrEWCQG1XS/owiKzxlfN
t7WIykYbx9Phlfmm9skQSAkQdbZlwIe+V+c7apiNkhOdhMtYTyEnYgHL16C/5FMnHAYniBu3d9zo
DpTR76kIJ+N2+pzA9555GqbD/wR1yfn3LavCIQjzg8bjlSR9EvwLuW0O9WPe16kGauvJFUMNIHfv
kl5v78ck/LQxNzdi4Oz3sTrR0nTNaKzGFvxs0s5T3jhnvqz9o2KusDMNDbHnkpSNDBJ7hzkF39YI
H9mr28Bp1J/JTKP5zICLlhlwPRjyv8V8ieBqn43klTlRAPtU8QRx8pty4MLL9NNze92adeXTEWzZ
63k8gUv0S90aviiKzEGtaVbs9tXfbcaTXEDgUlDiRqq/pW78YI50bURIE1T0vyleR5PoylVrk4Mh
/v9fd7/p/93Sc1gC7G8wMYwbdmSnEoXt7fRXCqr1uygkgcPlPo8A6k+hDwN3tIDhz8kKewDqqNFR
aNYAtNVTy404eL9JCHruEFRa/3B0iF29Lal29QgiT/d8C9DzIZuEfWrtUFzoEsom8Q7QXskxiAD2
Y0p2h52bKQ/BWeIgkoQMeJh/Dx+DhzslA0FeG7VZ1abisRNyXBEPTZKc6VUkiZozAb7x7oj9y2jd
cSp/zTlJCh8+GD6phHJYduXw+DYUJyEBvzjG+jqIILsDz1gWSvXkb+lsPcojBrjklWooSe8zUKiT
EsiYyRJlF4K0pC9DTMD+fCxg96rjC6uG4rqBiCfmUOUBxe37mNqzVIUzxR7Zvw4AG9EBc/mJtoxc
g5d2PHHBfMv7xOhwbIrE6bsDr3cTZpepNOjoV3vcN4uOzaDzi/FVOt/YyksbcQfIL7KavxO5XCqb
i+/oI31/E4U+2YpnSX42T1Xfos8ifh1+FJ0XbKAJz/Lo5UMuiD5oKUIaMqI1TLKv9Gk+CUU3YqmI
1Ya16/tTLcoZdCsy53ZKCGNLHyad0X7l25XGzcRXJWT1SaPbWF4t2DQBbg1cCBayJz5ZkccRIs+7
5KvsTHlv38Bb0z0MKQXTLYNc7mD6dMCLUoedWHk1B2Oqllin2j/ga5jtWq0r/sXRIutqgh+L/lAE
xVMko5Wb789VQpcNhYmb/nV8l/37U/Bd2qPowaqxOCzB4h1tB56yPDtQ/1CCJdYjRxcblCkpMjGj
aWvzg25B2wTKgGLDgFYmzJKpXNyvdy0nvD5hWWPNogGqt+KUZmQ/o0mb8xiLYa7pPOb0PyZQSLv2
WiKQFWn09yBNfTfpbaaAFshF/abf44bVn/UdxanKFcsZTpboI54UWbNLIJfnCk4dMcsMIiU1mjfj
KRNvbVLzpyviufmoHzU4egw9PdEWla0kFVvwYfTTd4u4cJfd/qi3Hm7tQgsWPceco+SfuWPoTILZ
UNvsXHH3bqrjpnDeaOD3F46FPhQrvB4H/jUYasx7R3+r8K+ervn7mT74nAb3S3uPMdtk2SaJtiLG
OAgkQScPbGKQCwPH9HYF/AL5L6M+aOzUOcSgAuAPEMWPwLrcFUCjO4tJcOgUJu3j7w9uRJT/wrGo
ABVdGdCeu06S3PTJJL5+5qPiwudXKXrFACq6FX/9TZ2nyemj1JfjvV2zJVErv7WbOChHtIuIWH4+
pvLp/2u66FXjfbOHhVc9Y+JnawKjWse8rf1fTIr3VKWwyqhP3wA8OjWDRS2kq4cbfgjARG+o24Po
quDGKr1fXorUf+DMzL29zAzusGq8EcjiY893UwZVvEoYex5f3RNJ09pytU+R/spgPieEaMDZmtnw
IIRuBCUCe4R8IncTNpih+sTXvGYb8rW09HFsTSe9HQkOh1wzQMUggZDpuB5KfInW7GpxUSmgJ3gp
4ix+gNvXTTZZXCSGbkOKWAquUjOQKqM/9e8Qy1WHlFH+paJtfXpBeTF4RjN19RiTflBm97arfMxR
LH55U9XSjGQOpWsgaW2hjix+TwJU8v1Iako6aRkVQquT98CjTVE7GIOA3A4vNcJF+OnTxlHe4Nqh
8dzlFH/JlLiY6gh4oNka3tz/gwIpnP3hAZ8FweRRr7qiYP6jUM2tkatxn3vqF+Xq0G7BbUZJJMKX
tW05afeTNCG/61liKFRxDBRNamA3l135gxPe3K2PknjuBDCXlTct9pDjuASfmDd9u997/+KokugJ
gIwWHWXxCIzXVApRrqHnAf0Rqknh6GXgtMao46uAlASOU6ODOVrKEFSf5eKogioxSqBbVglCam+u
xdLmsaDp8SmeVgkcNxM0HWM9BanLzS1o21VtLl7chPNw6Zj7fVK0OtKFDQnVCeVmYC/ZxDvHaKe3
RGhZLNXYf8eM43RZbpFivSBcu/JGd6ger47HHLpWvOujQrglvaowAjUynuOgy8r+B+yhwZ12YUgV
XR0eUVUPgsTuTv6HWha2R7zbcfyMkdXD6OquW92Z9AisduMaDujDvUUQfcMUtmVWXwklyAKISEgQ
QWsfNvelOHtWzLAnkNZe2fLDCiHscR8l19AcPidYYmUj47YPLuZwTxvHxYcIaMr3WiNVrh/IOK8N
cri8P2GVRBO+oX+Tm5stBqMtM74QdLa++0n+UksBB6bo9fhrXYiuI960EZlEaRtU1HH/SC7qsfNt
jV7voaMTN8DIn4DBysks8/bw1HnmD4AB9DkANQf8P/ERVdgI0O2SiVBIDx9m8Gz+3xij12CHhyPP
5IqU6zRXIs6pwqMiwmgtwbDSrZZIpuPL7AQLaRkdqUzBUt9TJA2uyMllk/Ai0zunnlLaE2knLo9G
KWhomL49giuwVG1tl5VASC5OyZoXdMDyaGDTvQxCrmQEtjYxFRxmf43RoFVtbQq3gqnx13r+I5yg
MiCXIOSyOk4yi8C/7aWWRfA5/vsvPqZPLXK5Xz+5aikjxKJx7l2YlQArUMXrmNXHMasGL9mjfZ0/
MYBNn/hwZUl8T1Dc1X9kKzSwiwd4wylYnAKkJiCWZBICn3fWMO6uOUEsR8PuYv6D9pMqOMyMHXpr
AntnfzPpjbcopjemUan0ve/hk97+2h+3AK+rkUdvAEaJxHxPegvZZYrNbCzDkrB/hpU1W1WfPli7
ddJiTp90soA/xLE4ZrLgVz3QUIslfDYTISZScyovCjWeWz5ER3yrulCMoK5bp6thJJZjpaYEVxku
uT5mX+fMr50RdkGVJScyhm3/ldIFow6M1vgaPGzfpup/dkBZpR6f1428/UGMisZ6m5OCKPo0z/FK
hzTN6BzbLuy2dHKs+EzFaUAFHFV41g2nzcrAOVZDY0XrxOisuBuF3dHN4MctQ1bA2YLvL/ehMlhU
TzpR9Glu8KhEi+mCj7Oltfdv5aSh6KhhXicKALHUsNlTsGB8VTVpICf9GK08B9WdouNXZ2qTppjX
wYKvlEWr6kY/yiT62yrARM6cu+IeuHOazGw401QlRAKuGkZK7HDVSebJMIpI6fmHQpjKWrEA18cL
ga7cUyrUXCnLd55Zlf8WDI5Efc06FOgpbV4iZ/FR2R6+pHq4nhzf4WpxmCl+YwM0/MG1kwsE4O5D
RQ1rswv/MRz/FhB2YG/NWMN+oxfWhRpe1BT28tshBDfx4c3Vg3PSbDYWfUWHaW6CLAzOVcFgxa4J
MG0pYvEHs9ClRZlzWiryaXqRZI1tTuHhn/W/L9z+V/qyDbxfqytFK6/YND8EUN7GdfSsVPldZkhA
6AMGTQlGch/0+ecst6eG/uUZRR6B6b9RYf+QmJ3eZuWNQecN8LxMl9klm5Jol7EJRNiHbBo5pHhx
gGhpdMilaVoVnu2pRXebAz1QSWIUyP+nqdTQcGYQlQJ8lQwErhjZGKnfduxeFesGU9eJh60KHOzM
9oqJqI6l9aGt+8n8Dk5gcc14MpgKNCHq/0QZ4+HBWZ1xtPyQ0IFSo1k3Elgz9E6csVSOgYFR2Qoy
Mv4Ot6ZV/pcUYsJ87c991RpzpbWgG/0Nyfj+wfQmAgEN3eCWxrp8Dq5OYBTlvRwNrxaDD8fTqN9v
IPyt7FHtuqS8IJG3Qib9KW3HwyKaqwkP0Jbz1/cwE+oa2UHiT7H/+fbh6Q+D4VidEdXse2inJYDL
LE1b3IFEUVqAmjBnPOUDp4s8PBnzgs202vzuWX2zfdV+DVhSm/zwkh7wNghH3JM1zBAhyg8okQvE
EztVEAmfzMjOf/npnXy9FqBI1Uqz52mwaANUGGgU3Xyw+3wpmAbLuMnkKlNJ1fgMMixqHzKUyRMi
nPyOAzLIxicIh/grdEIMN5e9e4/5tVvs4bOWrnYbv2tffuHgFDwKA0CQjpeeIpZ15V1SpC2W8mF9
QDBZ8g1t3sieynoEuBRtIn88wna7hKzuIs4g2UlegRhzBUCzPG1mEaPXiBQWT2XwuqbGyaSoCoce
JyE3s6qOT2e0aRdSklc1id/ggXvWEsuT9xFr74DKeO+dlK3rpgtEug/St7LkdNEZ66ba68erB+lL
qej5AIbHdEN7EN6sWFQFlTzW+qYHlNaVC5asS2NnnsuUxSLjPSvox8Vn1lWuVTWlV3cwcqMnmdkB
2JbHmr/Eg77K3a31jj6lzwIYOSoGUb76Cngm03v/zno03TeQE0ecT0OOK3/HZFxlIEmps4OtjiSr
8YQG96RfZcDKZtveteGdGW1jnvf+JWCtIX6FCFs7jPuCMkn/msV6aPeZ5QcwryvKu3pIAFuwHD/o
JY73YkBX6L2jWaxhhpCK7X3tNjB0PMthoZ1QWA1kQ4Mme0VtSep3HYJkC0EKQB1Zrzino8oe+FgS
Cc3PWBY2dneFK1luNWoqW/W1U2ny02z70N9kLkg/pyzgQM3wNUOrnLaHfTpyPKDVXjoBZwFe1R2t
NbqZQsec6k++szPPlMI9MkbVyykOE3BDpxzpz6GZ430788+NweHoWnNWkAOP16joDXPOXUYb+SDQ
iPGjbHEd22Y0vNTl1hrifqNHQU8FQrLyTXF15sHLNUOZM5n991L6tlHDBTnB6kHpw4z4542CvS1k
gZ/3EsD8FBGeGbidCPbljOgPy+H6q8PepHXxdstMKf1zgR46oAsUXVdcCJwCaE5WLFhPOXy/gcGv
tTQ+0A8Q9kCe5fESNbqZcbfYqsUq1oFrUgeAQoHg4JcwLHeQHJ6jzP4ueBMfCWFVq00Vm9ZQuGj1
AYLJ5zkHhXBZRV9jKKOCBV7GQzKu0aXnN8kae4OMJeiZsvTI/+ro8/okRHYi0FeBmyQAWA0VFI32
YAT8B8et6KZUH1VcCui8iFzcpUt2JgSrsHegiLpy2JmnJiPgpO4FODGxeFUxlherpWblnCjfurJ+
CwiNEE7/2jCukcZQnP0fSYFo/GtDLOpZ5czQmdU7dehKiDPOlT8BB4PnhHJtc8D1ZA7S51EBIEr3
6CXbZTaCPaCfNxWquEYuf+91V9oZVSaQLV43nx6378pTONUgPvmVcYAz72ecDUw5VOppLBgRZzKj
WNrY1GpaiTDYD44Ovr7/650Ias71zh7tiaJ7IjHJJP4yfb0bC6oiQN8e/FzecXfpmM/GOrFwC3/e
e8tkWqhkdwy6a/z8VGKLu9+3Cn2WnqMB0MP2lC2FeMM+rTTUd4H+9mU3KhxqHidviSEM0uxYyjXw
iRUsNsgFqZYPuOd19UnOzg2V6H0kHxjs5mJUU0APa0yMkQEKIQ1qUdCqK9Z9RC0m8b45KiQhrIwg
8+Xpb5JHarX3RKps1cE/ER9VefWyD2qQokczDXTAfp30AMgQBNCtvgbfrDWJg5IJ5aPad22gRoGP
lokKQCn2BfPfA/vU6SoMJQyavlQ8d3+xGSGovvlBsfIRhGYfw2HYtTqKLlQAW9gEK7+K3zFXp3nM
p303TdS72tpR/v5e73nW/xTCBnm1XygeR2YWxnx9dqR7NFJjJ+mu6honEd1GhQbyGvCgrXGXqomd
S6RSxjhD7bx9LzTW+CtkxTS702uodcjiZuVsq618TEaU3+d+RMhYtmMCwv32y8RqGnFfwTUFjGzK
VZXqJ4/r+Bebwsy8LeWB2f9YIH5f+IHlfzbZlXUjPlZtNzQJnwd2kvvLOADAK41xhfFnbnSstkvD
bn7r5fzRn9tyOPXG5rQRXIhnCLyE46qWjTG7PS8y0qBQJMjPzLrH+Tu4bkxKV/6G6dHSbsvDL46C
E9haTcY8UPUZ0hdwcLt1Q0HVpRw+OPzvZQztQXQLGiia53XMpMlt1/XWUc35jq6IfTP9nyQsWJYj
kTw5Uu5nVqqOTcBdeFcjs13lAzyPr+YjCBwsXjp/E7WZR8P20OgXSWPOF2uNf42q/a5vKsEEGT9Q
Jz/LcTDxrTlcqhcfMFF2mcZjLw0I96b67eBH59Ywbxkol1+zLdtW/ob1XTnKHThdLkfynxldVmVv
ovgGq4O32UpFNGGe2juRRNMkc9vkubWO6+QUUKkXMRV14edGP1b4tllN5w07gxcbmeZ8Sv+yh9kG
aK/EQKYs9PYvUUajc78Oohz3T7WWCEkZnWdyYU9tCrQqNkHKnRIlS49dFTOzWNXTL/+nF595oXQc
KI3Tc8+o8xn0SrLWwzl/62rWRspGoQfP6LlbFmOTma6mPvr/f0+B33W6T4CJVacM0oAbeEPZaQpV
TPdIm74fOeOlqkzb8sSxNxSHOIAYTHdXK4mz2zykkViWenQ5D4xe+I8bsh0oGK7EQmmy94UwvsI9
8bfwdmvtFPBH3f3bK/wn9sbOMaptG8ede63oaizkhSUf4bKOQzWRmIeWM5gVTerkfdTq+x5Xix2F
Kfx1FGtCO6lc+gyYpOKR/7JgC5Hms7ZzjaAReLngFFZFuxMNV3ME1nKM59ByUPeDEChgl5G2bkVy
zJwgOkBAQEniuZ6G/YM9yKpW9D7GfP9b5zHvrYgTzwqt1KUvosiE5+xQG0XoFGJ7UUAwqnynlCgw
bn3HlbOkJEIUyWTkgPYThLmG58aphHxoYRg/U9hbsAmXRHD/GoJnezjpjopCxXYhD90aMWAnXcv2
rqubvLtvU6gTeQLEq66HAh9V49EZi/dpmcbdRhz52FQepHekmvTdhbUYWIsLuhow6T8cVkMUn0hm
rYMwu8hna3EQyiKYC8kX6KKh2H5GnJdw9zxgu0wMx+gbYJ2yq6mPULl9AYl80hch99b7n8yUW7Hf
f0Vetpla1TZpyvzsLFlRx8wCe16OZaKWT5bLU55HIn46RWcIMw6xHDy4IIj9D5YLxYATGU7sltNj
YuFOwDceazpcW2HxgJPYh/SokU4fS78TGQCvDbLzFEk7RUxK38C/TJ2NsZ392Yk5Qk7C3766SDvs
xwVM1CEHVV7LcwEd0mdMnbjqqZPbRQNt3V/3DDz8znmBoQ+HTzcGCDSKoSAo436H7oI7ouhOO5pd
N2Qv5+pvvZGZdfRn3J9laa5suJradpluvonQUC2W7Bt+3JXIZZvdYGM14oK+eAALB7vvJoPqJ3un
eSN6ggYL8O9bYJy9TjQ9TloWSvMNclyQPER1qWcIeXVO8i0/XE5BVeRzuuQUKw0y863mRa0KFnuD
EFJXXcapRMbV2PkcjpcM5v8xRetXVELh5uxdR0FS+vfW4lnoRMNZfdTVdi/LsqquwCz5UZqKZwTI
nSnnI/FEbEE5I3nRLeCsNytuWoCfWJPoEAiG4Yz1Ga7DzIZLOmCRuAYr3Wyt/PQQa7/8+enzg7Xs
IS8QoNCOL07dTwkkdzW/DIDqnXoaO4XYv60gvMJqpnES4OMMsSeuc4BgcQYyes73zwUtyrEsZdEh
E/vFhyniml5loxUMPkMF3gH7YRkq4zul07AZkw5mTVzwxvxx3RWftCaozJ4QrNSHEMZWGOCgkDET
No8WFokbK+F9+cLAF697r7GkjO46jW3d23OrekN10ZCgZExS73ShKzg8yeT+CA39he7J33TC7F0F
vQJTIOakFGZDAO4O8UeIWtGX2xFTdjzhLNnXesr66Zha1clp6Wi46A3LLO8/IZ1QMMnK1cIxw7ss
MQnwUXoeVkb+hJ3/MF9kWbgAMFFYrrYaV0FrKQxAEw1VSjKYteZv7exsNI36ycbONmFSTJIkvCPt
6WqHNN0zRKg+4wbS/kqylFwq88B27873yRFDccG3PARyQekxJgxzUEP8ivdCNVt0l+wCqwtGTRQG
ucgrZ7llScZoCJMfRx5HBUFfrDE7Lr6CXsvhyS5A4LglH90P1WmD6XrZD4u8O4Lbh8R0pYMoxS+I
n+FPUW2dCjH6VWo8IyNFXKVPkisRHQkNzBDzv9kzlWwkDPPXtQvz/T+3Z6hbptxtjcd3ghxgNmqG
dfR1ZMjD/3QFy9AQC/OvmY16LliNJwexgvhoZNwENp7suLDEYr1y5ddiTuEasPdxxZ0SXkBWLtKy
SH5BsMIqeYzsn5PCkjPlDnCtGxg2u0ac/Y38QmApgATpU9UVqyHUledLP1cu8/N4JBQZQZJHa8ny
dQwpXaviyrnzas7hruMhW1WwXe92uCrM6GXepAWbAzRLQ2QKHPmcfEY5OegrT/EA1qFpWz7O/gn/
tE6gWAI54Ba+YVTUUnwyfppRh2mhIJVftzAFnlfBcbP4jDKB1ih10R2rPDhXbFlws5cEEng7TuJH
a0pcmMzbOFNJEw2iSv5w1BPosXsMfwYD0xhJgG9z8ZiUufWUXLdSWqsKzrrmGMNgVosa+ujFV6Uw
/O2U2GSQLaaWKl57cgiEld2WXPus3cwFhgJsFNksH2xaWYdY51IBkaDrXG+Enu4HumDBPS8NMmx9
0NHODERXFAL176Yvdk7cuDU7ieheQJDifmc4wTz629zj5t33PgHYPdtzurroXEpYtMAfCRpeiSci
/gHf3jXLoYSVlv9D98ao50ExTqDmPyMG9yOsyOUcN4S/VZh+9zzMWaphOH8wJU/0lWY2893geW1b
7orXR5nxRR/9yybIcBADb8lo0gLJFZickjg8rVChHhIdMmruvBxieh9yOKEiyXPVhZf+ARjkdKx7
zPmkjglqvo68oZ9dUEOzVT+SB/wDAyF67H/9y9DQkf3Bit9At1tHIbVlPZ3bGtEtmZw/55I/xO7T
2uhq7MBRttuhNmUQ+Fmuf5yNGdqKTg5wd9LjEktkA4YrVomOaTps8mTSN+pYB1j9YTBxe8OImtxj
SMVD94TWaIELfS/1D4JAymCC8gzMxIuiaxIZ6juhmC2yXJW241MqvRS37Fnd9ZCwnWIdCVKn7MPI
skbuZ/kGDKqDwAFEGgl7fVbw4PO8LrgBMLOt+VL6xruiArxkj8R8sClEVrGjcYirRG9KySQyg7fG
1cMU0TRFES4hi/OFmjCUZe9838CY0aPkXMSgnPAWVLPxBQ4Yc9WQMXB+RZ8YfU97LU0MXE9fyJ+n
b6dA8TATU07nCi0qCIIZUDxHLrhiGf7JSjYP+WgpUbdj5KpYoClKRspbFA9CIKWYLwN9hYawaqwf
Jh61GdaCNLGBfw6vJoXe5XQihMIVreGS79NlBJPt75DNzcVRytPPJ5X87Jvw/tWRFd5ljA6iqxmv
ztJcKj/1UthpZ7zjbih16OeXdLhCefh8ZGD7Dw8Dh9sXSGkb31abqGSTqZLghvyS7EFjhMr9LlkH
/rvlXrAbmw3b+ihKq1EN9JmnUcrJqcrj9mAAW7RusxXd855Ca/lhqLBd3EvDwXW0M33xb2CF4FSi
M1tZeBdmXqkGgGyGPD/uRpQOXN1LxVsNCgQtv8zF+6rA5hSvjaJjAgwH7CkWCbz2EtpixiuXj8fw
AvNwk3R0Ic9z+rLloEgGNn6drfQ5eLkaEtKaEX47x+LXOE34hm2ReFsb4Mil+9wkfjLJ8u930zNY
G3u2zntYz3ruhYRkamtV8HUQ67S+S1kf/OT+SCW92/rG72Av7QImlDuyBJpBbSEL9KSrpjtd9aB6
E6YyXbE7zLFp4TQSfKb8H0FL0MEMZrg48Yb4DJD8X/9m+90IDViK9m3uT2Joi7iLoZphYok8v+wA
wbunQRHsLAb0yH2o4iTJg1z/t5R/IIHyPx6hWQbFrX1mpYuDzegHssTUYGhyCVbCfn+4b5V3Y8xS
Cb2Ada+4QCx/l4Rdn/dX7SBETC+9Ytm5G06mAKEQEcVjxmhSpsnHpENj5bjv9xz8Id5YxXex9C+9
F/x56r74VhVKpaV4xWY0fgJUKLod9wgJ7w7dXd5hLC3xEozpqlU5XHcItfeKMXyUpHKCHDOy23v/
4/IXeCikovyFGS+NueKeiTm8M5kad3YFTJ44KEfh+E7Ip/b1dvTSfQy61WSRIdcEThPHuEK2UV2n
CpW1W08PftLM5PVCL73itf2M7oTireaVlO/eveS5ik8GLzpVcaN1nT689xBle1Mt6UfYsoznsdrP
Qd9taP88kM8St+wSOXaqZFxpQlrFk/0j/0BHskBCacDyF6NIsXPGw/uci0C1v2TKa2dLrwS+ZICW
N65a3ybVbqWY+h84RK3IbgE45DmssuQJZRmGtYH8mgD24K693XUKQ4SLxKNBkMV6xky8MuIgzn8r
P+CGdKbnWTtlHOb/DusYfURA6WsydgQATRhjAgPOErvjffUs9ci8gPPMbVLiDImWlVin3twm/oZV
6UHrMAdqWr9YmB2eo74ZEWYfWt9yxxVUQPjHp4CVGZP5/8JM6BNBeOB/Psy/DjHobw5IdLEZeMr0
Avwx/1SvGPYXYy+Ge9CaiOwVYKcflYbrHjI9qbegddwKw9IAHfod0C/ZY2GcymiCfHTYKcX05CVO
y9Kl56KJMotDxme8h513wnZzZ/ToR2FCyjZak8PiDZc2oMs70MlGD5O7VTLktD04+5Ouso7yogFd
ka1kVylzi09yVjTsmnKU2dor9CJq3/M16txCtzy4sUP2WD6Awxa1uX+hIjFiyV/zJkzuUMNHgmvq
T2mc+X+gTmH7oLhWflq99E+dSLfrkVCr/5ly70NcLOPy98kfnSdF30u/aObMRODw7vhBk2DXNt0x
C3ZpAwzt9JEKfvzQItyhBls0eVKMQLV510LnHr/vhVeOjaTTnr8DY8FS66beh+77T/g+iUTCG6fT
S4ZpGGvVJ1stbhhWr6VWKyeal+Mo7s+q9zBDEiM7QAFC1XTzQ5ik5k8jPwX6nyih8pHvrD7nNVgA
HpAAt1NIdq3tBw3FTVm4yAFOVKt7l4jvq11rnzKajtOJOhSgGYwLfiQYw2933TlA1n3aJm/eh5Ne
xMPtC3KXunnW+eLjqleJR66mA3j89j+KXRtDUR+OW6WxnZptvJeWmRF3dtfoxzaXgldyDGu4WTCN
4IKTxRx5tyq7QYRFCvhGFMpe3waDwmomQ2O9mKXahC4k7w7i8DNYgZM+YCbpVmoONdSFkK8iXelv
k76XIkqGRntDbvUukP6Dchnf4y4AWCD0fX80ZcdJPJWKVnJlyJepx+69orPD3WJs7D67wDAStnjQ
uqa/GtEIkEl11zlyFXu9+Pb0ChEfaTbmiDw02XgoMiuclwB43iuAUbS9tpkW8aNGh+uLmFUuOub/
cqB+putbTUDEC/x1PmeJpDvXSLwsQsI4/32VA2rkJsY17F3XW/HLM/JgaOOGcYfQ931k4qOu4Iyc
TLFp5KugsJ1TXbsNiKqJt+5cAaq38TbUrDf1VmO7X/SKfZknbPYthYLcsz4gs9ALgInEJHDc0H+y
Ut8T+Tj/BgXksc+yVWJEbAFCeK7mfznJ7Efxb4hr6HA+LD2NqHcecWza0zIeO4wNvPrDghBIvO7Z
lFx1ViL8nW1+R7TOxc/B3bdcC/PfcC/+mNsyHAQt9TGFUVH8QSgksGecAHJJSyXepK2k0beDJlks
LiNxTUbMBEvRgv0SedYvn4ewFl1uc1sabzl2pnTlN8JhEn+5TRAAPqZeiP/rlpgxGNmC9nbV3wBw
dMvqyFVOd/q8VtaC65xv5zz3DX97Xsg3HYPVwSX7IPww2nUw3fK4kfl/qtkQ39jBGc9oR2IMVJZK
ldImuT1jSQGR2k/u2R+mCuZ9U2runFjklDdWKot64VeOlcYj104PZ0OqxWVC5HWs8OH91kCzlR69
HfOH81+aaMQTmurVzX6GgKCZZaFm30J6TA7GZ0xLQL9uoT40TJyQayx0PCLvUCkw8IPSQOv08jS0
adc1PUhxjhAifkw8J5I0X0zRUyz5nOQR1jPJF2JlLTLn12f5kzsA9/vj0CL5POGQ4ib4Nd76dpQ0
vY4OGbLi4KTIbXG76dJRCidR5loZI6+WwF6M6WfWVK4No3Fx3WZ3qeSo0ka5hla5pk6Xy/BUlF+z
/wXCOACnsydRdJY1QXip+1XwrheVz+zKrXPkKnA5d55Z5ZP2bfrBPaEHI5IYnctPwCHsHcRGF/6f
NDnaMsiV2DeczpRGyHv9XraDtKWbBh/flEjA97suWM/LrZOuXdZaxlQaE5ItatlWFvF3ZvRJnKqR
vA1aKPIFoWJnKeMtuO0VTNdD1FV6JgPQxRih8c7GgRcqnCYCmhoWKADC8cRwACLyM7/v09gmdS4W
hAdsHPsOIWp5sZJZlh5if3sgQkh/4V1pSf54pAVRKBwGbcS3i/++roH1vZvTAewdIW0pu51U4lVt
no1XNU+EkOWrL67cUKMI2C4vKRINmsmmXMJDNVKiOnJpwEcJcXy3J+Zla3Gs69irfZ6cBsUNErrC
Yhg6IqiafDJHaawvOzKi8MaUqkYmd10SrQ2uh0NlZnbuVWyZwBnj5sUCtNa/nFDRtBcq8P1VGYJ5
xK4LsXi08+G8wBwVeTgPc9Omp0qCBxpeyPYBAt8I5UeEzVY32BFaeAIXCuMI9V6qB84R2Uk6Ckjb
dcCeaLQSpGfJ/JqTf50AsK+HKS9/0WwGZ9+9zUaz5tZ9qbVKdnvKJRn7lXweDj7tq+2oL2RHpHrH
GhizYWl0nBSKBB7X1a8sjGfB0kP/7AOcLj/1FwYdwAbKFrRQqgUubF9dcCAceXzjrHxnAXhXIRj+
py+dKAkYnGkzgIlD1/smgctfI7uGOGP+6WosyeCC9FVNnx7IIGYq3MEBLY/sFaur6z3Rff6kU3t4
33uYxLfovp65Fe+8wJQR7c6KSSmDpBvRM0e+EZODVvsx/cZUdu6jAWPdgoJY0Nq57Uo4Sgbrx1tD
ktvFksHkIJ+Tln+6p/UENQ17Y2dsAWTOYAaIC6WF5vwq0ELfm6fLaBOWt9pFscRz6O59X4OpxXVD
mpJRum1l8ug1mMRloBem7SxJD26Dl55RkakavXCcoEUaFVN43I+VUpUEZXglzeUImknCS0z7CO0m
KA5PaBGhIGbmwThob/hCj9ZVfbMZ7oaUFFMHLEppPVb51h+DSMVeIToI+K3fPi6Ii9wyO7TE/S7G
btdEUpkBX5e/5Djnt+rXv37rtOiUUKrjS42zAudpreY6PVi3+sBd9f6sYBWiSBqIlJDoPYMPh8LY
J2WuuZMTJXyHKJmv3MijTCj1rIvzEeFzRbFmXD5IJfJFQXBHdxoxD/gTfuCoBQOLJeYxdyYGnBM9
EZLw6M5u0z+EDuXP32aGgI05lZqpOK8+K98almiV1ODbzksvCZBlg9noJK+f9WzKc+430sX6LZ2U
zw25kZMXDTM4Yh3rcywxpG1c6NFSu2o2hX6/TtqbxPRC9gh2yh009fPbIFZbtpb3qVRXtg8ojx3c
rUisy8CFcYtf0nXMP7YtEmwFSv44KWEEQdjku7MHP4w1QofpvlsTFI4okNJBu1oqNZd1x4h+vjDz
t31fm0tpIFVhbfjHnw4/jQdnR8xPvHzSHpRjdFFzVcrHKlFmk2Hjg/npukHUk4/vCIvOyhxgo5Jn
WmohOi4rYCBiUWoKCRnIwhD+g1xpVslY9EuP8TpGxJScsXUdRTTkxnHtJZULpMCIDv6NOi9xvhUk
vAg160bqMjTWFBCLMOJ/usbv4l9DKy4JBnBY5lQV7+hEwec54PLroFp5HSZkC4MjFRmm98Jxn2Sf
N3J1rkan6CUMGpBBfMZQZOwmPpwW/aIoU+rKGO6a64QsMUzO5GFSmAcdzbc21M9Y2P3hhFzmRQIZ
C00NQEc0pCHhLO09qdNl56ndyFfENhFSBoFQLlb6vSx1HkHNPqHNlcQ/s1RznxUHmiNfYa2QbM1N
/mnPfyHn7lK9O1dAwUGmfRpkVwEilgINh1dqP1IBYojfm8JURDD76oHyWmVWMlsjzBdqAYzRKHhg
zsFT9pDDrHSS1nChN2TNwcA8XNIG2hjNBQlTaBchmP18AOnEGBx2kC8vk8WHHwZrc3j5jA6VHYml
mTQGwHC7y21wlWWAdugIpVx6Ou0rUBWoeQHNpJZ0cgT6Gt9V3yD4QfCfZ8NmMF/84HIqwB17bz3R
sRDMZo9RoKj2XNdZRRQ6Z0XLLMqRpdovVfSZJdRfvDFu36oQ2UDQpgd7r0DmIg0Nj+njdiZj1NSv
boysUZJHrLJ2EjhwYmGS4VlJrUg03ZmiyvmdD/aCLcJvvxt7zZVL9cdGFirT53kIrxp+kjdtKrBv
DUrz5RUzQgwnCknzBNTe1qTYdVWNzME5kRFLQDFrMAfMwvudeUzSRyr3ltv2oJyP9mkdrRWoLuyR
UqXelUrcw6ZS0QAs4Bba+9ocPkykO+qASLVr4Hd2hn0vCoAqPUO0zHyOewvU3rKI5Kxn+yHIZd4t
xc4MfTgsgiGcW9AzzDjnPEDX6+4vFQJrMI4Q/AFYYgxNSF4nRemKkMgumPd18CrG1j3awzZGEhiG
KiVglpgog27IHlRYGTrq/ZMTLj3hKc51KkD41uRg9Jur9cxtopd7VmLhhwsr2EHy3lGGUCzbKut7
7EzVmwlyiwI/obL3CBfk7GUr/nuq4049Ts0DtosWVhG917WVldoFCJHOGYWWkLuUur0vO3xn6C6K
0SHwMc1nLQJAt+cK6rZLhZNd6dWT0g/0xv0K2TVAppMKQuyGqQc6B8EEuXVcVOtFQsrNbeZJotdL
FjGdIhIx8p7VbkpXnEzYYFN12E0kRfOgMgyBdCRCS1XL0avqbADfyHeVaLGypPjYthDOdtU9/K1S
tg9CixFp5pZFgBIdq4btDtQNfQqadovfR0aZrEWOShfrHO95NVWlwH4XI1ueB5u/CTyYbwWo6RQF
Q4vXBL/Vryq7e4+5idj0mPKyL4p6azpr1aD2fWbzjl4pwTefoutj2NYNFRFssRXsuqCkb5qlwCy/
dHnnUlK4QXOOY4wUw4ILUXpxo2jInZFkoK30/2wSnJkcjf4dIBYPKSV6mg/qJ7/5bhp+3+HOoUbj
8oBQT38ot3ZyYC5TxD0/IyEu112JyUGZoClh5XrIDxjGVKG9ZCzi5mVdcCXS+rcmmCAsTKH6kuFJ
GTEaj78ndvQ5AQElw+XxZK3Ibd2Wki8Oyypot5+pybwQIp6ZD8WG+LC6tFgf2P0gSm393nOoXotB
fiVEe3g6O/ri7ChHt03X4xs/NzxXFGXGpA5+slLytYY3EkYYOgl9WDkpfj2FJB6Dj4s0Mq+DvfRV
VpyFgshqy53O5XGquNxFbfitRNPxa9HJtXoNOR2s3m2kAj0cVsknKAH+EtEnDtXbNheX6R3WGDJ6
Tjk877mz/zVVHnSMrVkbGw9Hn08fqJC0jB/HZEcguMpcIIQVJ2cAGCw1/5qEIEsuXKldGB6Ss8zV
Cv1d1Z1ccQRAr+aLjWKdn+peUGLmWrOWTCAKzhQ1J+iotj8u94mxIFJHr3HUw+ls0h2QE8jVAP5O
Tj9HG98lSzkEiJaP8dFqex8dKY0SOop4iUZK+i/7ZcNdgpkfdcyGYhaJWj9mCiwjAW7Hd2NfJ6O8
KI22RCEEoawmF23A3dpp1Nmh8MmML+3X2OXxuL65PEqUfbXHO02PmTzDQ+rGZJ0Y9MK+PnKARM7A
SX2z7IA0R1U2CPNKHtqCDssvZgYf8dh+iW0SOENkfm0lZEUDFFcdNdUg2B/b0l8WZZso7xxCZwjN
poz9LsyVYYlntW6hdk2bF6V3S8Rqj6q+XvWOCka0RuhRpXrcNIFve4vB0Um8M8+anu064VQSU6yZ
jTosIrj5ZnXbGOmUQcE5bptCvYoeVLpJ/8pcmzn4czybuivWQ1lzfg7h4Dp4XH/tHVmHTPVgdWv+
M53AlGmaEZ2TJDOzuN+S9vNVQfv53hoSe0UhuA3lXkK8EW3jT/jaDR/bZeTeWAld5tIeqfJr2eI9
ME6CEjpmfWIDSg9zZrVpPeQrhW+Hhi81Yx2U2ph/ue3Apn0jbuyxQL6uFAmMDPZFtvWP2YWl2uMc
kWxkFjsCnyHTiD9Qt19PSK3iR8bzdlW8p3A1FieEzsJwsrARoYWowog2lZ9UjOLziDEjWxuI56Md
DoTTzBEtBG0kk1GX/xUZieMznun6/KaiDB1dkQHEDW27dWbr6q5sbed3jxhLiGqKiHZgZC4F2DDy
T35+pI6hDjgExA44oHzSJBnK1EkwVH/86nKX8Vx00PTA8sspwRns4ryOnK0tS+9U0bxLkOh1XfxM
3R87fajcDeLiguJoNbh/QOrAeBLxcdVJV5XjTcaLjxMlzyu8kuSHIO+EIRSoPECDxVSTCTgu2zkO
cw8sSXg9HDl1WV94uO7h6MLJsI6nFG1DCfJnKIt0QiBxKwTRGuK2XJGYjlE43jgZEElu1iKfQUdg
XgExo4bZ6eto6t25Mk2XbQYnZQoxrfA880Ay8wl/ulsj1IuhxITl/2WFd25SPjnNHiMk5uCBnIEp
YOMcmyNaoPl64ZqkZ4uwWqxMPxg1eYxQECOysGPkL9ACVzw7I56xJvS6UfhaG1eRFll5gdTaP9XR
Ca629lSDKp4ioCaOaB0X8ch+GtCMYtnw8lkflCywXQ8K0+rk0Gn6ksg2HjL2vhgj1ulu4u4OJtq+
aFFno0gVIeavy8awwcfk/uEqzlJffWbrFVgBQIIW/fdtf4CUTWPnjpkD1TguhQ5avUSvNfGFVw4s
rynsHI7Nh5CiAlxlCt3rIBFFlIycHIjugiLl/n1mXzTNGi/Y0y4Am+35yfaff+ZotipDK7P8D51T
WMdO/vc1gTor6Qct8QZLi38rCfhUn8K8f49kJlCHhjrhxzJwC98Blvi8vfR0QtpOlUWrTlncCKgg
1mTIVuKZ+oa8U8V8HUILMNdMuo+uwVsxRB+yjwbO9otUdmeseSZs/EAPobN1L2woXw/xA3k5vk5s
3RPJLbKhhcO0i0hs5hvQ5TNLeXoD1pqgMn7qfDwzyxH3Lz6t8ThMVfuTPgOKMyYDvMN/k52Fudln
15R+NFTP8Q2Dqb+hTwmUgewPRCPGui0VlNs9QGKM2x2214/g+aH/8L0VV9VTMioaISUdatYPpcAT
NMGi20nB52LmzcsT94SPiAk2DtSF2QIpVVFjgMs/XrS5MQYZF98D20KWBBZTppFWJAUz5ShK+m+G
FLHTC0n88ieyYsulHzOWt3FBoWORqIiEdJ8yWuK0dX8nKpJ+XOwzHQVAx8mzc5tblx0pxVsSK5jC
hTfb0IKWdcUgvEiPo1OZqMTOrZdk28FQl9omYbErlDPGJwopsEp1ssV97+AtaCgXd1EOmjBqKVec
/xyk90nNhX5vSYzSVja8Is0TX4DKF/plajfeoG7NW/OAzCfzf6BvmnmGVXcPRpSyFAbUgN6zkuxr
E9LJZRDLI9d+eLAgI79yRJmCvbtZCbhBrAOqTsmhItfw/NPKff2szBYYNqM+KBPRsX/nPra9JQm7
UGnyGK2WgpEstzNU17MpW9qvVx/sLAJfjVsLALF2VfUsZSIo/KTIt8GHTIEuITa0hd52OcMj2X+R
3zOi6R7W05mGj7fq3dabCyxaFdBthlJGuNT9o13lV82WxcIHSJuh20FaRRg6fVgw8pMiRbYDerwd
dZ3mD8DLil4eZeOL01rXGAwkoVVhqbxAd6RAa7398uVjt2msC+Eu8Sq5tatFDoyPxzfc/dDp0fFM
R67PYgg+pxS8FRrVGhKNiw/ap3LEaambUv6SpNfu6HFsVqsHTFb3vRLqYJXYLKx/t5qwyDhGnDM9
/sJOnXk4H/ExSLX5t2Lh/k677tuqhEcOL0uJyAFUQrVqI7Kl3CFLvf3K7UAZgh8/D40euocKcuVd
Qe+ChXNpZpDxlsMy4hd0hWsMPPDpm/cImi3Ckwgj06al2kUfOsMHYzXbiCsMp4aNP1xGBPFn4C/l
qSCOPRhQSQFXBk+pU22kV2wVmCe9S/NQELIrjcsnepjB1rdjKWCU4DUzJp4mcaC+97wMud26zu9J
C1bulYppiO+KX30oh6h9qryi4zUwaPwj0YzFBAJ3vYCvuBwVcDPKUyEKS2xkZS5uR0VulWtJIoox
otNrFaGI2MVYcHxRb5TqJZjXlHKaT0cXJS/784f+uygRWJYpQD7jSDCpOvGE/bEiZwqtlpkvAlYJ
08ggG8vcoS2IpY8jgVJpZX/Atx8i3OmsPXF6SdqlfxyoJhFYzddBkaXrF5GfW3woeA79qrrDl1vm
c7gvl/9SYsYeureHeVzJIoNTIQHhMRzgiWKc1l0ALM5PVz+5Pg4g9y9Rt4gBnO0I4pUINvHtO8X2
2XaSa55Wl1YB+bCNs+tAT6IL54IWnFeOzuKyuVcoa7WM9CLbqVHpuIsKODuif+GmoZH2h7PiToDC
CsGDlWUY3qlBrrxqRFaKVgJBTTJspJn0rhp3MeIrEh6ZKbIXGlqX7WoSkFCDlOYSHVg4XYq98W2D
RA7jTjacv5o5PCzG4aUmBJURo3+t4Pexsh571jUdLDIKXtLOhRL4EmmHcThCnPi/QnfVD5rWVnoJ
cNiLlmlOBRAEW33zOTpyVmX5ouhSamwGLM2w5PsMvPiGw1AT5xkh3jiqCv8KiA7om9qNWMpFyuLT
2betOKROeio7VtQ/JHs/b2s6V5xFPrlv7u6IANCgZfMWQbjGCoouobdPL6TSetYIB+ftqV3xvfIx
VeNhOEzgqKkOyzKFiFoPy2gDdYk81sqnvCb1OboWamhYjuoZfiEk2fHuiXoOHUn/3n8+JWpd2RS2
C1cjQCNtHKSJ4QnF+fZdpV56UBu7ptZsPDAxL/ITmKHJV+DQfRLVEvJy3gdyUoxMnkt++mtdIqRO
WaQ6KtIVN0E9kTU/IIxhvU7LpivXjnknclCRdbIP3zXEdT2S0og/Pj7oX0JQHTFyRkywJr0iDDKp
+Wzb7wChxoRpR+DlVYJJSKQsnrQCLSVq/8nUS3wtrQHtzuYGlHY9jtiapXKnwGeLe3hxplgJbT3T
096nKWDlSwBHGoQQoOvZxsxQbtcf0hKIb/MKbX1mv//6+IhqCRQM4EOXNJrvb5mh0leHUUffjjV/
6/GVRL7yPYbstFy+8jPwOZoRYdD5KKWyNDoUe8XtXadFggh0xyedMR2VEIU93ZpH/L4n7sDkQaAb
Tq1x7/lVaP2uRJHZUTWctEP2Qd1rJlPVw4JRoqoYYx9b20Nih3WbcFozAuI3u7SkceR26dWupUy1
VqXUoNJ4njnOyn/dttHYqg1PMiaSKDEJh78ezPY7bj4ltpKp1+RpGlY9NBBPmvaZwHAg3CE+1t8j
+fvhISjhb4IAtaogO2p/Y5Py14ubOpqq9wCZVFFuhPikHwRRm8qjMoSdPsW3G53boFezmaparvPW
8oKs/o4/iYsKJY5Jb5Uhq40ZOx11OBvTbd4Ku0N8TVq8cUGuZwOTYCM5ls17NQwqQLR9eOVcnz1P
KCfF7sYk/gq2sM1TJGe30vF5gPDvDdY8CU1krERsW36atSMvDHeDiszwqVD7A5WUFoT3lfStgwo6
UlM1zRmC4T68GIxW7LhDXJfR4BOGamEcV50gn2OEtliLfftJ2su2OBOxz6ZcwcJCkccm2hPWExMI
aq62fqYq0C+6EnIuKPSo2mne+eMEhlpE1Z2lALj01MG5Qukr6tUhYpXhDcM3gT7qMOzSWS6TcW9J
V7Jaxf4SI6ZB9C1v+YCfyfyaiVI4hccKD+KVUhNsXLPwuefZvSu6/F3jGD0XmsLsAtSz5crmp5Zy
vPSoW3eiarMrbcY01Su9Qt9ljsFAo7DpsYcTde6K6L9lYWFuxPCaNAKWb3koHza4U8z4HbJNRvnw
M4P4fb+SqgLnvPd/wR0+eWfp0mgR0cZCxoUWdTMVxk+ax3z3QelnZG5okYdp4yPBCWlABtSus6xl
g5BVi/UJeRw6yU7ZQz9LH+isTm0Xj02mY18iRy3vQqQrjnhqegayYT4Nxk4ZVsPNQeKsHY3e1SIm
xGoGpeUHlGY3MBCqrf+u8KCpW9b/xxyTGSmJNtRsh9OpmiZzQ0cA9vqZA6MAB4nVSSS1jFNYld4C
MXmkinx/4SmlvG7W10XfKmMI9wc0ZS5qAu7ST0pHIFrx9xiHD6uGZ56DDfedVPVjHHnl77mKWZb8
amwqjTwgvTv7TMnqtuUqFqazS37CnmGdFjOFRB7nYGqBEX3+yhACJbgcdjhMYrUxULdx+K/izR9K
kBl6H4aOaqedyyV16SWInz1v61z9KmvfPS8EKrVvRDa6vQLJQyWmrk8y50kfBvOIYxvbQ8Bgk96s
RktdvzQqGIkZCj1NkOt8pxkBopxg2qiPn3DFiVppFqXfQ4pJ2HQlL2s2EPyWJJHXB+hV85yUZ5kz
is5pRZl4783/Do6sDT02BT2t28HG71TC/fJjwyRi1F+pQz9CiJZScO/LqX56Y/jqVWIs4p1t7yxR
KeQ17W9CVF7qCGQpr6q8TGXrigNruGWyc0qdaECk+IggViwUCwsqOqgKNR+YFDI5tDArlOWjsCAu
uFSIa2CadvgWzMiIrV28BiS3Xu9dOZsUEvrkhRs62BsmF+4gCWn9NxIHtIkI6T5FA5KKPoGeocg0
EZST6IPqdVtKRek8kxRaHr+KwxTOenWhGbVI3eVaQmiFVFc1R9QwXzLLf4YepRH1cu8hskFif2po
A8iuHCcK5kilo5Q5vF2R0Ho/IavgukuDTJQ8OS0Mrei0CxNtemwGpVGNT4ZPkxkOJSpENN6OPwPj
xH7KH1Gf1CWUKtcX8H5siEisaVTChDO/nA1sxEYg+6l4rkEyGHo7c3NLD5aqWscw9BKUdD2g7XMB
fbgPEirzbxvP4V/16QQTGisxkB+bmonV586hK4vzXZI5LrkVoUa3yczciG7uORtsZVvRRwLvD+hK
S/guxCftfkbDMM7C9kqLhXUxJ9wA/qEyuJ50ua93u+TjRUP7J2RxIZeYcGLf1C6XiMxXkinRQNny
Bnxb2cho+OmeXxZIWNmg/NwSr6r2QbY3UzS1KCrxY2Ox/I49aCmVPzaTGBpNHNQhvpiinKQ/QzFI
k6SluhsDxgarwayJ/LYhne3tyAPpu4058FBTo7CoyfZXBXC9ZeZnGq2cnO8+l79LmRNyH+jODIl5
FS8AinvlsSJGQ0DkfLyulZ2B/261deoxyC/e6y76B4DjsQXYwNaNfdsj88348smHD2YJL/N76psl
88ZgZ48jB/ZVBQTw47K72ulcYPyzvya5cm3XNXXggXYxtSlv30OaUlYdUeVL/Mr1tsOXg/gaLBMD
Ee0pJ82gxu1EbWyUpi+U0Xs8X+vO1iU2YxOjYXiz8kIgiIFBly94OWFgvGMHhdeEK3xs6PlASl3W
AtEDiS6INY6i1O/vo4MQBHFM/FDDKL1yaMPbhdAlvNbCEZj98FcT2qTj4sJDO3aj1k0eNxfJ9R+x
rJgKV2CyfKC5FOf4YdZe5kyYEW3UpLbuqR5rM8Uk8R0KkdR0I8o6QxFHA7WcRNwsPo7OiclJ/BLM
bSLIlsmZ+30nqlg6JVYbX0vnw1xUTNDtcp8xPlDJqbb8SBWPiVNGGBWzNehmTKC+laoJ++7trK8h
yNvKlwOhJEsi8Zdlchhc0q607xBg8JDDzNzH8cBm9Ru8nvoP+X8jkn3xND0hakn1OPxhNh7efJ+9
T06e4In9ZMaMkbq0fAwwVfw6s5bp4se4bm1LwLjEec/fFFsWm8Y7YmNMvNRhIG1JNu7yN25L+CLY
l6P6bRXjhxxpb9DMZ9k7V5WTJ3WzNP6OonHIAMjYrspJiTsEUtvYjllr3KYm9U/3XQQqcre27+C/
MBBze5CoaiDyO1qOuOUkJZT3HDQTa33m32A2TQNpWPvpCl3hCcVYm7mR1EkITbcVQO9SOlA4xCr3
LkZFkWoMDAXiE6wOqOxMQ2+5jWTsCqw6a+o+1bhOaMTFgaHQ+cltFpqBaQb5X7rvYEg68dPTScKS
HCPHgkQdwjPTSqTHOanWPCklpO4zKvM4401kRNwVqfuoP/ewz6RrD+bLrXxiec5W/fDEDPGD3dtV
ScgQlFAsWgwaPMZbORUO5mec3KvozsQsg4GK8/tJUlrfOs+P7dVRTQF7CaYK00AzgTAcobAnKp4/
P2N5B/HOoaCptx3HTuTq3ep5cSq4H3OVwglYSlqjGdNeOLlY/kkuMEH6agbl3/zL+7CfeloLLMcN
z66SqMsBY58rP2nW7afNedH2Ne4MGLC6E2Ph04AmdnpJEsvHGc+l2DehFD2zIL2wWSx0uHdTq6nO
qz/0MedD6BgakJb0KMl+3ddVkhW9r4/BFsADHWTAFQ7g4ncyTCLFpmdKQLCshozOCbAMRyknRtxb
bSdJyrlkeSMZiAgHVVJDrcz64aebJwYPNJ7shWPevKWIva1HAYBTexR7B10cYq7EwVZ7jFGcE+3U
PYuQnGyzNVblnOwuMMZTGTEqXQFkSr540wM5KOhymAzbG3hmE9KWLvHmVB6ULMDRlxbdmWLMj8l1
OZ9RLJ7bfKVpQNsknmEQQfqTeAwRLIhZ4Ik+fqL2hEh1wvmo85ycAPxoNT+vuAmVmA3yPrZwf/kW
nesVE3LUNHMwDa+r4DQ0Whb3DptFSSdz3jQsqKfLuCVNnIgjlikXPY4BvMXqc4OKfjHXsb6Sn0Zk
RCJSJ2R+OA2FBPiYQya7dgz8iTErT7GyTul+rx0dP3fjG9W0ukKQ0wXXoeB0Rj+Gv7rFwH5Cbinh
i9kN32lQNC2pOhJd9A+DcdCJBs6nYABG38ASfTemprZBuQVbyXq1Pxf31djr9BHi60CKPK5Fj6qp
xEnyrSFQ05/Wq/K04oDFyWwggI6+grvPVPXKe71I3UHoXrm67Ou+pFIOoxFinyavY2pUzUWHweNe
QsBc6hA8rocKWDoXIBpKuO4WGLNxQhgzaC3GF94upwlgaYEUOqBq44OJ5fsIZ54W8Zn9bINuZ5Dj
OO4uEiOdvA8SVFTyNV+LgKwfyg+sZsaaSWAabTDzFtrh9thFri80tY7f358bVD9+1ieY/On8gWxq
R/lGU0gVrWtJWCU/hcm+mc6/u5mFspAP5JBxjm1Fa9Ru8qx9l+JboQFnxNSbgit3jKwnIXbo8c8P
3fNKPrOglhroXg15VpSWgEoAnmGr79jEPXU6zyYlbRnLGokqN8jHGQs8yQyUEqE4gEUU+1SQ8zrv
FCHKUHhxAkJATlj6OQcgSQpMqCmsQYXxg73xohVKi6yuWyN2txSFcF+dFYhyWuCfoOmse8ji1tPO
A0fGZ/7GgdgVCoNQhr9jUSN52N5Xoj/i4/FJ8uJ9CdpvpnsWrhQO2paSGQzoF+xaAU31EdbhBoK6
xp6vsYfw/dPJidW93g5QpEnfhEAxrhEmYvIF26mB8M1LfqVg0MYywUqhHEzDK4/T/hVi85/0/k/+
o61evSHAyN4A9JZSEzTRds5sFubI7c1yg91WPQspkSJI0H9wuLmgS0V6mWOsT52kzQvbjPu+XvD6
AczBoy74PZY6ziacEQAAcDvxitZDh7fzHMQGObjy0mlxdx0ow+prpmR8lVBIXVpKkVA0mq8HGNfv
mvvq/RRwRVqorcpDqo6V4Y4fi2R/wlD+/VlnwgdKDH59055HppaFDCmwNrMdh8o8XzTnAeMpK/4z
NYQwW17Oyvdl5mg4QbzKtkq1lmshuDZRhvAsGkmGKFoGpbn9rLuAL3rGjle0kh0dZfLlRluX/Jew
LVex1h8uFz43MWn7xNlHpP6Pmc4h75ue+WFdzPuVDyURVZwxcaOp38uaCYGWOJnFPuWGRfO3dIQE
0cdfuXIFKYRmVItFtSD2XQ+n6AX9umMyVbVeJduVyFzGfgYdkw9ubsZJqvuW3sdrCA4OQO5Mw4LK
jD54GLgP7N+ME7g2pC2R5d7WbLkVjMEaOEr/5kQoN/I/EW4MserGQIMp4dqmYO/mricTQJE49Rg4
H/w9GEAIvDY+IFajqaA2SuOSlPuzJFR8Wlqfa3TUok9y7VaLYJtxuYkAscVNqg36wtRffHmmyV8l
xro5xvR0zW4vsTgoqyphAreGStQLMyIJkLvvELsWJy/TAuTPLoRBL35WECP/BIaxipDhhGqpKecX
upaVAc13Zh6aDu5EfUiebgX/VnWFzIDrEPB7CTrHEb71GytMHqOZch1eAho1BD2czvJ8Jn1YGtyt
Qj/hhZ3RPyqbvjs8TkcRAmmSwZcC4qo/eNur55YWnTI1cVQFKOB5LWXwpN2uGB80JyEMtZ0sQaei
5ihZRN4DTvbKRlpi7UhHV/I/Z1IXcosvfoLfKZE9EdVSJ/l3v6pkHx6rtPB4LDHwDTP3nZTPzaf8
hITicM48RuhHc16eICl+FQXSg5A3lLcmaky1sj/KRPmD7hD0Qx7zfwnIMXZ0lmG5XOrwm2HbOFix
mMkCHVQ/CC8DG7I0GKNew8pKGgriN90XEEnGWz+udyIVAiwiXbSa7M3BKfMoDl8tU/64wCVknyVC
s/+84AxAgm4MLrba5A1++mtnLdjkYF4SGt/VTgYowchbS850sChYMt/+xnvstirEcxoODau6oMud
EpAlHKZNGFm3bcEpBSDzDCuHqMI6TuuumvQSfYhQXOl+dQ4efYpIz+W4G0miJ2ugMXehYKwLrIS3
pzlx4IsCehcnhvabrwLsFmC/k6bTD3reVpABNyXUNgWwqPomuqpYLuMOFU+47Gfx6vT37fhHSbyC
b+mHE8ViOFoj8hFO/qcpcDiXIB6rcqoGAHRs4/+1DwdvE+ouis+s2Ceay4U122ATep+kwV9lpsAv
xYKYg65nMPdT+su9oXvEg2CgW5ldCakw0osw1PWHXRy63Tq4JoVCBXC9HlRV0NWO19cvLG9b3Mlz
N90KBD5KqvVq36sC4YvzTcwwKbCdP/klci56O18CQPT/QUELrwNNIcM36Pcn1uwq6ONRBi4QW+cS
xGmNkQMZ9sNHcocyRqOyukQc91dhNL+fGDoH50RpGGYeWJKk1fNJ9v8b1agbI/3iZuStY+34ScBM
GcO1ZDH7NOPjg8b/p+EwDdRIvAvD27OU1N6lSvRMbauHzqIjqEWYQe/m+1LSmVjYWq6sy2X1IS4/
gIHmrKsCwt4bq3gvP8qP6BrSWDVv1ci6F2V0uvq0Re94amXTTiOQI7L5bq0zXATpM4YEA+9qtLH4
7xwsnBccv61MkKkgCvdWECIT3RGnEkAGX/8JTecKfXNe7jZEa0XrxlJt5CJi5yk9dj/RFJjk0n8r
ov6/IIUn29dF20Js++pi+wbyNOVMB94VY2CCdwtK7Jbi9Z9SAKDmDco6smVnjGtdNNUFuahXXw+j
GGh4wF0hNOuRPBF3jYfyD1Ylsw/45clKpO6RGQFdEkGuASS9A2lsWU3zxuuXoMPY1nGz90UDmKn/
zfsCMlhoyaxXPJ5+ulbB281jyTBSNrtfn6eTrz9WtWUQ3UTryxwHTCzePcwBwshvEhmnCeqNUN6B
blqNMrjdl1FxOW4m+v9KzLMBnmZ8TokDZPj7gdae1GMhBMxbQHc2N/Zej+r+b1AM+gUm3FNB7YNJ
oqobYPbH3nRPVx0Js2X+yXzIZKW4BCg0wjsMrREmA2FvJqyKDr+3TZtr9vszdsBqY7xMcXvUUgUF
v0oYzGDfRi1GoZex4dZwLYO3n86w/RgdReiQndPKNI/Y/+zOs4uQ36+8V4N6q703KfBwZoAhMppL
Stg1bMHmrY2pFYEa1yUT8+kwjtLFlCe7u/e2yHlE4iHalTmfEbdQPFnvB4MSp6FQNxxPwv69F2FZ
7z7CEcQEeJ3LUlmr342yUwX46gYZ4bL6S501CnoRXkAhYUQxIotlwyM4bsJ9MeMbbdufRHENXuct
0Iv4il5b6vDmm1nlRrF/9D1nSAh0E8B9o1I+SG/IeX142Q81wfrPlEVQqDs/eDN1bePVkSgiYaXZ
wXv9p85BIpkm/m4SA1X9Z58Jrt84T5wUlYL6mLwqx/FTSsJpGkYdGNZnOiZDuILkKyz1FzQbov8t
Bz5bO3jMuzWMWSJRL+29tEq8v36BNuMCVJbWNqNYEi8T1w4xCb+YVAKfh2O/FEEqXwGBJ8Db3bSu
Qb/cWCZ4oHywVjZqA8dh77aCi70Q0omyUkyqMWnON/Lw47jpY0K9xf8ZqV+YHaak6lghUyq+JeT7
X3Fn87lNHe49UFigqj7DyqGAmaRyu0E0SaqT6uSwW6jAXo2RakQT7LzHUYauEnlKL/eBmNy+G1ql
JaLeCjQ5vfsDRhzazfax328LGBZ1UonfkeaFIU36R1jztFwACb4o79xVjuslgGEL5AjMjPHoN59I
OULPVdx7oWXfxEUBkFvkBKYO450HFzcHiZIHelM5KtboDmMIJETm3bXBEVDdSQTEBRaGPFXgImyt
5V4kMbLKs0GkBaZkh1PDCOcv4Y8zRB2P8bitTq1Owpvww29HtbEy/8udaypKUhD5Y8nfIEEEjQDw
4O9TapnwL7qG3KS5JnGts9VaiLypMJY1l6dVtWGigdLmgU2zcLk0wk72A+FAeon3+/u54kdtt11U
/r/KZJukPIw38UTuRHbPiim2xQN8lTDt64KonQ8qnHD9ty8ZK/LXEng814amQLFN11MgLwYV2L+f
yd1DC4WiqbnNUiTS69nFcxHKM2tyTZVdcuF1UMJQvcVA83nxHq3kuKu1r6vAEecQAJMcv/ubEloq
sUvYQuzwotdNEwsQJWWHPfy4Nj+0iFqkvvvPh0g6ceKaz6zDErcP2VlDM6SyTwfkly+1eRpgxbzu
R6a3qk9T3/IJIEpFo4Hq2pdV9iHKyso/xRQM6EAZLUswuPjRYLk80P/iMMKZ/FpQOgTQqGcueLSL
KvGXx6rVVaQXgIQMNxyuQ7N2ssGNreFL0JYQcnskHt4lgpf33S71Gs51plkAA84E6XYoDAZgLcPQ
4uDXS3fDM43S0TSJTS9jSTPpHM1GIzkLbwSi7pQX71pjDmWFFwG6jb1BhGZB+mYfe10+AYVX2qjB
L36jOakz4BOL3rq+wL4xtofRMOC+/q3nsrkT9gIEm+yGGuc1ieEx1vQhHV6UQqbfb4Pt15XRA7wP
kJZy0hHe7DBIT0UNd/ao5Dzg34VlseR3bL/rYhKd+O31UBA/4bYTJgAWhBnmZwBFw0kk8H7ZHkvc
CDGeKY1XIHtkTQqe1WJlG115Jr3bGPDMv2lhnFkoY0JT+Z+kjuDUCbDp8CWDum+KwiEogMzBrO09
CdOtcWSpGQ1BmIZo/6KZQotRnygaD6G+hJX07u624HkDLwCwMqqlbmmaOxpQgdbTYLHpcVTXrp4Z
hQDusExRiZ5C4QAzIMf4lyk3gVMN55j4kQGyWJBFylf7M/vI/kz/Vnwc9eETik8ZxM56cfUXWxEm
BXKZssJ4h82t2XPehpFNUVA8A4U/whQwzO4XzYV/c9cCWz8+zaV9xL2ekqW6gAnXWFmPLhSpS7lk
hOnMKs2It4Md4cLeST6mGOTw1EbVlGAmrSvctcR2zFuwAWdkLRw0DAMNX0JFAIbr3ziq82PlogCL
iVaEiakOculVChIam1v8Wj9d2+Cu66U4JZIthWaYDz0qTYJ7HYoHxt/NMRcC9rcyHFuvYPbxNNRa
XPxKTCwyb9nyPf4XIrdtVqXzaXiEYhFCqrDQKs3Makt0o/lVJykYG95o9FFqz0AQu8ilPwOlQXDR
AUhFQDxbaCIEGfIT7ICby8vYfLEp+8bFJawEwx5j91LXNLC/bFOY7Pm8+IsJhm6gkQ9BDOacV7mq
EkAJYsAMAzJfhHkTifMjkvKaHb0FqPFKDr+rROyargJsPcluREKKmcWpVAWS93XvEre4NLp68mC6
NJ30tsWvab7yd4pr2mVhmSSsUomj7UXOGxQrKKHBa1GjI4R08Ws58ojRfHNUvUrzoLn/EL4Zl9ma
8/UTz97jTPJv4R21XKp3U/b5zCbQvfQX92Cgu3tqzHZvWphAmGIMzW06Ed/E8ZnLaSy8J5vAbAjr
BW/VzsWdit4whsmcTO15NRBwqvgxzjH8pnhBSoOi1yYk8UOa1PJM4VdRlKXKoKlTjAqCUZkVkHdH
U/N8tth6wJOBmU7gIsZKNkqnC1l25g8qhYDYiVp63LsUSOvTv9j7B9qTM8CD0hCSopHU6MwL5IWm
n6w+A8qhT1dSg9M8rHdY2XTvpDJTRg0eI7uMdxSO0fgcOzX/zXfOPRBVxw2T6BnS3V2JcD1aSsqu
WWiFl4VbQnYHI7VrnnAbOJd4jC58HWuo/Xre4QKcPJ6DCMMd1/NJVJuYai2iree9uutQB0k+j5TZ
e72tb7DDuT6ggnY29FkBBBdBm3UPy5UQrhWZkVt5ed4dW5k+Baf0RkRzp7YRyTqWuKIYR9dCKzTr
xaq+aY27X/q6pdN7Kj3qTe1ZD1jRd4TaUzixRTyCw3rhugxrC3MiLNpD4GM7eafhQ4yL3MZuwfeL
7QEcajyhD6HT/cn0PEL+k7ZIr/y5dVu7iJHmTkMyKgpCfL93qWzkYGeOEJrYcol0yQLLXzOY4tUJ
Ijpba8a6UeKSfOyhq7sA8rTgJZLbGiQGwLsBkD+e/iXifLpnBCUOM0tpTikZZ7f62qZeds18YtsN
5GIZ890/tF7GD+ANKpPqZ2wqvKz/At/yOJfrLcdPUlwjs6agCtqCC/CsnV9UJc2ZIReBGsCUO7uo
GckeXls2IZZOx5vn2miQxMvD22wiNLfrFki4EChM4db/Zv+6Xj+ynpeJKK0KhnBFNYcOByez908I
2gpiTuHDU4h/aKQba+SJUAiP6hQonIjfaWU4e8SIHjkFCZvjjtKgu80jzA9oeFgS8k7GaETjnRzp
GbHQiUK9yNSVboSvi+T2ErL1dFyU/W6mj32AVSSCaKZhR1AfUKgDYsV1K7hFoAEV0MBJRKysvnXN
yqiPCp22HaoAlp03zJonP/SpZ06Zki7DpkELxKb/Fg6mKTRueUUoMpwnRe0SIARP6Af/xHbCfcXg
3/fyMgCX0pYhrFb4rbK2lWRR67RzU3r444TStkFB6kAax9VNyrRiSXT2DAKpAyxT90YYyoEubbjj
MK9W4mBDlOpQ6GBh2p0VVs4LLEPih1OcsNtmLeQgeAKddwf3Aaswx9ykdIXPacRpESlrZKOqEI6k
b16mFFLJ/O1mWbXWrSr/hQGULZzUP7Ys4HX7pqES4rloo2euHkL7ynycBhAR1I7K7Xgzz61cFdjY
3lQFpA3nfbV/pHisBi/pAU0XKiYFq3dVAXwihH62oSy4Jhb/cr/OsKmGIECSvKFLgc4AcKnMbLoW
nx5eheOu8fxG90KYELLi76ID3l8P16+QUeNK55QT7HzttS7wtDDOPElhFtJ2VRzHJ6sTurZLersL
GSyJjnvgMmGxaf+3jmxbB6eK9fe6bZNxjgY4lMZeuLV1fWaaW2fa0cYqQjGAde5EztEl8rfprMp8
2Cgnpmua0+AyTm+GpZy1I6GleWO1VdH+/4RrN+QUmfkR5WRafj9pk9GM8qO5B7i4GClEgYodFk3T
u8jy4cy3U08WpgPKcHsszXza7/HMhWFvWWnWHoRckZ5djsEsmOycotIEMd/D/b0w3vMOLbdwT5wC
O9Nwgc7S9jRLbD/YnceWTaWOKDtNjn1+JqESHS+Z0c+eo4CtcF2eLYN5MRHn8Hpwk2BUkiDJNP3F
YOetFaHWXBtBz5uYQjPPUS2Dvnx/0H+QMOgGS2JWZjmst2Z4Na1ZZhR37MjJws2cjWeyMxfNlZNP
CcG1LvH4iQfC3eSp2Z6WD8SpRkqDahMAlMSmhv6O3jhucAP/YeY+m9WE45pEf1qtIb1fiCcm0+Kr
zOGbH/VkRHVNznWeRuwNw/PoTV38QNRcOhJ3QrH82uQHeoR7zl1bHN3ad99Kf8X+/DRJ2wvNbABQ
+VW1eYZzQ4cMN+FyKhF/XjhtpUprghTzcuTHlcxsrZsHKBMz2bdJ0hIisuGAWFojFd6eydRo3b8q
a2E1mZiCCNW+AgE1LfXv0R1GGorPZbSmBSYPKyPu1TdRNgyfRof1EcEiIQTmiWFWa1TBMtS6TXoO
JBJMYRplbkZ8h6D4857ixBh08YckqqgrW9ZP4FGIq90W1Tes+BvTGGzUPnVArNSYq3CDKgLEBmAe
9JhxoywGqk//KDw5MYrbTSQwjYFi597iB4RNZyTRC0J1HDdFp7yS8ShEUeNDv4Fhl5eDHdUsRNjz
FCTMsxhLVI7YjHV83TesqOU67Niwo1zVV/tq+86ex3Dlx3WolNn+AD0kDMT3LC4/yOe25oE6Y71E
onpU2zgtfmNgdD1cW9D2Nfienl3R74nQTmFSE14r5JU1jv6laI6iQ0ooQV1q54IhBSVnH+bTSi98
O0ZROdjMVBgXFmaZpe9141pcFLiV3GPNhzq+I/uQHDTr4LUSHXxlYCswLWBOLsedUuiCWLaCZfpE
NmxsrZtVtIs8fbUrPCFaKa9ah7WmM2LyO5NtMb5IH8khPfl2gkmsJ6F5pYzsG94bxCSAv4n1w1aj
FyYfR8Rg8rbH2X6qcZTSQzpAB5JheYxDEcwEE/HFguPwWMs7gyvJf+bATJ2ondHx/xnn+Ajtc2XN
YIMHA5BXQhhtRm8pW0FPsP/pu8cv6MTZXEqSf3KET7115wamQDYq2LMR7c1SvpEnU7S027lbJjV5
YX9QgZ+/ECOopMvt7FP/7VcGH4YUn0YXbIptTq1+ERS26ooNxp6PFBNtHF1gOXazeUcod/DsXipr
/3OBSYoEfOifNBiXwcQvQMVtP59Fd/3Y/NGqHctnndKFQRxQLSjzojs69zljRhcG6ygirTiKUDqb
BQSF+s3AE1VfTWqZtnOAc2ckQDOJYcaxHSkzwwBShCYl7qXt/xUtbfuB3xeT+gK1xBQV6LBsIWd+
4Yq3civ7El/uPyA7A2hvNYzIQL7uqGDnDqzXFKdfWecRsLtU4YsjJNh2hEUKGWJj2hOVzfuF5ci5
HU3ZhY1XVEyjhWPtAe5kYL0hggfibcEVIdTu8+4kkPb2bLcqTug3e93Hz+Y/yP6P4SWL+gi0X31D
EHwyN/BdIJPtlM2yFFP0cVV7DC6/PogRM1YKLUDkKIHu6LLKyeY6h+zMvvSpya38S+AmxS7ftXUv
HX+8AsyiDfV7psoTPRc4tIC7LdEdpjl11wB2fRi1J6FPdayejRamPRRqjK1i3xKJyibimEEFCOTR
EbNBrt7SwgME51IvDejU6Okby6QqG1BLoCXiyObDf8dyYNMk7i80d7VGKOroORMQxwnUwQwf7a7H
td+27RM4lC+E//Cz+ENOAo03QzCO2W0/q6izBLUdCNkuigmZ3y42dllXTWPTAXf2n07Bq8xe+HXG
cpUtJss2ONGPHh2pmPTMoruW+6909uE1eJjFCdC9h7t1q4K/KwXQnutShWeY0LTk1GmFYNjjWdzo
trUd5JWWdgWUT2MXw98cpwhJAZ3PJfgBdVBYvUvYh/wDV+A83E9ynHU2yv7RLtvT4sZ4RUFgjxHz
oMplllVqSehu5VTTDebexNiweWXUuB1IVUaCT0x1r7OSVbgHrH3LI/TUBq35SodQ7FwGsF5lojCJ
UHvQO5V9h6UjpSp32R38QtwrrD4T+wYFXG2AsrK1v4kxtdZ6pk3Fx4QtqO8WmLA84r7yLrCfrhp9
b228NefgjJ54q7nKQkB/4iJfaPvMVAS/cn4TZKsHWTBX33EeauE59n79ZFyVkUKQS+bMuqejn8Tt
nC6ybcXcHVAe8kmKfVvX/RlEI6BPQVSvl9o8OUuuR/Fn1cnvUjBeGqXyLs14BLl1G7Qu58uX3Y9y
evv0VDnhlBIw2wphYstX0K7CcgoBc2fUTfO/y0Mw62mHWkoQToxgBosqDY9nU2+Vp/1vAirqsmPj
9qOpuX8ibUVxiODaiEwuywrCHJUNoDlSYKu67c4t1dbIELydxzdtWe35EdvU/Yi9CJyATn4+u6Lr
4FbUBLaQRll2dV4ZPqVvR0bcSX9DyecFp7+tbEMh7U2HcYejK+6I4wyGl9tLVgklEh2thNfZMhEX
lm1UyNa6Xp8TYNiJRt9OoT2RDkPtk5c794zidl/PBcseTLz4LWJzkS8gLUU35JqNWkU+Zxoxe/1l
O7FnKgoS5xLJ/bF6xpcFHBjxnBbM4Wz3moNsUnNyup8+/V7dKARGCKImt5oRLAhH0C/qheIZe30S
LezbWAM2NPWjW2G7xKpg1X+1zNtnuTTeMOR4P5YrmpRBBRvaGVClnm6Pn1iNL/pur25nYK/8AAKQ
Jcg+ARDVmDOI+YzSkXM6bMPKYKLK3wudLS0K7yhlxz/V3XxCRGn3ZLHVgd2QQJWMSCswFoX3f7Fk
A8sU4/smJlp5+KSj+0StYP4S+LPYC6QEIm2Dtt5YOjW/D7RJN4d7i3Cf6kGQq0YDUNXuCGW7NEiE
oEVMj023lYllDLBUMVW5Cp5OVUu7QazPP6hMdaPotKNk0X5GLrBNfeiFFSvMtAj2rSPWrapVTzsv
r8OqqtqLya6kry8fQVvqSGCR+l/V7w4UC8LlwazVxCfr/Ev5I2ty1vv1ZzJMUKvZWtAR22kxTrEt
Wru2QsaI22nBhzkzmeKY6WldlmOCBOiAJHbDbyA0uMvePwT+/nQm774MKIADVX6fFW49NxPCekS+
hrXVuEM9qygToZuMeDVcnBHlZGecmLUT41YGQLf/8gY+HBZVHEzYHFStHUWVa6oTeB6KtUXo16xd
KqKVw538eh2ZFR/eYJuaEvgZ/XHBWwlMKeZyAcvh5XjVibVgOiCEpDK6LHd2ra8YpMX8T3Rx0CLP
YGhf2Rw1IB8EdEmfQwhDCU/oaH1Vz6sEDLxHmHc/qb/tvSiIvcwucqWzAIciaytTZiwH3CsDbcvs
moXzNYe05ijc0jdoJx+mQyHuJI2xjnz7qi+Mkw/H4t9at18iZYSvy3h1JyQBhJhhbaZ+AdHvHwJ0
RppeXhQwwCQDS1Ue6Yol/PZTaPauptNgiHvddcwpwh7bADpoNNeP4JFc4wTE+qE8ltobeRYclL7e
d8rY7DXggYhDQfpoyEL9odtqC3YtMnuXqbN3EAiDgOWogiQi+PVBG9ZpYTu8GxNH5b9N0whTQWtO
X8swNmLLroETkitlMOnceFFz9udMRmYtwpti8vNsYJK3zn8rtwgt2w87MSG3ewvCC35voYUj9Mh5
nd8OUnRreEei76TgghhRqYlQoWjFlrr1hKB8amDsMh5AT0xprIRGOighXLDCKcnZuMfS/nwbAKhj
idCRWFJKopJ65QWK9sjWbS5qUhTQf8ZHAleiNZpCe/ORBZiIb07wl0XqkQ5G3tg41XgvEtUKN6dx
mjYezcPzzBMlJ8gFZm6NI85Nwt5c73ZN8mjm3B5ie7TiLOuASV6BFjf+ZOJ0BJ00+9cyltqsmErQ
FGXNNHESMElQY/+I1oIIkbmBxQKLMGLbdCZ6GTaetXONhed33ShJqdu4rGdTOJyZ+WbJYnPsB4g7
S/9qdSR8KWrFrA8fcYUxqsQhflBI87aC2WjWJcYGClpzS4X1KVZEzIaQcy793NEU359+lNGmtg55
4wG+LQq0kY6soYqvgU1LdGKryc2cpJ2pcHLaiYpzF9evlgDCXkHQujkT/m2i6c9w7+qhLqsOOSDH
aNQxOMEC6DlJyila2OOv29IiB1yUDW+8euMNY2NbNM7xC0ewLnQgT8JmU/LA/0kGYCw8lNsFjZnB
tMkngeqBFJKOL2oIYvXFPQDGIwjyq9gmOeNPwVV726xusoeNkG4LKizs01htinAnrRgwTqu1gu+V
nTMarM4koK79bJAHfRnqcZO+1ttPnohYWKW7S6z1zjQ9R9hcQ28kn/Dk5DDKZHB+0NzYhCzslunD
OgImg14pxukkgMYRvKqnbSWwRBKaJZbEMlRQL6Lf7wbyrfHfUPvipQuQMgl8YqB2V+gqklCcID4P
h2djFqE5oQs/qnm0WqEd7IdtR+gyUSxU345H6A2shs5yjbgq7kFaxsUs/Vs5KERRsPOJzZhQSrm7
cBbRnWu/pSm+7FFaq3/822/4RhnOzgQFNpQgbNzdUIrOs5qFYIORhIehkwpU7dS2W32SsBUcQciu
QHFvnpeyd7riYyYrkKYJ3AjoItht9qvtrV4egoohVH10rm7JQM/dlF1IelX/alCWtIATVnB8lB0p
6tuUjcbS1DF4XWwaH+Q4rXcH0FY9iU2Vvz9BaqzLETCxr2g5dYJ51gKkQRsPzCAwawoeTiePiXvV
gPAuBVgv4HrfEjDqBkXBmeeyDA1S2m1CeLrbAiabI/av5qwsb1b/VFZU6Co8oWWzZtRXMj01QUqV
t+Wv9KkVF2xS9lPEiFLTmPIldOLIGXaKejHeMqA3F3SG6ipefc4dzdeMudEwktgxqRfxsgCrAqTq
Mol/37RHsDOvMMv+VYV4fJAJCRsNeyHYsVIfm+QFPsS9/kC3ujsaDIc3UBc5JJba9WUnWW4sBtBw
RZf53/UyiiCeJ4JcoDKJGue38IqyOF9o+bwPFaLHLCxbakYdqxMCjBLoigu09DNXb+Ws4dIA+05Y
byoTRspLmzpFtZBDEvIR9LqkEoyxs4BE6vsjnb71EHsoVxwhvEY6wIWLaSUqvzI+xE04TuujsNW8
v3E2BZV79Beh63JbARZghbbqd2hYbUverkM73zeoZEtPrh8/iOkUtgF41MeUkbhxu7Dur0dT8Tb3
AFaeoELcx6eD9F7q5xEU1+fxNWiJ2qljp2F+p8CJ1KcTJ2a58xlagYmKcraDRvlM7q28GfzlY3+J
oo2rwaZ5YYd0JcDuNjK/2rh4BeAL7agS5NzqKFn8IWg5y8JUmTmmWMqoyE9Ozw9lJwDg4Q0wVnwd
4IlFEngX4DsAlXeQNi4D9ehzMxi0Sx5hOdqw4+VoQMg8jxUF6prGkbiqQJT2CUsyA8OjFxHhchZO
d4CmsNFP0l0IfroGerQBwwsEHh8r6R5Ie//7e/+x+gSUhroVvJc4fe2AjouO6Mh9YUJrI5krU91b
YNzS/SK43Q5Rp4cC9us5YEL4NVm37oOxcVwUZWyQyFM0X+YZbiuDYveP05TR36Hy+bS3NlEv65z7
GEzVkP8IeJnnrcoBXWouVpcnecHtXNNP0PC1PjeXXWY98UGUu99bz15LNioxc2FyE3NdJhayiI30
mib7rApXz+mMpCCw568UfY0KZYWA5e+6ZH+OTxv+IDw4XGhmk4TArbMKBg4vwrmcps0WsHSazG7/
t8C9i4vMlbAEqEGhLBNrtr7uu5mZzx90IBuP9/HeM16pBaSObzphJ3c3ppp0qUg7C/eJ2vzL6VVs
nhcoYFI3IvnjO1QiqVV5fN7/AKeLmxx8ap+s58gZYCPbZeRuo1mxNo30QCq6c82IC/BfYTmabHc1
hNBuVqd9NXGUljOcgPoDTOVWRi7fGpQLvNO2sN3qeQa2w9TW/MZw1lUgpWTw2EbgJdmQe4LJPmdM
CvgTvCm8jZiL+ucsAPvbB2+BMXA778Wa9SAAI34Fv+AqYG2UHqpCoCjeQ1axHnPjItB1FFYbIwVo
rrSLnRiRgXmNv/5DQzC10zR0ciYDZmzY5v//BJ3JG/lAfu0WrCeX+5Ka+zxC+E1A2szEwslKZwaT
u/9mbeyKGXRopk34mLpSdJBuXBnfwU+Q5yW5ysLr+URNFIcdBesDkXHhBnCROGZA8uyCUC8vEVn9
E4SgMx60X9CbguWiQ5/E0hLkjZS/Adc4/wsi9Dryafs5pFTgiwzD0x++y8E/LOYqJ3dQFsHPNtn0
7eU/fM0ARkQ+K/mIDKY1nGrj1Vct0EvecMKgXgXo6NMDmsuTKOLoL3mVmpqHJHc4OYOct4ioqgW/
U3zpk3zVooqj9tDdTNhWp32n0KjeSj2xQE3p8t/5alqiDsB8j99XM6V8tZKnq7jsrvlWgYH8RMs3
9lQvEvhVbr8yUTNaxW4fcN/fU5JjA17+f3/NL+090OImn+7D74t9pdh+xQFEw4UX3Obi8GosLFeu
j6ui6yB0GolOQSd5PgQ7cJjZotIo1D7V0lZS40ckH2C1W3/QBrGZgD3AIwzU1KIwd4hZhNlhigKc
i1qeduV0sqRfplo1p4kPE0iv8QAwNdPnGovvOJZNnzcHbIie0TydKOFztU61Kx9DNkVegy/sckq2
5PQmda/0Qr2/U2fhl+04mdYLOmz8dYXnAUjWF2nrlTD2U1a4IDraArimknmvjuV269GpsLrKUTKI
zLNU/tUhiwBPdK0eMCK5JHBriQbzegbRcs+akBFSlJ92hByJ9soxCnVik7IqHoAW72xA8fQSbgMg
bPtlCK5VzPlXi9O2upXaV6D5dXdgIp1OSKV46y/w8kqQL0Dpvh6bMHjDGHuKTgNDcPmp71l2LAJk
ChM1dGNnaQKXRyzMIri1tlhP+hs+70WhiJBkk6vMb4m5K7djaKF4sgoq/wNFMG52OVblPm1vt+os
mhtuwbvJ5MZPoJmnc+ztfss2CkEkVYrHFhWiJEtOQh8GhwtleE5I6NO4ubbCrrteENukm9FbedRS
HzG5klSDA8H0kMZVxXsLfEEtWY+QGVh5kgZ9olWTyDfZUCdodPY1WlaaWvR6U60qNPATYYGkwGct
NqLVMqRcyBJxqsFr/rkDXmV8Byl60fcAi+cZwIRdGsSXpgX0R9pwbM0aB1Vmds4rgSm70wxDzslN
W6fgL/tkVfx5hriOkuR/bkptMq1K5DC+bWeZx8GjP9ZT8gWWCcq67G0ik3KsQSjKQPQWoEJh1r/g
zkYFDBqN5tN7IIDLxJppeW7tCwrNWNyvlqCiHpML/er1tzLe3dFRbnZAWP7yZTQ+s7WXmbnBYdl8
tYSXd3N951ugt5yxBLGpHm+O5nbYakeVulZZpy2cmt98ILFhAyAv9hl2yNfgxWfezqU+VUYjoAyW
sVcD0YS7Nz2UKCCZ0OBDYaj5qMk/vEoGiPC2jb2tbGyW8oFJyW/rM96xW4QZ4PV/P3DZswMH9ALg
0rOsDSh4T+4pERG1+8X3O6hQoejvoWEuumEx7hzLiWFjacxnWApNFX+MhpwnfqjWB4+Ftj1JjTaa
lQNROy5Cs5qnuakkcMRyzkomxjTaBP1prfEeMQDZtN5pCUirYW8TIPrV7srTPvXWj3SJvzgCwuYt
RqXSRJo7NGt5Id/toGB8ysUIwQJ27eV5mi1e0YWNg3D0zrBL2krKlMAhtaccPQ0rqCwJZIGTg+/u
yYA5I1pLYZqB+l9QWAV1CRLwVObzarUBzPFwtPofM5LhcLm+S44s28I5O2pN7Np74c1KmRrRwg2H
dQnFUOgaIIxxnSUENOtaicD8Y4FQhq1J0OXoKJv1/JpOIGeK58pqWXAWhRmqgpW78O8kf6l//4ze
XGYf7OZzI0AJoW3sQZA/fjies9hFaeU6IoS1invrwUken8G05+toiZwWZC/9y3SWMHMQQfE8e5Wv
ggrAAIeTKqugqs4SyqeHKhT6L6C+yBtkIFVLLDHGbzSfzEt0SV29/zHmkG7SiKxabt4rpJuw0dEX
sUCVC44uA/rk5coh52JuOxr2k/OOyaGrju9MnYfA4p5PiofgKZ1rLyvUcJJ6ioKXqI/KQRFKh+Xk
LeT9M3nko+X4BMjseUl+MjbRifAyUxG9glfaY3B8C+Ka3oYPzONms72+xEAbdlXUlikyABHdbGQd
eeKJArOppJrl3zcqX/VaEyHGYrD3mmZRoFGR59hNuKOqbHD2XjpUBZZjJ7yV4o2mKSzykN+S8VVq
CIjzSghj4pWwTHhrVyrKfJFvZJTIxBL6KrNBsMvlrMVdAftg+nH1rjxzt4OrLgP/83i8wEJdLuAU
ykPu6L6kaW0cOoFYc4hvt/OwFVIKLj+9fcBGxYyTMFPC3JMK+SfRV+tI1kctanpURILSxHraPVmg
lg4Kr9ctGXu/5+/CRP9n7KWMo2VIVbQp/LvXOGGtLyzwYtFN09IoJ2cQqJoXiCuPz7rKd6un49H6
8RL6CxcVkbIFK49tJirVirImzqnRqb/i4hw5ywJtpYruYwqX0afq17lqsqAGSXXWT+NfTXCQ58Gy
PKgjbrvmndWmm6f9Eg1cTOtzNl7csrTePIdskVpqziqCwUv1vM9k68XXBkoL6w9QZZiCFcQzVg8+
enUHYppSlFEso9LPS+hkozGoTlHtJFJkQlfEYo9ijJ3paqJYMND02PSMA3Wln4T0zJh1hzuNVtiD
I2HAcWkRZMUr3OzPHLqC5D18Jgzby02M7yZC4rvQEbzOVXhcc3l5b4sLBaOG1Ulz7hphtDaE6yh7
ewx/aeexhxS/Nkm/eW/zOeokKbXrJfLgccu3HW64hsaPcgA7mlK/rFJFVJXI1CAQXq3lcQaJhnnd
HbZtLRb4SSBlH9Zfc5vpZP8oW4SrzNeBscOBRNJmk2pnuUbh6xhQa89KhHaCsw8mPa4iEDa7/RwO
BTCcld30IQXLiOUC0O+UJAPDArrX4NJ5+TMqPtS8x/oaie3eZcb6ckPWbIgeKfHAr4IjQ6mPLJXS
bnpr15TUH00YVtM2JGNzhSiOi4KIRWQs/P0NWbCFV7imDjbj95KWYkp8BBuVolOEiADQYYbisfQh
9UyOWCAAGa7xv2lzCTpzFlgQ7zbnd9rQs3TBcGCX+AbE5fldDN8pOUub26ECzJaorv5UG4fl6RZj
Mqz1YnrjR74hibG00pp+o6v/oebMUPK/oB5zNyhze9uzdMx60mbbCUMiM2sHJsGD8Ho8qpXolW61
MyplvCEfWhKN1HHvniPMLYGrzpS8Ir+Fcc7j3YgWXb1g/THLtmZMHmCFylgvzTCgNdA57XCL/YVO
QCS9+itkUhtcjgMVNObP1KI7gKj8jZ/Jx1gC4tPFjs3Jx3N30MrP4aBG7MUhXYbLa0HCsV+zGw3l
p9ICR0u0VKG1I3pqJMr8Lb59O4CgyIFrwM8413nqzV5I4SYhvomlNolrkiguCHwzW2RQlIXyxCjy
YKjMcEDGzRV2gs+Dq9OAHz22Sf5VIePTo/bw+AgAh+niyI/e3pBFuGoq8qQc2TaKidZpxh/KR0w2
jLvOO/Ll2LpIqia2gVFlO9IzQj9gshXl5WZyw6aIj0jy7dJHqOZBxhnHmqbXtO+R8ExHpmaOIuj3
FX7QT6IILgzEerbszXsmVb4BS0YbS3Hpw/ICoE5/ayrIrKrH4Ccbh95TgR3V6UROR2HJ6iEBODvG
iS7PMHGRBMmws5FM/mpErQ6djYYJVnEpuzskEG+ZJ5aMQn40vdffzb4b9IeIiGiuOQjIFyp3g45G
kYLc/O4H+taWZeSp71OELlWoAgy6xpJf3dEQIqVZluZ6b3GwJ0wNKQ+ROApSizi1urfIykjk5SfA
zh7wUCqQe9GTIfbLyxAFw4BIYT2FtM94gWLC7LgQMpi900vgkzcECgIvLgk2pzV138NVtG6nNc82
Ra4O7/3Kx8eMh8xzCzgiKLja0QD5SZj2v+IMaX7xR0E5kI9pU6TXnTwXnA5WgtdP+cGvW89TA5Ln
xA3PG33bFgZ1XcQTLwlmLyYbNfhxIwc9zLfR/RA1Uoj4pAWy/xIYg42XZQ5HbeNUuLHKDcxzRmab
zZPRc875rbUWAE1aPfvRhOPtFQ6iTRXrGoKBbV5NuShWdriTtwU3mk9H/uhsGLjUwoQMcve2Olw8
h6V9mSSQfBa9CddBGfaSQz7tAuAT1p6yb0l3xyY5zcvEB9Se/k/T0mU8iBVwIDLp5jtCnEIlYACd
085nYMjFUGWI/7uUbNQYmCRREW/q6YDPwsuc/4FvGdORNA3FEHRkIIh6da46bWMeux9W6kVLM5pF
M7ZPX2dy8Kj01YvBy3z8JzTjWOOeIcqWGUjglqArU+rhdsL7nX42cAzpimJed0YHE78YyY2LtkBP
5vgFIvQBpguCgCVsMp3vcBQLBqDzRqHc9fK6bRmKC6PC+Mw0Ul8dA7knuQqO90VdDFKH1mVsqQRq
0BFVfoaTWr74XygupiP3+75Iyy9xlnCEhb7867wdfD0wtAojMgMDtJz99zu1/QneT059VebYcQbU
3aPxJO/P+2lxi/ExK5DMc8bLhBxR/JY3gKrwFAAYQntH2vf/80f81dS4gzIM589WW2xAd7L3RSpX
g3Fw1tl+ms4ruOvBhB+cXKvJnhPqO3QHgZIjnT54nYhBdIjQqMGOP4AyAi8AXXnUchmX48IqUN4E
WSmoP98lUQ2Lt+TGnA9JXbrM9vuT1KfL4Ng7HrtG7EX4HKsRXKQE0lZTJU/x29hxXudndoK5gj7T
7Ey8w/gR74WPWGVvNZK4QzmrJATX2Ef/8L2/pXgA7pHsTFyzLe6O0YekfpMFmPtONLciwZuvPs+h
omN9CXzCFYNKBV7nWulMukjtD6NTamoeKS1/8TvJSBIrkW74o7iIkYyfDwfB/JAo0I4M3s5x4QL1
diXofSsPfsbsdx9IkYH+NAqLyL1EfH0JNnP51Ld2EgjVdgaqK4KV65vofGxFqtNqJodRKmKQtPwR
Q6MPl1fGnTzE7gvwEPzk5OuqnE2Woh04GC9lwpPacNPNo+36Cs8yxRRu15Bp4y2QxYO14Nz3Nfcw
PKzTd1sz0PBDGlp22dtb5zSxOsVr90OWAsPORWjCcCKgaMazb92QjiVSrGWsayZqaJdA1PCZWQZ5
woujT00QRVgfsvYHOiBdAeTyUe825bQh2iizkKjI+UF/g4LwWI5qfWSq671zobs8bbsDlHVMGm4P
MOEFJmtoiN7FjLf4izQZzcv9A1FCupL0OQl0DHZWBRASXth9WSMmMT1PNgHIvMaaItsqa3v/3n1m
WWHjt0HNyuPm+1WbV3Uuif73PVAZubNrfaa4D/Vwfz94KGoTTN+f2NRmOPw9koP5Px4N1B8vhm6h
lR7TiAYmBemhbaTmOeIL00tJnS8FN1/xwanpfhe3Q9qsM6FXd6NgjWspmd5xsjtzhsSWG0agOpxE
kUJsxveKXtXSZNO6H+/tQO32FJLObu0ZJIwfVubippie4Vx4msAcaLknzyLdaDgpg5rPYRSAUhMh
Dwl8KAyY+rKCzo0P1ZpbwpHDpvo9PUnJwGNokH+Ces865CX7krEhJ7L3XCFQQuwID0SkaALibpAi
wYB7IDlPYkq49luMYz589cQgOj4lKnOO+kjSy4Qj1CJXohwqGmYi3EBZ/DUvsF+JzJc+HiqX51YR
T/WU3W8seWBCrA2cVSf/mGvPAEToIB5BbhVSRIGZolGcY89A8KcdDF+c294BQJNXf/RmjtlP8MoP
/VIm08ISStR4iygqudcQPFOvleYlzlMSSm+2xUdYEnpMq4Ges1OKRZbWiKa3S8aifszE3a5VuDKe
ocg79eOhYsJSrX9KblAQjj2FuNwpg9Dpf1+bnib/QwQ9xrGEWCZhBJtrTjMMJy5F8mV3KaSl02lT
L/hp4Sg/Np8ZWixPo4ce2y0TQxUUst82jaUxuIksOj0XZQQYLkadYRZXWBmDhOaaUWzVy7HDQvIh
UBSSzNSAnbp5tkLY1gM6PRzxjK5fAYNjoE+2z/409y0P3aOFwxkhe042Z/q1fg4VMpKT8qjziDDF
hEq05HrUIV4iNk2uAftglTRmTDu8sJOuP9oHm3sQSJYU9Wl7uSCZkQxwG/tQNaFCwRAuhLRs1bVU
WxoilaaMYFV1vi6cXO+miOUpNFT62gmUnQ+1voxj+WCCk/aReXrl5wQjit2iAp1babUXD70dv6pN
fTKd0+mH4ZpngQ+kYOw7RYI+FJmMHjQ6zisuJdzifWl7VxL3EdiAdBGECQ7N4k6QT/OK7YcUCYMN
QuF2iuWJAOXQ0GsYFfQ2lBenoXFiRB8Mz/y8Sa9e/Gd393UPkcvZG2zCHVWwqq3r7rAsWdhyIeLF
MCI/HFpo6BkXM5TMtz0D/rpTNZCZoWBa5t0DZ43f0lSZzeROrsdLW0ZzT8hy66tuehc3bVfihNu+
itwLprzopdKh/4arAFd9oB/b/ulsjMI18jW3KLOZ6o3Ye2OB948XhfhvEs8yRYQNQr5b1povM2vr
dm7L4Qe8wzw8e8aZfh+9SSrx9RG3DlQoDcdSmySwCTs+UpnGvbuu47HJ6Q8kJ/3O++w8OmrY8wFj
9Vv/vmmw6tOHme44dRFf2CpuOS91XLozA11CcCvNEPOBb9Ep1l6iAxAiI4t/lWIcAKDnbY2XEgpQ
J29IdMARv+q5tzx/UltYeMYryGNf1CHsFVJN8dLWErNV16Gx6GrOfX8861XL4j0NpsKcMh/nZC+O
dZ9EiQ2dfItC9GQ2ghBlbxTdm33Plb2AA8qM+SnrHc4WeAXAQ8K6AgQg3H++HnIcnti75c7V2TwM
xq1RggdLBazcBKKyJD1/SPdx5KW6lB/iZwNdMN9aC0aaAV821t4VnL6pdP6TbYUm2i+GTjkniFcH
u3Fran0dDwp/1adRDI5VdXcJ6xpVOPsJAzL+oUG/CmXU2BO2L8DihLT1aiqGoWX44SgXBBaeWEca
hAsA6S2qcFksTF2OFL+6oIxLmFC9H2WfWni0N0ow2wX+72ru3gxV88Li4QOFmLjSxtnj5xr9+ZWB
wzAhJcRZbFUd/7TEBNmRg+bxD+sYJfKy7KKbW4dWvATEqJ4fPM3e1E+ujv1T05IQPkaQ5zJItKZa
KGnvWM7epP9nhhiqpJ3TI0ZpGN6tAUfzTSZnAW6vDGDb23mJZz48OMCsfseOmqsDNzOAA825NBTx
MQtfYSvtjstXB4cePHR5F1zbLLJTjPpa+8edsv6WPLO59EtD9qwEbTDbTd2W0d0zHG4wDLqyIfTR
6Z8AZqwFrtuxdUe1PmkqRgQ/S5rFSXHXeeKKCN6EeYve3CxLjFuqtc5Vf0Efnax8pOoqAwrZpsFT
qxCieGBujZBkowKObExU1+v/jrzN1lRnq2P/Fx+5pY9au8zdBO8duEH+mdzunspAWXXzBUiXLCcC
4Q0oo8jA7MCsuNGC+KH/TlnBBB1TSasSA+7VWq+x6Z9YMPvAOoeyEbqkxMFCfQi2oNG18lxfTcaA
OetRic/xbLKscMgj+pleiNvuh2IaQ8c60tzq7vFLQSRYLjC+adaTb4OJ3Kctj/TEnV0kLAETlZe+
fV0DVT+/A+rADMQGzyQ5DTQSPCZzoGLOW4wDOhOdfI+hIPB/bULRnUbFN1Jx0qvxINGuWVIo0+ff
C0+FTvaJucurhbXAiy1GSQ1xwePu86lVgPXULVvQLveEOFC4XQWoYQvmKOZPEB52TLSKVdRZ2VA2
BSd/c4wtTrpz5VxV8ApX9TYeUuvuZXliLBoW352EFxRq8pOAK0PBhqRrvrMouVppWDvWrxcC1l0e
onUBu44m5ioRCyIW4hGK6/ykEIa4Z2wRSr2Jf7KKOXkgmMpCsrDtsJBIZBYtNb7AWRYVjWIhv0zl
DX13F0y9Sj/OqZPemjQZzPmTT5hUuMD0wH8KViXnJE2ObPJEkobVYOYPhdckt14MtAIxC6Ed8NQQ
1oPB6L+KQ/GzDBjAGWXnhbY6wz17Rr5gDmyHyjoCg4uXhFIwoFa/wUOOMPFAjEnxLc1pFF0CTAOP
ijPkA8Iek7hoASWyM9Ay71aM4dZjsX4FN4cPS4DLTaYH5GH76plsK2IfyMtAX5F3byXO9QNTDXyK
OMVOyLNtnMWneqoXYQX2QqpJdd3dAqPKVBD7+P1DNsnHySNEryO8GA3G/5GA7c39rJx8TpZiaW0T
l4OOuJh0fQ6ysEJqKd9oitOwfjcbzui9b39TO2rflLpGqLJ8ve/o967LuE71ccuIP6EhzvGvevIP
jLjZNTpDxOXNh02+vPhBvB2OmUts+KJnTqWelpT9+qf6oy26DGiq9UtE2Chylogiu1SYxISFMJWK
tQOy/ju7/6OHjim7lM5FPZBeMLi8V23DRZvWesp/6DIq3TxLErSSpdB3GqFVDlhe6dia/+IohizW
Q9pRNqoxHs7pRTZONBdmtjnlk0B/oBsw6i/s9iiLZiI9zvm2IW3hKHkg73xfCrP0nEpFMdrhg/vc
q2ENSztZAAPC0rU9b680YdHhTUuxW8GsUexjLxiGfz0MdmPhBdb4ru0wrif4ATuagpxv6kxXhd7m
X/KqRN8Ax0MxgcuUBUStHee07n/rFr1UFplwTNxDndPhzY9P/cqY+moJHRSkkvjo5jKF1VJvZuVy
0FQsFtPekgzwqoM3s5R9ZeHbK2qJjOWPh02Snhj0I62iUXhmGZWlozofyhsxkTPzT8czG4RU8DDl
NKfB4tRbY7tXzfgzZldThUfL+WvNMz0hlAD1kPQYiwvS3+zdWVJVDAqjDCGXtbryRo9Eu7yHbL68
GUoHe1njxd+ogzN1GoDFwK9oAiGHVGXP8fTpPDd9Uzww++5rib69EqKGws+DegMQbMYgRpubWWhf
6soCRG/EtDliVcYExbJ+GT6SKSBMVaS1VDTVKljq9Gs5wgrUS9IuIhi/Ijrw2cvTTJp8Qof4GL68
07DDgtdA5nz1wGQSoASF3kkkV/pl04nUsROmrzeXagF/ZVSeSFeoQ4yZEPgyx8OXFo6oYp9ohguJ
2j2GHHXMDJOQ7NbLZJmdd5G+hdcuQaBR3BohkYDkbmzzY8Edel6s8t5CGzMGMnXBEE3qTdCaiBiB
MqEo/iNWoMkzE5biPjV/ShGJEI+SZ6BiF9TCpnvQHaYkmdGGUFjMo/pIFaQYwN+mUMOg2BJgfXuN
Klh1/d817v28mZHzPrw3EyAaSoJTyWB8G5mXA2vtuwbZty4PZSjRMuNQxit9o85SNcrSicR/YcTH
C3sa9ziZJeMPFHpmEenqjJZGvSK6ETtl5zEZFSjrxx6BdVbB/E7kYLqbyOFcIcrPhsqyOh5A4M3P
Nt4P6CrZ5dGuE6hZed3IWQASxqrnhRoQl2Cv2AG0jdxl+ory56GXLHna5pviyxL5rAezf7GTuYad
zKh8ojdRrDXYcTy0JVMAUvGXUn0dWnyDiALHivWjux/kKLr3AovzwG+h+pKpWubn1h+TytuhtNAm
bhX0Ti5OghCzSI0vIM8ZNY9GE19tcdu9nvyFdN4Jm6+K0Aa0MCOC/jTdoBo7D3UL7SobralG7LCW
4IAyewirgasMRh3CcwgrGeFBdiHSV3MjG4MdT+4e8zLJ65F3GeguGY2FppugXjhlh6vjLwwzNtrQ
FEAXGuHAzBX6tyZS6QzJeQFVYZELDq29zrMn5gmvpf/Jypg+hXQeJAR1nY8NMXnOcfwGZPz7XfM3
jfWeixGLXPNjmY/a3P/P00lL+mlWoS03ANQaAcA+ksN1dhQfEr35Gg6txxBGB13Cpn42rIFia0BF
0CqeaI2hP61mWw4KI5Q6g+ydd4Cg8/l58N5NbokpbuB6X+y6ma1+2QGYglBYN2zz521H/YaCvMoT
IsurYTa6M5mMXAarzwtSxud3vCEeCUosIPYfvMnHCke9aWZiKUI3WizDmWD7biiwdiAR1N9RJFRQ
+3HU1nPt+KvrKTGi8EPrpLr96UkCAjsoiJTi15gI5TUyFUnT8alU82UECqw+PpbHSNhcEsTiXJlR
bUrqqN0SQ52ScKP8hK6ljAFaiS58pkjKG099JgYhfPrv61GkYv9lrOKRAcyJkeQCW40csWWN97Tf
oyqU4fgUjQTbgBZ7d9opV2u7jxb3f29xr9suQkEHtMZUNCHMxLbhsqZX7Rp/EECG7HamXHqledzT
O4Ehq/FgrH+uQFdeCEu6N1aoyai/S6UrAltPkXEcX3gk+FilUSbcY4IJrhzFokPmDJU6HMAYu1J6
mmnWLMj3Eq0gs4w1Xd5vVNUD3Qkg1hQkS0HjmZ3RWg4Xu7JUcvbZ9O/lj5HMWAoKaBtp5sSSbiHT
dMlKUUPvzFJJ/EEIEQVbjlG3BIG6Ld+BhzqZiLQuC0XxPzPNTWbJ57K4hjjrESN+L80seURXk2Ix
6IcjZTKehc8htoEq8hwcooVadRdHCOauhGT5Gxz/hSucfgoYVoD5ftlichXQHAJv8PPd8evD+Ks7
ilXbRHe6/POTkk2XjzKrHJjJ8zk4lPFYOm5x4byZpCidTTHGDNQhRYYaaKE5et9lOkgykERpYUmS
wQt5UfMualAzXYMNA7+1swZ8vQSVq1ObHpCC2BDMZjU5/yyYB2wsYcsPl8Hop1llV/i6l7DbAagJ
MDZoBr5iEtZsFilm/rOMGbpQ5GgbJG6kMyw2fSoWx0DFQVW+FPWMTDpm0wbAOObz/+V0vSa6hLXc
8mCSYxUBZs7TNwrKyC8FSOzhA09+FSiQ1g8hK3JKpIfnPM9RG1ypb2qeU9n8wcUaCKoPfvm8PJzk
bm7E4V0wpvK4qzomGgrPL0NY7qIsHx99/tQjc8ewHOAtzG1XQvKB0A+7pZUh9C0AgaNVTYCQJajF
3bpUmO68z+ndfSyvrF78IyO66Drr1hhCUfP2aaTGL1AwwWWivrs/pA5aGt23Mn4KPyqVOgSZib+F
wtASXr6j9qZu1APi4lDm9ujFvM1SHqdX8LjnVkGFVCVwRYOTFHV3kuGa4U5zeuks50KqLbd/CTN/
6kYhaL0V4JsidgnbXfXkwD/KnpagjpM3MjSzP5eNbg8xaC1Y76FaycwG0IWsRtxNivSkYDstBBE/
xxE8tEIwwL7XQ/KqmF5DID5HaF5/5qaXN9+aGZKWs6YN6gcr4P/p2+fJxxatqQMqn1+ZyzGAGdYt
Aukj6xBe21wx9X6ARTBQTI/ymHgT2Xfqv5LmzDITQYcWPPxSLRt5UkEot0lH4ago7QpdVJXLYm2f
OW8JxFWxGk07oQe7RzkL9oX8tRGIMA324GVd+irbRgtJnbyYEDT1H3uXEyby1/OL25mqtWHmPQ+5
VLcmXoNclhpu33ZNYKsqPGVev2m0GclJWzkG5eD8nB6qb9JLAECUUXuUjaVYiEXjDeIgDsx9kZHr
DP3EeE0FQJuJbExNSm0b9fUlnMs/sDiI+VAt1E0vuvxvAwCwyuoIOCkykrLYuqzIo6BdtlWMsp11
WTdip1SJjdsIIUxHQ7/gpfw93/w5PcllTX9UG9f1g7lPkXYwB4+KViq09rsRucIAP4dnLmb0LPeE
k2KuaCCNOghN9VDNUeFwJngTdn1eWEUIsxkmurZFGLT5L09O+qJOB0uZ+t0kxYD/xvqk2C3/4Wlq
s98z6FCFHrBNiokfD5OiHerlzC5jUi6Fj0Y1mto2i51QAs2ttU2lZUExWOZdpXgu5s2IHtb0oO8c
xYHiWTdVaPJtd8zhWLMWn+k9ExtPfAm6VV6C+9o+AQuRUaxgfENSj1o1qFJNv7v1qZN8NoO4FO6G
e3CxoQZzVF8ForwjrEmnn7dZc70YQDjYKySrR1c48H0Jfc3O7BrKIo/2bKh1nb4orRqSw4ErR9ka
elYrmvLrmQM6xajy1W7q//JJatuJiJLcQvD2zn3HsAaxQ6TrK5lZbfRul/BsbEX1fn4fxrtg98Tf
bVps/H73mnQKtKhU85SppvVNyI6PVou0NGOUZQCxON2N3SUZLv1d2owKScDfpNCSn84WZ1GbQUzA
vNXd04+jn6126riZjKM7juuASsxtWhDpW5r/hzSa3TYrCnmzncTUVtDIkdrEjAHSPTrUWOCd8YJd
j25Un4upGxsDaf2uKE3SEaPAybRvGMnDAz//qT9rybGziFyDWQgEuVF6tp0oS81cWxd36OmwsKAc
A8tbRARalSWJJ+y1OUowrn5r5CgzMp69Y1Hjp7BqoQynNyImrapG+Y8IMJP0K6tSemLaEQ6MlZkK
loKWBA32gmS9VasP72eTZCxOuCkdp6N/ArxfauErAo2Fs68rY25XDg6ALMOAbEaYLium6XvIaUyy
aFVXvPK//96QV3SoO7Jh/HyyFZuB6TV2FPbeJDhmPxN33hBMFufjeUw1WyEwpBY84aTQIaM+vZwl
jLQNnqUhz/Zrn9a5ubMnpHBOH9NXV85L7lCCWegewJx4kwmNn9+Qt2WeI3K/RDP/IRT2fDtSFSsp
c04zPUblkVYEtZhSVqgpfNNw12XAskhuU/9Z8Db8cqEkuug+etx8vlEkR9xcJTGA/s6TF7zZyxs4
Clahf0lHfzorN9KcoEkmILKYBWF/KAVFMuXQ22RN3t2Rl10DdiYZZZwIfEfCd6GmnzgZTWLapFVY
StQTwwgMLsicYlDtDtSfXAztflNObFuUANQRYFggdhPdHDs+n+PMhqW7GNjZqBnRbZynq8uFXBNw
G9qU5dmQrto1n8UEUyZxxQBnvH6eWcxtz/kO+rGTwJzBpEKtUqjurOqYzq30azMPpy4fZheFckBY
mtTzB3xx2PcCP0CRNVH+jnHiTQb/wjhrLCiypqmxC7BUmByTJ5jYPJK5ez8Gz6Lrwd9Uvm0sc+k4
oaVs08ob86j6mQ0tXvIwDOGOMMaveJstXOuozIYpuKUgnpvXJ39Xf7NFSGTII5duFO6wzB/ryTtH
aIuJsoi1HSwaOC16DAAUIrIXmrWN7kvMpfkzkT5/Xp6UcEIMrJqk08Mp6x84lVsHOyR1UGm/YqqA
sCJfDY47b1xYp6VZ3PwXRYAEI9y8TftaKdHxrC9Kg8lVNCYZsUQWDzzPVP8NNhf8/suW6Qc/mWNB
BokK/qj4FWFn1ggf6eirO18Y9yvayP/+588lqSqqFGi70zXZ0jvynvf0qBTpJftNfAgZvQFAtJmP
9KzozGo0tWPTbhjkEIVLCt3Apyhc1kMN5mhDqeHtHfMvC0EzdOk6nhrp3PESG79H1y6lC52plN23
PZrhCKS5gdOGzExhzYbsEWHGsLnx4VBGLEFqmTXx0dK/yiKtTxJ2Voa9bayEb9/mhH3ICq33lg+/
LNVSheOp/wEQ0UddHxoXyXgL7izQRKrzDnCDmy2f8emi5Efqn/CJ+z//kB/8/yV12Fy5jB9c8pWs
nh+F+haBjrlH9hxklmrD2q8ZGujRiCg6c0dJ+wCX40MGl5nSu6R+xi8QW6K+P5Rs3uG7nNkfHaFd
BLh9lSNjnZeaEk/6YkvOvvIKIdHSfarve9qtxtDRiqZnVgcBrIVMmNdKxngU1kvsTOYcwj3u4yeX
xbJ7ovYkheEiyE2x7ogZvAkp9WcdVEUH5fnit8KJZkFgx00JOQYAhuWd87dQEKwpEEU4fKkdTxIx
adxDmhP2z9BdsX617oBXqNjHlFazxuxTBNDCHFYWPsjSeSUwubvZ4go7FXxUrpDGBd5V2FRyRsAr
e8eZHCtieL4a3bBib0e7CV/dp8UBM0lRUwZggtMlziYS8MRDcN3xEaZ/j7Vdyk76Kuc4osbdS6kr
9XD8ym8VZ0ommo7/+usKr9FTeMQt4V5p640cQF28n+toZ/ONqhF6uDMotgJJM76YjAAaGcRHjAAS
V09ET7pFBLlRZNWtTETUWnp96Nsg3VRG2LoJArZ1WWvnKZ7Yj+GHbpkCdNzw2fun/gCEJZ7vwuEw
Pk2IIw9G1yccu7UFVad6WaFPwZP9vPt777eXpQwvFz+sQsgQdFjzeFffXDcFbjV1XAmUSxeMumQf
waurQSim/HvCEovoJYud3lzJLamle43FNFu10bGroKONA1FPp5h0iIi2zGV5qR9d4VYQa/2mrNq3
JxxyU3nG/LFOF/SLL0CzJxb4SeOR0M1MXN25cG7qHQ6ACn5SYw485AIgimZRy/hc6putS147kOWB
rgNwgWXmaXcROCAY4LGamAowgxpDvU8euiNI4MMtoHldwuPn1g2wJRfoWJs+AgkOf+8kYJitwgsc
s22MWuhgRYAlnp8GYQrsjittBtwhdzJXw+a2BS9xJkNpjBSLDQyGGTdT9ylSQ32dyoBlGnbMhM8m
2ye/a05EDT2FSANlfZdmhKWC2KGcGqgpziFHwL40zPhorkdYF4Bhbhvhu2ALtMR8DHJ3AdCC2aUx
v9Fi+/DyQHssoxhsB2pqfcXoifm9fl9CIbdM1Kny72dAgMvUlcdFDM6JirASWRWFEajqyh3uzrXR
Bc0OGFgR3RTR3w1rC/HLA/7JMema51P6x9BJTeZ+30vvrceiYS6VThYaGcOhglFwh2R5f0Zor1o/
iNXuGKF5Js9f9o1FaHu5799IR43ZvHtiTNXig77qnwtUPNUfP2EZFrhwqK84Skbl36ZR5sanEFJT
dBeb04jV1ULzGbCDoRUCgC4nBdnS5Hl685bX/SnKohVtmPz944n2Y2ydCIv2a7RekHNIEz/VVeMD
IE9aqQwQWAhUng7hWiu7r1QS5/7f1umvGi5Nx5gtNORNTYA0al/GZwlagTpD8Zb1KtjuHOQRoI7m
6+58blgf7H/ybqCJnHl/vV7qeJEDGZuDYzvP4rKYg2W8pn+lNUwZsnYEyO8lilSXB8FaT4ManVUg
QqofGBeilus/3MG27K5iyWDs2RR8nsgh/gOiBh0P4Q8BpmEdEW8kRMFStSdqeKUkKbWxddjmIBLB
CAoYQm0YkqVkNRLlCN3kkX785NS1V5H/QKLpT67/zcEnFr3XFpMND0482LtWOC4nCMLz2HXiyLnp
VAI8oKgSE8bJfDBjmdcBzsa12PxfMk1Km+NqrKiPRp0laRrBbblOvplR1ZZzAClz5fUIPS6OZAU6
WNuQmxqI2iKMTmDxik/9qeg4SH3nvMDl+Uf9hBSSQmnQGTJ9FYq4kx9WnUxuTq+8DljL+uLpLvG1
GN+Bu5s2nSadSwxRVF0uczlLWGUjVkpTeNGX7y0Kl4kMeqfWkSXmBcxlOVhzMkmXx6MuqAMgTIdv
lh+i+R26GC7TzJXxV5zGvIhy7qCILcU7f+VodWCRiQBwd/XKMVP8W2bxaybLlzBVctbikPIazVX8
fAzp0nXRTgt3S5uodurvIxEjgPz1tqaLO4BKav3a74X/BMn63btW4XuTIc0p/6QVAer83/v0YIor
dm0QkwzfF0hZdYEthXJ/uwk2fZ++4bIHF5S4ZR5YFaoqhu/L2pilI8jxg5lzi4FhqCK3CGCEKwgD
vNGYyIkrzzkRPA/LmEjaGA0XiPOLLIyktqM/XtcLEEbgL4hPv7H7bINQggMokAU/Pcy57wlUhS6B
NAVgPikymtl7tikE6SxdFFNxE/TYpyut7/Y9cHlsjXH/TA6x6ikiq+m+tvcusPfRtl/4nYk7E/LG
Jyt7AIoT4daJINk/dFTV/cPYQgcOsSf+aoRsrXQGGW+eff4NX6dyQDj9GfFNC7+SRxhybcMMWtbN
43/B/VUgDf3mAO/JpRpsMzPFb5fpEHrT3J62BvEMATPRteuZM0ZZ9g63QAqm7/mSKZkX5YCq2FZ6
9jmq5G0FQtGhqc6mSKVCKNBsFglR6FoS9oSjq+o227qdIhOoogv5mgyEGi5MB6G/eL69ZE0SfLzh
LQY8A+NlH45vOQWGUfsRihaIFepq0Pl0aRbxPMAX4YOdm8LkBN/4qx00KztNg4Sg7yoyhpRaL7W5
BwHaOCK78YDzsHaYaxVB69MV2QbjVWoZcFJcv6p+/QpEgaiNUdPuvpI490ElUbGuzrrurLlhUXxm
slgRm3dr+fCm+U4EDSQSyYcZZQn62Vdq7bsku/ddnlcWASnwbCoFcxNifutCGn1gYFXF0fM0zK7K
aAoQt2ojb4IjWg8rW0XytYMlT4hF0Vd4db4VatMOWykjLcbkOeEnvwJPCXgPhx7J5cd9hEL4oNDZ
iidX8EAqPp/rZ0jQ0tkCNYcK9tkF09YdQPbeXlHrvMAa/hDoI/GKbO6kjjT+7Iuhd/XuQTU6KXK8
bkc11ZC9rqYBSyP5/9D1uuiyafSGRU82O4NH9SubfKkyWaIPDUIrOYDTbcQioGgEIi3GgMXsKyD+
oXhlhwiU1Y11C6x80WGBCwr3aBcYe7rTMqsMz4SabnF6Ywb6P53rc2Miax5lyg+Dhxzt3NXi90BK
HppjyM+gqmvQHI9otmnTUw2/6qTUTOlkHClcQ/geoPRKq3UZvTRqpxQpux3GBcYPdV5ZgYCZ4qp9
tcK9j/thdpyrIwkUHlk8pkTJf6dXdKto/jnl8FLbN9QSSoVJ6X1984j/oxLz1KFUx19LtzQLTD5F
ve5QKrE3I4bJrf3O3vV+uOFwA6LYk1yiRdfiP3EeE06sQiLnLAxGufTNrmKWpX6IFYIj/nvOB2e+
upYlrx+CHGvMYy7JwQIJpEAhYMlaLlt3W7CjhXN6t+XKTTkE2OZJmgaHrBt7Ww0h2KOmmlUFQSB6
JJxO7nQ9I2ADFVwEclkS+oelDWuWjwquWSsHTpkX7ep7bvOL0L1fRpW1FiY/yomQK8Vvp8Qjvk1w
x9sviCvyeJtTBTiJHyKxqIQ4nLgtqH7SOBe8oRKfXHPIM4uBoKgdpb1O3CUxHyQ1S2xSwfeWNIyL
xehXtD1NvMnc4mskl/FcCwhYnU6HbZRbMph6BRE4m2oAvNVOMuiQ2jBhlw3gzNDOiLqk1fIfeyBa
LTaTG3FpfGmzGaUS+i4omt5KCEj94xVgJAmVnJW1Pz/9xJZXf7pD9unLO3TseOhN3lZbB5KURG+q
dEWO4+kJEuNnbMHYDRDLr4+iaYxKx5S/98dL8G9tmrlxdwNACzGtdpcO0/StycaZoAHoQ9jhxi7o
JL80DRPDewgS6oAy0emokB8VFt5NAHp0j9Qf3ihnuoHePQn/pOjpnOTHFrOpHnefylLK26cuNPcm
xFtUNN/tg7oILW2EJ4WQaApySKPaQEPclc/QOAYh6ZZ0kKnTrQDWjY+9wgX/2ZTMLU01TFB5rAxn
+PbGCb31WoMRNpIAuDtQkSdaydKGTERtDqDnZk7Ucigoq9WCoavKBPXGx8O37E4bnjsp8OoiWC41
7PkO9fQ9MbiGOlyyjEjH3f58IGKu0IMTijoR7SgIBY+k0cI+oJoc4etjFEWQdfTu3WXeE/PdNhXj
G/9PyFFsRPX/tQoSfrNHmVwOcqXgrOQIUFaY/qEILPP/uZVwZy6fGdNjp7WcEwIbC1BgfEdmOXZl
XldZupCONeqjfidIZLfx7AJpe5HEYQ+c4QEIZtUgACv15Ukqijphk2nXIKwcxO9Z2QfahzcN9Fsv
G4Xjx1LJ+iIY47X3zmaWMa8L2O6c56If0W7UnSheBJAGzvyu323sHrV92GYD5yO8ul8360CtxWVe
5/RxZ909qLt/ZfB0X9OwuTnFxIaiQQAUiXA01ZD72KzM8V3/xplIloFFlRuTPZFhyZHUrVnO3oFg
LtHfg/FFLXpF1pCiZfhgWcCpmpd/aRsgjhewARiQo+VANim4aZRdcmycCGL9qqgtn0BArbKZupOA
7OHAUU5InS+iVtgVF72isBA9jbX+YWmdV7g2D0IZrNgUXAxE1+L4IQnRrHKPY3ePUpQlr5wbVS+i
kWBKQD3bwLSYRk/+G808z1iEMAoBWTbp28vUSf7JRCA9Qa9b3Au8RYQAwl9z/MKtAp636cV3z83/
Pha1tuJsJ5Us1a9BeNNYr3f/I8AlVLr9RMGThhcdC3yZ9Pw94nkOBanxUgfK3UQprDd6bLugr6+G
ClIdZQYjHz36clyplmjUZj6NDLD1CaAZEVupiQK0ZC4P5YXT980pRym0/nJRhKQzlvUDvsZyh6z8
asccmA+cZB4OpKeVGpKAXJjBCuM4naLdWzFQ2K901QSje5N3dqclYg4rnY8j2M1iHeFBj02HPcvI
2jW/sj2DjNxUQzH154I1OG3KvSd0pMiyWtdy9aYP9KqScrbhFzgdu5nC6Z4KtdQkmzeKt2V2laXq
4TzgJhQtp8pohlhLLmdRt2yHzFQeaCWnTCCrkaHLf/KAryZCvbfZ4UPXHPj92ABIkcSofdf5evgM
920QwDXa3zVNuF6wEiksJd9D3f8xJlb5ZNaK2gMR+7BgwfOn3dzqy7gz9uW2hlVWovVtANDZxqrz
YjoryW/+nZUSSZg34pgBAiSmfiw00DRIIoOM4BBb7KPVqwFtd3nBXe6F+TBU08y5WDtWGi9gjbZl
YQBTu2mH0DDETcms7hnbReMJ6gt3WI5eKZCT6i0k6q1n1eBc5jHGyadIcykiRJDsjeE/00FExKDn
+UDd8NghS2k1ChOrGhVHfcNlj54O/oRIMYR3f/UrWXgtN2LdigSxLq9SHvQkT+/7IMmbAFIBmI55
N+CcyPz2BTgADSTFD5fVKR2kztoeGJ9quntNH1sboVQ6k65cTvGGHzJLPjwDYpoJCVsOSGUGVrDg
7w9NSGB4JPryIKFhKLjTGtCI6sebgOHQ5rVH08pBmFQQeaU3ORLAbmM+AiaslLRXIOamZwovA418
WvCeZdLDk6mIRiWh/SBbT7AGFWvqF7ovlDSm/r/WOpNTA3CG/VrSeFMyknguKvEJBE/bHYO3QOLP
BM31ry993XhQJzjY7tbmhcUfvlTNRxF8NbMnIIp8FGaUX8pYFtCkXIA8WOPtb6bqndy/S1Fse7Dt
ioVzo9sWPstR/BRC5HnAAqRKcKLUw9fi504RP7KsIUxI/V5wXtKi9ZZOxoF7JfvGb6ih7ffQXLlI
SrcrKz1DZJ/rSR0torsYz7G4hxryaCwo7OICfnib365IXfTSNW4N41mAJxWbzanHTBCINN5DKm8l
NAYx275P1L2OdKAtSqJl/cdje3HcbaHFOKkT+hkD3iW7L66cE7dRwahPtK6Wa9TH2ACdW9SN54uO
oaeHPheuAceBatvA1EDLKvjWLXpUt4CQUviQzv3GSvBrfIJa+vIQc0rSq8F2U08mVBPVs7uCKhQm
Ge0kEwbapzDD5PbYgIKhJiQTT8u4Wls1/xWNKx1OyaKnQP+QA4j+6R9MFF+KzCsYCl2ZDqh5/4Gt
mpRgeHha53cRweOrMPUaUKDFJSoTZ+6lJSHzOXsJxr6IfTxmQ+POIAxLfyLuI+YBRqvnMMKFQ0ZF
cWT0ed6E9IkFxx9Ifv1cXAt9lTu6o8GegP13A1aLBYQRnwDX6Cj4IwA56xDQYIMszTMNap/iaV/5
n6PTtsfmlZm13DtcwWBnRZWYnZ8WGEtNPFtU2FuUCvM8+l3QQEx/W6bBAEWckuH23qPk1biUQvzU
8a4UgYMGXTNefxiyEJeUlP//FYr+nwHkHSZiWaeGh7Gukx6Eg/fwQH8I0zx1bxHgxbF1fxVgPUtA
4WcW9czbZgle/6+uWN7QPQ0dlvlX6QPiYo6WrmUW6JfEMGJ8qMn1npDtJSCydemmLT5GasqR/AZ0
0P6YtMlQnL05EnRWPzkKIItRjjYp7NBTsa2nTGgPVDLy9PxkBjMH8dxRrdjDDq8ZVqBCPyvt9pxi
5/PW05XdM3lyg2mkLULg5138ALR1dj/HU1RS4h7chYFTroHrguQRYypHzm/+JB/GBRcqBBD2IMNu
25P3x0JOW4ujv1g6IqyhDuMcesHn5Bfp0UgYAdrvJljhbO6bQ/6srb4J3HYgIdbJx7ZKumbWAyMx
1bCN8j7qDo5CYauTxQEhPr3U32It3MMzYjiFurLsvB7xpRgia80caOtOtxj6iKF4wETfNjzDg1Ux
dPxn98RhmNQJzjsapyCa+35Ghsoyv8WC182+j/x1l/M9j+WCooHXBmDLX0iJy42PwmMtC2n8Saan
7eqgWlOe9f3OKmojGjGEqSBpTqZ7RcJPPkcOB8INImISfl/DRzeA2Y+G4/dt3OjEguy19dVrkPbd
OoLZvcyEMOsyC2OWotOqxhXwrKCuW5MTvA0f5eAJFShkFWiMpALGjFBTUSvXu/cL+IsfDINqfxIb
GR4MAWavYCAK+oSOpKyNCSMrSnOMGTUbK9OYaxXgoTICMob01102I8GSfFj0PpSRNQG93ECG6Kew
gd/8CBCGagtCkZqiUGsFyca+g+VJKFzaetWdWOy1Eh8JmXxzseQ+EWcdrV0lKrSx0MepCB55ygFY
oCfKLT1Cm4ITe7q7iZ1RYUsZV6ogGgsIaPX6KnMnHSu2oYT5W0fXnHGtPOhlOqXagZY8Y8WIPuXU
kfuSOoEwSL3ZMNuDsYPlf7O8iEp0VNj3hZ9goig/VhHrSYlS28qAP9AWjIb/o88V+HOLIWDEZ5Fi
rrNoJtfn/vWFrTXB2ohJFwcpBX1OUij+PILE01id3aHMuDqpydRiwn5zSVA9DK+5gYt3JVw7cMLy
a+7ppFaNfFWgUX+IhOol8CQ9lUgkxhCCC/Iwm4vwuXucFQybK48AybpmQQkIYi5iia3WI9IQ9K+v
GPezyXe9wyRSoFdVPZpdqAPJvn4vf/EU20guLnvjWLO9yA77U/AYJiiZKGM1TQyVGm1yePJTl41f
mrNJpLscLObR8TH6eLbK/lvkKf9LZ6+Uph7AH7d9c3KlYgtD2DPmiMznnueKyVRaUdFmaUpuavAN
upqTZn1sALqj8sw/AHS4PFpViHPpWWvtsW3UZGhGaf7ihJL/2sk6lDp2meGtwN8L8rxPim+2Tfw3
L15QM9AYrfvHJuAgfpf7Oj/GXDntP6GfhPRsY+UdlJcg5edZP5iuS8Qu6xkQP0cRoRk+WDQtcwf7
a8/vJlFfCf8f1i9yG0T2RJxUYT58/V9/triY/HophpYNDdFvHHBPzuiTFNjBgyMIA7iNt3f8Zahq
zSVfNiwZPZwknOIosnFRs2OGjNlnP8Jd1DLd2bxNplcbMwnGvbiFfRSl3RfRcaP0dddH/2sG1QVi
wwyG7ZOvRJRTlcuh+JrToz/pwSYY9q/L6UBlXudJzXqvIMAwPZ0TF5z/CfwJxoG2sCybNRPBA93W
0B1E9aP5Z3GYuLW5MSxkuhFb9RuWVtPvyr8QQKbhH5sTjCoDOnJT4rC9dXW1gY1n+6PHPdXxKeDe
z5UN1qLFWBnNKm3UDuGO0ripk3723xg++D/kD2L8p4jt9yCm8e7kR6j2PxagtM5olZQRCfJR6ky5
sahCqwzf6Ho2hGcUn9z15P2u8eZjTj/ENuy9wS1lVkBmuVcuWg3gAUbE9A4q0GLKZ+nbmcK5kXvz
LHFCUSrvWnlviGLOWe76vQXVlORWlrUZV49Wggae1soHLFW869OaQy78AWefbTaWuQV4yAiZXsVj
yvF1oThBKAWGKqiA6H4az4UxgSakA/GuHHnMiT5Ld4FYozijUs45N/O+rAxblm0DxuPDoe4nCdqS
N2cA1Nsj5qJYM2ybtiNoRvIkJSD8gxeeykqciGPyFa81HvM46BNdYuvK7TPfKao89rlJ3/+ww4wk
NV6cugPBE132ily1kDQjTQMMaTBR3h28A62Hg0KPfRwK9FoOCgaX8sE3UirxeEdUS3NiE4zIijF7
XeExGp66ByUpzxwBlxs75b1osSdOaHJE6CqZxlzuZUJOsnJ5Z/2p2ZEuk8FhI7CWBipL7eblAB8b
8eeCLVFS2yZ7t4XMrQ13aPfCz9wXUTKFeUBfs92FlN3IY92NzImiCYGTzfvAj6Iwgui5KoGgiWfx
aAdeDh3bH2QM0fQWr8UDlGwRX5h70Uu1V92YOmG/btgrp878D/lywYmieHEtB6vuSU6JwNMUdbcd
DctZQSBH3+d65WKvd1mPQxYX0bIUee9O4bY4J4aUTVG2gO1QTXb7aXyesblMGDSrSyNIKem1qEFH
OjNnF1lPluRtqqUJMYcup58w16tnEEzO7AwKoDDysyKeWfOJjuEr3Pon3zwHQeicDNCQrBS4EGxb
NwxmoBevRYqZDIp3GY5nzUxZX4qd66Hvs+yFf1H5Og2dK7RhKKG0mrI6o8uFhUa2HA9Kpqah74SZ
axec1rsWdoXYCE4TNrpeX7xGR9fUHFrj87/PXdCeVqFHvN75h+G3dHCfRr9W+YlG4pzvimatv6oT
qW0ZoTh0ZelrQdoLQ6xxsVO1fvWlyPCL/ucY3WPWeUSJG2fdLV09iFLvyOeDwUmGxLlkpZOrCxnZ
UzATqBa/Jra1gqeOqGdL+CqMXZnc1l4h3jndBwacFZr/9F6t9/lBB2UumVCAtWUoGcPP9vOPxuxR
ggthOdXR47jwGa/y3zfWcBbYt87Tqcug+OjNqK2bCBX+ov/Q9TDumk2zpD+Lq34qK4TBxbYXz5sG
nb8qKbjRLrKF5roPxtT+qlNswqO+iGUj9FzVkxwfJgxXuHVlmgwxwqraRkh+lEmkXGFgc9jtbjxZ
HnSztAsKD6uxzHj0+Ew6NI0UftWXXjYQR0zXgXeAfg3k62KdH8+3LrDlPxf7vlZJoZYA3dUQUNt8
1xBsSVPDcihC0+urWMTCVd6Rn+moG0lSS3zO/XopCfXuADKIDGJBUuKYerYE+gkEOvTa5VKOHVqf
tXujwVRN4Zpm5m74NHd1rg71mGdHHmqNguDk9Mtt/imf8dhsaDV9CitQ9A/zEGzBeaWwx5O7AoOd
3++f6r96kk32L4nPBLRBPATpNT+S3z3s5FgLn1LmU2m3Jjwrm2IGrMdonZceucT85AMunl/VoEDf
zK7L/z30hnVdjFkj90d0HPTmPYs8pOEaB51jKoflcttQy4KgspYiItRdb63nEaMr0RnaBTjh305d
ueMIQkoOIHueHyDsNfN0o+WeahceWbisuv8LO7P8A6CR+dhs90b/eIPpHing58hk6nixuqOOuIpg
m+BgQp8PdNnkuTugnIXfRC6EfIj8cIUofaLkuVEhbNaDZEfA6SGjLMNKAS9LMuQC7iD+QtzIgN6Q
gFUg4HIBAFkBfYuHIgWyVOOrIXKyAmur7S/YjUoU9fSfqjLN9kcO6WCTzC0vfWyIMuVweBeremIp
sCYgB3oV7Ozv/n/SXXBBOkQDQ3BEUhYxYzS7TW+a2CqqdZlRtrOtz00A3vW7qT6ib/y/GLxWsI/P
aoGj5K/fjNlyCQjnqFzKaQR38ZrlHQjG/wHfPr+6iX7e3f9QAREm7frxV1Te/f/Ub8wFc/tjhl3I
PeVJUI5WHitrjk4b73OyutOPtAyoNTmSt61OY1Mhj6FI4ZqV6Wig+459VcZ8q78fsyKzpnMBLrPO
+cUeoMQRz/dgCgaMCZaOw6oGRCEF6s3nG3tXHNJKecvPz4kGP/UMROQevSnDiltV0gE41bo4TkeC
4c2XUEGiRi3fu/gxyZcq9kUzmp5HThizIbbMoHu7ErQ6tQ3nXFrgM2295PAWLeZEaqWh/2WKyURl
oQ3NB5vL1gmNxkxC5tP3pFlOwGAepXcc1FKtAno8kWOQfoXa53Vzlzi6pSfLHnXQ0pDvhKhRhzQw
a84TNErGXFoiR1mxLxuD0qOt1CV5wpt7cwX8jQTzVm5onorwPE36RNBcb9rYdLNirykkpOuEYWkm
9D864zVzWQiQfdGPYRcydEYSfZTBNeomhZSbycJNlylx9fQ+5F5uOZ8KksvLs8hzPQA50A9ASo0B
uvJdjWx1syYTow6q1JGTb7/XAHZiOvvumhF84fvdkDW9UzbfkQvsTEagVmRPjJ+6fbWrCZFirD5f
RfEV/SaVgn8lZDFzGYBUALcl19QtLGjS+iLx2JuybHyQ6kzU2XULy70yh7bt5Ybtj52SgCBG/crU
Ca2kksvtwhUPpPoqrbTfCuYAXaA2NQYWC44CjlD5DaPmE9L24uTdhMavUSXr+V/XP28kUaMNX/dA
P5DNBs3geZQ/GarPirshnicuTd70URdkrOLeWjt77ADVvoQ0Kynxo9uGsZQMD24eDhEJuYlMyUuw
jA6S/ySka8hjoCrUEU3fXPUOIDK9dzr7hn7lVs0vXZsHzN81cZogv3RSt7w7PSnQVYu0+1FriPQU
b3/Sz4nOE+agqSAZMiXvFh0IVtNFHUmA1e2ZmPb5B6dueyopSiXN82BOFF98NuuXHk7fC7ocM6bh
uILBHKPzpowveWQNUXkV17dQovNZo5PeaRWCAJ5Spt96rQknw9Vfpq0st5wYCbRLJobGR+aZlKGp
UccRilbrRanGio6DlmqXXZoClSFLviIVxsEpJZKOHhSq45Gyn+uMPWveqxiG+1FGUEs0xI3693a4
0bA9eNLjFom5ZmPHepiFhwQsTHk25KL6qm2v354g6065JobE65tIoFVWo9RRWYwXwCpslsY8HJ9+
lERYGwxS1uuwbTrTGMz/5ztFxVHaZAGKhWKRDQARC+hKQhoXfFxOPseEFBxAMuS4FdR0zD7AOXXB
1YNc3t7pezt4sh1zt7NjO08uOQ9OqrOSVJDwRSLqNH6TRL+9SCABUq0cLOKbYYaCAnWlc2Bd7Ma/
TEPENWAKJtY2/fC1rh3meJT5vWN2gpfYSUHvTWkyfTfczNzaQOFe/mYVKBEx8dNTduBCyN4jitJF
r/B2H433Yi8BCR6qWKaZ2WvnWVs0R1ya1d2mZk++JKsRLOuIAG5rEKA0/HV3saqT19ODJ+CHPEOV
l+iKwWgJzn6uGXUg7DoMGdQIsoxeQ7TBOcVh1Sa/Q547PxEBtjj+CAG5RYsYOOeYMdL4bdFpFCny
c8l7vIPhzYq7M837LkqoXuDAPeF/a/AVtXTUzFkZfFdKOewIMyCbPEK4l1YfXPLLHn9UcLj9G0/j
QIOJtfTkZYRZTaZoDUp0cCZfbSMK0zo2qUGk+GiPy+94iN9pZFKWws+0ZGUY1Lz7VkZPLczLnzNr
xSAGWLP+MJUzf7mLzelzcM2ASI4ujdu9OIsLLR3JDLhHBN1/RsFwec1YEpvh4Eq8XAcg8PaEvh/m
1qip57/K91p3fwbHikEE9rVJgRelAZR6jQ+xdi2Zn5Sy9XV13TvJ/7PV+/irywwjR5JxvlIfiRqL
bJGfRabHR658KzEmnBwKonI+RPbF1B2iET4iA/5thTPkIl01ctHV1p1pJuwfme8K9Xn7daVodJwJ
PIUKmivxkmkZRXa3frnpUO470PPAt+IwX0MxZ7xSRLJKWEKJLxjAalLYLy5dh88JpeomRPm1uwsC
qZNWdwOS42PAgAk/vq9UtFHg+3wi2cKWiM+cY9wOkLAN4KMqNVV6G3EE1Vc76wf2nij8eJSQNqVz
69lx+TzJwjwNAF77Me0uONz+d94/zEzTKS397vN/PArkCy7V4xoKnbRKvrS8BYc1TBLueKFfbKNr
Bf285PScsVLe1lvUBdRJWQBRtwZr7LMSvE37FxtAdlyqsoB0mg7slGz4aKEyrZzi/dU1oskLHLRI
8VqOuA6Fctaa5BYjgksW1qzNTBNoIZwGsBwazi0z3krsTPtNWB48bknIL+ZrIyWPfmKWCrXhIRQB
ALZ97TOFAKNogt7C4rFRDcHwRa47e0tPESfzjJq5LY+KKb55/BK1GJVUILSGb3ganjelsvH+uftq
cyD36qOwa7nAdH1Z99KwWk70yXadvKKAbVM81iYCj86oFuMjl+UPjiekMNi1W4MsMQWEEzCudXZB
prONx53h8W58CT4OwSkSUxq6Nr77eJdk+UjCE7FHVyhkG86bF90gSryLWPpAGVZoSfXMUhF7Bo7h
P3yVsaX72mDzczIAh9+WS5fgBRviR6nggtPDSy4O/CwPZyeKA53AbPRUhiloOHoVqRZO8oHGKPAu
yFZhBc+TUd8LSNWeQSxO75rwQYpn1aWkwPHac3bwIa6drz/eeR6+Pil6nxM/MKgLETTvGn/pbqtQ
653JNjnJUeWVIc6m4dPHbKio53e3MdJPOJ2R4kWTqxGlgDvA90LZFu4kzs0sZtvaRPNJ2FcyzaDq
OnZgrTpf0HcdF0o9fQc6TRu+aoI1S+cUaU9Myo2QPxRUV8sA1osYvGH7vBVWByeA10/dLK53Ggws
TtUnUA4zhAvX4MTh2ivOVbzkrZ3OY3vb0Ggcivtwjlw0GdRXdFf+ucAYVQ8xw2sarng7roOoOPqY
jumZlId3sFSQBuQnM3RmqrmNdIWuhekIiC8NzhL9qw2Mego2lJOnGkVBqsG6R5gsQqnAjr99h2Hy
/oezIZjwKImUilj+wnclp1DxIPIMzNsbRyXRm5Xap/293FGOVuR1Q2Uk2xWByGnNBwylNy0GYoXW
cA6m+ilMc9LeZazvcE2j6sc0Izef0GjEOhXxDRLwIsT+aNZmIG5tJuqfUAk7MV1fiNm/CdJTvqOq
UQsAWlqQUPwXtQOCYuTYepdjz1xK0XekEwaurTdt9sICN7/Giq1bbk39dK/5hUCz3/9lfYEhHuqJ
ldktDr4ZEWpNn5WRwFA1uw0mWogtDOexjE4FGAFIFnrtOWyActlWsZPM76Fl8/8FJu9xON3h2Xue
HbtZVShnXX25RZyE9Owkk6htguBAS56tGDsMA6axgrSkeuYkBoYXkrDafGRmGDx7AYSGIXe31UwR
3o43cPsrNST3ITiJHb0AC4qj8FslJqstZkbdhfGYCYJ5Ccy5viX4HOg555ojidv2JvIbksbJ6Nhs
CmdlszK0jbep7LBfq4jdYqKySMXSjcNsedOWHePurFxGiiYr1lVB0IySTpv4NsVpvfk28Zpu3F7H
/zcQhYYSAQQMeCDKLhlPAmxwF1rvsprI+C3YMfL0trpOn/82wpKW+pZ6ysM3prznJzhAqgyFYmwO
Vgn/kXATVdGf8+xjyXeue3TJBtX6LNFlyd2UGkmwbVGg2aCUJpGP0gPRW6WMvFaBxAbhvLUtoRdt
lrAzWkcD7aFD/eU94CrhF/ZUxmAO+ijtE2cY481s2nXxvVtBjDnzP+6YUxy4XOKfB9fVPQ5qOf/T
Ny2wks8ajfjJHR9h+RxGPOMd0Hf0VMafXvPALNimHPKwCaVkUgX3r0t00bBOcAOeDRA3qHiGxYnd
UW0rGadcfiwv/2eyLoh/F6Qqh/6g+TWEXur63QErkEDl8Vn9I+AtEVcVZVDAFx4nU73cRHP+jyO2
okgatY53HyyEFXb0PLOT8WQt7e/AQZrsSySBkRf39cdPDZSyQ7rX8jZ/rMSBGm2H8+K7i/qjFMyu
R+jX8sRdCbl0NV/rW4x0B2R+NLISAO/GPOUlTdZBQVs3GWFYLJHkamhjwZ6/96yEULh4Oz2PKjkE
vFNC/8hKD5bNZ5Cb4R6vsx2Lnv0OT69vOdX0XLzYDi7bIY0AJejDG11NCExSV3Ukc7QSvSNOtTc5
HBgW7COs8Ss5kCgAtsvHO4E2SxD8pZvKQHHTZ242VUesIh0CGGVAGGQiXLtPWhyV7OIiL525IPrX
BB0u/JtiFeUAp/5ib87Yo4f7Yh2rX81jSDeHkyeSpTm9aU+wmpepK0nS+IS0fhlxdoGtNhOzm7Dk
cQb5xMm9uF1GHnhalFCg8Lp+HldOi0Sg5RrsMJaabp6eYOLXTjdyRT4uTXEU3PbFYzUk4iSHJpTc
D61GeqbPz0IgbknI8RDJNKPRlQE8IVhVZoULiJu02MY4YBE5CNqrxtUYgp1cLz7iEZnf4NwXVp40
Va5yO0WIZ1i/yNC9je0eNHpe8xP80HU6G8n2fSih5sH16NcoPbIWjLizCniC5mWDevW88rABF1p0
G9+/X2IJD1J1uMKgfHLZ4epIA6M7bFKBoqV/7HMl0qaBkrMPb+jS0O58jbi/twQ5u6VQpnplGmwD
vtYHKeOXbBXLUCvjTl66oTehF2pDjiD9FzGsyJqCJDrmrNblyF/KaoYniIzcnK1XKhtlS4NgLz8n
hupiDV+ov59B27dgG8N+BBZEGxYdyXCRV1NTAIlBrh3tVqYHsJtMhUvE7SPBhxYU8N7n9l6Fh+tj
EUITWp6Hl/T9C4a1M/7J0nJ9rKBKFkI0L5ABDgrmb5IfVUmxrK9uyfOC5vE5oQ2UPvlP8kd8bTOO
IUNeYWsajDzbsFzYFAK9DRM2tg1jh+jmcO5XDjoPWqJ8X1ZKrcnsqeuC7ytFoSuMiyIC/hAZkS8U
4WgJulPVHk8eGtVmJAFp58sf6ztM5iWjuADfi94dxxp66opnl0yw9nCTj9Fya0ZuFZd0U/FpjOWD
Okrb737kmlq7wfoS1XcbDxhSw+ieSYvMuT18WWCUI+Fwfk+SeJyMusRotTsNSgK96jyPFgAZMWhT
f1viRFS1NfDXlCoDO3W8HB7XMry7CS8MoLH8wTei4G8Bo5SyMes15g+KgGqIQLrrB+KW5PLlS6Vj
glT4Em1xqPado6n3aKxuCSCnnse1nAUqM9szGv745bqnQcW8oshALULWfZc+nOh5xFGUzLFoS6W2
lHau8myouieNSl11K9TQncdGABMMU5EOfZQYlyIR2kBRjTSxXJ6/BBBk/nmuW0xbxqBEKlu1Z7pn
q/fWrFhQ6DqGv8mif/w3+YzWgdp/a3ZD/cx91oeAURAmsY8TCKth4BqJE+nbTSNHlo1C6eWtOWpl
Xu1rR1GoKhFZKE1JwhZtkAfuDMy+C9V0+v4ppvlN+iPHX3uepJo/fJUoNYwsGWhLXaK7606cqL6e
IM5cDHLX4kMyauSpTlDYlGjkmF21LxV8Q0fJU1k5dN9OW7lWYlVsxoPhEBoNLnqPp+vpY8kLnDIC
brMprmqylWNV2nH3wAue9a7xPvr0zimYOgxwwTkY1CkQ24lfdKwFQsTrF3wi6mzffV7jDaS9PtMj
dXWq57n6fxI9Gdm/3ZwSGKFPS4j/V2oA9GTUvSgPUy7iQWku9rdlWXlr0roV9NYrCedClnog5nWX
U5e6aVyEPfiLSluF/pyg4wRIDjp4x+xfdT614DUPoPNE8D1juaV04z7FywWZMxyLhSe1Rl/Sxvlu
U5O+USgmRUvudqGiNJ5JIHx0Se6DOVsd89MCtfyN2btGqAqY5ZghMPqt8U0QJZ/PDPucOC3VounR
1tEyyOCMpP9ys9IVBQdP2NdDyEj+Sz2i4Rny3s9do7jDmwsmfK6UsmqAmhznxCayP3vVgxRaljAj
TpSjPFQM8Ix4qWXHJ6pYX9kcWY0+PyU8a5a5wRU/KTvOCXsBDQl/bvN836pEOwnzM8F6Sztg82Xm
wjX19F+zSJPP0eQyORn2pelx8YTu32xm9yuiNCSv+3B9UCbobzqAiuNiHtqz8P8F2INo5QcIMreZ
tTYy1X+BUhtej5VpGrAqi8r0qebVxFzIm7f8EjAi3CbnFYLcmajUYExPXkW/Z3M2Wj6mQx9R3WDt
QSE/cEBz9izJ0hkOlLsSMLZfCzMHiZndiXe5o0xKTvD6pqxgKc8AevCSLreaJ50gP514p7i1R+x6
PkSdLrdc3IXw1cH2ZiIJmnmjYbypIrkA+FwPTH4BpAKp0HlTgNEFTQFfkdrhtnYfdxlMlNhPfPzf
Oin3wxM/HqzM+6/37FAQbdcVDET+c4KbVamrSIulOcOTg9plD9gG9aLuzFBQqxwCPNO0UkDagIpc
bKEV958K13b1ZHmKaHkFa1JxXa+B5+5LHTGwC/seTDX+2MyK173wNrzNXhbxfmYPT/EwjYFDPkOc
7k9mGZdT5s+7e7/lBRFXvO4yX8Sx4V/wbOm71R1DirioFsfSEQj+jyB8j/MbHqiWk0SS+tPdWWQj
Z5b+5gH2TAQO2veAvrn31nHr/vj2fu6k7xPRw102LfUfBoQFIX3KJLf5QSpw/J8ygZtpSScqITJ9
fDKd+LcVEOUvZWBDSSAQ/Uulrvyn3Yy8qrqjwryZb1NE7N/YF2HPSysf5V2/rUEEZTBly8X/tkDG
5VTYTgG95k0Gzz8CovZhtwoqBFhCecFO9Gi8CZX2YPVIZQrbWapUsTChsy00aIjzIceRw3/UmDBE
WUgAlJaltrzODB9P6bvJXXOELPBeJSXv32aL6XpuiEpICoSrCq2P+u5tk6wlZre+Nng0JzFBmSDU
Y0MZsonxfIk3QRPPlQe77n+0NzSY1BQsYDZl8QUMc5/cbr0HR3UgLMtkLMd0bgsqVBsGu5JtTNQ7
Nx+rX7sHKX4k+sczijhPbXeWCCu0U4LUlK/0BWc0pjV1c1Su5AibpJSoyQwt/o3aVZKWW5gcj0ST
K9XUCL0vC4Swn9N6AX/RahP7CqnU8v+Bw3AWqxw7lsu/I0mkOzKq2KRQA7qmEmlrEuYnCHdWBJPu
vx162Xng7fK+xZzNxzO1NLx9hAUOAs1hitrcTO/EDzAJEEe0S/GXO4NAEOIYKG6VMGuTPkT2PlS4
qaUrG3akf8rAtsBbP9ltnOqdqmM9FCHqse8A6orx5X8Sbt/qTiwuehXEikeOxGuOPCHouCHtPGAs
Jz0r50hfOP5iJ2G2m9o93ZjJ9PNDVEBhSES/n+A39Kku3bqIsWiXhoK8ayRKRLTcgbwo09rRMkhu
WoweH7oAeQ6RY1EDs6KFnDzXfUc60Wm9YuQKx/QCMVq+xH2eeaIDDwrLAcJ1j5iVFakYZyle85o1
2Y+t3y9tSeWDkA5VoGhrhGxpRgMV5AR9akHa8UQK5JKhhr1LFY8Koj+vOAkPonPScIMSLiahIlJx
/534ucGEAEOoajIKHz1JFcAn4Ew17MsRN+OicaNaIg773jCOfDe6zOcP+4yra5hfZ8I9KXFqZjUm
wjNOw7U6Ki80HmEpl7ErebAJWnBWmBr7ySOjTY67CQthx46R7miVMyyXPFXUqYbKGqUoskrcDS30
82WZmOpQrWd1lSEdemv04kIPEdiJS7D58m7npF3/X0AA4HquIul49gukr4ThpxjO7QRdNwr9/2er
R21MhTaCL9+kv+ZjISwTObHlDLUAk0P4TvJ/gadIypWm5EY+K7D51xHldmyvyw+eIPps3CPe4s6w
xRM+1Pa9KtNtb9PEBDvkDuRqtudpSasaYdcbRZVU1MnvBcm1GXwuq4uq7gh9nEcszSzSqIyrk+8I
9LY6GVwleM86lTbW/nkEhz6NlMUs7sYEFzJyNXZ3rDpB+BFCUaXFyyUmwiORxNx+lfuWpNboxajN
CF4vkKmhbmeEanz6aTZnVBSMpQrl9b1fMoJ3Xxt2bcMoaiRZ+l7i0NeVB79UkpKTbwaiKfTlITej
IACI440cOiAi8WLUMpj3/ReT+RojwHTEHBjVFrT892zD4rw0zswZS8MWABjmzas471DJgoKxHd5g
l8VkLCcdD6xC/gP/cfjDZnMvsZUlluaEIoqnBiYhYEpwgpL1wn+ar5xr/gj868T3bF+w5Q3ViBhL
xjpMfxItslZnKFDZe5UAAeEfE+dC8wBdQuqvXp5L+1/dhUJTA6p3CcAyCgie1CcrLnlDYYCGZpVI
+WmHQ+Nvq0kTSku8cGQMOn1WVeK1Z/AzRWZlVpyKe9yTgKHZk8erfwlpiFZvaqbp+ak7v5kabmBJ
IQUVpxb6i4TPN5tG2rLbh1Ljiua/f8NTCz7oRaUIArsRedbt0O5ASCOOf4e7+S5jKDDCVpTEZuYN
+hWq3S3LyaLvAycBN6TKqBDr34vk7rJ+WW3PqRz5sMHGiLXxTEagY7QfQL8XWEnAAmksq1FW9/5o
+/FWlFyAvw8VzxzHeg0VwUhjjpZfrnlCfbN04q7VpSLjz/LGoj+iRDfAlFQuKM8sFszZCsLwCZs7
FDls4Yyd2VccpoU9Q6qQMVyt57Hr7OnkmCHMwTA/+l0dOXudQT+Wd0VIimipEgufgVAalp4ZL7kj
CRGXR352eX/DIHyB6SMCxHxWPwUf0VRla3YuNxXBiG/slevrsgWO9ryGuxlvsxmwDzCSYY6P7T0H
kh9jyUVdmdhmhi1cdgIOxSx+jx3dcith9qPxamQunmUd5wuxaFtTBZQWDfR8MYc+Vn+VrEZOcld4
jHfsSuI1R76cSj8w6grswC/KpMilpRsluJ+uiJFJwxUmSoub1P14aAkkViqPbKb4HwsGJtoBSDq1
BK2vvoOCQvcRuKOig69htzEvVytSh5M2/2gt3zc/mFOB1xzSWsa8jCbGdwZJFXMBChtl615psLDJ
r/g39nf4pJ3GWjdmVR8LBX8gN1uUMcTV2c4PjwXGabFOpWUEUAsocx/uhaPp5H089EE0KjWI7upZ
2Vs8hELUAT7fM3ky9z8EHLSJg8U/cS32JKaCNE2uoRWKNQ//Dg4daILVD+Amw6Pakb+hgIyB4AKS
j+8M5B6sbZD02TddFeLunwKY6uIKYzTva5fv8cNhyanUZU8az8Ms9PXIX2q3xonatdgoKzuQQc2E
XJmMnoBJtosOFl6OpbAzZqcrQQkpwQaWoPeDpxtnp6aVKTVumSxuBicWc9IIdTJ9S/Ezf/l+l451
8n8dHRKQs/Mu38EwCtKDqBhYnycUr1SRAHwSouzG5b2LTD5Z4VemWkuLdiZFfuBEa3YWN2YhE/9t
20H0YLWtb7L6F+SY/fOjebXSwBdqB5w17yDZsAwdi7kL5oLsFtiGeg9kahLVFRsNF/UJUHR4uvvf
VewohfthvNNpO/LFhqoRJ1sMj2TmPVIkVK4e24GtxGB7e3leFfO4YptRVavyVpB6QLr+0MQB2Qm2
v57Dz14e0fZwsSfacNq0dlQqaHaMS/cYaFybKPBTSilfr20wyfyPyntwYUz2DrLfl5zn16LYjVff
tVT8WmGeGqQtl7Vrq/ob2Ik6dKEjFBMoYmdREbIQ+IkjFjMQvFj7Ws2Giy+NtID/aExrtZO5ImrM
YKK0YsSEz6YLPHl3sBupNr2K8pr5iMKetvxlivycXKLNciT6ByOAi1z1LgW4WNNV35l1RyJaIHFU
pFMmEgmWWWmoKr8ZX1DJ0lRcxjTwUNHIukZnwaMqwOVz/bxyfKbUVfevYZ/SG7smgRZqTLyLVnjL
aG36HPcdRjolp8MQ2166xug9xnKjFuYIrqS27tFwUV9ADkOoCYx4t7S/xOeBrf3y0VsWYVNg722I
BuewC+jHwISRZgyP2qpfN95cwoUyfACZNxBwWjZEGF7YZF6sPYB4dwYDf/ses5xBJadAcwReok8v
u0qk6W6AmAPAPwCVUoNXfyi4asV3NrLOTKLvlRLzEJRLQ1OWfS98CuNZNhEqyum0cYFIOU1TIEDf
EKjnCzN1CRK7pVzf0tvXx6PGtmvVyZY3W1EIb79tqk+GDSbev+VY7U/H99+XfC6+KbghWlxSCyiH
ISW2ZgqIbW9LMGeN5MCDQkeTa/yiQhBq1Ddyiu4H8SOUI7D3O4CJaZoLYkTMvYsb91+Po8cSM3kP
qmJUZ0e1JvavF/17v5W2oLp4zrQBV/kKOmoRSfd3SmhQr3je5T5WShil4MmCkRL2WAn+2L7vSeQR
ODiSND4gwKGZc6iiZpz1EDsWpfoEcVlXiEY1ZThiSKxiGfC1LZknHbgotkqPy80+PIv84lraaOky
TOrJfVpcjkYsz+lhAnDTarN0C7cPLjrfowwg9yX7ng+JQtFgLl/hdBexN5rTsqBB9PAWMrP2fD//
xYLUqYD18hkwOxXqyqnTW0/aEZn3dgAOd6W8uZCOgOM3mwrv15vYV9WBKdbyP/lVFmA7P9D1NdOP
5/bZHHagNOf3NnLGqU9lM8QQT7FI7lTMaPb37lkBZJd2rB5Bt/mIztto5uuIzMb8J7aJaohr0EhN
tJyLKuv+6Lv9bP0zorDwtemm/2piLpI63nhCz5hsciWw5vNdSdt3BEtoTTI2xmCj3VfJFpuCnsbb
mE2/Q3TmBtsMMEcaxDrZc2BHc51EcWc5s2KqA2mC3ZIILhV2rOilYSSXNrmurS8yR/MchA7Oi/bm
0wK+vDcqyRaKghgOoE7YNfGQNnu625pokb/F+gBMLotcAktyenWV4MIdyo9CbfjopDdDCaV6YUAd
+1VA9KGjeWpwTY5eQW75eaSvz9pOpPem4MxD/ObLZ1x5WHmlNx961f1ayEsQp/fq8Bfr9FyB6KxY
4LaJs+Kkz+Qqj/iANqkqdtN25umQstUHwu5J3lHuBMo58KsKIcps4EYAhbrszw79TvfPYso8nQQs
iK/DzrhoyBP1SJzs5wamK0R0+Q2BVP04/qlF6LiGEmHJmGONogrK6BNriMfbON1Ss71p6KPyegBc
BsXZ6eHTZf+/fYxE80LpjJV0jXXSprrRH3L5SdPWGc1m9wfp93dEP20fxrAdqwLTe6L4/xt7NJrI
7YHSAHCRtde4rSUJXSDm0gtd91v4+1PsIqJe1CBlWy91kWaNLIvjZUUkCMu7ASZO0D+p7sYJBc2C
0MUswYxE9HteI8hZ9B4XSUUUGurQLmqiNmki02IZJe3K1XwDzPcIhk30KCUkaOOcrMzNDstl0iEu
b2dqCVCamyL96I3FdREPMn55WnUaRSIOnHhWjKLQkQdgVnLPG3Bn/WvfNr0uo0d0qSlIgzbRoHVQ
qb0bm+HxDAvahW0J2IRySFhLAErpsKDjL/ZFlSDAk7EQPl40pS8R2+G9qmT+JmYSEPXquX9+5Oxa
kv1fD8V7HbaMuy6TXyOUwAdtOMIGZ3/LCmWALceMPRxGUqJg/Vuc3D8Ev4BhU4tLc9zHUvMSQefe
knfzcbCDEiW6/sOIYCsy+avsAUDd8an7Ws5DN2f5tlKJ0OLlv+3/p/GiSHbEf85d9IMZmWWcbe8q
w/DFF1r/yPWPnKnr3IJeVSswq/imWqhRJfWtjTBA6VSSiGKfMJUXQWU6OOtdRWxaLe2TtJmQdO3z
Co1gnKb/d6ZY4oQN2JWXeADWimvlKiwRM1rEZE4MlnMCFPQpRr40MGsCvi+WQElYB47CFYcOxWxC
QKGRkz5oeSh5ULEAO9gMYcXFmLDk1wlX5hX1rW6pooGVf4SeCMnE6N7DyqL+c9PsEFH+nX02Vm0F
WynYliOAgxRHkQxz4DDfNhm8/8vZAP/uSjsykTv7mMgBU1kb52NdKbKYJ3tnVu6MR3Puxtei35ye
Jh+qLMpqHYIu6qg9af+7yXdPwg0eL/tRBOGRaCPkEIEZ00jKdDHjT8WbksVYOVCmtaaOIknu7t4y
VZb/XxlLwzK5k3IwkF0e3YTDgQ+x1skvj7Aspd5e0J/lxicho14MTB6VGt3V213O20sIkAqebFi3
uMvlRDvtjt5OPUtrLV0zaPX85dCIKaxOVwDtq6PaSCj+E3Z4IiFm2O9yUEor4BPMahTlcYFziqkC
YJKc/PkbS58wh6WhoOB+Sv8QkGEDAncEPAn4LFmN5OitNh1VYtZF1J9h5qpmqboT+kcUblg8uVC7
84RUHF3DbEtho+HeJ336oIL0nhggJdFGgqNwp6Q6UxCuMNhCCIPoMm2sl5cNsY3HDMdUzcgP0Bw7
76cu7tf9+0bltMqGGoktgIM6WSpH2sNgSHlzxPkaxZfselkMA5F15iAMR4Z91Q/FRC9slCkqllWp
K1P1Zha/LeyQRGFloM0LWbTutgJZUSQJIXViUtS1nc503O3FH0Hhu8CaL5Ea1Ww6oKKcR/ZgCyFw
M+nGUqhxKVFdXHkxAxa0wIMsrtrvFTmAOjgrPh8Ya4SkfnKoRTVBPyHqH+IzbT4qEkrNqE0VGhVT
XtyFD4nHoJqoQk68Fd+nYmXri3sDWTh5Ncbq5zUrxamDElrk1KnLpaM+ti46te8YD+2Lr4DGTXdN
AWFieop1Zxga2UbnpnLk/KdC2bfCbjlBVq2ZWfnfNKYvBm0aQrhNrRpEMTPpbJsEJMDNlwoUXFJw
d9/mWrOo68WlaLAr4fvarg3FCNIrN6RlxlvJvBHVfit8rktUjLBWiUhokFK13Oyc3GHqpz4QPOJx
EAnFGyH+zSWya2FciWC5JceDavrKJLBh0fXbnz6wkTZSIdduPwZ0xTYeg0MkJi2XPyae6e60JCP9
LcVaIJTxYWGKHumfzBavUb60FhEO9/rbKJF1/SEuyCaRPgWLLjlDm6DEpPZ6GDuPfZwbloe5w6Kf
XDW3SEOGeQnMewPKuJHaXjrY8Ba5cisFnbiYNythW2w9oSuzL2AuRhAJ+GtVf/P5JfTBxiesExJq
gSP5HIpnSy1hB9vlB93Vj5z3drjq4AXCtvrLue7BK4spcAcmu19ZkFnRUt11HNkPLbnF0p933eHe
teIkikf6kugo7yD0t9WToZAwi3Huuu3oWccdd8NtqApkP1XkSkjL841+GnkqtNv9/Nma8A2Nlciy
4bwv9vi0nWXt3nlv6MTK3+aIJQ7CZVQB92fUl3pGngWd1a4aG4j97J1PkXeEFJTXS3COfez3T/89
lirg+J2s7b479a/Uv8XXLv/X34IfDSzRD7b0Gb+FvcQlohGZCwUfXDurD1UT2yOdmBT55uHka9k3
0+v9GtroqvAFO8ZxMsSMt2dME4GnKV6zuKotprxalYz6vW3R128xGEvgRx4f0tboOkFDIu0DpEd6
TS705r3WCOYkNskxraWRfnJg61kI5380eLFqJjfmZii8AcR8vxXWddLJVxYiF6SYqA8bTsa0navG
XPY0JeO2Mn+1KYLPMn5tYo0pKmt8cM1Mjp0EgjG5Gy7NdlznhemWTvVOgWxxUkWGSAyZHchsvTDd
RTZGD1N8ovBJy9AICHzvpp/Dp1atXRHyZONjR0ShVpci8z6vmOokV+DiF2fXagGBiMNWtBpeP2hK
JYxqwPombt54kW4S60TxSsHJonnrF8D95x708ljgNZBu0JX1/Pe129B8N9YCr2OtJfaOK5/NrAyv
DzwB0XEOeQRmPpDPnogOakg7mtFvPbAf2TLZbYfDJXGh69Ewpk6tybVFjceSjau/GcAof5w2qW5r
tx5pLSgUA3NZVN9QuHLiCx7S+5C5KaeE2UpsReBocQ36OAM8wmy9ueIAeb1s8a3D5hHP911a6ZFg
5vum5zafDRVCNzarFapxpc17FNTorMCL/4TBdxdK42sivK2z89SdnNKxtWaq4fo102FYO4QoK1wU
XCpv4yx/bYHBlVauIY2j7DPfQefoE5Z1q+N4eGRnuXqBvBTp9ENz7ZgDGMzHcde1UnsM23XPMPdU
+0N3jN9KZoOVs9Taea05mSGoP9FcntUGiKNqPpZ1z+ThsB4jwdK3woKDfsgmEIM2ycKbBgIysRuM
BFow5Q3/XXhM9S9PiU1ZCcODpItShwnWKbiyKkv0SVhe6V0Z0ir5CDw+XCQkmCaC9m1hfqVrGNcZ
eiNMJX/gnis8zkHd1xvGZZm0WI63tcH4grqB1c+FtZyMATQMI9F22htniACze3JxHh6D12MjVnys
cNYA+IKflmEO4y+AJXbE8JvYQIDXtQ/AXQQudjhMuvUwQ8cMKRvlhUNa0rn3vxmaCLuHam1ZQ8FZ
GD3BPQEB8oce7s3k2610ISQGeesgSyHHgG1+GRxfYMr42I99AJOUrIeV+0d+7QaHxzyMugJQsnJl
y4GQUFGet0sxPiOIS3//COZHyJdRMUMVoTo0aiu+ucGaO3zkf/9W8u9UvmIB71JKNiVRwj3F6Z8S
YaG1QS0B2hlfg24w/n61TKkELOU267MerR8p0pdi/NXMGcBEq9i6NJbAqtKGowCcTel/1bOdyr8j
e80r8dtPGIS31RoF0Ld6y18ccXmi+HTfVU2A2y6o6k5o7jehdxR9nfbl6hUBWwe5vX7gwJXla6Xg
XD30go9dgInHQyUe7S2jKq3EnDweQGuni9gwwJrtQ57LMuXIuXDjywgtcBeuGCWtAug9pdcQ5CSH
1EEAw0xrWd7e0I9+RG+hxFfzupX56zcxeDAc6TdBcLs2qKyH6vaXg7Aj+ekmDWW2GL4nhnEqbhy+
ShuQnW+Bbq/18NwFbYCfbC6ZllhHwVkVM9gzCn+HamTSO4cv9KYUHQ6DpijlFlEhXZEcXLBMCQvt
GRpO/3i+Awpxwd6u7I9AxVr707R7U3HdjXlIdCyx2DG/dx0w8pkjIkRTmHOa2vwbaksOqXrvzhMH
XXLDD9viR3SkqqgJQKW5qO8C/3oahQyQOjc7HcPOEJo4pJ8aJp2PprHXQEqs8Te1x3RkmoFIPkZC
GcgS+wFmRB1DLDUdEF6TZnZ10ii6For9XTMS58mOARVpt7J5/Qv6MfJBy9fyeQXvn5lrGJhqWH8t
25Z5cqk0VzolvpMpmO3AbzfcLOT3LpxOQaAheWCMF+J8HENkI7V16IeWb1WwzGKoLMgav2BO+5Pt
oLO+tNwlkrM3IT+OMZnkV/IRgwplG+LOGNnnP/0cWTTVa8pWiZgYF8OImXuhWT6IvUAXHuY6Hf20
7dpst3NjSRqh7f5dFmnpOgEI9FAsnW1+Gk8iABHRqRipcnvLes0qc1VuvMrYOFJXBZAI4fKORunv
XDZnAaC+Q24KZhYS7LConzj+RK8BREAiBuA5080QTLaGDqy2mfx+qpy/A+/OmtIzYXJPoztKMZh5
cJACQPd/X0vGTvvShVHha9LkSKjkgMX3GEv3a80f4FlNgvlb6gsohqZTjmnE6HJjWAiu/BCyKF3h
NmFQ21ROwKX/yO0P0Y7tHOGVxgSxvVIB7rvafUjah40YABTOUZU/SDX+qpxHFivKLCnxk4bZRb/3
s/PYk9pBzgHHOoiGoI2MQwqamAGSIaMotMePy/5QYA84eUfEkXCwUTXiJQ9MiZEMMWf1NObxBTW5
GD/4N7i/cFwJPCS6hiBUo2mmp2UQ9VDqs2+RLNFGux0nwYZ/tef6IGZl4On/hp2VjCAkmYcno6wq
8E4/Buchi13HVNGHhJ0O5s8dHpH6TX7mZtgPjiiuUKMYXOFludjiRU97q+8dAOdyrtH9yVA/s4y8
Y23TotEOPDZ5VHdC1P6WnCNZoyo2FNdyF6AzVyZlYHyuQIu8s5kX/2BIPSlRtLTW+c5Ij3jHQgie
6XZMdY/turlNeIAJTjs13zZt88GFF8WXDxg3rV55UvvpYf79Nu8P3y+DpIwG4BamI48Xc/4senmV
A9EOO9qJjoh2cZ5iKYrH+vqoNP5O3EiOrd5uYz6YvaGNiFmfHsJx7/0hStBnU5lScYghyD7p2tML
t+cbXmfBw0jSZUfcbxfwmTJ8PYUIbU/XCIAGkqxQd+1GExVYoNAYVo1qgELN+4dVsy22O/ggwL9G
Hl1YrmS/PpzEYZMmjww53BQqhhVw6QEvnFM4Uq8LTsoXQpd9kRT+4gotmDNy1gnJtyoUOixBuy5U
oMBiqCRWtARQRiIrbf8Grf2jzCOVT8FwGtfNQStYeKjNY4QD8IZcoAp8wqAeUA5lbveWGRaen7Jd
FoQFrVEpWw/xKBbKd5hL896ozp3HNiQ6cGjj43QmdPB0eaQh17VQt1B+jSGNDS/PmtY/4F5TEjHi
zSWpPxKzQ6fMi5wnnMpeEXxCreEkeyWanU6tzs9HYk/jqAfOFWxrDlUge4Z97XqMjBfyAeYjsyZN
vGqwyQTCtikGm00hE4eNWW9XqTgO1J7OwGvt9uwDc+QtkhCKOevSGJS5dsxEhkG/MbwQX6nL9uu7
3jyDYsXbfxk/dNUKA4yjSqnuk3efDdpF5vVSo7+oi7nRCiXW1g2oc4YlfUozR8U6uPLdfaq6kSAg
YObiJfAX/U0bxz4OYXTzTbyfeESvvsbK+wDjfHMRQq2lwd4mq5d/Fx9x6Afv2QuczfCanQzM6uD3
2ybmR/ZUIwI1CdWz/GAyox8cr3vT7KX9yJXDBxJ+fvKNJGsLTZmq7my531yglfB0clQF04wFZqUa
q8D5z9LNcryqEH/HtbyPrjVR43uOwca3+XzSurEm8rPQUYSxzextQvj8Sfm3rh+PzUPr8l3b1QSh
uLqxYU0l5qLKoVQ6TceGQtAj3VJ8yCIiSk+if82QDAZJXMFTSoSjaIuf0dN+VeZfvh/QQKJm6jHA
H4sTTrF/dr5+TxFeCdHZAaVwFHH127vsAzHjZoidbjAxMOWugNZHqMo6hR92HivyGaL1cQkm6jga
T2LOKZVAwmWX9/3UdG97Upvwh/+ccTZiWGz+crTGOlEV1TgshNhV12o3amJq9a6sjB6SI7D7Rr2y
lTcVr5jWzcLUPI26vVLgA/oeE9ZEuJ2GCQLwwjonGhbrYTgRaNPfBWHvDfY1knWT8JPP39FAbPl9
f7Wa8Xizxd5bw/TIm2ZB7draLlPntDqUOUZaGxBXdq7G7uY9mRB2PcTA/hVc+wyUssmHK6vbQr4w
GE17EnmEhBoPyxmWkiKlDMTi2mceSitYbOlgkt9YaJRco1SMT78/6JDFfnPRCqnLiCuuSQ2RvzVQ
fBjMERwhtAcf+1pqg9sc/8sfFga/EYGlaqWnBaMMm1G+maEC5GtQMIUuiCrNiO2VEc2t13TSFSb6
z3gw5IlUpvq+PcV+uHv2UUAxuVg5TzQg0iUZaR/uU2oWQgwR4zegUIUIDSKJOjVbM1MB4zSrOWzE
tt6W1WVYOnwkSrQw5wYVXza8zxSjJZ2Qo/Yp/SgqZ+UQUhONVexlmOzRlDvE25hevul+eeeUq942
+TSD7kznST5L1tqGwaYVM8H4i/spL3pDHjw7hE10qZBw9zZ1qIfJEQyNJJH1MNW3XRXv8Pi0gece
io3DWMHeD88lgP1rcXc6K6sohfkVro+hSNVYXx07bh9wNjoV/9bpRd4gIYKGkmKYCys2ttv1Ihbr
5GSWFLmmD6DZs5/21m+gsPiCrv3uJXijuAbK40wyPyuOwm/hA43PE0Mos721vWBKFDmYwcvUDLZq
IHfs//2eZ2rBKIIe3qqAIetUYeM0na/HEAsG7/xTIfdnHGQ0c/0hDjjzreCQMLAIcdZZhl98ZMn9
xxkD5QVvvKj0wN9S/29sdFfJXcDB/l07Vnl5+AuE7eFX7fDJ1uUX2ZN8KsDMKDuGHIxTNaoDKRt+
NZKoQXge9zcYpFvJt+3XnN7gQ2KLHbycVIgET8SmNsCcJ6wsKL/cFrb3YIsrld90yu7+IlWeKNEv
qSA+chA87ZPvBdPtnXzNg2KhS4AZovZ7whXU+FGhVFYcz6xIlkXRqRinrDaneaOmS0OglEwXpu8A
fQQF3ZkJKvxMJ16LYPP2E7monVm3tD0iLzvc5abnzrVFlsjV2O/BAGvywJY0Gx9JG9cWLI1ziDfH
bVhnGjIc4K24h70J2hD+jBRm05KdmnBzPukWvR/zterPf0tysA5DLS20NIueXEH8XEStLhE1pNCp
YvTTVh6G4/tyfnf1Xq3F1kQubeBjuovsaERoHdoVrBGLqoTjPJSadK46amvs+S7Rc4jkb5iIZYRe
oKnFmpgGTYPvCSWO2jB4RgBe6ukLmZmX+Bzj7YUAV+yuuyg2Q1FXJMr5FuCzuWKzSI8Z28wsN3Id
XVf38ztrb1nb4okQJiYqGcFi5+RMKi1qUOdDJJ1VQQFXZoFvFgAaXXbQA762Ngaca6PGUQ05he8r
i7GNvMvC8FUTvK25gLKOUggyaSHbq0ZPUm816vvrnzvwJz+D3qBG+KPdSwrIUUadvYDoD5xbrpuc
jbpuMkjoflTCAqejN26O/1GY6FHDb5egwLeUREhDEcGF4uInrFKyJGpAVcT0fGRIEIjEsNMxi8H7
/n7kZGcfrFP8NKhljY9U6TXhEXACFrq4CxhCh+6VyJGrTpieOjJMacKFv07QCkJ2ql9XFs03cuLz
5DOhDCIIHQpm5mvsHGXcJ4WtAbK8qaHk8tvA0KVtJWTuZPAvIqDWOnbZwYWEf4Eu2hcwVq/q5pHJ
5HGkXsS91sb52aKTgHNDPjc0OEacooQANqbhTKJUKcokUembkZaqcrdQTg1pjn5J4I4bOoaFDrA9
N6Bu5hN5FwCJQ8Y8UV6y4JIN6vgG/w/H+5WypC+hgbxDsEDAlC6TWougwVGoPLBAuH08QH4LPRrb
+oD4VKLSJneaMeXZqqJNHjoVQvjg+hlPK9sLSyBBp8OhNEVl6t1mfdVoatAXYV3GakeA68K2L2yL
S28Lms7fHW0Qz5/NI+07H0CV8/ShogmETXZwwibnvXVHeC7rkEkuXpUYUTw08lEu8Uc7vx1pAvU1
ENoFQufQd+/pHPJSApI4VmE+60RU9SpecG7Dq/Xn1PcyyrB1JPhRqefqvE7QgtgBCWu70yB9FeRc
PJKcqiVmMazJKJqwfnSB4Jej6BgxTKQBEvo5b8ilaLXjBTPaJLlW2LagNW+Vlhb3ZwdapNVGvpu8
UXb50CkiYRb0lGyswbWrWc4WCZ+2MajSNKQxlh4xOVEy89FP9RlhCf5EexGdYIugbjAekwqBmKlG
NCVmx7jS9icQtuOMH5IIat+lMD9zk8vpgiS6lu7DwXl9YHlKCHDSPNxCwdEeFzsn5URJaf8cAEZu
GzyDzlxyxS4YaZilWlSccfg8smdsjOGSWHKPhhMuzCc1mbHIxj8IE/nOxazK4AIn1pC4QIL0pc6j
/Ska4S1GJ6G4iKu/8RYSOTsBhMPjwuGD98n4kp95sCCk48aClxnR95+X+3xPCQO5VQKj3ny+R9jA
aOJA2j0sjnQQb5e5wbBv5f6i7ACG9dUMj6YryFtaNSWZyd0pyesZITnjqwxQqA7FMBesc4Vp3Gz8
XvdUwT4AauUTh7Pec/8cmux9nVkLMNwMizxswiRYRV8eN1hZLvzYm+TBq7pJkU/kv0SvLgqGL4ih
GmfOlgxP75u3EC0gvMLVMb/T5HPUSeUspLMp7ypnArm8YdEN+nV4u/7k8vywEoTuioyCbjXUJ9Ec
vjwQ5yUfhPY8VMZoKDoKGe+wBwV1Upi2jPclVa36Rm+dwDnpZ8XYxMcdJp/DZfhnZkBVmw4q1GoF
xfpQKNb9tHALBPdER9OCFuyKs81/rhv266DcEAJ9Dicew/52wDCf0LVFNTKpJccnbMd2P5ApShGw
qqmZ5pc7LlsdRhwWG2RSA2Ca7vMlHILaeRPp3Kr1sou6pPggUc/GV/05kihnxcskWLdoBBJHIepN
z/5CLQtxs3/fQR/8HmyuMh94TjHv+Mz5T6o04gJt/a9fy7eg4VlJ5qYCTQLoMBpSePXHCgrxs8ms
FPpQxb6gp78+gNZjw0HNuYE9O6Yvm1IA/S9ndKQ4SEcdHJMsBFFzxztcx6BfIVqT5249dtugcQ1u
C+F9JfN3KH2Sdv5Wo/6vui/ZJQBt2SGPm5GhA2sUkjTwYMKOwMDTgq2RuhyegdA7PkO/nLNAlbzk
789odnNm88QJnJ7vX6sN+JZXEFxPx7AsLtHeDACFtlbqBYjmEfKORm6khViIR2g4Q0CfmV68+WBD
XaLGTz7q4MJ+Qs8Kqjv2QI9vxAWK314QyThcXJkQDae8DeutWVm+yjkZRiCZhkMrDH8VS/C18rtm
slt/YW9RPvy3E9UiPc1LolFE857Yyi5dCzPlRh8hzGJzv+rfSeZP/K3PNZ/Uy24GtEtFV+X0wDT/
sZRwO7Un4g7fxrf3uQFZCfM/5YVtHI3i3OskAJuOKV1pg6pc8Qv7JH0XbleNY/OWBqAu07XX/kl2
cvqkfiK0XhFlpPZLwabwC7k3sk9qPqPUyDCtuwuxDPY4x8WxTRgoCJtAkJILy87xoGY46HBPzsQL
Tq7+07SpL76JzSRsV34/Lm2P/0kBDOfOpx9v3pIY5qgQTZm9qdSVSuumOof2j7hQs0Bcdk6FLpKy
+jRARkeSYgLgG8ueb4+NVHn+eozWIUDbDKhmZDjxbVAbbwpkADHa4/4p3zCETGpkvhkoEHWk/sMT
E8etttQfyGRsH19JVAPzFfG1BCmec4axZtZsFOekvFfQVbdibKLAVuGpz13F923U01NTEVVoIp9r
FsBBnKQdqcPWZBaTMhgKWWEyONOQxuA6bNyAvDf45ALtU+LsMFlZ442QUQzH/jUjITJ8iCWIG8xy
XQWmBydKc0SMz0PSJE9rpocHyqYvmaze01Af5NMCf3jXVdFVMYKELF1xBaW8TfrY+mFbT2Issqts
w154VvtRe0eVzqvPlA7foTzgfvu/ytDhckj+XTtudJaqvdGu5sDENOY4cvVXUdogo99nNCfymKui
HnzdKbP3KMjjwFpuwU6m1MgEgh1Gw09s1zTtlJjiE5GtSsbv7l1expsMUr+aUDPiJ7N0eEzzpQG0
N8ZUu28c28Ou24+LagT60mtHrV9jex3FaFl+qLDQLQ+59o2JTBN0XeQ/LQJ8aYC6mBNbrACc/Mpi
0a1TZGWiXTG2KbB52DGp9H6VvBWiMfC/4GSr5i6o3qSC7MxrwLj/XIjROgOKiYzjTHB9W0+VzAK+
1V266UQRDK0V2p1ZQIjjp/AYOFypv/dOt50lhKIfOVElUIm2pIMG3ThGng4ztFS2VBAsLsdImXVm
jG3X7VJkx51T2JUNPi8QamDgv38lkqOZ7Ih1PoIIuF0ruOgyeIxL7BDAsHQHWM7nE3U8kfKDNp/Q
9y5DlHuMpd+wo5Hz+6fH64IbYK6yhYL6k/niFjRoMhS3xXNxex6v4Iev5/3JRnF9GeSPyUxtKE71
IXluuwSAEYGKuRXWid3JzS8F01WsC0d6+aSkP+THGTeOR1vcnIdBnnaEAa+66jizMx+RF8JA5bAd
EkgqlujUyXc4KjB7OezdsXFxgJdglZ+YJ8gDzsCpi5L8+Mz93V+kMU8LthaYwxrXEq3AlVR/L4A6
CkgsT7f5kmmtjHMjpuUyaHeUbXfY8c2Whp6TgeoePOSD+N2pOCZg8p5isgREyLVb0E/GoQSEf/+3
fd4UwP+zWVEa/fG6JnqK72t9UOfSLxuEnbcgYhWNFvQQPhmuT6a83yhX7Ec1FUgFnDfinxmCBM/p
GL7xgJnredb0urDwBYtq/S7bTY0kGsRrByvV4WrbvrGH/9jqU+RmewuYmnPKpV4rFjfXbd2iy2Q8
HUiw4P3tbZJ5Qeq25CLr3CS0EOCRCXvjX7RVJZJoC47IAZJg0nXwNHKCX0BFExcEckJ3Ms/OU8CB
27/Mg3UjUpq3verpNK39IBBkBnDVM0Ym4uKfYDfu6F6bikJU2CznNWYjqoA9LQBoIck+jv3XENU7
EmSW2yC/gLnB8S4JDhiPAO46faRPgUR9oA9c8cQ2nbdDIuxmsimtgHfnenJK8dXvASvIiIltdHRI
2BgVCA8fopb3C/pFrKapTDjLZuo+JTk/N7d55cMm6ySIvQs6Kh1qMaUcpKNbYWCvxQ7TYVUX0MD4
Az/89nFn+jsTEwgU57nBGGlhWYBV+j+sPSwT6jPIgC2Si+El3IxfDBb955MvVevlyb2To0hYU3yK
Z3NDv2F8pN0B/VTXtahndmIIdZDyVM8rMvj+d/mTSUru8saGwwOwG4vhnAmZXW5mIgDrhGxHDIEY
rlLBoSaEbCVZ6S14Q1KzmEX9cJzSXLDcQ4BS1OHn1N17JjvA2fvRB+uSq+z2MU9kj7IfB8cqAGLu
S5xjjlb+jtjU7NFJDrJnPGKPuIQ9um0jnTRY8AC7+FN8jm6pFOvr3jkIv78CmlSCw21KVzjREhi8
NPxWLKCfMuhAXnd5eN1EMkkat682fVRZndSwB00ALYqTOXWUdhg6BPkAd+f70nPvPsev2Ogu6gcY
dHH2LRuaVN2KVkHI8q7VLsHXe4BfrZLJLqbZxr52I01SYn/tPNjuRLeFSiiABt0mgpzEOpzFJwUy
+zAbET2j8agr+F2qeznnrJz+I6wSvv/KxyNR9v/NZYgy7Nl9k7M/Lu+RiRx40WlqmqCIbmQQ0ZLE
WkH29LpITXaGmdKne5mdjcpVbL8egQomAKOFpiyKgq17lxVrFFRwubPH4MlDjCp01GlGwiDXJGWL
a7RpDYYoaHjICnb9yBtzMLbUDMT0e93FvnFoXRyYZA2ayM5qQWuJzzpWQ3oWqOZT36Saxm6VYYod
Ra2iq1DmY02cnMORTXSIbA5dOEnNM4g/HOtA8xqpVtid6lnl7pNCkYJQjz9snY9lB1DsrfySKw70
vNj6P0G79SCPObD7jaAs3cyzoZy+4gsDScdhvqePsISaS0SaU75WnLsbaEZPgJt2wQRk4osrkLxp
OeQ8RYLGMeJfK6PSRQlMCenAAOapmeSihmGQ7vXvq8gGtDHEq8uDgmF+LZCm4fhdE9Hq9/rrKTPF
trqLpf/QDCEVY0PnPjWYnfF+nx2wq6Q84Dm8ZAFxjPlRX67uf/77UID9MgwEhpIFvWY7oqaFd+Cr
1VFHDSKhsJR+u2OLL+9JdZcThus6JnQwwHlilwPtM8LCj2ZZrNZfaPZ/gWaamXaKkZkszOv7H/w+
bnpd/e6f8jViAcP3AI0Tho6D2X3upohaVqIYPVS/b4mRNfnsWMLMRso8wF+ODAB8ZlVkhWAJ3bF3
+c1roIIbpYuMs1CaGGbXiykCSEV0ic4NB9GOaNsu1OBdY+sbzPVRjlRm3U4HbXEBsIXohoDi2m5+
5Dy+fbpkqYMfEydTS9VVhOOO0Vsae41xYS5GqnMPcLpQbFYtBU1JmHn2fADC0qyL/pJNzXniqTX3
e1yT6qODziLhICEGqvP4WBIszIykGw1FBtba8PhSCFellgNuNZi7Q0YAk056QGZcvkOKEMhHhQOY
C6itEkfTgx/4k1V+VBvPTfm+uE/5MMWGM6CBeiML7LemDTr04KIR/F1wQKu6ue6LORj1quhNid26
/NuTJ5No4QxPYReOPtodYfPzf3MvprM6uLo5qkHVxUSafJmlAbO2RBEIZIvywhhvb/AqvbjrgbsD
SXaGLCRv65GnEVy+vqWblJhKEblrqiHFifqKGFT1C6dsPuZyjSHCAqNt9tDrd0lEIsZrNDuzy65q
aMRAD2sMmFDbNmm6CgJBlflaHaSUK2PLuz7lQQey3ZJWBVmJ8386Wpx6YBVx3Jz2FJ38LnRryn+m
02rf6T11MMiRlCsUEYk8C3Lgl/xk/UiUkElL5I/NPCSeYcabDQPtPR6//ZcyUWxcJqGhxExglAq2
EIH59V9m5+1l3kD4PUIaoHGMzO022xTVt5Zb511yyi1JGfSJPMcAuiXlOR3vIbi31HyQF/w3y2o6
U90kqVA5E/sRgO9Efvkb+yBuWoozWm5IJ78vYoubRYtM0ekRf6tIjAK5KrpAL2cwpZvdwWYyn72w
uniJIv+Hnl8ARz+ZY5QGpg3SwKBDdruNEsIslU8LSbfnZyyB3aA1AcmO39AVeAQRn6TNudFRxhzq
9gUb5IFQ/k7/iiyaJ296ezLtKdzvod9ZaN7XSrJ7RgpNtgcc1eXEyPP2V5YUahhcbVNlN2r72HF8
uQOkNt1sxCpRdbySE2OhB1PrAFqs66xhie0slolhYBRhMKfMBHM/15hVItFawKnAyOQ3VQ8Y/4rJ
eaHFhoI9DiU8/hUh4r6BOUWBytzyGSRUWPz3MSYRVM8LgEIY5oHDmUGlrYzqxS6BeyFsf8jF+kPF
dJM3uRcw0j8/HOgJ48g+2y6zdhfQLFW9tpgcuAF5bNS+uDotRhpk8856Aa0OEZdCuRGlxaC9Dc89
NzGnrQAz/XnUu8dWSriwzdEQkyxcap7QCYGaGzoIMsY55Y46QTl0E4qrUc73iaeRtDEc8sSRrg9u
XiNitHLm5LL3/AgCk7MflwntS+Me+xfhNGF5pMvG4S1cyQOpr5Dmm+F60E1AVjH5s0bvo5lFszh8
4C44wxP6C+NvMqGjYUnxhWNNG6W39aiiMOtUMYVLsTDYCkpaPOMJgVw20hcRpuZh+U7Tu1HTWsl0
T4xZq4X5SZujAU9mrXc+Un5TkX6hJBGZ9+3Xxi7N39NoUxJhOdSA8+44Uw1j5mvlzOMzMOs3m4RS
3F8v30bzCHolxTHa1pRVMX7vkD9/dbu/sTDxQgKnFDqBaWyqaYpZAAjwnvuNBsGQyX+YuLUm0RoB
/kn20MT4EdeFsJD5xnvX/6rAjLD5zowmIs8WDnKga76pUkObiBUTqY7j9kL/SABBDobjjDxHiMc6
Lj5tSe4ygV5di68xioQlMwYXN86BSH3T5MhwVf41UfB/NLEbZutKG5tqthUhaHWUt35CSnS9OPIW
J2KR0dMQzRh219L9Y47vLgQjwZf3OpgxJmzbym+MkglbDHskTUCY6tG+Mc4ZTdRuMIohzuGajpXR
UdaD5QBJpR/C/XTbxU8NCVLONyD/Blcl/enfvyIXpwNN8YWY8c6L6qlr5uEj8oWW7k8lqW/PB4+I
IuOXW+FAqjeGi6zykko/L2cJizil3AU0OwTM07KqVFyEtcazvzmvM9tbyOYzumg1x01D/9Fnq1lm
ExSlSSsLOQqUWIZ1LUUBB/3ZxroIz5TNgn+wkByowzRHWTCjbcXHoQACSg/o5focaNm9Jwy2i5pz
TKG+mm00zXRWDFooj9nMnIdtpRMy/2ZRUzkrhDOidihqvMqY9s/OgWmsLgbD6CEr+w6dD13kmq38
xzZamo4OWOhi5sJ/rPoBFTy7U1vrwRt0/Kznq1BjTu+TTPH7deQ75XDAWGsds6tc+WsspKN5NRnS
2nN6wGHkKNTWqNuEK8rgFYqz6f0PJqF3Cxoy4aZJv3vjmlqGdNAgsq0QL50W5mmxGeSYoO7kIgbo
60RYDD5y0Qpugaaux4bsrtsu6lNZK4rx7JpyqiPovBz547UZ5GIcY2F08uEwA7QiasK8MxdKTtxW
VA8EPGmqe3xggrzRx0tz39NxtBlFADGhryZ2STkvEnFXEcAqv8PadgM6vX5AcbTNB9Iq7zhBBVVh
iC1lyaSFubnIDdrufxWUHpKqUZ0GUBNieHSmjE1gwlo8z1o7oPasKMZU2ofMVqhfI9jVWqgRlbxM
icgdV6KnJ9EthedpS/k0dWurcRN8dVCH8iAZ8fLZsoxmCgO4HuP6JzmcCvgKQWDSXix5RUTODyWY
c+dfAb2A5FgqOAaa55N6gHfFACrLBhNRnt9bqEOCaz6ydXustIRHPeX4MzZwEYy+M3niZF9fezma
9mjCRuNtSR/gN/iFQWvOlXD/YcQTy3x43uX4W21keTU1dI9zx9QI8ALyXCDT+L1P78EspCa2xPLU
q9ntnBT7qHkT1BS+8YQprGIri8vzIyHlLsCUKwGQ/3lyyhB0XPyUp3SOJbqFjzL8IqO7EveSzYPK
9bdPQ5bnAKrF4sV2XKq7Y9uoVzVkQ4+snVYlopXtddRqKakV9NKtriO/swrMA2kT5jAvT+BZQOaY
THaA0raN/eBisgmiQHBs8kmh/Cnw5C2llf9KSwhhbkINBKPJuPOVp9FHAUPSglO81RMlKiw2BF6o
R5cokttK7X2KXbzgQKlK/nR94LkOGZV0EUPmFSa8fcCu6AxZ+YnTVjlhUL73a7y1KcNAMvY9oGY1
2kKsMe0vpnP/uIGbbVbhzPgylqZRTDJ0PITDDXR1W+tDWVy1opkEsLY8DjIHH1sW6lEXISjprgMR
rkCYm6DPE+QFM8uMFr1oBhiddZO40yzqwdrMpfFcn4cJGNv8+d4nxqW8srdyLfUrO/vyRys7mmFs
IsQ4kplQkVusy2Oa8y6rdhP2g6+m8HPGTCb/f4sGkbhGGdEVa+flgKkjPnl95hmqi/WUPLAnikyE
H/JJ1Ten9PjYehgJ7GTuzcxuCwHc5zMdflWnLmwi6IMVvaYweyetPxN994F3iyLb0jo2AweagHVQ
tkNC0K62NofuX/HvWk6rRs5L2VD6WAMVjbVudXkEg/sQbUBFRo+UFNped75q6yZ9Cu6TqnUW4Pzk
Ity6Bo1XOxOsavWmnGT7aTP8244aYV39erTW7L4HVSwNgqCHio3g1oEZag3KrEBzhj5kyV3tCcOP
8UlCJkp9GPUzMuuGzSZt332NoO4KD3ZVaxIjLNsG+M3VK2rpit7GoF7LFNxLjSXfAfB+szy3cYCX
/1gX5rUcahWjlxUjNwIOrF4DdIxxCa3oiHa9YMmxfCM8ILXZaulDNf6mQGEDv/wRDtJuFvv3rH8c
nA67xZwrKNAfC43BOHw1CRMCTjLFAbPUJRus2GseQs9/PkHR+TdmBLUwNfdbRGTM1U0yZO6lrrFU
22TexEd1HLJQn+FOUy85arZDoaeN3s+WjBM5miXhFlPdQ2NfFLB2sQoGzGo4Xm/5lHSwrb7Qz1PJ
+U6x/f2Tn+8KXE1gByTqdlWZYlawxUL3gkFYsXjaywC7vGt8xoJ65heIE4nQATlgbWgpHJS58h63
xA/f9dBG4UDHAN3t2Zpn7tz3wtR+GQucNrYJVHWTMdflirEyFTfsDWrFjzAQHi/FZkge3vyfj8C0
1UesgBSgwUgYSAnMZK8hUA1ooXf5mdNkTv6hVGO7hXfdeL1JmAajdHj0ESuvXVdX5plnNTJLgO4f
BPMMnH7MIkApIrYQqBP6Lwown/jbRxMoTNULvZpqGkPUrH0HnGbwn2cNuPwdCoNkp2G5epM5q5Gj
GIlZSjU0SAI/KpUsbnTvndjQiISKA/Vx+PO1i6vhR/CM2SJpCCslyjw/doccEQ7kR+A3o3ObD3/G
dzUYZbith4WlQ1aUnvmYkLAq2UzLYYc9P3MoA7KjHnNOiE4hqVqsgMLAG0Y7oCMYYJDuegj2/X32
ZiWkyWAoM5/oc5uJ8seEPdUIFYeURFskmotTdC865Xj8Jaxd55XuHw2Zv2xUd8cfwjS7gLg2KjeH
uf3ddA+hymsPuuuMuneRzRIAhTH1sEfxWamu1EoCKk0GSa2fWPO9PnPujavkiITYlpjXe5roE05o
xRiqS6koBWgKe0mDjA0waNsiMj70YZ5zdhDignxyAbhrWgxpHO3ljLK0iWiJ8Vb6pC7Kq8mEn25X
uIaYBH1r7mMIsk8rrBvlMEc1M17s/41iWUlwcp5ey8yaI4nNQJIYMyzXmCHwI0Bxzkv29/JeO/Ic
lHKD30/tzUtzJRu+uV/MSiVJqCWt9GjpBkQ2/uU043d/l0u7T5LqQb6l7WpAO9PCcsf2/RW3q645
pJprZqXDXT/ewnXRqUWELnVuKeN4j0frPYPjk4vYE6klhp4kcXXewCbyrsP8XeeclHzxkVuuPrWf
3ZDm1g598kxH75GDO10SOWDhtJC69EFx028s68xklI2HwQoswY+k0iTc6WN85WR1P0AaVSUxgHCi
4/zQe5lSxAtKu6MNjwFyLWU0h+er2DGv599yyN3FyqzkiZh3LYltEo6kTlpufpfQvqxgIuzqYNkt
UIRkMv52lkuv0q5qlpPuvGau6uGdmSb0P1LYi8MwkkCeURD9gd1QQ+n3BdGgv/hKvwYvDXiXVEzo
09StYAvIGHzLytbUvlX1g/j9rJ1JBI8+6bXVUC2+LV8UTPr63LrZgK67dTJnD2lCbsi8BFrZyMLF
nLFbXb3zUBKi30r+SQsb9SlA7F93NrSoSORL1MuDyqrVpx2K/ZWH9977hUYJAysh7G/3RicBisj7
t8x7kLzMCEOoyXf7MX6+SUaIJYiFkuzsCI1QABt4RAYjAz84BZv0AjelQixeEe0FRgwYITMYMLOt
7/jjxQXYEiB49Pfu6TNpdku9BJza9Jgpzo4IbsjyHEaR5ULnGKTyOKc958BWsfa0grEFmw024q7m
zFK9cJykJP2dLf/Cl9Gh1VIrIG98Mqljvj8T6asYdlFZRY27pXs6ZS3s1nf8XohhBCgSeEDzJo70
/iRmS3qHSOYn0TU+W4I47jCRGDSogrY/395LaBGrTR1KeTQsMMCRmkAbpdEf7wgPNVUhGMcfKOzG
tsKnJGWcldlgrSwL+SK63L7PRZLV8jBkl+TuH00MenZSXdj9sk6zioHcdbdibHPGOCg4Ne1lrDSx
XAyhNIWyxYl7hsTBL2qrOr3/xTpLxqcjvrpPcELaUPcZHfdw/lm/JyLawF505WFJbTGTuCGCnhoV
Jjt0AlJiuQH//96Oyll7XFXWMhqXjNLq+rph2KSAkV25eV05OKyNv0bY2AbGlJe76LLW3+Rk8nAA
iTxegHEL5pGFB8NAobf+VvlAUXUglTZiNk2XNRhFKxZ/CrZiibOIkjamV7eXSSxo+zukhWoMmFGi
z1y3R7CcA9V0Pb4VuQS6NOSLmOs4V6+rOsOXsreIrDk6K3fLtll/LK9qJgbuVS7ulRgJYm5aXst4
+zXEOl9fcUjbIY8egAGvDALhQ/0NuoJ+Czcg0MIOu+WN1S9//glDAnXx8KgOKQdFmulE+RGNGn8l
jjJ6yNCSV8PfyBINyqsVYQ49KpN3q0mqDHCWiKltlxElrg5DJSw2l3aOPDlZO/+punfPuEWxi0qa
7GVjhdTnu2aUdYfVY+3fy8qvyyRfS9ovpK3oRJiHyJ5zRW1R/g42LuQXZcuqzt2s75slNlPPR9cz
RgY42+idY5ZheNTqZVuB5ACAWO0su8xn5mIbou6XwLldSFAt/RO2VK/k42lvCklo+cNIfQodqWzc
/otg41GU+HChIqEAt04n2ui8h45BXVhcjz4l6loA2ln0SCn3Y7Jz4md2xLG3hvgTp10g+5Vr8xuo
44vHbm+IneFnPnNYRQMeOCymUf/70Go0Y4W/9SyD5XAy0F+2/CNOujOR49FJJ/WZXW5gcw3Z9xlX
XVO54rIh/NKX2JfDlBaiOIUvxObWprJtfXQwSpROk5aUYDufzXj51u04keP3PRuVHT7rt3gxV8RA
qRLXeT87FvisZJJM2iiRQn1fRMwn5ekcDGuY3kUUY5QXScoxtAQUFYmqssiqWJWYSbSGH1qvYVCf
qy6AXaVcTlURZPlYB8pfgwmD3Sr7Qtp0fH/BzV6/yr7+oQBmCLVXYiQ25N1tVfKFju0MTYxIkK0s
kQQywpP4VbIHdhn/Q5zz8Vx94jpDQ+VHawX9Xu2OUDVIa4AhvPN5AIiWz5jDAM+IUL3T8BvvLlCY
vddCgYv9qHNUw2yYSgQxg9CSA6TOdBlyfrkofB2K3Y8a5U5EwOHsoFIsvHdcW+dTv4wPZHvXrNk3
KJhlB0xYJktvDL2IAadZaLVSduupmOijfHoXoVtdWWZDI0VPkCQcg8QbNUS+ijcTVY9ZJNGgPwYM
7FOtx6JRg8OpKpKI06Dv1mmzkWSiIBxgGXeA/5HNy36uqE5sA6CswxAyJv/5EEHwuraPH4hjYo86
Xo2YXiBwhBUl4TepNaBWRL0QFJPxlPRApg5RJsVSNKccA6s/WXFweiRHy/0WHg4oAAbQl9Ghd7pz
/d34ImIdJ7V+yixH3WF8CJHT4BfeF21GH31eqrmgZzq/3TYuzfuR9+Y01cb4dpHQXigqMpNcEOZZ
wjulLMadipNHu+Llc3nVzTs4wAs8eabpCoD1/2mqcGQqA8NFWCEV7xKIqq/c93jlBF1qDSPNiZ4w
KfhIF3K0HDhjw6/A0DYlHTkOUwxZ25djtu5cEvfy6RsZYnhpTIsgoK8fBE2Muv+x47Ao6NVh5e4w
qnX5Y6WS8t8yO7Ac/B/3uSg5D9pdfE9iNMfC/qlT0sHbTxFXyuTQBmzaBG1gE7EVv8jH7eaVaqIy
TSXcZLDeGHfFmGJ0EmVx9YQcfqP1WsySs6Wb8cLdev5CNXCRPfqU3AYFig2k/FUiwFOTQ7KvpArq
/Zfnx5H0yySYxVPwdrNQD90Q3DAiocsJ3kMvQLOx52AfrLJRDSEehS9PzzKg7mchhRF30mHHW/Ru
g65zC0UpptFfi7BHHs+edy/77GJJA/k1G+b9xY3toleXoyD0pCLyPEhQeuCnkRNF5iAJIkQcnYvl
d7netL3mXThPMem2TY7jwyhRgrNfrcO4u89o8HwbuxN4yxUMpneNw1gFKEUPAvViCW4wkN/xUXpG
fWiz3WrLJNKTE8+Oz1tVVZTBKTKVwxhwvSzzb7tX5J8Q43vvnmN4ee+2ChBv0xrkKZ2jWUa911Xz
vLQpLo8uplmTElBhM4yoMCTAWTGGMfQ07pBDTs/OeeJBVDI42mbIf7PbQKq8tfhYrQSVGZoYjZrH
gNlHXC/EsT+whm61Gpw9+UyhhODugP1X0FwTIeqIqVAxLCYzQcEEFpM+6Y+Tkkr9/I9M/cpiIkDX
1E4BPxIyGAGJgY+QxdIBi9LRnlE9uvF061ra6Sq7FQKuIsX800LC59pDhWi4A/Zq/Q/BYpLrWARt
zuLKiHuPofdjuv+kVy+rhUMfrb/9kYs5Z3UyRH/mBNJXEy000CP/IK4Ey2oLJzwAApztEgoqQ9PU
I5zystYqmAHJIEquidyvS+MMHUfJLGyWIabs3TGQ4/qjlg2EXXkNOFsWv5rpQs0Bu3ayvbQLTQr/
qcyNhXf9MlhC+xnBRfHEAuNRDB72gBb5jn6ui9vAbvmjP11SRNUTcmWHJ1Mg2LKCXp3/WVuXGOCQ
NQLiALpOO5mbqn+SGeiUr19ksGHSX8hYafgUxVDIdx8pK6Spnjt1A2tNKbMqR6YyQyc610Ru17vt
M4vek4PyivfPNcciMRY2N4fsOXv/rh/Jy0CCeIdpK7g8YtLFnX2A4STbi2Ti+EMX5VPjJHXPnBUc
qMn/JKYV+iHbs2FR5vIBr+Xuj/O6Z/pineG6ZJbbyXjwdL5483y6TLXe1YyLOBg9idLbX7/AFc4A
vOa8Mf0/7dhI3OL0hBcX7LLKK27LnK0qY9UdVyXxAFaLaq007fq2gOE9ErwCBZK2kU1IijHrmNX8
HqV/1yUtn7h1OOEGFD+X70ZlvYtH/jL7G5DE3vPViJ9XwmfOgVk5f+9Zz3N/QYBFfIh2EpgaU7sf
tzE4GAbkpbkWTNe9mSrXkNxZE2Z8FBjqSYVIDdtLb6oSqyK+PpkmRI8pzgT0KSc2iO1DQKQKOvng
fHTiy0Oy3e+rAlHABT9ZwI+ox4XHnWmgV55KLOeCcYD1rc5pK88bkV8ZoAo539LwcUgrxjYEwTTC
eW2GbIu+3K866UMh6tyFRs3JrcDm4bDUqN8PSa/uoq/gXqOgkehrOSm8QHzqN6wabtjMI8Bsd2K+
WsKOzthsfM/BvN5pkoy0Q9rOzVgKkhAXsEDuQMksEhxSGi5NepqjzaBycCfxSdHEgfZHLAa0kn1F
d7tnGVynQZ9npuBkJJi79afgEM4x4ufzSYPfaqCjz/ZbPl11q8xX/+dPkosmRCj2kBwC1bcyV51Q
zZbhN9bNKPhgeiArp4wiJwMLtfCUN3aSnggaVJQk+ev/fpjRGibuxybeYX7Nnmw1SmndyIfw5vER
JbBlYsdFZKxwatu/caqiGz2LRFG+kZVtepBnyHu8zDCzx/28U76X/jxaL6VO3WjP1hye3VLcCN+U
+dyZ8Esnu6KK64hiJFViS9mhMMbAJmtUR2/tm8FeL60k32tfWYXWiQ74S9i383810z+sDnXAohyV
ILYq79kZdvp59Lr297xvehfN0RigktoR7rQ2wwlzNUjD3GEHYOl3bVGEXwvRvIqeBYjnnzez3goA
eXpxK1pcO+NeIGdbsRyBz6No73ArsNcKwC/JQ6NyutSHIeOZ2eIm+OssZs7pDvrvz3qz4Lt3FHfm
IdU1rzp0QyxdqSGJMsArCPX1a7Om0drp88/yffBv8NMpL/XfRozHAJo9F6IgM3cadEHCNuhm7ain
K6V/me2nmthV323RcL7kJWdUxPrVSn/+kEEDYedv+iPZWqWSlnRHcQYS1fmWqujkruSbu0iz5xxC
1w9kijY58wpawpFPlSwL8vbNsIaudx7rnG9NHemm0sstg74t1S5fV58usM2AiEztAARqDS/MtpCQ
EIVHCrYCURIJXZl/8MPZVfRnIIIIGlIobiuR5RsnEWXOuih1okBouxEz2ErnlvemE49d1aCqQWoo
UcFhTlXqwFQXjpaS5Pc8RBsuSMf0qnTsBXiXFq+CWrzvDHVlCGwVCMaV5rrqLdVEwI72Q49djHEk
kP15+YpBn59XxGzEtHQFupR2dF5ElIIO2QRXdeRh0VG/ZlRt5SDSPyDMqXJgOJrcY8WkLrpZmPKv
PmrF2zbcZoClmhJX6ycFMAtGD+1o3EVbGhklBfwjQuEp88/DhykCf0EwvBKcumFZHLTZZ0pYeAnb
yenPvsE+fTEn3a+gdvdJ4cnKkr8CmcOMvExQPnvGwoVxhSTC2M4FH+a8lqFd6669qRgvOTM29Xw9
Mxz4Xti5bNxI6xlCa/9OiOOog9CNtX96wRIfp022mYNBoixIe79C18bR/Bm2iYfGKlwpkGAmVQ4l
ZIvx2h9bPgssPbE62xfZJndIvsiUP6/K4mlcB3LMrcV3XUF7UaVWkueOgJaxKSUrAseCqmX8MDO7
eWbRi7uRHKmQM/zaq2whEY8qagcs4SXeHBcq0TN8iYuNIgPF8KVX8QQhoiycbFHT01HdvG6a8C4/
+7KFE+f7pHIZFILQFpW6UxobjSrM1pimwTFx9L5fFAfLAQ7Ih8yAq7UeYw1ZaKe60FPMXyft6yu3
Yo1JKh1P4q7solSL4eoUs7f5xypCKT4AGZBW7hCNvDlg85NyJYUNL/cJ+ujdWcgaE7uZBoR/hHWK
pg/tyrSRvif5GHRQ8KrW9iL8PUtfJZ/kU54Nl/KG81zUNrRqXutXWfXjoK47fyL1ID5emBD2Pt53
LEjzu2eN3djWAs3cdQf40MMpT9+XfVLb6ZMMteMltzdy8Fg1/RBmIykqFDRB+LEBNnd9rzsDQ+cb
bvAv9LDb1Y6x/35Lr/OeKfny/CNfnssplPSLfVUCdbHR7qDATsZUK6haIxqky0E10T/aFuOW5b/T
H0OV4oTk6XLjB4kao268CVSoRQwEuSFxkeOtSEqjV/MaavxY9R4X4Ys2f7klC7PCQHHy8LUVRBm8
m+8naUNqXRjHJmgGvQNCRiIoEo3eW9hN1tqjHBf/b4vdIjQsuna3ZP0x2WP6/IxMVldJ8C43E/Ds
jGwxYeYiJ63G8m+k/QfCoTAQFnwyc4tL2Eg6wL0lK/Mbu5bobjKQLYoHDXUjylxnvIS2nuBf+1aC
T2oTT+78l6OT1P+eQ+otlR3Je1dEsVy1eNDH2vUzBkfBUBekLIxudUXsowuDU1DANhiuthjI2ikS
KFsAsjXuz83pL3ofZv2FN9+Nt2k5pi5KQXUfgwEDVvW5V74LBQhUjXytwYgl6omvFoT+y7vU968A
D9scoGAdRG5G63TzeK1zwnAcNsV4L5R/P8kRDro4uOxWDNs2h8qqtEQjUFiT8rbHs1mq0ul6bqM+
uYLMd4OtT2CREHCT+23OfJvF7M4mCjzYdJBP6YBPVQkHOqERpbiTT7xfPxkTB0Cdj8LesOTAtyDO
+fJW7AoTutm3zqsSugsLEXHCg9dZcVdib6tkCh7aXgLuWRFI/fzkaIHt055+RuLtxCl0k/bkG3xh
JvyPRC6EsD+cfrlAatJz/6bTQ6Yh00zujNBt27WLA1xHRB/h1ICwgeaZYVxFAAWk1vV6U52V98K1
93b/7R+x/Jb6gftyaHoMxwDwO5nbbeCtNU0k07yv/TcxsiPTo8wz8aXWFnJ4B+9GehLxn3rkhO1h
DeebAjRKcexgCJXnyK8+D3pbXSUiZPmlIbZJdCfLQZwOifRECoGWoI/CVdTWDmnt/MTHU/nC4P6S
2E1/uXo3PRsnXOCkMNsibF91zt9BN5rQCnlQALYRtSkeQGT5NeKgnI0OojuYx31YDaiq7iYyhl0j
SmNeY4uPy5wA+uhH8jNSUhrKh6mvjgLGIEU/1aJivYBvvSUbCzDFz/PsI1X3srPB0LHrWUxRbg7j
Lvj63KlsZHmG5Pr9qHwyM82/vBWfJXQDFsSS4Qp/iXWwSze+d5x8qREwt6hOB3IFOqibhmdXvACw
FMsgeLJTZiQZvMSPPd94AU+RZqpcod9b3+eah4m+Uo+RSixY0a5zjp1+DmeZ+LChbCurtO8r31Zf
IkjW0Ock4XbZHRxEhj8n+V1QmhNAlc7BKV01Xklf7YHXucVI+Uuh5AjBIm8pIxog91WFKVpA4sHL
ONxHEYuEzwJBfYKiTyIESssDLXaohmDaHYNdVnOapPuLxmfsuqbB/EceOpQwbHVOTcyf16Qaj5/O
Sfbg3/Yyxv65TUYEwIRCYUyoP/h0ndhMRbUV59/p/30E0iBW77NN/h+uk4x7zQYLQCDHKInUeEwQ
KOeSGTuul4rNr9JqXFXytdHr2Ta1ptr1UJrYWToXZvTYEn2IXvkA/SGPp6vDjjXb4mP0xsJSXORi
kBkUlZL20NG9x6PRGQS7dlsZZjQKdY+9ETIkLf1BqxjpW0lIxS6VGJgEFFDjvD7o8Hj0A6kPeyAX
UnTFcHaJF0AJZXadULSdfb5V4FKrzAQ/npy8Cy3XNIAtdJvdmNmdP1b5xf7M3bqT5WkVgbUQZv8t
nv0O2OaFPhpGZLJoveNsViGlNVl7w+0N6hJDRANELRo6K5EHVEcyq6NsHInoHwGZ7cp9YubATF69
m7+lTjLz7GM+O4ZUTLpEfcbybGqYScdpEI0D+9Kf0XSt/DGMfjLC1M8Vh1kK7Bu7jy2bsVBzbW+R
YkQRDnvqRfiYVabWhM3Xc9NtBnFcn16ZUTPejD7i6Ro38pxIH1f0ChpZq9ixDhyWi3WsGa1JshcB
ab93TCNo/Fo95nTCIQleoDuva5WfyIFOzcek1rZdJXaL6bemzxN/5FOGz0V/bVF49WeDAdR8Kr0p
BByvGKOegdlpAsvuzjxD7JFLAI/m+vMDOAh3V/+J5ouIZZS4+TuMbLVwG2mUps1+S1YXfc18kmOl
ygWrnXkK/pyc2xXCs0ELvBZyPStP2vcc832/w4FmM2RSGWvxhcC7C117dsM1zqZ8VGoOskKQcs2w
cN2Bkl2nTjY6el4bMGTls9oCJDGp8+2DpJDvj/OwMloxNESKgLeZvO2lix2/i20DEVIxjKW2lAIW
n4Dz8gWCsmnlEbCJshjIwGIWk27EqzfBtcPmJGYNdDCuvRItuJB4RKNwknjWLwoBTR8KvhuZPipm
iVpY5gWt2h0N841/U61NTbhP/L+rZREuhzhzHMD89m4GbS4AVmnkIyCWoz5YAO+IGwd9wX4suWzv
6hvhrbB9eyDi3EXxQDFoIVQYJ+fnPCXKQDpbGYjs+buem1mxuIhyjuJtIvAQONJMNPlbEhZbX5+L
FBDxFO/TDqtzZFlzFXHuBV+jL62Oi52QWUpSZU8Ni2hbF96eI8X8l/tyLRdS4rOgZzKDpGU1hkgt
x5kBK7XULhVKlG50KWwNbjBEPe02fv6SBvjQwyitukBFD6YA71OskqoGyLcmXjmEW5z2Ld2AAfwQ
Oo6iP3Xchj6vcx9VFbxBbA5jL74+oOF5LLBeD/3YbNpaFann0G8ka9yqPLG5ItZ0Gnmu4ffjYpPN
Juyn7vi5E70PMZ8SStKVrlZjd5hdt+D0REkJ+fZYYIEaDGSEqNEk5X6TJTzyuKbIgZwebcDyB3pf
S2Zo7o6bfzOrkEmOAHAY1c0eazFh45aSEo1FXAgnaRhUeOOliVwNvFWbIpWZMmYf/gQUnOvpMmW8
NU3ZJN6tZ2puU20XQ9/gpKEwLPYvIJ03QxJ79/ah3WbwvjFZg9QyyHBMYtT0F1ITSEMB3U0DW3pg
Lc1PVBYBDYg7C5HKrSchF9tdwqHoj5dh3471WTIsas72Dp2ESOtM2M2+wVdYXfLiHAchb5+pjA8t
dzUVeiLtfeh2rJRqCygIlyo3XlirRwucL+vNTXOnJ2iAgVU1GFclSQ3bXJZV6jpzycyBtfOq760V
7dZeA8FTcyZr9RmZFaJRsYYLz64EuZj/c9HEulw4wVIvXWjEycrIVYkwMK2mDqR+VqG58/wYqVHX
h+FDtZRia7jmXEnRVSDtQrLGlAQvqowtCqy7s/FY4ktSpjgP61qYzRE2bPkboVvsCVeAXYHThYfG
wGpJX97RCblsqQMvwuexHjfDIVerSYo/dXJuOFW9PJgQgYrbQvyHN1eBhCyl2x7//mkBWJM4fgcC
DIHOK21/No7wmkrj7tp62XYPkWYkMcxPsDNQUw4tBCeOLO8f6FKND9m/jNY7/pjC/Jo8rADRn4YC
ifBmtbcrMKerX5FtBs1oDTz9FNJhqnNXPjWk08WR5ZmZ+zvLknSfaPOsC/5Bw5voY56OPESVCVNy
ItU1GDF1sDoovf9oxE/6pOFNyu8erhQd5QnHPp0uF5SsEcfj2X8dvMJiwGjxfTiEwfoTyjVCfwYb
oe6IU30Ue2DIMhLJ5A4ScAUQZVPTl8O1EpjmHLV19lLZB8SzW53Om6ERUjwHol24YhN8AkoJit74
8itidA+vj/68JSk9pv0jan8ItGTzYqlp+wTLkTBgumgjEN5tOevRX2GT8hH7t0pLt4+Dlv2rp8qS
PSS3uLukDSrTvbNVOIera3rYKTO+KHPw2pEVklcs3+vZ47M5kA0GFe5UZnQFPw4IJ81mFDwwrIZy
8AZaiUd2/tDvC6ry3wTyRhXSd2eLR51pdGUYZue2VJdq51et9HiqbIcsaWJcaWHcESyUSOKXb6jd
rRz8zx4NyUIA++z9b1ox98jrmK13H2+PaItplkW58HFDWr98Q3a8fow0hvmZ6rn8uB2KVBJ9vDoR
CPgIkV2c2c93/R2irTtzmGdxLjffc9iBVYzAyvH8jjuB4/RK4D3+7wwSPQ/I17mQgNRBWtFda97B
ZWN+HWUik9lHzUtuRBcNi+6CMZnszOxvuNjMd3+uzfqocvK5NQh2T8IdlhJDIEILqQIbQwXrNe9N
FIs0qrJQaqXGlqxAJ+ePtThvbO4gEknYsnVoLggNubKsfFjSk7jKLeQnZor/E1fbz6E4iwkGIbe/
r3aOAF7vcNBKTJl94Re10mfJMPk12zb7tZcQVXcdSpCDz5TwPgIt5T/NtgKSipRCtg4wHekkwF5x
P0sQYGNb1mw+86KNqoP9tC3gh6GuPg/pePJ9ox9EYm275lGOZbk8GXi3GQB1HpREqr8pSM1q3OtD
pHFq5cDLxgb3U5OcEAHqT4ULq4oDyRFa6w6OnHA4igowrhh2LARx0ndhmHTEEC4mTn8sGoON1ims
tenwwlB2+kb0vkBF/GeoYoRay9pG3rpkOEQaUq0iY4Vs4y38YW+GgdI2P2ilaaeZmaloI1pgkUeq
tOpWNXukmGbE28q441aqnbIyHRkWCU6T2cRwpQOoW1dvAx6TTAktr8xpl5SV84lKk0SoA8LLna1b
/pGLJHZVdLo8TsMqxYsw2ingHFSWRxnmtnpIfD7LVCaB21m1H2ebCQVqZgB7i1vro4B/WUwbmAwj
3gBC8ho1PrTlb7ac6eCk0W4oZoxmjz1XvSB0Tb1iGZcliHWfx/jLYUyiACWgWVg7LPe6FGnf1lFx
pNZrO9n7s3VdU3/H/+ZMjwtxF8cwzsNhvb23pID6Npccm+Aub+8OHzKljIha0On4nrI4hGkH0P7m
Cr5vphOYr5olg/BrvP71NtFXlGl/aT4EDGPSq+rhQXHH09CkA34f43gh3cj2xMKTbf6xzqlxRk3Y
efHJo2zKcFLaZZ3arIC+bIwdaVdb1Z++rP/9UBxOzDJIkIgVkC97rFC9+hEwlNRMzaxs70LYgIv3
bTuBMB+1dmYStHj1RCvQ8VOq6acUvfTOxoKESn3QGcOcDf1l3mS+9XMPKqHe9HR9hPBSswyBIhjh
6BeyBKs4TEyA5IqVenFeZqkE5KoLVigQDkSF++bxHJw67+OiBNGPk2MXzG1RIYLYbfDvbWP50DvT
H/JKKOZOBF5KKIaVu3RQeFgI/Jh/VIrBwUrsQEKBuaXbLhL1zCxH/ES6aVCbM9vGCiGV/3F+RclK
nfznRbdq/samXkWhv944xh2YhSRNBcXC2OaZLC3x+W/TQBmcF9dh3Yg9z4kaNw0XkSUJ3pTr8+bb
NBK3LYX7Q29G7ddExA/YmKSXKODimZ8nu+gcQ8U7GP5kP0LtyiqHshKFeBKlKH/86s4/JosKcgOn
CQsy5Hh0B1BoCnlqWi6gE+nvZlGBmNQ5K7YQ2jOv0NPVV6Ip54VQySzhB5YJnRkS2LwW+3JVROhh
hJe/EAlWEeBOUxu6pffY0tGt+Ny88u9UYPSnbiuFwZB9JMbIudye8xso3nKr9Vu02NSEEnRr1qNr
tFlG+AxQkrS+1MYE0D13vrPL1qVEnCzlXaFUxCNNqQh1T7NcVOgddI1UDH7DlbbYBEo4xMxYBAnL
565MfysnAwmXDASzqaSPiegvpNHC+c2vqvV3PkmVukBdf0OP/mESZ3HeFRo5IpmzAkqeEIg3BvYd
KZKtAEeFC+8EAjknS14oj0af5GisucjBAJXk3mow50oL91iBgtrTmXoLGz8TvVEjLwqwpYJEigYq
BpF4KYlG8NYjF340hS6OOXlLc85PWnhr2H7vfY5lMAA8tmhXyH+us9kP7XT3Dt49ZvQ294TYXMj2
YROPdam0J+b0H6kd8XmtKDkbijRHUB6u0JoCqi5Rf5Ui6f8Ok26DCye/S8HSMrn/Znd+w/YCw78S
tpbJ2SwEv1Kk33egn/cjH3uHk4iQIgOPjwwpLfZucM2nSbIGh0Wx6sLbXd2AH1R6FxV33I3GbGyC
xFk8Q1m6kniEjwnBoMZZY61E/B24e/407YYk3W9Wz+Bui20yuOf1bFK1TuVobOFqFY7TswD42YZI
posjb9AkFz9kohx3KDTgjKC7FTuRG+xDXsLRY9+ZQ54+U+xVzvpwka0p2RVXP/U/9u2s0NtVVV1j
nwk5M9fQJwotRVxn0OcC/AoVAaSkoIB93OtLYhi0JWcyDdLlbwLMsbyG4HSW1x+uU0cNMifkaHXJ
rRa8dY8mlG7k4mOcmI7RMtlax8n/dyA/rY2PozJZYUDQFTgGsSd2orr6cynYv6COcRZiffN0D6y2
hnqjxp3Z+x4zdqZMdsQZRBblDhpAOTJK3H/xZRMHk9heMYPirT+ZeTP6Bbcd9rf3F8hqINb0qajx
oweQDGiH24wpcUrCrADAGtqZbZmvxenulY5ZIneUuh6sqQUd+dhU99j4GSnmaafI+Qr+wKcExdvX
hone+S1M7M8Gz5NNb7OascwH+6LZaIgZpHEUHW8WYrbPjg67TorIcAw8TlfU2cP3n6Lw85hSy26s
qVigadtLO1h6U0VN5iM9i3Elgt09PvRFCjGmidMM2MH7DPP2Yjd/UuH4zA/kQCb1QKV6mqOL/LZr
EwrIhZj2QGl2huOa8G+4j8OlNEC45XiA65cHptQv7J8aDKMs5Km+uffIZEoFcyej/gGGTv9YiCsM
v6IRkK7JN5vyY8WODQG21jRnHxNfj8kELmcuz8DbrAqQbzja0Ml3Q1LxdkL5y9grYyn000c20NHU
YmWCrVc2yejPIiIFhNzrtwGr/2t3GTPljDAprBqJua9UHwYHQxwalYB7spwTZb2Bh31uRsFn7EU7
DD3I9AvvmXBjLOYzHBHLNmWzfT2/80vlbYfVSqiHBicFr5zKkpfWz1vz8D0gLcnByRmvqxR8bPeh
sKMaujogffd6oAqM5wYnvYqep1U9MoX/qTlvdh6ppsdfFGqGFiyJWjM3FPUT2du8gIOKnkRSjbir
oAEvHppXFBW7IaKFNV6Js+1wF1uAsIbmoBkxFpm7A7GZOdQFGf4i1TNCvna35x9FRyYSJeT6+/rH
S/ovTEXQWrhQDAcGe/7rKhl7LqXT72lkPJuyolgoTU4zLpK+Kovqws8jrl7KSXJWJpR3Ezdk8Wyq
urHJe8S+rlI4FMLFW9sDleWjBTrz7FZAEAOwBUtA+iSGxEqBB1y1yALZRIrWqySPusG1y16uJx2S
rHW6r2eZ7EIEHMu1BB2tcPOWEueYvYleVYYePwFKPXik6rH18oO4XSF6hIuREdNZ99xJgFRXxsa2
7IASfoUrdqXlT/g50wqc1cCOkqrreffx93nvUgoe9UF564w/wCR04BqnC84MMhLnVnigMwfIqaTo
7xaPmmTNxY8I1rUI8bY2RzWui3f5TKCaDCqniwtNfC8/5pZQJTR6PjHQ2dipim4qVwHSaa4stGsD
4JbdVRlxqK/JsUvkes4rhNfts/hYZrK9YNIMHtwZR0cuH9Em1gL2pQwQTCTV7hsVwN/KO1uzxb92
TnBoRb8mn0k5IJ0xqo0IbZhcm5N3dBji++SornH64nbWQ6YrkfZ9yu7KDGhlNomc6aEDprTtPmEb
4EeTA9cU0kFRNbCjTNLzmF5dI6Yhx5PwYzCPhWnKWFcCeopc6PsnbqbL9yp87JMGMNE0vBX3iNtx
y6zBJ+p5RKt4ykCkjCZmj/wNEYUBLyRNAwGcRHmDxI2cQZip8GTfIUO0VVw+i88L5Pn0I0GR/tnv
7qjccxzmmhCAO2/E5T3wVuxG3geg8DYtlht80iu+kFafakpR5r6aOWxRIrsZF/VMZGs2XIQCmyNO
2uczG3iIgsWHoJy88r4qDetq310TfEke281QEMwdJUZXSkk6zI0oHEJDMfuOuYMOtcCFPowJzdqd
iV17rtscFOmq6E1WSLWgSKribgZqctyYY8GaMLLfckJLafyurc6u0YEokcKGTza9QrRA09m6akdj
3KHvg9KuN32WKuaHq8TjfsF03anyjHpTiGtrNuQ9JUuxEEzzHNDnKnMTzw+0NKg8kh60838iLaw3
TISYL3CZz+jIcl+WQb2BrtaNb/6EeciItJyIL8yxnJuQtzwlBlzazCVxyi2woEHIZbe8Aw7snO+Q
Ui3OwhQ4GkIDwL//zR0rBu9a7jQdLzzVNObsXNDx8C5WbCG4zSnrXsJADALcKwNw+B+a4cfVOmO2
R1bPRHr2g4JBdAasmhonu24HPdcboGtwA+HSY6Vp1Vcbrsw7xHSqpRnJ5LD3t5BTzGK9KtvsxgdH
0xg3az5HctLTxG6h1RSLXI0x1OLsvMQBGMNYHaeCHHcoX7/2tF4uilH+IR1/vMspsg/AcxC5ykyP
/MgCGClSSFHpEasDFNPu5NDIK8mfPFnv9kk4kalvt6tPJTQYtkk3U0RpOaXcIfCrG3DEpqSZEwMG
TxCTLlbHqPwKD1VTgcAflgeVSt/rpXWl5SnwAKTuXojbckUojb8oR3vGnnCK86jDCWj2B4qmCe9J
4kpozD7GmNpv/D7xe8nCd7id3oD1sKg4mGusBj8IZ4drpoJKoVxzTGnSPtPcmByA4xxpQz9Co0vu
K/l7spH0j7VbVOfE7dcnUHIM7Ds3+C1wjreQFz31HtJSvBVUV0XaA+eSeWtr0ytMh6zkyat4o+Hr
ll5riC2cOEfQOBpMu2r+6KZ08w6lfz9kzQRBRHHYNd3bkXMxofotYEsG3KFRlkdMHIJzBrA3FgIk
q2vu0vlhy8nhGfBtt+M62CWBdmfya1oNta6SUBmPBKaivmL5NHIR33T4YzCQSe/lGnSgjMVJ9FzV
DMnsAxb4HsBjcFdZU7QRJr8eRdJFOh8ow6kAVBFNwz4kJ82h1m0aXGeS7OoysB0/95dJ1EEYk0Je
tKzxnPJgVDu5iKZiVsLHuCMUPhYv6I7JDxHC9FUS+uNycUv4Lcs2E+le6ju0bUPgitdDwrX+kI5F
bWE49/DMJomQzw2akJhLtomMOQNpJxp2WT8Twb1dfH6/55tdxJ+7vnoSVSvIIWSQnmYxEdRNuPBE
kcLROZv6I/UGzyjOfwKP0IRgrhIRX4X9xAnfVfYpbqnTj2GfmdKmQk3kJRRujqkweot+Vs/J00DQ
DOuRM2WNME6+HtTMmlUe2B6i4Vx9xmqBnNj5X0NecNaVQzwQv17G8baS8bZWW2QHOOVIUK/i7c3B
/FBGluO04YhO8twqNAIh/8tnCvQgOsXrRrQcff2d1Ma2hxGIkEcLHwMt2nDd3oj38zKbG/dQCEIr
eOutRsVLZ5XG8QzyJcCJMIZlGdW81x9JIo2UfEHcQ7vhL3eg6scGjXi4JE+mcSs6/fmR8xTQDS6e
8bMov3tlLX2LzBiezK1H0W7L/WKCX575yQ7R1lRUrnG+b35frpMJ3sqKMdrciOFU/fJJZRLIh90L
0s/Mt9AV3O/m8VSIcqqm7ASKv4SvcsG7DehGUtp+fodo3n9N3lg7Bzdec5yuqKcClyE6uF1eyhMD
Zglc3MZ6qupUsEZutEjZ9SewUYen5Buv0H/thDGFilyXci/x+2fWXVRHTx+qLN1rS/44UIBeby6E
stUlGI1vD6qIetnEjLT3xioxyJGpcjFsXaK3wCu3SJM0DQ3ze59LkgDPP6MATV5eqpWxHTc4yMol
Mkj5ag2NDZ3eVuSap47cuuT0W+8/ps/J4WxjERFM91f+AFYzEYWsmbytvjIFatTxxLFRyMqQHYRO
cjm0xKybF7hOsOLr06saqHfWXa3cdtHl/N1ipFJp6W7pVwUONhrMx88ZEjiGDB57cvJmqs8MnvUh
GzEeCCe7Mrzd6Z0G6ZJ6kcEoruRgj+A82hKSgHwiUn0ogPUouB9DMWoQZWBJJROGHcMKzKKHSVfR
2WOQWWxINOmctOir3XadK0Ez1PG7y6f4df/w8daEk9UMb+1cUAAOf/WnjIRrfGwTOhbmGnpHf0Eb
wo9wRMi6rLSx58SCYl8Qgpab43gCC5KU7krZkNCqsFKljjrjGdaGsH34PUxTN6uD4K+gGnnnvRIs
tkeCvr+qWbzGmeZVWxPq2kFtJLF7a51LgWMoBbqdhAg1WdvFdOKWTP786bUlktiGdtPrcNTf3jlr
r5wTI8U+3Vz0JvHXCKzjQe/yYdLUKsQ0g9XFiyPSAfrUHb7LibmdG0LUBx8bAwP3oH7Q86XUWijw
zppM7sLFQN7A3T0TwDWgHzB+GPdr3TWWn1Cqa5rAPLzoKgj71i6npRT9wJ1GVOpbuW1ZWcxIVstM
MyyzKJy26ptAtC/+xWfLAeH0YsD/YbYa36FwNKLgFVyLjh+72RB1YvevE/ObRvPOT0TB+ZZsfF78
7kG4bZApwPk50l/5G49ZadbFqtmnjk3/K6nCLOLlRZyuK/208KoomTDREDNVRE8pDm+in3ENI2ES
E3gqKLvJZKc5c9dCs1thC4IXDcHmjxOtBJH5E5fYM7fEPudxIbgzfBbxbjlBrY65NxZAnAjjs2gG
bi85gb7lRm8R8mSOq/55GNrISVeE2il2J9whFCnhOLg0vtzmQlQYLxs55+CzQIpPukAi51jtxqES
zZKQtc9yFIiECiQUNUeNIE9EC04LKqPMlXrUPoojVHdwq+Lwvic63wSwexh1R+P8bZPmZgiFfo3t
HPQaVnDEnpa3S8H8NCV+FT7WyKjbYgv1bQPR2KK/9RVViXeXqZooRlq53fLKpJTwJTjHg3HZqIDi
N7d2+/TpyPOvBUvw/CkAa4V1ODsIj5Y8AnqtQ/4J4m17iYim5Bp884LtwAs1vwkoGm5RPTgX1XC5
yzRxa3ysBhj5R7X0rlGmdPSk6IM+ByH9LQEIUTJXxXyq9Y3aGbHwWckOtz5RkCGajyvOEZt04uVz
F/2fEadDoLs33EyGrl9+xXcjZR9tKxKeB2c+l/2dyxSVIc7FC62cxiDXPB1L1PXlw7HsPDq9nNj9
SnuYgAks4Vh+PlySF0jNaUgKdu1omWLo3fHCw4zVwrO0IUbfRXVft+X61bPEP1H4TshYloyLFngD
Uypm639vK70CPSLMmwHxWmV7T1CcUglcKmqmeex4AkP4jmZiI6GrEaY9VSNjoX760Hgs8tnoP5rT
SnjtFnzTF3Te1Zth6uCadP31wHoUsz74yoMeNdfEGlUhI2VJsqhu0qArXCORl0V0HmA6RjYE7HOc
97kUkjj5BI5RivzOJd5D1+jMz7FIskVgVhV5fWiDzVH7hg9YXUr8pjFtM0nEWlCkn4u/06Yf+xvJ
TqJtm0bItLv5zhZT31wh4BhPUNT4Qi3tJ7oIno0hYgJI0WSexvb6R/J81ZFa1rpMlDTM/aMDut8F
D2Ai8QBg4pmpcJ552KQsBUNl/FdEx02wiDZFZnRFaXUkw31jPaVcv6EQbRkFGIMhTwURwgbVKJyz
WZ67DKwh/K0o13/BJzb+koYGBsSD/IQHjw4hhbeMuz0L9qUbBACHvxO8riDy/YKOqwUZkRudwZAM
7Gref/JtsEPKkchG+db3Asn2Z2vKT+Z/PrmOfQcUNjOHbMh4gExYOGe3rcJfO8YzVbATHnXDcVeH
FPdGk7QGIYA8PPXqPcZkF3i++nvpRq6VsRpW66vn5pqJYraVotQziI6iuqWTxC4ta2foNC5ZFMLp
F1SvDq/nD3Z6R/EYuuS+vH+d/cwipnoEMpc0Y863lYERmoNRRcoY5YwVWHjJxx3MKwhjmw+2CHig
Fo9y9NiHXZpi+O73cxMqTMvTpTXlt3zZRUj+7JKj+64ym3kpsJsLT/baquQHPaZnHErRQ/iGQaz6
eJQiGo06JpKnsOBicXWAnC1kUmQ3iDjoB/Hgx5TdXQZPd+cy/p2fc47XKDv2uoC3IRRniJHQZGEt
jXUQzsToeg46WXYqd12MITRDTy3NbVOVnUiYwFOrQYDL4ZE7m5US3KKtjoUeOjwepFUsdUTjkLMJ
fy+WvPCzazNjWON8u+UXXb5nUFKea+w+69Yy/3FUcb4WpNvm3ef6IGrmwG+GNkbzeQd5QnMCzR8i
7/ucrxqvAJKiaX4L+kQFGjuAVTfnQAKw9entBDRYaqVC5lnQI0+xyGo3AGpTIrvRj+daOc03t7Dq
At+a3+BHKE90vtGc5dIDrLElRsmI7Ltrfgcz44d3YRnadarEEeJXLD1WXdMQ3jKdW360XVzXrWbE
sIWZC2R/PtsKCh1N5iWU6rJjmfrdsquFKbMjPLDrH2IHkN5ePj9PAv3qmd/4TwBYl+LTff6rGLRw
C7tjPF3Fwceng/XdfaImpwV2kFUuG1IFxK4IVCU2XCOkfX7g1iWMeM0GjZLyf5I3BPv4Y+XPYR5d
sYSSfaPOLi3bjz4b1BLHWfDmARJh3e/wGyGwyFhp2/eEiWICk//PG3+nZAS9vRWmhzerKgcOwt1d
K2aR+Z6T/k/8+sccy3UCWIe3e7zGt+rVyIuhTxm84n2O7+ppJw82qn/ZNHRLeywyfypu8AL/ejYJ
xEyQnakaGE0TL4Is1twnfqzYC7tBhWlKOgtT0uXCNk5f0fUBFHNxI0a6A1f3qw0euUZlfWsQ1fH7
Xse2ofD4QlkxzliKSc7+VjgU/kqtbNs1FAWRkZGarf6MC5Uj3Tn0CNDfxoY1TXuou0Wq3xwHQbB2
D/aD+sV879HveVRbo4cyrGeRrB48g6EAlybehpI/pinfNcp7z83kEoAYT5jJ2KBJbLGgMyOwuu49
jOgRgmguZrDIwo0R3OXlrx5L0g0D2uWllAIa+uaCBMbrBNvuxS+ZKhZk2elymyItHdJiiD3iNLc6
3liX3m9uSIV9KzBz2lzoVW5FFWC5vPm78hfk6a6szwNJBaSZCHmXvBsE9/eGdTEIoOhzWwCIdmzY
7YFWQiTbCE/t7lj0Mrm7Prvho6wG3aQ7K65LX+mFG2gbu6JzwWqXO+JQk6OEu8b5X1+9caMNlzXX
uBWzGRQN80Lh6S2qdsJr+2uMtbu5lgnPPVaeuRTxR3TlzFYzf6ZNqSc5eRmBkq3Z8TW+mphQK3Az
Q1Y+bDQWQdTAVp2JbqA4oYhrHVNHR7K/+cRFnjD28cL2oaePBZ0wuw0eaDrx5hcm7T9Wa6LYeI3E
/gWUa11TP4n6bPWUjFmFZqWkQ016iw9OZAgb7hWCIg+AcRt1Dtlp6WRakxpgr7gxG2mRrDuDb4qU
52zuuZFlqRKTk9so3V2C629XjUHbLufbO/TuWpC9qO2hhSUWPfbeCkwiIUHEGda9nduDuqWxj1dT
9SuFRwWbXNqAFirqBZ2m/iJ+MFo3G5ZcN1LtiIau8vtwlM8Kt2+7WMeuL0cFJk9W1WHlvacAXY70
qwcAyjMHvqsqJLMatWDykQ+uZf7bofk5pilvo6Q1ohUmrBu5cnLNSfbdNLMYVCjar/NS+5QlO+24
aS7BEDeVYDY2NeWQqGeztzMQedqK2H+p03A+14yYs0PVQ+gKFE0zrCO0EWo9ei9NFmJL/+sUy2hc
PVEuQHgkDigxfGyNCRqmEwvDp8eO8Nd5O7ST5JXhcevrZlGIUT337MQu9f/Tcq2yXwc3oGreG68Y
l8w7qVuul+gB+HawlDPtB6SqM2x4Y94xmgpYsU/+EINBgvnNlT1pKQyxQ45V1WFi+Q1SnXSqm5k0
rEH3fbIM+2D49DhpkozZUW5snTLO6Vz9Oc5eQfrqDQXdePoe2Cq6WLaNGSz8HHLwiSkxaaEvplRO
TNfs+h09yfLhlh8onubd11tWIwRI5C093jF+0ra93rG8JnrjLsMHEdkFKcjGQkXJW4v01DghX42X
GPQr7yi23rGS4s/jIcp/1DBZqv6r1ZhcNzaYYl9yTBS2Qw/SMJ6NFtr/iEL6ZE+PKjCmORSsRbm+
5pSKvTDPMiRXypRBAthpEFp/8CkuAMRCzAALlXsfBrg1hYA55u5MU/RWkpGTbo7o9gUeVZ8b1wH/
vTT6Lm2/zr0ZgRXsciW6eKZHZJZGG19qMnd8Ux/YpijHMr28lcwEJQc6SlH7eoTxrK5fYQUfWutO
hlFcPkaT4wUnP4ymkBP/IoHtqIlb0jldrOCN5OTB6Of1ZmOF8NvXgwsV46jqSfJExvq0OV3vybtw
owODA1Rk78xeQ/2aaNvlSrILwbYcFNvocFA4uRlpUIT0CMoxZj7zHgE1qUHu6KRM4RVyStnQdH5a
9InFjuy7PGOJjlspbdNASRiFlGyb3gzPxweEgiiyN31OhR5hVoBEBq+kKB118RMoiEJ25U69Z5dN
8WW2yB7+q5Xaz8Ls0IXHCp1WzMMjs1s3WI439LxYci47JXZJ86bdAelDbO7r26dYTuPepfV/zCLN
qhv9/3tPI+j205J75Qg3ddnLLfiTcaQGcgseds7Lr8d1mcev610sr0D04Wb2Fr7Lrr+/CohLHSyS
NLbWGj6LqcSU8MFt2ZfocmkKaShqMbM8zKFIV7odHcAY8f0koLgOCJLYt+vJ/cElfpxQ2m7dEFAt
PrHM9KMY3ozfc/i6c0ZO4BnCJMx5A/OkWkZnt/A3uUezF2b+yMakTNij+1cNIILxhKAYZ1GvUn/d
pY7DgDwSpyljOUvT0YgVLzS04ofV+V1+n0f8XSUrR0IkbXZbMCDFaOVuWF7Cpa+05ucrBiwZWYCH
48Ey3TeMpzEPjGaCVi0rS9kMAnCtsdqD+ZfiHCIRQVfVRTWHYz4pmwKgF15n1i3fMs+VX0flbD8x
KrZ0oXssKantBr1hg6pcClBggn7UG7JJUdoAYBtXJT4XSQ9HtFiVV4nLcoYURyF3adwq4P+ZfgR8
JEb5XpqXN0D5k9CsKVsrxvlv0R9GzYjvppR8ICrEiQ05c6xPi9A9T53dvvD/vKzsOif4Bms5Tn/T
2zDpxNjrpKVBeFoBgkyutdkdFB7m01erZTFw0iky8LdF78eQD83gSkZth7zbS0dx5E2ja51ToiHU
9wCK4dqyerHGLh0eaIec5HfIABwrMsa8Xb7RA6PzS0mx5hQkEl3D+Zt/K8K9TKTfKmOpfl6TAocd
XIeh2sjt4RiztuMb1EzhzIPjlORQaqS1un7YVMMcHHaJrd78LtLX3QDSs1Dro4iU7VAS1l3rdbHQ
9WGWE2UytehbacFWF5gKvWx3IWOO95dGwNRlzwNHzh/1Quml4VNjDPFdcFnnqGz8nD0qT1CK1oKM
tN57llGyv4/ovFdSLVnwqSweJEdSNnnqYZNkGGs8RwpBeEwYVPDMAvo5zEGhV0wR+Gz+wo8BpsdG
7SnkUIed8SrcsN0yVGYj+Mmfqjj2emDqxkOkNxv2YuG8xsgxy4fgqAGoEYhZZ7bwUkjGbP7FLGqm
pa5BAHXYrvr9EH1y532KmJc5L1Vc8f8t87koW6OLwai09NIoMnsOYslzZ6yZVRIoIlYJI2bbd5Y5
y+6jtw7z+A1gayR+0aJ72LTBLSTjGRi5kBdqnubpvkQ0e+I2LzBuzUgYUaj5roEgZ7yHNatDkmlJ
M/h2Cb+74cuMjNNHRLKFwrdwonpSVOhbspW463mgou/jqr8br2NuvDvf9hJlIjP4tKYb9GyhEoTp
iTsGPsCuy0JNnOIPA/4FijFhXabeS26t/wDmX1igC75xBqlEKoOPa1K+X13iAnRb2qnZ0LJ8254v
RdMf4N6WDGGjCy7nxdZPEfw/qeZp/Jl1XHB7xZigZHUjiffOo5oURkYGN4hXPw0jOkv68PqNBIGd
lnKZtD/ITqyFH1wA5yY0ojeBfLRIfbKoC9Qb8pH8SeU3vnUlfyZxBllodZhvvWBpx8IcD9+dm30J
I1vx8k/djaD7sTL5kOJO6RRdhA9pLbu1exCuaFaN0n82OiXOPKeH7Nq+xDom1syhyR8exvBBIPMi
0pdfYuVr1adFK7K3K9419kUzZ/0kXM26U0ekL8GSi24tfsLbyXEYydobpIQvXDIPNyqtjnjfqVAU
+o2MWI840Vv4uxhIv7Vp3K+vTDahTV2MCy0mU8Hi8ofSUXlwhEWKwGe5wVr7KbBlaISzCktOKDuT
qsXHyDQ+ljYVPx4xOk/Qdct6rg/YcLJZKoQk7U3NpiEgpQbz6dILfa2iT/cs2d3QsNe9Cmwem1rc
beA40qT+DjR2iXfm9bmOlhw0KpMUE9zgChgjueDWqDft2KRdZEQnw4FJ5XouG6E1RIuDHhI8P07E
WOhjN+0Mn/oAWsvAsBsxW92GSLEQLRvUm2FPtCR1QI+cnKFAQ3w84HlFwUP+OnqZtoQ9PJCoWdUk
hZ3Bx9BxC9wx4DfpcNMhAKE9UCgIdUrjyy5LIRVwYMxcO2ejROKANKNVoHqraBLgQttaP1tKzJEF
WQo1gsleQpCymDxbfDYCIvaORxaYoixsig+M4mBgdpkLK7CTTTv1whVHQtZcRLt00pl1MjW+rP86
c7jyOwLJkzSNyoaGhd6OZeN+LS9xMVyODL5q3xmAdsESC13iakVtkik1ZTbOR8sceQ842b8A00YW
Dx9u+esojZiYsCfCbR2MCb7Uc+g0aeI4d7ZjrDmc185OUyMY9fhkQoKxhHFM7KUYV/FZ++wI/nsx
5g0yxIukUKAKpjCkm0/k5vgbQBZy6nxe5vfp0WzeZWflt27ZWkB8H/MuO3kzWhz9JNP7gyvcSq5i
fxo0gSA9eY6m22xZQ/z9joErmRWkrGqnTcLkI6t+veX0BCmDCJiAvaj58cjsAbGVc9Bo0B5Mm/kr
DRIxbYQr5+Pjdb+JEdC8u5f+pav6WJY0cvBZLLLJeO8lLNmVwRQFU+nkWZTpvFornTLVSeA8L1wl
WP8vDT6OcCCf4Roc8NcoqsWjTBSsoWonxgR1hFO4K6Fiiu+k2qVDv5SfRZKUXOlfbQUVl78/W58r
klha+T/e/1TU7qum3r7StiQEiQv8Ldi9rcEnBaB/kMiauLEYC42xX8j19sC6Sw0H6Wk2VleLaBeu
IR8sM9d3eyGa77rcx3AjuRTrVjDFIwGcL4+fAYnpuVbuzI+VlHlYKV+exJLqIwITXA+7BekJILK8
yqMcdqpoY7A1aF2QNFvxYg75lA2AV+SWD9KwnDtCGEg22+xYSz+gKXvPqnUXFut4+UlMWTUvr5p8
uTwqtI0IZ/XlaaVpgPQ0W4OJGymYMLXoYHkKWxuwkyF3iYE7d4rRnTaqPy9U40DsWPTJVFwiv7nw
Bd9H02EKsQmvZYSlfhAegPRm2rzOWnd8suCgUUZ5hcATBEqqJIIkHM3mB/FZqP7YoJqXe7wILJ1q
kU1mmtuRAcvDgCUXlGgkbWyOa7f73RdvZdL5ytLtAEpDFzFBdNNUd1iXkStRhQ8SvIajSUGOWFZF
Pjh8Ijg6DAsFHSVTJuUQ12q5Y5whBt5bCmv9/Sh0xrJL77ZhO3vYZ7F5I5EYm47bs45MHUfIDb90
vJiHhNsiH/+FIgRA+mgdgFx+7DmtO80H1X3ogjYrDTXxpJNwREW5DcBlPayZvF3bJWqXgL3wubmU
tCrPrOnXmEQtP+B/MvIQmYOQFwtEYGJ+kx6m6zcKekhuCewdr4ARV+ERBxBBtMyUZow4SVYfSR6y
ZiDVUmw47nhN8wEwPGvIauCDsTt/4Ybr4UWlWxSYlLX5FdcOPXSSfADSvwg/kBjIAgMy8tZ0N6r2
fZykQUDPt3xdfho7OULBVHOCFL2hm8Jw03Yt950osMSbGJfRw4Xga78+0oPdw7usq+CGK0vXzL9+
93YD8lrJ+beX5KKEw/TXfafTc6eY1Een4eCla2q63SfIuk6ZOPH6dJjASa3xp6lJyjPX7m3FhoV7
U51AHNIQmnbTVSzCCaq+hFhWeC4WTuVPaogywJ/ghsYlKVeazdX3zliWipf3YhlMJW1/yOkrOXXY
eMvNcDISiy7/ZY5EQrM07ERyf4qzFAGIHCfQnGwfN47apmaXlxO10pznTQGfpE6cfYJSc3DTv0Zh
gHYVwGAxogenVyP45JIIgR6PJDPF4oFNkL9w3lFeaOc8xZUKifKLuzOt4zGpixqW0+vzfZ62T6sY
aK8mZTV6tpiWaGCZGFXBDN33IIdn/Bx553DUX9o6g4/PBH7b7SN04JB0Xe3rkfQ0QdlxXvzqc99h
97fouNn+D1/uQbT7HwsnStkysz+Xmc/HMNILU3A/vwvFpGI3U2g2bhbGKrxKEUS/espV2fr/579u
MlND2gLad837+hGViqDyJ+AOzLeU9nPHzLHMAKmdcSVrzHCwSiR3uzU2DAp8U3gG0SLZeZK9Oq97
1FnEpbGUYHKMT0rBk1S0MsVWDa/AZHzbQistxmlob6LJQjuNW0K0mLSgGsVvOkO6vVbXtwNqQJIL
FksVLzsqvEOYyp7HA1+yVWyOGJN3GrhSPFfROQ1jmgGmF6zzObigHsEuwjDYz73ZS2pIG9DxClpH
DJajBh9OjA7exw+QwtSAVSY1P82qkJhgLsvlOZYfBRg8eXd3nOFmv6SObB6gAvlxfnV0xGQsu1Vm
TN/N0Ljwri9tQ8jxc04XgZNEUwRkqjFd6WCMLnmxellxEhyWYWGXmLUy1KYl26bt2Wp+dib16AZb
U1zROhUv3nC2T4kclsL2GHMWL3z+oW1KUkgvbbSX10pM7yLtJG1mpARUNgEYpiWXcSUc16il8bpf
FeNQHAKQxQmWECuLO8ZpxmeVaG/uBNCn5KR/1fi5yGuX43xPy7wb7LuhtBYUM05witCooamK8A2a
KtOiamxNksYM5h4Rtp67DghEJIcZLNS+4oY/AkT/UaPYouFHO8N5FSYn4oHcXI/WG4H88eVejuQz
/cHal1lcXBgBG5LmYsDLIVfwp/pu4gxag5CPvIZgVNMLw21BWcbYi2CsJA/rt9eHQWbv9Fdd3hDZ
eVowPSeKwgZ74cjpMxEjjh7nZQ4hRzzftfp24uQknN/uJxlkO2M16ZlMfBAI9sxoSopZyFK0vHn1
zW0MjsFz0e+UAUE5emRE7JdHbQ66RddrYVT4Mb3lO60uHcj60yGZZoJJJpL+YsCOCwoBu8cqU9TA
K2Zm/lmoelZY5DIMDp7M7706qDc19ouoKK3dKmAgmbvIrMYa6p8TXD2ryMwAjAhmlfaR1h81sys/
1MzAkRYIiDxN7Uh05fCY2CpT3XbN+3tZ/FLX+sSVSfK642xY31THZzYsp+FW8Boy/lC/VK98xeks
CPixhfm2oyiLUIGTE2HIJiArSxJXBUpjq1jGH0elsTLjKKiJAdYrsJHIO6ODxzpLDtzN4B0F6JSB
ueDxw33jNdqMYU9WDGjSeAqRInb5a1PuTqnKThrMy79FmHvYxTKgT38S63EUSSwNhUX+IHCo7OX/
CbCly/+pHvIZy49lgjYsIR4fNu0KSsFfPJ8QbeuXLS6JG88x64Lc/qV7UjuGysnbF0vHJmae5xYl
jaDvS1TUq2YGteQYnARBLc27T4NLf9c+bCaSH2C6Ybj1AgFv9aG+omfbFVOXZ3/HgKbLW1Z5ukF6
Y12xl+9W/67grfJLfBZ/pMzenVl5t7zSs1rz85ywlfVKxvL1TWTWrf7oDy/Atl3w6gZoBGwjTtQk
9YzB7gCPYM6DfTgUQtsXdQxAMjquDWUFK0t2NfUsRNAj5Av4lJhzOFPOR7JLbPcBLHt/t1iDrrby
wgwVy5cC1AdjX5T8j/ch4lYl44RcAbOhZhJfTd0dHyYpusAq90LYvG1Q+IgU7YuN0KZTaSOIAzwW
3gOQWIBBe96djOVxNSrbdxG8/lW6NVv7LJDKm8Ka3USKpk/r2jSWdY1FZXvxWXWeFUx34NoIjjGO
qWnCjV3g9wezpyladLMktt1l5VZld0LFhFGxCKVmjFHR/g2ZOp0tLDK/LZe1CiRjPp59iXA4duYc
XLEPFvPpO29rzyERvMt66Sqcdr4Q2aV0z8mJRE9r953rBZSjvzVCGBT9kT79gtUlOJ3ePNVkaKON
zy5+IqWtB1THO/fiauuUrJ++KB5vzJxab8ERoyqVgE7EqnVGs1nRmrrjnX0ReqBPtDnRwrTamJ4F
OfTztyy2Q+/azQDAED5ObdUfgWSk7AYVNp0eCPHjXl4qk64k6SZ7t3S9CIFv4xSzOhbxg6DM4UQX
n77UMSAhOwbV2imXMUBzMhNmlrXPHVUYe7zvVe34uJfcaQwTsTfGja7pR52kivGvCz3zeKuT+QXv
4bpyMNbxUc14geGHtUtt4mJeAOOV/WL+nyf3PNjpz0B2vXaIa4tigkR11pkOSRZfIWAVQ3hOLOyX
TFcS5ozk5f1Hiss8O78+7HXJBLewSneBjkFLromDvC6jAzxcLyX3pwDML6GlMlmfyhudXQKi5hsZ
xsECuy3tRrWUajmFsqpH+lEcnLAIXh50d2Ga7KtNnrJFIogw612MJJhN91+I5xTWNd1ewQPOfQYi
wHla4UVpyE5ZClpqPQr59pg+sHptrRlJqFWFQMFlAJMuCIzfbc412LknpCRiyot8yqAj1ACpdiYs
sMPUxwkH4ghq7HaagjHWHfhQUEIGj/YmEHxXgI3ePmsuvWRGISyjY+nLzcqXchroIgQqARJvkz9J
s7RVL5vGK2LjRCQ71QTOgUkEh2y5fWPDJJ8m3HORhhvF7zUEM9MLepvLXX7TBzO54HS5+CS5x3t7
o9KiKPZLiB0uVkmsRHueCHwamvB7yreXC8oF9eEXaO2/Y/LFa9U35YxkKgA06ho3Z7//5I0L2D87
AkJyE+/AwottzZs5zrqYrlOpG4OznhDn2TwzO2VDg1WkxADSM8ngsHgw691p35Bt7tDLU5Zxm+It
xIDkP6vNBm0jESlOK1IvHawmhnH5x/S1+Eh778/thfJLN6CTzUW8qwzge4AhVojGmf1q6hQYE2uq
zfqcjUuCLY2kNo+Qmac8EIJj/nZN7HBL7WYFCwGMTfEc/okhJ87noN/L8CrfqO04FjFgDX7pSNM+
UCid97wHdM4jeuoTeHB/waEN4lZ9e9gf0DfvHuBQ29GntgxGQiehfzM++MeMIL2sOu5e629vaXc2
t6Zfl48RE7rSiFtPMj2djDPHVefngZQpCrM1Do8U9zwDDLTzPR4OyiAabz5iQlw7iF/yjx3z2pbO
IvVsffYGy3VNNmhJtFh7lShs/JSD2aEBYnCGzm4rDjf2tfTMPqnxHTfPs5nNbg4Wq5epLl4O7L15
8Bbp3f0IdRFrH+J/Wimwr5LTTx1L/7mt2lTerofsVAMVix2qYX/CZT3myJuLj94EpuCc/W4pN235
aI80USLWnHF4mkjjpPlxm+a+wM0UBqacHedfv8N5iVRhKw4ro0+QwFQtEsreetb2bRjT16AxJJIO
RqvqgCnPNA+9/Qc38RBxHbCBL88X8Azo23XrD+6N++W83Bj81ZEsCeeTaTXwHpz6+pexpIN+yS26
yvMYTm0UuSvHd7l7vAM0njSz53bjUylyQNK6ZPrK5lzf+jD1NHgbS0Djt4LYhVYDKFpeYSmQap5I
/94IbwiFwVxJT2cuFKQ6euqxOKgdmgb26qxYSaWgnYkDKO3t84TjnVUo9J8C88OEPDWij5Jry/Y2
OFRv7myAXv1F7LX2iAPQsxXj0MD1o+SUBkQGp4+tPqJpfvG5SL7IxfuFcHDN6eI9LkqyA2p4ioG9
1VKPTzoYa0bLMXFzLzAtLbbtnfy/k508637Ndx4OKWaAUr+ej+G3bJtk8Du5g2JhmPoDEsQJIFVr
JIL1h88QHCUy/4TI4LzW9oX1sLYAXfE9vLO1D2IqniH9x8QgjrKSa+8L3UMIta2hStV9DzEQP9Aj
Hed0b4UsXQPVq9k/9wRilDni4VtCV8LqNz19yDAEEpI52t96BCtRv3PCrGQlMmIlbYCzmwOaamP0
dVzOo9qEiWx1j0F5KBO9WLUjv/L8vSowNSH06oPBpZeMpxhe+g6a/cuMSnqmBdT+PcmIts//mWc4
WBX1aMCgaCqCdufpIwsXR+uOx41CwEd+EQ8SePF7plc25ZV5OzEj2s07poLmafnj5jgUzIudkC5K
9JZmV2n3Wa7WzsAw/SP9SVhuwEIQkMoE5dkZDlrnXZZYbLGbv9kfdBTHvlJxHJBTGSERuhZehi3S
1Su1XkhlXh3fyKWwzzBJ+EILo1xYIfUmBIIAzzctDrDellioAKtNUj7YqAGFHW0PtUJYHjZGSywi
ZON5KKKpPnmLAiSMjL1qBp4bny7Uap9C5HuqUC3GZIZ+u3HW1P8fYTzxxBnvr/lLjWtFln8oE0Ww
xVwO01Xhw6mlOMPDLo7mJEDxStELu2M8miXx/m3kRIHpOm69miionnZL0624MkrhaNy5npXwDFui
4FG3ThiRxU2OEptnnDI4oOmgNYlx6nbGOSxeA+pmbIP6YY8tZMPnnDfvPATo2GiWDIS4PV6oKteP
7YL0bupcP8VDhRa43HjvqgV0qWpSgOgEKJz7GkIlWvulfUMiCEcx/wuJ4dPR0J+vHTh0KisDyu8z
UNdK9NssoxngKD4xqAd3oqQIXy40254NDGokYdPW24ELjpPj9bpGZilpMKvfuoKzQpNiHGp75WBB
s1Kkrr+gAzG+g0hS03EkJdOhwsaK6yUixbK+KPazeJjRwqN5j119HNbc2T468Uh9/pmX6JtbwON3
vpCvc7VjJEcnBhdlc6+JfCqOYrFD8mPaNguvWsn5wHMX9I9kmlueUs5VbKHCr/4NwTJUL0mkaXU5
W0AOTM7G6OKcz06r+ONezdu7W2A5Za9QtFcINpyQ1oGbJPQxH6kvxaLJNybJe6/A+GldiXg+bWn1
zJs9QmtmXsnQJFbH4nXf/Povg2O5M1OGX5qtansKvmswqE1SjcLNj3SVY7hu97qR6Sav+YvaBRjL
zC4bVSRm1z4OZlcr6Jj+WbUHGigNm8Hb/oYADltzyCtASCp75n5wGR7Rll8m2MAoOGoiHuHsgHjt
0JQvTWoSY7EgZkCeMfqQ87wtG44evTPj4tB6O7Bck+/bzmLDuBXxc2XibtTygzBQXUh6BjZujKiy
eXCK6ZZgPQcyoDagawgg3irKgb+hcErXx09d+1Txtj7LZO+T20jq6V8tSw8XWhHhCO2OezSSGpR1
kDc5jBB25vOndq8IR/Ewuq7bndZjRdSHgT7Zfwo13fIsMnlniuWLPiUwSVY+iGjMKlhjQ3rVzdkd
lW+2SHmxi7SfASdDTPh1hbNPS6piK0tG2LJHyJz4i4hi9l6sJ/CX4dQXQiw9blNTM3CTB2QCkQZr
n8Er5nbrnZ4WH0m2DSSTUu2QralcY+0i72oJuPlzUDxMzl9GltNb+WfzsL01E0gheUTx4gUJD+do
/BoP65xyUIGUvf1NXGiPgbNQ873xd3gbsu4Hmoi8tNgsj8OYjQfyIMSR11Q5rDfalJHaOYM2hmLU
YfN84k0+s39OTra3LaqKweIVLqMDmlt+g4AS2g5gbCKVEAZ6stUba4bpCZr2iy9SyeAUNLSpLl11
p1+ferrG5kGA6ucS8ro0wkfG9l7Ml/NSQDjyRAYNtDBU5f4j22VrPv74aFIQY7dn95oNKLh/uXEl
Vnn78NCbjoPeqo7jS2nvxxtSDA4CGdGVJPyggGcHyu02d9EUlz6Mx/9vq4o/l+BbGv8GqcOgocQO
i02nbG3UUYsgQQr0pfy6VusV3npxAKwQJOlBxkZRnmzg0a4QmGgFGvSi6TlRf7Ffr+Icg1COjgKf
7Ty/z90+wXR4rPDx4HbFjQ1Urxu6cnXw29cL2E6FFdpHaGRGZ6ZswEoFN0xbZTTj4kjF8trRHNyM
FAfsxoEsqTtdS2ZMVABdF534w/vxAE/+LyPRIv9DSmIW5anQhyd6+BzbvRynuybRurR3DtOn3FL8
6PAQyw2XKKPWTNc0bJCEwqgqWSGjNgC+Wyiplw/Vk1fMZydg2Ju0jOphBzMbad7Vqn21zbFgI4m3
qSQydHYD1tpfyMusTjNMZg6CP1CEsGB99vakOHk5kOHToytjcaca4kcvY72xfNPdk3K0u3fkwBqq
hC7z8SFmDRkfccoeM+XQgsbTobgoU5ben3dOuIKFvNj2fZyH56MjIdhdAbvlgHddqsAuHip509Gm
1lQjx+JwYwJWjD5XZ2fEa4XtR7I/piKjq1/ZAuajMoyydZIkNLtBu+sP8k/umTFxCPk1h6kGOrS5
d3rJw15OWEenRg+nIdAsQ18I818mkAUjdl3GKBN1sA4Hw+Lxt9z8W1KOI7SjmFd8WUxJJSKlONhT
aYd4MSycULY9tVU7QnmLPUUOJa2k5pXBklk8FZ6e2wNNUq7hEb2yaQ97CE+4BOZEqipPslXbkJOZ
HQUzuYbWv7qubKVp0aEu66HEGH8UGB2So0M5oTf2DK7FC2RkRE+r+a8foMdPERJpz9VjQx3pepT5
LzJagCOW3FSJtgIm9Vq3XIUoE76AOnyfTy4h/4+j2Vjcge2Aw53qMcl93dvf/FE3Psjf/q2OWDI3
E8Helak7ln0IdmQY3oxXq72IIKrSIa78NaXkC7MuKZ4CpCfPacVBEyhkTcWHcNhxUbOL2zmsX4F3
grHdo8LB1huJR/f+/nhnp29Ksp5B4VqW/9igOtvXRcujKwObgJd1JKCW/eoejjz5qsh3QrBfjPgP
UDDkiyMdED+w3Xd3TyENk3ULMv+S0FP/7t8H2WilqSm2cibQgwjei/AFibILsz9N7pRCiKtQ0nTM
w5ihr3zPyS3S/5kq7ZunHP9W7LlxGbrRz22w+9sOKOFBlNYbUP1PYeCwWlu77XwF1hY2ijeY5H12
J1pFfEpHE9PNICEa3uEcc6LxyOIA3NzgqJpoREElhcjkt93syz1VRLIUZx1HTfy/wDBsGGnhpBQb
CJ6gUh3UD4g1+0TiRaqkwWtByQ4Q6Nq7nOTO7qOAkBMVT9x/+8Iau1cvXhwgUFGYgHKmUilYSSIZ
yDXjVqBrOTnE0JU0f1NDgHvJVzYRWDdw4tKHZya/zqYpbK99MP6qNPHTt26XxcD0idCJkyMMNSZ/
RlvZPdaaXWa2yw7kxPR+a+gtEUJfbO21E393LGvA/0Qsx7B/2KUpnZ+paTtGJq8UtlyWII4SUtmr
TAijq2WHLOb0zv8EXajcL6rhvFJg7D7PZd0twCEDwShSQfTw76e53pf4LxyUefXuil51VmYaWeBu
oOr4+0czTMf16NbmTS8S/Obo+HDTwq6xkPiPLBotIqv2uCNjdt7Um4aaByxsV58r6ibBn0Am1lkL
QrT3oSKRDNLy4Tjs/SGmql6Rk13+Xd/KIXAGKnZVL8LEOD87x6t/JyL10QLu+3g4JaXDrBbVAxcR
FtYLdzSsJCdGSjnaHYLfeVbH706xnvVc2A8ReNqzq8JNKb7Ai6Uw3Nv40Joz7MFGpy7ENdmvMMew
lUBwDd4Gtl6Tzh9yWOFefT3TSLfgxMwErZ9IL0/Q2u4Zed415q4Y8GYcBgwo0CHDX2VGCOECMgTZ
0P91UkSXJ0xCPDocBUQDIIRid4GjcC6so5dnpNu2jcysAVOEruqrC2E9ULnCXOIRgUr/t4LZph6A
8SPvstD+jac5K/BDvwjyQ+7f5t5onIAgrP96no9OvG7f34KtInEwUvVHS91ufbi600knYSbzgHaF
6i0JUWTTP6wI7F3gaG+TNl5SHE8VIpf47TRWz22cAq2LhIYkL0cMTC0QLaLKyGO3O8pGyL6f5XLg
esO54+QYh2NbsQV4bYILlNApSqkdQ/fNuJKMgHqBnRn6ayrTFmT1ZqDggKII/1snI4Ollu5jt8+T
SSE3w+7yqSWBwqF2itsa5AEVWsDeq0Csq+GGxrPBj5NWVzJegjFcj0zpynEX3T6AbyY9/Vb/9Njv
xOcDx6fkATLbdazis00hi63OKQ7TcPfwZh3enSDoB6p3AYk3e5FCZNMTtwwMb9fKJSvHc+x23glW
wxj68ewhGeBkW/yzyTkmrO1JS/mek25vsW8kNR0JkbJmXq/6+aInrIekr4iqmTQcC02UCbUBHz0P
FGc4evj+XMIXQUTE9Gthr+k1EAEoMthlv+fJZAG+BdsbocQ7Wg5U5djCd3WK29cJ4Eaph6w14bU0
wzWPg/NuXA9EjklkzYXZ2ibZqnIXasHb9/auenUoiKHBczKuw9+C/qMtBnjWN34r0+It6IXFHFvJ
zFlODKgVCwvOvttlUItttgcn/eHLObQG7wdVD9eX45DMr9OCKqtd8dcJinMUes96k1U0RiZrBqxS
uP6HfRPS0wl22gV0KwXuk7FAQvgbKKeDwZFqVS6+NvulhCS5kMpsRfHzGpBF6+2da+jbjbIXklU+
Imt0NiSCESETfoInWXg7Z1oeIvMmBUrkgF3vWe6BQReHeCzgahesodGvH7jd3DvMfFdMteASoLHy
S8l6M3Q9DESWIFa7UTzLWFaKSsS0Q593TNADXhYePLA2tmbQR9qIxoxBC1a3Mll9bkthbHwVXAMj
2EqRhvfUs2ha/BqZRcxdMFbIuItpTJnl9PpRMvhcIZc6EK9Vd+wk8iYA4F+IknA9hlzI+EgHKWSr
HWpxRGondls8XHLrngsFa6gQWtrDWG11bWZeH9Ql2ydFwo+k4SiAgB1wmlKS7v1Z/lCwtRVbUtAW
WNWDfjSX5pwK5sFKqzZhunSn4h74xsoHO+zl3D+6k3FDWCCgckWKnMkQUTgii6t69Wj6w9Y0i8w8
rEv1xu6xvsDoqgLP0Nu9f2XiLsE5ZWbLDxIc3i1UHgnn/HnGoFO61hU+qccnaPpugYChfNI6Fo1a
TwQ7fXel+47Lqgk4UhyBhL589jOPYVk7k1itTTIcqIz30HObRZxPRwTwK5M7M9X0XC7kjNx8JT4v
3lhgLjtlRKAYQS2A8JL9wApbPBI/s+JREKRvF8uCHCPj6yCiKoZpXCsGzse1gyViCso+o2hEI+px
svN7vhvpTnoXGHj+aVBjR/9pip9zeiQLVrM+QUBsjWJmTHmtZ6U9dSIIKEtHGGNuoKQBWJd8pveq
EffEw+RPwrYnGcJZOIwZgPtGz4LilhwzgJFE5eETlgu7gdsrBQW7xLQAiDlyd8iq4IIFEfFC1BsH
iB+k2iuSk4F19T6iPw6VXOBGL4ZZp8dgjxOt+/zbdRfVrNLGzV6QjUE4Ocuyefb7zo5VvVr4vgyt
b/osSuhPnJ4NyHsLmrVyzt2mwwARfksujJtb+UvjG/skzYoQgvMp910xSFggMKCbjncnXsXlGSpL
FMwAp8CXo8lQd8tNkRVAH1dXxiZx+IG5iVNzahtkDvgW30B3Low+XcJoWL32Uo90Di6youb/SQqM
hZi1niOJaObq4Odbheyd02voulOKLGfJY0SgGkWqpGVgRfv+JWcoB5Q1WB2T2jHkGCE5yA8cs74O
a3/O/pd9HrOpwYAvSo76Ctdh1jsEIHlfTE2wK74VzCgoqyNo1wZ3sLUhYFGWs10m0xZnasXNMXHi
zoS61gVfLqAAKilOmZr6Awbx3OrtKGvY2nFW39+fPLln+ho4r99c5z+y3Cd5AE0lJhX468/U/6nM
bPlyyfjjgz5yT8JGb1HQyxG/i6FWpA5oqjF7fHLWHkE+N/RzoNmjzveayBFX0uwcd59Ho7DzbmFU
Z3DkbVzaRaS6zMMx3po7GpejH8chc3zsun8HwftIvMW6kwt2ThYYzl3T2EWToVuzDohLzhsiPv6d
py+RenlAScOKLT+pxGxoR3CC7/1A2EjlfJIXWWSUtlm7goA8/UHtsflNZFWypWHk1RldHjpOXH5F
uq+wOs0cs1gS9V9g8mCYirg9sOC87ZTSU1Ny+DU/38DRQFh+2shkFFA9h1DDpxIAMmIo28xw3RTb
PGHDQCngQy8nOlyJ7CpmxIr9Fc5gJINVGRJixAWIJTnQ2IEjATzYMg8lhTHO96HMtI5hvQmKjlaS
16d3zZisc3JnnthEiKjsHZb/j9nE4JIYQ3Ezeab52i0vJbXDF5+aPniuJXNliYbHa9P4XaPfKSj4
DV7Uo/v5TWLEnRWzCikTNt3Iibpxx98gPWzV20DNFJlwgGXJeqxbhpxY/BQmLP4UiGciHWncqyDA
SHR+HZpzm5aQYCANlrIQ8Wz6p0nZqAFG0qQZRm0UFKpwrTX7LU58/yfxxJi4aPQp+CMp+tbYvjtP
06ck5jxtgHj1tPqmukXtcxn8egcPu6gh7lP6Nu3xcLocz0wCm2ptAuWwTXCjN4RGqhsFDH6nMOgR
hbiaoNq7X1xWH2tdpt8h6vsGYVJyLIs8S0QipClWGYVgG/9guhrAwmNiUq98EAkNDKzKkkLYh98v
COSGS5N/InKFfATB5Nm6H/53muzVcWGAMC1D3tTYDcp6Yw1RqkGtwXmWANkVoLn6zgP/YQjMCveF
eONeuKux7WXstRrlRdXJf+QiHLq1fWJk5rH3tAsk2TiV/uYYQwsDFEhiLg7bxc50gjvqBXSBiX9U
ow+e9URWNZSpRJY7grfoqvub7qAykKzvK8VsXKEfar60/xtJNshZADku4/A/ViUJuxsypR8CJtWd
TJelX0QSCcFSp+eS0N+LVVBXDRVjREIhomyZLjezmEPbHRS2XE5RegJwcDiexzSSJiO3Kyxcx1C1
wI4rjRmB/JjZuab2J10USxFxW2P73IPv83D+tQpjhJ5iYldKTDhwZ3m8X9Bz2enLtY9bRTdu/1vV
ejWNxjDlZjNThOt5oIWv47MB1uctDprwFxpETjsiKtXbgmmI3uizTxDcx410Y26Kl2pfK1099eU3
DMxWayiM7R77QtAJLNjZz1ngGy0rLWr16Dpjzd2GF4UpK9HPHUIdeFxXSitmoqzpfP07WsYK/2B3
o53EUiNEQa5AG3r0heNh86dPat26RqfTTko9r9Q18007sxmMmhIoKAqZ6klV4mySNtxH+FtJJTft
xeygGZ5a8ec8QqpgZI4H9saMXDGYGdPmrqrA3f4cPHedEvdMKz05zkhTmMIkXzRlOdPZZY0rDLa+
8LqUnEOey4vcrQW5PgLQ+816eM1kNqcKX+bs1Twfyr5eoX7Bj+3qrjJLX0jIk00Vq96/fa8gmzE1
KRaCltCvK7sqYLg4sEcS0Kd7JslqEU5qkfO6FkhhiEXKslbbnue66JVDq597VhAMeF6E14ST9JCU
bfbrzf2acj14WCCDeERqRFVT7/VMiBGWVC71iKF8jYs5ZRlRRVVUrGDw8LOoxHJiMom17QuIZQ1e
Dy8FwTPkL88BFJcmndxpeTk26f8jhFt4vTmOUO+52i9RytViW7/AXf0E9SMZvydjVLKYf67B41f1
cWbDAuU4cXnRZaCEnfIgjKdSbuBt+4DEV47QaTF8fjnrTgn6BT9ECR7xZWobQYVXHSBZgoIyYJTu
ySplut1ut/oSX6yxf1ncxpOWzIZUE5wsM6DfkHxb9Jc+4KaEZpKiFCSoU6tG0HXeZ1NWpRaumklS
UKD7LaDHo+/u+zai3eWPiQ/QVcUBFvWmYB4Xg0nY5g8JwmwZkfm1dsKoejE+fMEYdUQcKvRsdFlr
v28ECoxzc4MAtnskqqDNgGOauVtC3qHAIi5OIlzBdY4XzegYz5ugWwT5V985Ixmv+Co9sTBidJp8
HMongnnBQBt7xCl8NkUcATiXK5g9px8wtkhm01Q71DaNPjsQA8D//M5EvfmpUGJTVdH3mFCXxPIw
kIjHdlDH2VdZ8IqPBAAwmL9GdSmoCZFhwObUUuEr1EFJ4LTo+znBIvPeBnnkKtdiUPTNkyBIBJyq
x/Nef55z/AAD/KcFEsIhOlcuHqK+9CgzzN3/h9SzYEitKZUFyZMJjXkG8XgBRzcEHTs6y1jIJ4i9
c9pMgHO+oLPoVJlOJpUEQp7sSvL3YZaTQOnmpxip2+ZiSgYZP122SVB9vKV/RKJvYJ6alJs5PWlU
oR8UOir9gDhBIBpwEHv4P9tHa7tF+Eexl6+MZpKcD4XzHRlx4R2y9zZXjjj9qdo4XPBWwbYi6Ffc
GrqrRxTRS6DcEuScXAFnwCiob3xziExVnDdFaqYKB/SpirMg9cOG5b8WcgIxUye3AzXht2yHkPlu
ImuW0zpCr9uaOqNYFVvDrd0bUH8bTRN2yDm+I8GFxViB0xO2DuL7a7oC2OC0sR+MM1QweTlY2S4A
JHO8x6k/0Q62D+GNCppy0lkVz2AZ9TaLjWO5n4blSBzjTp/Fc/Mi9p/NoXhbrV7SfbTeOTO7qX5E
HsHYRkScU0NRDeQ7Ff+gmxN3hQi3+Fn36exrPtXjypsjrGHGWPKyd5GT/VmFOwKxjAWcvhj5nZ27
p4dVcyxz6mS6Fx4VnPuogDb2Gvg2QXv2hs2F+9Tioqh1OQAV8bA7l16uxQGTFq6fqlCydSLNqCrN
0RafZ+022h+7PeoHAHqfXcU3VdE3FdAMfNhlwa+7sK1WcLDtSUjEvn5Ch6QAvHPD/qXcSvGqaAJx
QIeWpAaUa8dv9/ZMzS1Du+BHtZhd8z0oPLQ3EmdoXHIVk+1uGs89G18zgsVVdTC8zmx9JvK7c0sp
MB2M8alqHuIHW9uiyklyt073+eUi9j1JrZxs1xiWdQbBoloUfFdIR5Lw0BUA1PK4kP23SRDYUw3u
jXSU5S2Z3K8Wbak0Xf9TQ3LuMK0lIbNSEVZQWYa9BkbiV5NDsAgRpKdZbzvRtm7Bvpw+S4EnnZaN
8N8isghToRfQpAtRvpiUn6mBklVfx3g2koRLeffkyOr5osrvPETdedyHlI+/jYEXug3M7yFzEGqo
RkaFy+DB8wFeU1meF18u6whMROlJNCxCHEEMOC/mUazx/kx44oQeaazQKRfcmLiSCksNGSUtin+N
1b9yOzUJHO1Dxst7Yt75LKe3aNIS7vZirfdimATJDXr8Res5TnhWFsn7xYGWmM1bxXDIool58YEA
1PnI/kGvUXs2ouSl+/fL8i/c4ZX81fdLxje4qACAptRz9MXFD3WdVDsl1D0Nnf5ckD9ybmJLfDt2
GKVUa5CMNW2cv5t5UfGod7YkWzsvIisSYWJsurrrc0smWI3XrN2Ss4aYkKMJr+y64ShFF8V6HeZY
zSzsAcKleN+yxyJ2/z8e8NvnLCHoDfBF7YFxc+1dhmxtT/LqzEW0r7VnqoAYpHaSuoaYiH033tyI
jxwR2qp9tIAoloGuf6f1iB2Yyvh0BKWFAxlXoba0jsNmN3I3qy38ivF3jiFsSDrAxAYAZ0ZBSf81
io/MtYJzjqZtKQwfe8utb93y6/QFAKnkCh3yHgSO32bRn3XKCbrrxgdbvkoTfKPg/p2eoUFz+oPd
Zyq8+Egm4NWUrR98BT9ELVnNxZpHMyC829700vf+s80unyU5MGq+EajhWNbRf9zi1Dm+nzKCaoYa
PIK50G1MgZou2iCejn4AvOpvLVlj+bD9Re+HuGUYbKeCJhhNnhjuo9ymQshUEbHDyEtH6w8fBr6x
6uPDaOzIB7IiNJ/O7zljZ8O2LOuCiPI50WJejMot8r504/vbfrmDhTjYNzhla57nw+Lk880dYt3q
BUSQ6Qfqd2imNQqvkeT5FnecTrAmloFUJRKZLh/tpbbPONaDvzA2ltTPvI924TtwAvtRCCobMHuu
RS7+/j1R/O/IBg5oRDGKGUnyO1LlI+GJ2ljkFrjmH6BcG7KKl0zjvnUPRcYTBCjssA8dqUranqy/
XUffHWCchEPUPGLUuo7fIrAHGTNl55cdmnjlpDqPaSa0kYuFh0jzQPb8NTfJ8rSYpm6kvAH0g9dJ
5B41kHrM3YcRBVRI7ej87S0Bhci8hXCqnm7nEH19q3hXBN+UDM0Kex0FU85qROlydxQrqrxDwiWo
p81giH1Ap1seryUWCQIDocT2KhymyrMR44vSwAFlWgPDsVJK4h92TzotWqs3wEA5e2LgRUXO0SW0
IB7cBahaEj8gVvqyvht3IVgMq+VtaS1M+mBLVVlWspFm73XYjOZcA7rL8Z9knRgCkOLu9Ec+SCC4
0gmaVpykmyxEfkGh2aP4+fb/TErc03cPLCb7s/7XDhA9tyWZNOD/1xFW1wUwTlJBThomxeswmZQx
kNSATDjB/POPVbz7QfB1Evcyv7h2eXER6lAxEsjeNZ5IOdkwVg4ZGSphw1nkYJhnyoS3NUqff8HM
E401up4ePPARIQON15J2d/o5hRCWMKxFAYkYdAnfK5IXeuNvF/69bS7rkDFiPapJ3RAcvsJzcbor
PG1uW1ys/GpZ91sD36F7z6pjlhXIz1j/k1Ndt/MzV7RBQeyzvkwgVooixO/4drljBJcvvFQ6uEnM
UyBAN/SUyyGHQmXDBW8B8q0bhZsHuUS6FEO0/obvrMWI790VLSorNUiGfjn7chymbXV+ZF6rqwan
hfz2INBW0CRQDugvSE1PhXgYe71/QnwVW36s8sNKnQhHHuZPTaLUK+uXX0k1N0vzTik4qFlLGOrs
k6srlYyNFOwH6mToEimoGoP1oR3pD2+P1D6qiWCnwdT2NH90YMckQo1fL/87NoAfTye1Z/tFodEX
f/LabiwrV2rhq3YpqOVZ1VwdM3mqWxJ2O4XBj9ecg9UOUIpmgscDzRf04n7MV8freGm7xvVg+eKO
q7lBvnGf1/TB/dcyeYSmm9TvVTrDOLA0IfOlM5D9t1du9YqiTlXNFUFMSQle0MDqTnnvXCKY14I9
tyoglZZvyQllk9BGq6zvKzCPoPNXQJh4SwceWCiBibzZRfChzkVRMhQns4I+N378C2UtbTuCm4o9
jV84176S3Hyx1eVgaG81fID0nmCMqIFxfVV/3HYxCr4D2e5Pl2U0kpFZ8oq6KXfI8k83P8LW57ng
QFKGHUzPYpFPtPgqSXc3wKvF+FaeG//N6ezzvBAPnZDv292jdy5CWRYU7Nblicg7QFC/vtufFgwE
eqmXi6y9HVx8ix4nZ/pH2vyYhaMkE5NPX+J0UO8xZJ8HN/rjRIIX6V8tYAzL4k9JIKQC6w7kryTT
tSVY6Fj77yUJgg3Q+h2+XDaACLCluhnJ1VQIKOqTnV6ehdr2NBxix0qruDUZukNYIlp5rgF9/mRD
f/SzXDONeL+DdAeTNEXbCQ5x03caE9Qa5qMr9yInSceJqib0CyYYPHpA/TGWapIVXeTyqODb8xPO
0kmRMR6FzsmxrYZAWGRH8z13GwtXVnRfTSVLudaizcJn7wNHT9puXqqNx+CuVbop0E9vO07qYfEj
uGei9qwv+vC2h1+QTiAU5RJEF/iX3XrNVlJTecOMEp4yVMwAW/fecA2jSm5gmc6S0LCd3iAMWO6T
FZYc54uI89Q2AC/aJ7gQ12o2nwoxfEQ+UNhbduA2NE9Eoiu6hF+k9bt1cKbEuJd07U5T7A2qgzzG
qGd+IVeMlrJ1G3NnQAHvKcMzqxKqIHXYPgmg91KJQO6uI1cYPLipwrE2Y+Z1BzUNW+lU8LIkbK++
x9tSDUdAyOyb1Ippr/Sn4OmbOoSzcqg1vaLAS4Chfy87ocd9WlvKRZU97Hb/HmXcYDM9YBPCGqDb
I4zbVziZo84YDeP+mDORN4mXYzL7m46eBXcIlt/bEw/mYktNe3mnBBLobw0lEMX7kXI0iULs7MNC
BOKmvUA2k38IrAdiVXQTYM1RuVvWQOfM1G+L8Aj119iQcKiZaC/Meh3qwBZczJKq9MJ13ONsYPAF
QX6CuPQ0ZlHD0p6Yy4zoJFj94KGVONP/GRauSNpom3/L0yLu3fSnJLzmeUvy02FtdsgFCQTFfaaD
BGdZtVmxamtI1Z4NeTz0uOXCg7IHcFN4O7HpKeZriYKeJCRo75a+RKHQzDcsOgQ7+enMey87jFCc
TSto7RIlfC1EpGNauKMH6sP3jHr6JaLPyTdcaN8fGl53k/dhmcuwE8Ur+bv5slFS2V0ISwsj0hW+
dm2MkEO/A4VuDcHnF5dTNoufbymBo+hTpJjuRgizayeKRafLStTk2LNDYboPaSO5HGBBHyF+w+Yi
9HxwCpfwj5ElZimxfojh3stEr7BV9LoukhgK+CViWYy6zCVp4C7OD/XjXQCf/cOKi0TNLcovmWKP
BgABxmhth7RT54y9j3VzJvyAFxmv/UT9H/7yfz7BfyljL+kWjiprwTWVCtJsT/lBzpK8OXxolVae
c7j4/xzlFPGVFThxRIo7B55hG/0FVGtAieSLDZAt+/u8HoBSlASePJxHNm3tB2ndiy47nMrNjCoZ
raZ9WylTXAXiSgp/3COxKINTCs8xJEIOfEnfuoCW+j19rjuSuhpD1iryZmt+TyYlPxKICV9KVYnB
7SNebBHqbbE8kKw+9/2ZIjdMzOgHo6Y7TbLV16aIJ/tnwNDTdt316Nab6P1UchZoVdN+J8uvU0hu
nsFFvGlFt8TKRBqmdKeRvvzcf2jsOOlBoElqvaXSVOZaIGo5ZPypY8wIDfK4ceKyZXzZrRJcFaBS
ozDuVEG/JK+qsrTIIxMykWvJB92LkPp5dtwG2Zu51FBRuSKGgOCGTVcCrqah0MkiguEQPffrW16/
uqmPtYb9uXX+lujz1awtimeBdiCV+GpcSAL2NxvtKfKWulpFLGpkP2vof7EtbraG0rODrHxsHlYu
ZM75qhOxXlncKGquKlbdQBm1kEvxbShwLT+cXTczvEwJhFTEbsgPPkduB2r1EytfPKjXsr9OxSL3
jLYe0go7izP77QmjgiFrwP8GWbSAEaH1VEm/fzXkNAZOn6zL7nCKpEZ9p+hRz1Psut42ejBBGEVv
pE6Q9ve6jtIToxXmD7CXi0TxOBxpd2lBEke+1vEOVa5L4YMnim+4ZCaxEgA1Gj200PXYTVNM4v9J
jsWJ8BETKqTiRQS5r7siVbBZCnHc1h+lGURoh4hgWSRENuy8mQe4LTceajyxUWW0CqekwkTCVin3
8SKOURnnURDztyiVCU3WwrAD5P8G9Zot/CJIWRmYE9BtoGA5tdwy1PpuPfW0EGgXoQAicUWqjHKh
LISDe0r2hT0amM4wCxXS4al+nm9uP5FVhHHYFVnVDC5lVBq2Jo86HxwrXR052eLA9MY50Or1b149
Mj9flRBGdEdFA7OJQ/y19sN5++euoe8QUKdBduDHqVur3EAAXObo/jysdqsZXsh7EqLZ9Vz3pwqH
CcU2rz+iByBG3doBrZA3f3PUQd9jA2uLXTsvYB4JlM89ua01qZce7kUxzN3L8QiiE5VfaFXU4ZZu
e0P04AZccsBz/ZW+R1bZ2AzMM3cCLkwfildovvTyUAt+x9+/a8ZXZxWX5G8BUuA+11A3iD9ZnRcU
eaPFeY3NLJ92S1n2bNR4eBb6OYJ2x4JbX06FPaTr9rGlLOJOJyBRkTLKbQYis/a/5zSZ6tay7tGm
dXv0pGesDeczFsX/Kd6zaNZ25I0728beF/JD96YdOWlvr0qVefuLQjzTL5Jju9dVo0jektFSyGRn
I8WT3pUkbu6B1Gzhl//WhzEu9MbFlkiu8z8Wx3kJTCyQ4h29FWlNQ+dxp5xHCyYwGySQhhjWYdZ3
cn+k8WILu8wIPezlFJs84qT4b4a960mDl6oCYumYFgT6zmuwOYUl9QMEgWfhCJkKRd2XruDRJN7y
m0yV19uCVP8Sc5Wq/onPPRdder2fnvpy24PH0UBydLZzyf7NTUjavjA6LbN7sGHk4YHdWvnuwZ+m
CaYLWJfRwZoAYQxiIwXo+98dVVb8XtnUxINuSyXQoKbSCMt3dsFdLhky09ytiyc0LJcfpbHuEQ08
+/oYGCyUsBReYH8P59Bl07ynxHEYUs121lR5gvNTWJW5boT4xnjMfBDCrLOaqX8Us2Egzn67hTaR
ujMHE+Hfl6U/RirHCdKWBlmNNl9/phwE74xt8xJirUPB2dsJT0uVny35mijvQy84QPBmZLf5Z/vN
V0KzoLRCVJKIrBKKZWgJzKRCkVFGvszsQRDnVFEN9cXedlNowQFD7qEn23Df8tnbj94ezc9GO/N6
9jYBKIkbSfz+Z7GB/mGvXr1zR2K8+TODMQW4TIgwaBcdcbTQVR4+qamXBuW3TKohO+g8XNqhzc23
asWNVtM1rkdMwUS/K1WneMI7qzhuOeo8J0gHiYAaKrNWpiKWcjsT56LgwInlEQqRVvNFXWO2DIBk
enw82+lYAhK8QqtvFwBXTFPCtWm9GKMMO7nb8jaLd0oOGljONv1wzfVy3fjWp+5JYR3r4V6tXxxD
T7W8fuiufX55hWbyRGwsmzsPU/oxtzOJEpEaPhff1b5INhsP99SOMhmZ+5QObCH5W5VqarrliZo+
MQ4nltFxeQfOAOqDq8HDcYKjMsouJa8c6p2WTH+kr56BgS6BDiWhPWjPiS7UqqEL5/3fpC5jwwSv
6eD1o4SkE+QzQLMeMSP9RNx7g2mkYvk5Oac2ivPBf7KCTYKMc87vr2STG9c+wt2HlHuIxkQ1lmuP
mnP4sswQTd9p7IiwJN26shH/6zpVQiDMGnyLOKoHIVIpD5/6g6jr16Eoc97CimUm104lQ0G9oXaB
jh7iS9NrMGh80OmZNF2VOiOk/YBf6eCUYoU06Ol4Ysvjma7vNAR4hJTqb8wLjHX1mmsuAS0G7eQl
Bkzaiu8RbNKFjf9UaZfx9OXrIsGIv9pG8v2ZCAqvY3kzHic5gGN+FL1sO3mCzfVMcoHt+Ys5dTgO
a3S5eTLsJvIjPtxzD1X2F/l1px6cZ1LmwV8iTDMdrEXRtcomrtQKtSZD316TKWIOG4O46fh87Sm+
SVZD+t5VqwWJH+Xrk5VAOOyt5qGg9sKv+WtUt2Dl6ON/7vHzt12o4ggXGjAEt6DuXdGQY3Ji3L1o
YdEhsmH/WcLpMUgxEpopa0VfLFMhCC6riKNKGirl4Jiz6FvUUZ1GWVrblt+718OXSLD4SkHOc74X
AOpJ7liolosnVmaJAncuBhdTCcgI0bkQ2lE2rzJkDDkqPAGY7RVpwPXFnoFxlZvx7YcvC8x5THqO
vb6EkkoI4Q0HVxb2lTZ/+zzzpMzugh/8itL70TsIAPfPpabCqOXdggmm0IViQhiilGgPsUSvoXHj
iznPJYd6fWLdigvALv14l2C1z1mHRW2CTwjxPfh35bBsYm8MDKd79U/vlh4KABGo3rtkyJYX38Da
UZI9eE32Dvz8/Mm/0jqZfE8+2cCtSFcvoNnj9uKBkXaW3P5hiLe9Oe8YUcVSK9cypFPo6SSjx2jR
y51sue8c7CYxmqft45AWY83yjSL5bR5wmD3pmZkIPueDT6Yc/Pz35LGAVkjsU3nGlft4XUof+lTy
WY1P8Tk0GqpURqLoxJymvryKR5/KpMehysNf0jVveS2xL2tn0e9DrYDrIkPtP9U62WDy0+UzY46T
oFtZsSraQvwC5K9t5KXVyaMalN+cJ83Qs2yKFh2VKl49yUKIYXBXFf9+EAZRjiX5rNGewiR72FTo
MstoURKgmSElxfe8Ls0dz3sUbLveXCqxa7/1lAOBPN5dKUx5CuBmIAeE5beZvIqCmUG+TTShDlKT
cPEN9mJjujXuooeSs8h1Gd4N64k7MBYv84p81CEQgNeou4nqYq0iC0/kZ9fPfKmK30c/k4KTnWPa
D1NGcTAqyugxiGnqfvzJh7Q+8DAUp5M9bgFrfrz9PXEgKcDnQ2Er8V8qwayg88/oDl9tQ7jBpaCQ
4aODj/6WeW4ULm9drmyySC+d6z+7VP/coWdH9EoampFTXOvSEb/wcvw96EVsVWTKQ7VD9ADMiV3n
8gckbee5VdZsxQnHAwfQw8zYz4qpSUItJnrDJjQayKzrRjBtqaDqrW7F6ec8oJ/q1IMVqA3POvmg
kcIIF+dWUbQ00YI4k9OZAOsBC6hkDB3jZ+n3wWv0AxJreowcLR8zPODOAi3169PhdkkSdYS/aKR2
4MukE1kWfoZ6EQ4kg/vAvhxLnyKPjcD+PdFHqfTeQYRW3oUfJuz7QWzQJA7cr0em1R3D29C3cnO8
d0XfB4+4qGliqdQc7ukkTRcLE+2aVMfU1sOYYR8K1oyEassMRbP6rsOpDgdLBo2n1LuVLGsB9Ui5
M0djnSQR8LTfcqvNk16gew/SvDnh16xFpJSQJ8ZNZHxG46oJLQfIvR1TPuN7Vw1OkyGwD3NXRxM8
jcZpi2ueGB86UNxILVnWj1ZNiBUOy6QC2BTk7pdwPQ9Wcz1rroXwWGgwTEeH6BR/UJYOgo0VjYRl
cnkbxio3tlmLa0eLEP+J4FlsyyJmFqzs//XTFBLyQEEZxCIcr/7l4/CESvN9hKInEdE2zrBushzi
AfPUt2cF8M2dhH5Bd96VGNIykArq0wqLrI33DkFlPbaoxwVQCHQm9f1ufFakgau2X3wgtrir/u4/
4eepILUL4Jp6TbKVfqV1KUoIgT+R81fwpISOWIDdsobwv4sq3YxorTBtaQMi1W4NXCTbAg3t4P4a
vu27NlIxzffYdt620raOmwKWsAj2bZlysaILWcTVAd4+8ijWaCz7qzyRpKneENM7OIdM8ZuJrc88
4pmzwrL8+McAMdeAD9MychMOzVuDgVNYHAh8ga8uk7GSEvLk4JpycJHojL5fTWMbz60IFWbXDz94
uM6d+d01GYUKMenKwFpsoTRSzArhaKaozi3o2VsHYAzqcBrplxir0pUCt8ZQTHEBMB3gGdwtv8jy
Asl3bcd9Stxh6JTfjAW0qwTqBfaz2dOrwMyzm/VbBFyX6PIEImKvorgn3jeGqWPEyuu8BP1zkVHF
A6d84rcKwN83FoY3h1USDmboy17vhZwcxNujT+10D00EUOnGA2EiVo9ZzcNfooLTBLQuF8rWFNd0
nXJabjbMjIFWp0nI9CDCKZwX/YDOrcNWMi2FX21DB3H4fcoN0g6eGThnNMI1CaZCCelcPjVNTDA6
bI+72e73bD41ThINTH1eziQZ/u5TJzBE6n9I9MzVAsdJaYxDX3Q4hlv+sw5x/1nuFYxTYIl62sLU
UAXCdJc6kvlV8QEgTa/TScuZ5AQsAYgFKmIOc3HInOalQUeRouUSoHuPB6jawuaN/SxS4W5sCMxT
GA1KrWNlTlkEK8UAVkiNpK+pOeCfiXUyDNRGPmDpJ/3KuGGfqI4uc2pbTD9du5VJ+fDba+sRdSYV
A6fHWtZxcAE4XhpT2WDfxLB7l7jd0r0uyJzpqPWTHCR/ertHDvukh15PRasvTiikSkzZ1lxKBhH2
Tpmc297ZtPsWZCtMCZ5s4hV7MVO5Th0ighB7WekiD6XpzWQzoyimZ6Hn23661ezPJgPF40PszWPw
HhNIyt6Sq0zxWwTEE3Sd0AZVX9UnRwxDU7d6GfCtXhtWi5WRaWXEZ5KWh3/7bXfiZQHdFg7vluGY
K64QyQe2idoY/P6txI5oj58fgJfxPwmCANS7nma2h73bwWEmnFpqLhLRE5woi7lVCehU2xSFjghD
UDWp7xUPzUqDsKmt77jN29qEy/LRFQDnPEajA4EXav7HQ5p2Qvdk1FYsi64j6QYN+raSs6z8+EMQ
iKLKoQx8giflTBXjAYwbGtv3whyrTZ0CS5VCs1Fe+0TAwsW6M72MCj/0cWD1i6N8MCKiDFDYUlj1
/LnZM5PzY6tFqw1lDTnk/NG1AqxWZjTUn3SX9W/EmRxqV04byk8rn0YaProMS1Cp09lD4i0U+TIe
N4p22vpMolDma9oSHYBdAlR8lPqLcjEBv6mGZX1S21yKwRvOeSTSAbdI0gMwvbFXdFLZO6iRO82i
KLAUkMIWg/GL/5dGxnjX1uN0qhAXhZGStuilCUgM0/7cynx/vqzn8tBhpJXJkfP3bvWajjQGlGsV
VLbLpBDiDXTogMg+qLss3bNfxwISzZlJaCnT+8qjZThXaG5/oa5cPu+Uoy7zKbXO7M9AxObCZ4KD
P2evkJEcDtfGVzkayu19CdHKMYEsk7BZJKv7IQMwUnz9Da6hYn4kZoizbzYn+BXtS14C3OFC2+6Q
6PoEj4u4V3T35nDhcV+v2Jv4eFcO8Un6VqHdOh1UHAVBUK0D1H2RhGbtKXZOOcFJN+NkyUAp1W08
qP61l81W5knstrSVLK9M3Geu8z7DNYidUNQ0DudH2YPeoczm+JE7Tvvl5G5dlYi+JNJ+uioAeuex
IA8vpP/pMoqmpBKX0RTzuXQDP89VKrHWAvkfwukK5DlnDLvWH5ZpgwPEyfdC+274nPW0Q8M2yhfk
p3SKe1hqP8nNXG5EnWF8Y4AcZMalV3NyJP72+RC/grdIsqOmwh5GLIGOOv4XeyNnJFLeh3+qhEF7
jrIWDYxgtUl2WCB8K2biLvkCwENLon8jKXlkoqyCiNW2fsAMpgnEn6P5tc277e/6BTA1q5spT/YY
fM5ygQfB86XgCLgvlfw7TrLB+hzn4LF8cbzjRj9GeyrSbSDWtj6ul9RGCIo+OlL4rIWjRvlnMt3B
5HKUDYuGaUCcyWMrU9WXd4B7L7rlo/N4spSNsM9Y+wiODXTFmgWxpu0iRQRnEEBMZQrM29H6NmEj
qAhTIelkPrpNepdBCVt5A08oSrlJzPGHVRZYDKUb+FyT2DUpG6yC/GDNu1mTv8ddpDj1+CsoLMEg
KebkqB6bFiAjxHiKtrg+ClCC4CiBvFrp+rvHLGE2zrrrKnjoPhHNqxnYmte4n5ZqWKq8IIC2isb2
RfBtDcSnyslvZM5UQY2EZ9EQBrwfVYCBcgWB9/y4/wsqGJleWRHp7goJaFofKTi3Xgtf7ld+zbEn
Ow3Qwf8J9GleQG8FSxOydFZu61nyYt89cR6C4mkt18UqlzRb2GHA4z8AFZO25alkOp1zncO8Q3Ti
sHEkHjOpdu34LGRU97uwF5pNAdnu/3XF8WouHOyoIKcroxIYatR3b0IzI+CEyleRcOfiiicrHcdt
slJx2wEqLshMZv27CNEl9yzdFF/xqO4j9VRzHwFrD33OWzObUOXYqL4tsIwkd65meszRAjh+dfZ/
I/AQXOSrGQJPz1XogBS0oPSMBgKP2+P7Cvakj3WMZ39r6xEM3KQkPKaThB8vCO4Cj/7pcsw+836S
wJT6IUEyHP4PFCpbDd4fTa6f0d07v5e6UYl1jekNrxCR1s15Xew1udFzIKgsfCF+tF+cCs6/Q6Vi
KKlvUlwA2WMenOwhqM3BkKdCczxGCh1XtufSsAs5/VJcQ5Sp/hnpJt490IlbrW6DpWfOkwYvO+c8
VOy20x+gXxzeCZhkU7LBTDrOsrxDLmwk+kJb3jF/+bIddrfarYWZ8e4SKA0qX8VvHDCUwyJPxM35
gAooUGxoO7uEoKfA9EWkBWy1t43M5+XkkbiW3HPXH72tiwc4n8jSL/ekGGyHWqAfGSLG7247RKWg
fouJ5/PpbH6D+ZAdYXTYTjUNydhv77JdPPDlyoU4CfMbReLt0JGYSnZkzdLd5hHUPlACfE6BBxZW
Hag45FdncMfd+BDHWKZftdn74BzIYgMyBXPjNT1N+jEkW+yB60mNvBvJBIuDKS93bPaEE2DSc99d
8dKNpywg3zg0MK7WolXWDqfcsJNcbDGSRS+lZwaeO/3J9clMUPxbURDv3VEjf+480WqJ0vqnuIGb
5uI/cexze1PQApZT0sSkTMkXcwf7SIMr9pBEyhwr4Iu4/bqI/wlVf5swb7BsdfxNxxwO4h7L1Uud
h9uOSxZixGCf7HKgXFFug94wHM53XKppV2Osf5o9aXL37O2tJTxRCTo6ydzZDJEP/lXMeZaZ/Qsn
ywRUeQHPpSU6Xr5vlrPRQxLRpDUj44x8hmDSRiOPLeMSvd4wSu5h2nKn4bgQ7sNDH7zKJgj71FKz
9LpjRVqfYP2AAgMvWIkhqXSmxc7XN5LEavCY5WIRnMj4CevAqmE55NbOE7IAKMZNlY7wahmhXrz+
ixer0/G0ohSBfq43uo2owZnOIUffKz9SHlRGFoYlxUy50+p9y3qHolouaocxVestipwOoTx4nQj2
uJHpGwaKPhv1SksNs9+QnPk1LEPH4Rn0RVvSCDzstyXiBTf1B1CYzOvATEVR13U90RXZIOZ3C1qY
xR0zU2DpV/zmaycyIaeI4zk+Qy+fRRM8ppgxey2jCAFY9eFeYIvTwSD1RWkCbgNTs2xI/Nbgu5rH
lmu1qs1QtLaR227+6kS9SyhcsQENKGYzpQlLpnuiSttkUY22UsQhDDWk7ik3RQgO4hzCGHoNobji
N4BaZlRlAIYq3nQqaboOaBzfDxlyDe0ynuMQApDxbWFDUxrjnG6OOYN3i1771mPUawpB554zGpkA
LJcHegij0agSsHW1yGh5GN092974CGj91BFc7RTuKHxyTIa3laCVeBBbzead4rmRWYg/GW35k7wD
Rhx1hFuxkfmyC8L2mTBQ7kWj/T4/2SxyBl6hkg1ZyUAUOQfmT3EWoZ9r1GxJHTonoWNIAqLPQL7/
tu62iIfmCHwutKZKCCwg7xq5EE96kG/H44qsjlB5+06jCkuMGXFwMshSRHEbdAVvll51VX6JiEd7
wtdT3ZYChLlMZ8fyMK2HdHspGi3JgrqHhJPWbYDHHjF8+RrrjuNm5wv+pRjKiyeIl+pejYDd1TIF
6B2HAz7+UwsRYqj2RyfSqMzm1jsd0ca2TtumgeZayc6qRW+ptuj1Q92ENEdbztGfvavctpKzLoXU
KaC9Br7QSNhBWDcPLf/s4WPIAkm9mfGlIJKwYv1uFGvJ5gkT947pJLsHOKh1SolgSoC4KIVkxDUu
vp7otyuDUKwdnm0wWbN4xKjdQXldTBqDmmR7Qz91BW85lieERj5jz1rRoJc2Tw+gRvoMxrEkuq93
AkdRtiRH6QeqfqwOFBMtJIvqm+rt9RXT0dkHvQi3MVinN3wrJYfUgk/b4gAOvRMKbtBxXbjlEXDs
G1nLcVNxKR8TlvX2EJFWyeQ/2al7wIxmsiieiJHsoyU4L+Q2Egd+DCFDg72Cy1v1JTLB41M7nTdd
RWU157GIDIdTqBZdlu9+4g2s8oqSZeWq64A5mtDaxWRVQIfwKagUC9pia12OGirjDrX3diTnIAp6
QyQ5e86mA4m4zg0sFsVH8qguLQ+wPbiUpJd0hT4f9k+FBs44v4fxtGYWUYsGaiM4rkpxjyfyeE1N
aC1RFVdx/J6AygMwdXdYC88zDh6c2yjqeTb9GxdlVzKCi/Zg652qsX2CyuUE0oUKtzS3aCtg6brs
GoiiDq1WyPvkdqrc7UoExWnPK8hKqeebEcuGhZ/WrvLBKhfMjUYBsqVmnyexAqKsJNV3XXY8zsfO
1evOiRHiFs76pfOAvxpxcUp14Hi8fOCuSN5WtiD51aFXBcEo2oO1YtUdteQI/YfyemU9zwgZTbS2
gyJGfedmvCxsePQ6lqy8Qo173RF7R+b175SSfMgIsvklh9uGUUxexTt/5R32wJMK5jOZXswFXqAW
VEuIOiDRGbmc9/k/KWPXDuyiIdUmKlZyoy4airWiGHJofaWSkacJDdfNtd6Jo/V8CRhJVvK3pBUD
6mLktRWy/D72MiFh1PGxbuZifIg1ngIZUllPbeygO3meYMwGLb4HDkrIkgfiCvYeLIHc0qlDG/Qm
ZHBIg/nGsduf4Ppp8yOpR5WyE5P+v9jfw5g+8hj/4O901JjVfVK5zKh9327pOiOLN6nN/ubDQFnX
9XpcaUBlTF1QiHPTgo1DAAWJRWJhl56MyplNRPYPuUCXdJdxWwCjVs8VagKTL2C/x/k1PuHkmDwA
AcVkCGD6WNktOMXmzStJ0OB4lBaMG0cyUMCFJ6bgX9Rx36k7R6tIJuPNw4gke1DOadK653K2c6Rf
Te0ziHLFqCEls5U+vO6X/RSvHfxo7L0GYwSyVYZBA1lqtDGlzHnh6ZvOJMyI6lfFq5l+d3ppi4wr
+8Ngj9CsnO2P1MNG2avVwVgyUzWRzgMiRgQmqqQfAgdYViWS/0cW1fKlmqMW8ZPEecLBVtbCWVB4
QEhD1Ha3Ph3AGLGyX5lJsm8d8/bS5zv4VHjpwxfMdtNv3o6URB3HSD5UMOaAkBRCth8KVDY9ur59
z1y083zUD0x60JkQkRoTJDVcubochbEjDEp72n2w0N7bJi0iFyj8M3yzjy9K4zxh4tsItUwtuw79
D83djrlsjV03lAaaJMKcIeIKptEjYvLD67Hnrp+wF6wjpNgznjP5gLKRNCQjI+nc4BgGgXRLNAJN
RRGN1pVDQezDvuCNA3cBsCi87OG11EUBsjbCb/9r8mxFFVH38zaD+d24qMtN4EKv6bFw/rHZO+iQ
ZjOnrfvFaC0HLF8zScOku10sSMuMr6l55R2wF2iMHY4nxD91CO0PqsPubbuNiCHohagTsorH84VY
7CHJ+MOeL77stFUeYNfComOoPKq1rfQnveSBDvI4GCAjFAQ/+NiSIqM6FApJ6xlRfN8DMhV7NDkI
M7IQ2617c/8UgdOQ5ohsy5XC0EwxMpFtYo2RQx0L6zlxa1TrqBV1gZ1/oN1ElQdwQoge+gTHyMhH
ckEJqiLpfHcljn6SFkST8C2LB5xaqjr2ywQJOVvt3Bw61MDm9tQnRIT9XMrXHeSLJNoDT8UEOw19
XiOEshXZAHwoeqj7j2AoONNCg3fA/7U8oOQfbvIcAWz7Mj9Hgm4MytTSnOdUp1+yBfqjPD7vaMNf
JXF3OK7ZCaHZjxokjX6CKVVAeiIsFzW2jOR+CVveeSoJgstHz5Wu+1CpXXxywJzili33AgXw2PIT
e3LemcLsbaOEVnhDPFY1/A2HNlyCpTqe4kdrbfjqXXSCU5KyHVwjoh5tft+Ip+9tjba7lzzdtK4v
9NzH/yzadirJpUu2qpTNqVIyjRqjT1lV6Z/dhSHJccAkDxQYJHjbjRLWMRACw39AoXdCVw4F/cVb
dpIWEFfNTlcuXL5VY2xEEA4zlkV2FiPMdAQu4qrJabq5MKIaL/N6f3BsS5k1UsP0P5VSdwlr7UUa
lEfLrKzvCqCjvM3BZJfEMy+E5Cch2WFpSroiImbDg+vLmOzG3rH+LSBVYmoRH6OrO2AHgqdB4zMk
3qnelF2niTDd/T2OOpmZZDLyVHsAmcKVW71s/GFNvHfSjMoqQlWR6buHX8Ct3MqLuIGllUB51D2d
/XeH2E5IQUO8kSGG9wVA0HLspdQVSIkmQI6NO9T+Eb2kWUJVxIwl0OfJbZc1jTNSYTVePI2fDrV5
+b/eEGT3qCqTStRl5F/faLwIldgRWsju6HZTfdScR6noyqXMSQU07lWgTuuI3HONowOlcOYkK+Nn
80ZjWMVw2huSzPwyqEji6TB9hepEQg7YLdN0o249805IDahMfbTnhb/8WKSykx2h3HTLQ//untLb
igLLGPRzsPbSd6i9ucsfMVx8otEmJjLcUieQaNLdv68aUbNIGmXPOZlxtamuZhPvJ/Y1vRVhQ6Vi
NCULv+TEqhh03xwfPMZFMPqa3ollf/PzBLdjUcC7ohSMD8T7t/3LK9k5+aTFUYpH1tokkDjnlbC7
bch034LLV0cGk8y7P4J083PDqOUhpU25WKifemVlu66ZBVhc3QVSgKszvnJ8dsezVNUBmNZbDIhW
n4Nh/6UBFlz0rodAqISl0w9ujIPaDZu8PaNqx4fccbqKSG8eUcMzNeK+uWa4oOtSw1paXAYBzOXb
QMg7Ju0WJ2MNJvsuWHtOX0xR2VcJ1Q8k6175f+VCHw2789VjdJXHljEdqTIIckawNZIjDbup2fHf
+iFqIc5ojMPqHgqtRjt0I/5GoxSjr/KpA7333FTSXaCe6oo1fA0AovT7XWrpppHD1tA2WUpJ/p+z
9yiESZqjS7adRxAOok5OxHw66AXuiabgaFqQZujV2psCQe/4fBHQDt26DBiXqtcuBmw6TKAxTZjl
7Y97S25ZKYTsccw+hv3eyjJPBCvHD7ovVIkFhVVwXW38PeT6ML/3OLhL3LUwY/5YdGUADYh/d2Bi
mXeGmyJjH1A8EMml4yTnMQchVsgZg96050udYovDSFXIPRMff6W0giqd6GantaGTgQBdvg5D82hO
feq1Mxyk2MHxSkpm4FRRrMz9OAOu/6CRcbrJMVin/ghclpL+O18xlc8wTNFMRMBH+8y2VIvZND0l
AYlwW6AgW5ZQ5mTScvL5B4CUSAuprj6H2wqT1FknjQwvL/tD3ADdKFAH6Oa3BXBJEIjnw+rj3nEi
GMs1aGPotY6+x36y5fq0t7W2u2vqfIY1seRKdeUq9mzZE/A1VNwzXESDrBMaAz29vqQg9733L8hk
fhFmR3sCjJJPkj0ocuiljXZhHxOA7KCZ4pVfeRXGTsWRS5aHpmY0sNIwKmA8oItiH4EH/lA51/2L
YArNhZnw75WvFzOS+g3r0x2TKJ0zaAgI+sQJky1Xoy/QhXVbfjIcmXABkb3LrPkTBva537QDr1ku
w0FuV9lOaQfQctzudI7n3q542fuklUpfDJqJI0TO02zDuuEYXAK5/DsDWy6BnWxruPOwJvvLtbow
3J3XW3OLING2syj9ka29DKUDSYnLDR/LJ4K5lt3mpk34WJYYgaH1WDGd2psJMQyJ/qTFbD6bFURH
eX373ErITxsZVdQ2ap9TbzQBP/s9uwkzqLMmvSCTLFkF+plVCRMPhRs1jJVMZaZIruGKnj/1UTlX
Uzmdv5a8HCb37IXDIvZrV8QC5nMA6Xa8RLYZV+Yt64iMjrweL+3tFqXy07uhKzEX2g7olkaGYKBD
PV4URGMIQU7cZkfNmz6o1R8HeX/C5UZvsvjeMUZIo0Uzg5wtQ70IqMl7EMRDQL9Yx9mc9WnW9AqK
Ki3mz/K9KjqUkNxT9MuBjhxKIORe0rpyQ5WhHkH50J1A73j3+UMtnBo+mOnTdcSD5uEfhxe6Ds++
XXmc6KBgMQxUsm9yVKYN8Ysm6CmOkdyrkzXWYbKR7c8R6QweRkf0maf9mVCgvkQmlAc8dvEV8gT8
bKlov9zf+3/7AT6fF6fEiL7rKCJE1VMbNT/L84wetKyO49g7/sPFtNnMfwvbp3sZaKO5w3sUud78
8lqNa4AdxXzQxGNCvQIyjIy6wUJkxBzoE/b52dox+VvQhmLK5TStrC/Kh6NyI4GN51ywzNJPD1Jf
pKCCzpcSiLkQMt4GJNb228ILWggAAOAwdOl3Oe2q0af2eRhEs8NHnGcqsNcHaiYY1fvVYBfMMaJP
Kqt4EY2SfrhHs52lYfRtKJgha38i4nrmJhZehHIFPm42youBX4iF0QLQx14UMyRa2vR06XnNhGeX
/vmvLDAsPJEy1X6cPhSJ52bMgr2KG9O6O6qAX69TD6cBk8LwTtkFMqTLh5i+DNSFHf4smbEhEkUd
EoFkztntv4Fcs5ff9rgxCf0XaFsDgPGw/QOWN7RSL8/3MyL4QDVci746eqXlTXBAhneQFslF3Ixy
iUYZaJAHr2v3UW7hGfWquYEqtza+/2BrvQQHC9g3/MjsHvMKDup8vPNVjDz75kJngjLx/Na14kWL
8SbsEEw+OJJ44QpIUc1F50GNiO2SACnHjTWUiAcnfR9Dco+WTutPh6SEv3HsR695MqyF/FrvQkwQ
elIvSaf4ROZRu9RWQhvLyIdzZnIijeJy05uGTvdaVxYB4umm8PEwzS+dIJbdXY6MwWUxXKVVgywQ
AisGGaDytfusk/31xx4sG4uhhqP+oQgdgxz+4LE5IAzCEHZZotD3kLXqA6pmx0e/FQmW/p706uGE
HLED3Nv9R7VW8e8Tl9ZDXSaS8oN+7Zdp09eNd0hU6T8kXlqfFDPuvWLj6bzAPLknYs5QJCWvgNQF
sQ/4XA+QRLhSDlSXu0H0XdMysilnWQBXb6ve/FhPC31wqNcKYhoGwHCzrEPRm9culCedWAnpwEsy
vHDq26nAlcY3YIF40PXYlHgiM5mhMqzi4u9Xk/BZSiSVK5bycM6/miGFHRREhsM1RjqjJp6dfpjf
0TvQKfIS6qHp5uDMX2qXPuZ8Xir7BqNHqtAODghU+0lG54SmTWr7GzQPVW5KP7qAEAjFO45sJEr2
rlEf2ln1ggy4RUXrtCyQio28Fb0FbzqL/E7l3ktoJ9ulKBIocf5zQaIWqZVJsXGbzykop/5u+DS7
F+73Yh9PQLjMhyyZXOTK0s5P0Vh6xpHenGlbdUEB14k9kcte9X3uCx3tBv4P9ehC14sl9VNQA18t
aNtd/6Ov2buc/OKUnMVM7QbVZqxGyRmpmBrJcuTqQWboMYRLbAMkW9mFVeMaXqnWkfiBN3Mz9fM2
yuJ/m501qsdby0lMCOSS8SnyoOtKHv85YYWOOTpXB6DHUitaLBTsZVB1Xv0wZkyyHIwae6jE5kGH
bDVf4EjS1rv+eOxw+kLfuQ20n1vHs5TmCP0ql4Kdd7CgOLig2oWuAlaH9+oZbaMRWn8jxKcyUC5u
q8AkbhzrBxiKZTIarDZUV4l4k+rmfVF1oqqc8fCku8jB7c81P9MIq0BStUwLzhUer8PzUM+vYtMa
ls/8I+lSzGzKhkXYeZe0yLBSYFg7mIAkuRE/fVS5aNUlLpGS3zL/DzOif8JUbPS74iGdyIJt7LwB
YHAn4eDeuqx4zfh6JdCxZYM2yDWKRoEAQULCZJK2UAzPFX0gZ721Lpy839nBYWjNZCASrhiQuoEi
oppCJVGtNIPgHODN/Cgdk77N/gkDdFBNz2S/2OY4IA1PB/9qAeKXHFHhU1mvxbkLT0G9wi51rMuZ
XEg5I5KhYA3m09OmgHnoYstwmfdeoNP+BLPq6ui2jbpYF/Ph+uI1qLTnz/1TIcJBTsbbyViVeRT3
7Y4en/F/+Pv3Ceq8t6wtcK3KrQic8NVrk/aVt3FrQkBQGTm5iw5eyhyf7qPZ/H44Lo85gsNhM0Aa
EpHFfT8m2qQhFXb8k0eVuwKyDWuhm9tTY55vv6axMlS31XicIK1BXOZi15VXziJ67xeNktqxIBFn
4NiS7Mz7uItUkGPqwm6S8Ee9Z4luNL/5oTqZJgH4AlJoAGE2R8o27qbQAV5TpeGErDyuFdDZGoX3
Cg/0uZ/OjZR36uvdZF/mq5sQ9eB+n9RTaZoQcM6usK7nTWYP/xKVko19st9m2DwF3b2hTeuzeV9U
HtQjjkbuqh22AhXvt5S1+VVa2r6hz3S0+Y9lY3A6qkixY9guI6Qx2K/dJTMWtF7NhPto+QOaKRVY
EhLR3DJPAub+UsUPdk2UwJs6MwsKds53S+tffTsandmuQmSYXCuLR2BKMA68QH+2ZjHP5rKpX599
XelPNIzrrUVck7qH68GSkLKJzCMlf/fx8cAj3v5oeQzRJAV9qe+LZWmWMVoA/zpTJ9uGV/8UwsRd
xp1FFrX47L7FqUWNmn4kLtO5hRY3ihk70tvucmQrF7JrlNCxdA13q14vcdqIpOZ94yEMV/O8yetw
UIL3HlaJHJ8/Z9rpSy4vayLuusb6Bmc6a50K659Vp90Eg6Yvq32BvPQHaHOgUnAyJ2r3/68wHQ94
/ysA3Y1RwN6y9xM45tmmppWjWDc2Xfl6T5xt8dAGDUjN/I6LXOXkddPMvywcEltm2i1m9w5HqW/M
dmeZJq49T2KqzxzefV1yGbzNGxtTSluulmEd+UlMrHXSsgCvE/bBXSdnjAbflcsCVZLZLtaMO0jJ
J1NqUZQSsPE+RPypTDPgd7rcGlMbSDR7hfufiK0zzHCboD00MK2bbrmvalh7dKAPvDkWcouU05MY
LhgMIzYdhyrZnHaMaOI4Mn672FI4BVoQwO0jcx2Jv3fU2BNl7cRTlJL2g0DsyzMv1n1qNsgs2s0e
V7lCoSahC8PZJi1AorLEcKU9qkoCVIAbz8ibeP7vMEQ+6Y1VuWodJO2l53bqBfobYlH5yrFZVZfr
Wfm9Go9zIghoxq/TSoYeVza8bSyLsOSF80x7TAjnCJAQwlb8KmsUy809jlIOSlKK4ByIgGqCw3fP
6vHN+MuSfwg511/vTO7ZwePVz2h6yPp2Wrt652zFqTonOX6DFW3LvERq2kgDMxhYcX4ZJWCIxYRE
fxoAs43y3IT1pMcCCgwwv1oTKUAfEXtZEjiMqJNF3Rl/zINdzzhucPClcMCXHnKpBNS//AHO5jrQ
xEMjEDzr0BGma0i+zyeTGS1y2sqwguCy2L7F8NnVA0vl0LwMgOu6RQDQnIARML8PL6TZVoRJEurB
RyZyBYhuqMXoBflOx7eHhj2bnFnxY40dX9JBkdPaxaE/id6Xa8dKkKX33/5kbI4A5dcnC8VxSQ2V
05GNHMH7SRXPEP11U2zTW2dcu+cmoLWVJuXxpXXAMs8pehPxhFqdqxVzDJADX9DpkIaPpEKp8ua7
SCBIZ8ZlrKMd7g6xIGFLI8R0jkwf5UXp/tRr/BLDN9Jrzy9riVOt9RqyKxYbEa8l8eFmR58QrP3O
pEskOT4qTlNLE8HSHU8/UAqpD0NsxKr1mDhdn4RwQwsYRzvh5lZji8FqCryqGvXZYXwceUEzv6XN
7sKp6iI7THafb39BTcc/4KX9fOJGzxHrAfTYLlIYTIkrOVZyz7msQU2dUEDl7/RiRm7uLPI4fncu
cHJTRhqAThl8LJgqLkDKtLtOH+xyIg3GuJhnZxHCVotuRh/KLCSESJSj0dDN8NULHW6poAWTIcg2
pJyfLKhNLUJnaxJkEmW5a8Y9aSAB1HvzWvcyTX98jnDrpcM8w4VQEL9mcz9yYNdHxbbTnBohAwcT
asK8Vc1u9I/74tIInJgbBLMyIDYDTah/OanBYCfbsPJBevsT3ybpcP+hRm35GCOwA3S8xaTDctjP
JCbZhSBj5cluXI9AUYyPvIaiIpWRTCEXVz1hgKhbNTFeCKAsMjTz0WkH5TL3LTAcXBZeH+RPXRLT
EGDaeiMBdoDgs+kJSy5ivST9J87EJG4mdVrszfrvtIGPjdFN1ehPkrTUx6q6+4qRamtk9F/nF5xV
C/oBNAnSmb9PcAx8oi+/cjrcqR68twGP0nAjWcD6Es7NmjtpLWmwHpbNOYXnGlrqHy4v/Yl1S2pU
VsFROHut/ojPUvsCi5zzAAPwvUWHQVx/FPkP/ydiyRjGIMaRXv1ShkWSronfDN+xmzV/olFXOVLS
6VNZmnzlePPY0+RMwVuDhGmYQmSX5nSzj2XRq3bdqavqfJabSTkeaAmQ5v41BJ0JLtELkoVA5Yzf
De+0yHFBVg++7TAeTLx0iCFqnyBCQPcynJVHdPFvxinnVdClZZ5qK2yOrdHUhA+fDif0iXeLXOVa
GzudPOwVP8GqJyfp9hbgEY+YDRzVAJM/CvZoeRku3x1hR+aJj4JVuNbv/fPcik09dcblceVFO9Rh
szjW49YZ8OpRBQ3lvEZf55eP7WdRJkkNa+2RT5Fjla/TY81NXLNrH0xtpu/ZSym6zcgtpycdBHhz
AmqDqVvm3OaYbIVXzAepbq6P6DR5pYnls1ZipxOfhZf7FVe2OaTmdB2xt1aOm2B4nh1p1ImOGb+3
P7CKkobJTP52IVBi7c8JhhX6ldD9XjJQtP8WPcL9RavxFD+x3zaup/fseg4UOx5hdNQ9r5+pEVfp
6Kuz5jpJsiJw6TRK8yvSwURQLX3VUkZX5HXRQSx8eOcircWrxCMJjEDFJNiWv3CGvZ1482Up8Sfp
TgPZT6p8BDFGGY1IS2n+bv/x+wRcdGMNWqFv5vqLblP9y5FBgJEWGwO7fTl4C5pcodD3SsPoUFxq
b22noG0Ghfr2csgy99z0QqJIIpmxbe7ItJDJ7heuRapinB3NvWz49sZ1VTdymAFT6xu3VbFMD3Qs
eShmHXMIHJVhJVMTpmcR40tGYX1SkiGQdjn/4MPG8LYpxV34crsRwP/HS9OgEi4X7DMtpmVajct7
ajJQBO9sMw9eCg4NEJi/IW28N2vaZVQiL+9b7Bak8v09p6sjgnqR1OlmruuBJKM6+Ne4PTP42uHP
3QvYV8HcB4fY/+A37Cgj+88E/HPMXdhJ1hU5MXJd8S/a1q20aD1iyexllS4RqweY6cil4Vfy6tnR
srDNbEsdMK1TOhIYr4ROExs4qhbaAITDvzEJhamrN3MEaLijKf+r2PmLfR+1xS8nX38oVeTQVfY5
EPRrJM3geXpNcrhkq107IqZXHpWCjh/V219xybIJPPn0zdRUQKsZh0Toc8/i9yE68m9zEWM7RtzK
aFhdggBD/cSpj/xui4uLuzQ0B+ekfBJqIIZuPjWuTWbwuvfLAJDCCFl+N5+x+udmESROf42ckkt4
cHLH0Or/JvT/TRXAxFmwPF9+61QelLo2W4UTAc9pEnPq+8q23akRrpntM/D5ZgeEGdnJf/PGs4o2
clFqPX6GfBOSbKnOyBpJVyGwdz3ScnNZBRlWKF8b4dQXztNzU5xQAGgTF/VYdJN/OiMSGs/cdJ4K
xUOntCXrfJV3KVbdYfGWechCv+TAuSoh89WOVLtDWJ55R38rUTVB6LaJCurIGcs3RBeyoUZnJam9
EBKTObGly4e08MlKXZHAp8hRYLMxLaTwMhmOHuyBFf0zZ8+U8V0k73JhBLwpmo1VmWmTVhHqAPP1
QETrSxxoHW+Wpscg01D9TZaODv+WtOPn8lOrew6pgrV3g6PA6229u9XQXmZ63sDCgYQ9x3ehPI2N
evd1wvFOGu8QNUaZUY6UDTyW6pBloKKp3dlxjLx1EFMRigVrrnv0cRV6MZ//Q1CBz5GLYv5KpQLm
5u0bscRnAMSMBwFKauiI8nQUI2rfHUW+h28alTi1UBZWXC2tb42Wlmq5kwxcxcOPe8KzcAnCck2C
1ol83YlUXEns9YZ6mi9IA8eo5WWjA9ILB0vfpm6LvrDp6nHhzXExvBBY77xh06Pahs4LPAgi0ZQZ
3Z8QX/UDFCfH3+xPX7r33OqsFf56Qfgj7L1W0OScbOVDo6DNv6yfgTm2pbqOWSrSbTar3Fx4mkb1
ACBWEmyJF2DD3GjkloHQqKFeUXKy6VGnSX869sffWiprkUcgI5k3d/dRLW74rGWK211Vv5LVXgkJ
rAFqY7Nl43B5Y0NYcREXorIV5kqqv2LA4HM4YzqLqCRZQ8e53of5GZA1dcfOZdIUIJmCBD1wAlF/
Cid0xm9YKwt8yaHM6rauafCdTUl7klCsQJ7PjM38qaiObAeyoSzabRD2sQA+rWuBuO8O/aGWVLc/
zEhJyfXf5ZyJOpjIWX6WaS5x4vR/BwpJO/ntPeS4FHbEexyCm1yOMPxUoovl7uyWaf+bYaWgJxkO
rVepqNM5g6kmyQm0sunlyLNbPsKr76gZ/cRN6Oq3JQZyuE2+w+6vgLopVt0mctCAIcu1pKSiNRZf
4alSY1fWaLJtafH++ZvRwYglY/Itfy5vGuk7yxggt/kZqyikA46KUSyhE/NQGGhnk2efZZrh9ihW
setJ0AbgfH+QKPLqgp8rVZspSL8IZh7h03gOyFsZfFBa+U59CVl+Tk2/1r4AIY4ZqVsIGVMdMnJU
FjPVmO94w9xve/CweJh8Vihxnp8M0xnjmmuJkfr+9BmR+4j8r7VRVWoYwxgyE5ytlIgholfwH9sd
hUNHnqhii93sUbrXe9ymsmXr+//M9aguikpxH0GN70VIJPG16Eu5rT0hjTXjHTGwxJmoUpQCJ+5m
NwaviwT188djJsCUmatkokFHjR6O0/Z5La9sU1HdEdDryka1otiCdG3JdDlNjZtg1gDNTJsGMz50
+5d6KdutFUDPym4dIHWM61dzbWxQ6CRXXtj8DkdM9uY/dU+aR+d/bU9iVhxwohW69aRM3mSGVbAW
SBe0vN3xq5J6pcU5xGYwpFDClRnMfbxkBd1iHfmyCsGXd5nZ2TtVBqjssprJriFn6guVzkHBSBwh
M3ErU8SwjyA6SjXjHQJevwIWRo0AKPTwKmIJwkVwkptiOowc+f824Ox5fDLzIBz2AYYfLMYqE6SK
iZIH80LbChPeytWqSNR6RzJPIqu5rfJrVWM2Fq4TsE1osmwOQ78f1ddT9h8JzvpwB3kcJ10P9ItG
LOKdrxKFfyqxvd7qinCGjejchi2Uj02jnm4sYP1aQDPCHzD9JOgDZg21GC/TSIdx62+YejqK42Ig
tZBQVnviBv9b+YOEImc4wwvOh6Ynb4GbAAdwQaO9IKp9uJIyrHKj1IzXhlWULZtJH5nxBfzynKD/
ZDR8HlpWM0QnpF5wWW+oQ07dADcMd41uGvo0CPl2jlSJRgJvJLUyQOiMELq35MyqGYbZiilvwtHT
B7ZnXiA60YJ/kiyiEEjJCCx+ODIB1pSqYXjLjYq2/hg1aaYre6sglmH63T1Mpx9/Awf6npZqsyTb
tKsyf836BPP3QH/NmNDySQaps9UwyBUQCa3tY99XZ5ZE8OOHqGLW92ATdh6wj1UjlWoEl7qd5Zcr
F7rTSku5XJAsdluXL59EyqTen70MUi63IPXl++ZBJODK6osjXLmRJbHd9IO9aZEjBsHLtq5+g4EW
zDQXRuIJNt7QenbJErvdpWC4A4vVT3RWHUyOU3vG0UWen2s4RQzdf4UKMHXPamnoXwCeMhOL1EQt
RjCCttbuTN9QRIe7Yzc57NYv874d2rrLKWNjA+7mfneUDiOCgBNAYcOKoY14/H99/yWp43lgdIRp
MGRVuz4/2oy4ix8aW0bh75RrgcXne1V8S5vWD5QzC0yYfOeQj0BNZWyzyHAMhscfhL07N2TduY03
Q4CejFjB2PW9SK/rf9nDetA67iiXL7bJqY8Tj9XDo5evcRQ4DvKSknQVxWaGtGsFFCmXptpSJV/D
YhyIqoW/KmcfuovjsiP7ODQfyJ7EpUraAWOEAzb9I3bqq2HZ4nMe7/anoEdNy8a8Y4KV36S4E39f
U2zbkzlBaR9IIFauSfptoSIMt1rRS2E+vmLMdPx2BvAtC8IkRMkdZjdnV2b+iYHs6EnELkdnB/c7
helHUHGVbG4dWeBfQAU+XXZlDXZcVAU6FZBNNVzuXPCrFkUho66nTyXfeZbuRjhnHMu0ah044vp9
ugsQL4PekngB8PCtF93sorfUT4c/C2Q4h4wHcIGv/66Hsg3e4izlogzBiWJa35LpkMYgCr4FnP+0
8x/knXjNi1w4kGd6b8MYk0qO/gsy6pnO0zZ6QRFXOz0bfAnDlMWilsag355FVLvJ3e9TXsEXiVju
bCx2O+DEa4D6/VZuc3V/Zi4cBwtiC3fRMVVMfmMFFsJsCvVnwTAyofJyHU21gPLaiLUqYDeVgazf
8ERcvo7yWCZiLXqrKmU8ZvD5ExEJhXOYAsEF4yOCwTeAT2M0MAHqik4fsQkzOwrwSKVax5brgRSV
jAmcYcmLJcooCOfHGuRJK9wOs8VUtVWRKZJROeWexH8Nzbyr8wK2xIYod8XiwZlIbgTg3sr66cZB
GbrQS0x7+znSSulfz1CgogEPGKEcOfYyHzQ1KI2zTpCt02mTA8XqecRI/mSWZw1MLstEYzg27Z9+
MRNm8xG0LK/ty1ue82eF8Yuu6J/htTCu7KHJ3sKKFJkCAL1dqYc12dupvhYPhJPbLj2E0cb1qnRA
gOl6IGkcGxCvCNtn2Am/178e5Xr2OVyS9LYIPBbSIzCwY2ikiDWRSPTaLfdQdlj0HZuHUQdE7A+y
o2pkHK2/jbEskSzOyEbOclC8kvV6DeqPmItvH0FnnzX/IyeZyUFV4527T/bMXkCWX+rB4WD8iHwf
jdRNPwbZ7ZhnxZRBG9L1gqTN+2hcs4EVudhWC5Jn2LFbPWqPnMurE5Gu/LVGVJ0CwUKSAAriM8qe
odWdP0yVPRZeMXPQJex870G9sXJ8MgukBRKTrf/nOGCMuCEg72zrGC5TYzQ8xLdSmfgfuKW7w9ok
ag9MP7oXdh7zCGu5XpjQ/ErgobacmojnC/V4JC7I+D41eeADsxi2fFvfEz5I0mSxt2vhYX5rgpYt
YoisugJMZ7oMi5kk24Hb8RDgxU1FAMkyAOBsasJZl+A/fUcfFutkXYHgHMCuTytp8R0GSs6EMB2b
5JweWKA+keW2dr69ar1f7tL7Kt+YkntWWtx52HO9ZJPzKqQZYj5Z6RaID3dFEx3JdoB3LOhebEnQ
xg3Qj1pGqeOE1DO6fiu9Orl2aZlLO2swhYd8Pb+azDer2xaArAb7pHQrn8+w9QrGRqDDdp6CiSPQ
MgVN9J4YIkCxZdKr8ngQ/AeBgPJ26h9ofKl0OC/5TCImFMucJLtbIlQaE7u79VUXI8we7Ixwls+B
FOozs3VZCxWMDgMyVKokmjwMbNgd2xFso/2n3GmcIOHXe+/OBogOgPfxNP9itvAxGpB0JHpfr+s7
6Yo8m7uGrRJ+3/egrJrtxka0rkBKy/ACtz0FenX9LjPhpOnVupF0gtGRDH60DwtezxlKkjAZS5nB
OiF+nqS4NNMeIWZPn8d3AMISwojflJEdYBLNLDgDQgVEFnrP//mSnj7Ri6m2J99QiVOy+uVnMkcd
qJJH1dwBSDzqFnf8YKrjCEM+rALLTxn2DnaR8/+HrE+ztbLzUM/Fc64rJP6pk1LHTKMIy7T+D+I7
PJJ+8HGKo4Jblr5a5DW09Y/eiFImISd9pvj0s87Qo4+clfIcEyJepObyDLjm341LovJjSFp+W33B
gxGfzvV9fTArIVvI7dzUYtncm61KREBJpXN9l7v8q5dOOm2oEfr8+wlZccDqarDpItgvXhUOUFui
lZDWvPUOwvq8GY7ropyfcEnvqWcIiFVDC+MnyBqqipSn3ZRBT2KgtYX7ayXdW2V0BujNsfs5/2eC
3tipZ0HvpjA/Jdf6tnLPv1a+1r5emyprZpUHFt2pHTukbmaYO8l54RDU8Ebxkv6BzYzlh5af+kyA
UT96UKa12byKL2TMo2j/euTzHbwxFsHsNZyAFEdPUNPCH8J5Q2Feq0D0IeJ0YSMuuLt9vrSkuDMC
tJpWWzYPGmHVqU+esKubgPBeSf267p+uRkDVZQxIHlATx/igh37/K/mrNMMdt4BnlvF83xTKqkxQ
EUOGpiAVWTbHTiK2UtC6fOZKrSWfuNC4B3PGKU2T0pgWiE4ppXMxfJ7DBM/2023u3QiMPlp/NTJb
sk04NRaL7cerNFPP2uKC0LhtoJ8a0A0YvxKI360+DjoI2MagK4VdrR8AOnF5OkMj8i5ZUO2oB/42
9Fb6VhNIhxPw43twPrQPjTVryNoKTpGmHnrnHyEfH9wl1q8zSkD5umq3oxAQqH65qcQCymJ0FNoc
7dYGjgmmg30AdH8XH5PXrlRPp90BMB2YCmwSY/m2B4pv5S0D7dSjw+WS8I31isikBMeI85irIk0b
5rLUbFabKG8F/T9GBmEt6mMK4/e/KNcAGaR9jkxLD1zL43QfXfXyHSgLxvfhz1EU/OM79lhK4YQE
MNkC3UZDbC/v1ZduMFtYeOJrIrYKqC9ZGe+fD1I84E0yWeM13as640k4KuoceFLjBmATKtbW05Nv
8qNKSQg8gjXuMWMd6r7oQSrtBQ6Fer+hEzOazN0RAaKRerlpmXvYRZM9mURNKoC/PquninmwOymy
EHTGx5dK/tjOkCoUOmS9j6zotBsmZC+fvGJhGhgDc2LiGsGMHykzc96DYwF51tn6iA+9alEeZKtU
KXFFOR77b4zm43KXNID1TNgu5nIaPWFzXwBS780m2VSAxI3Ntef/T+zYR+Q+GWMBbGfZpMtNBMaT
Mk3jtDYmi6eIt1YKr00ZXCW5pc/A39JM4DQhXPLx/9RkX1fzJhcpcUq84ecz74uMJGhbjrNcgm6B
5xWWkMcmuwbSfQ0fbJRhLFhqL8jXcy1IllpFM7HlGMrJQopQbjJtBYUKtfkttEPsj/L5SCSsNWdC
tcZZWcqcNOm0kdUS+CB23KcpvQ1Eivvz9vSTJuf9wRpHw/7Ve6hg9kHb8ail1Zydo0yPTppq5NRV
c4XO94dZtQMTfE4stR/IMH6mAHSwnlKjPblnImfcNTayEytNOdtwJbb6LayMRBcyPXVZfvKgbdyf
c0zbF6ni0mYtFHPZMwwi752uyR+uzD8tKBJIyz/MdD9gV2aKCd3pRAVvUZCZpKugNiwseNYP+JdF
WUY1t2Ih6inAE93/CUtV3Zs6dsRvz9cttvBfDrZBElzJTPZeAAeSCDDoiGnH2r8NF36IFsH7ZZSq
RXnqn+SEsSw/ZmXI4Hc783G1yVC5/I9TjYkHiO+QG0yp+EC0dIIo/qDDRoJzN3PA9mTlvIdoeafx
QJNAGoHuv2oYSwm7IwsD7KRMzCd3Evb9smkryj/LJ1DTLXYLQcgFQN6gIv/lqVYGOHT/i/sq8Ws7
KTp/vXTafdhIiFVoxlzUar0YMn9YaJcp+7OVDWAMPrls9zFAy6NXwQzJWcjfgd2OhVXGuVPNOQIn
Ua7TGEWgIHt/YK0+OI3S1qOFttT3gjR0KbAgtuljGMIUQ/ChMYTX7uiH+8iWTzcd3ui1ZL5Jath8
JtcadcRxUYl+8UD/elAOueiu53aN3Iqkba/yxd1uS844G4TYQfFOBRluvYmqh705oQBQdCVrcmz2
Byx9RzI9QXQl251IwYHm1R2Z0QSQdnGkOcghWW6UMXimV1iU2ilq6NaWl3sJDquSYwULtoD8hWvB
2asT6+Vu4x3xDOs4nr03ZbjplNP8Hu9afnX7mBU5CR8O8Ptm0J+K6o9+ZgwcONXEVj2DFAaHBrWG
zdlXBRudEBokUgF1BsYCU3qzEUmCkpaiEH6YGxXTimCzjB41o3jpYlYPiupOdrPgZvk9suIkiRwb
ZHJeSY6rN4RtnQu10gtMKKIjDd7cREwsLppd+XFg5oPRkZYCe2tRxuV7ERx28xrEhG6vlMrqx71E
yIpAIBerzHtPbeWhgpa7+URIsY2vFzL9tGwFk+92VB+4bNKFUoZZUYVtbCJmSem1e0I+iUiJmG+S
QL+yUrgKokNozvqI3/zEEmdNetFolDq2G74O71WvcO6cXDUOvgQKWAvgQtk9rRWpn/zWW6u7WoQ3
o3rf1caOc5oWF+WJHTsHYPvQUBqtwWIygdNs3gDaiGyrRZeYEwdHr8MjLFYYjjX4qd24JGnGdaAX
Io+xGuxuTdOlNLYQke0IMYRa3ziTqFTGxM3ybWB35nRokxqFJq0rXC3Mqd11mifY2bcaVw2X0pnw
l88eRRVuqsuw/coME3A1f5sO8/acNRjttPR4lJs/m4dZmy9COHwHBWFzrKXHXdhqyrQDAdPffWv5
06SFBF86lfVr3f8WEWjKS4/nz95HyUNSJn1sD8g4YCzvJvPJFghKbZZjeKLCQumMBIf4yRyS3XLC
dpjAEM6qew9VKu19A7kXKY6Lmb096bCc4WFHTlAJ7rkGYewAbtd+qTtb4JWeBY9hChG1VxDYDgbi
n4SVSRbdWHHMBzgQ7YsfawGpWMQMW5GP3mTDPn7ganmRMTyAWPv4qh8/zfBOgiO1hibOAN4UecFU
iq95Sr5NjjTHtC5GCg0fkd+6lp3uhBJCGWhJijp5RA/RUesMU+6oV+WKMLAVnIi9TmN8jcbSwvFA
JPEBZL55MtILPZkysgU5KPrziQvos9wpRU1zSz66EMFL/BvWrMyjDlhQHyJuhtMpd+4suoe5yslO
U6Jrl5PGcVMcyazcEZYLJjRLExBGi+x46ON93U8aWDldc+WXyDi/s2HH/p1K/OSgb0RMrHmDGAHi
TCQ9/50DqMJGbnYFZ+EfBNbUeIDYaZH9LBwaBktAUHyBts9iFJpyNcP2yqCGDeDozJhvFWBDuGV8
p3sKOjj5aJqnX4XC1GK6fsTe4vCNO+i13QXFNseGUifg+805SG+jHmS6ZW6fIMWqrctkNDHfcJTK
0NcLAmUTZ65YmY+imOhCo984Tbz8twvhpNKJM3fV4QkalEVdaFSofKNGbCth7CPOovwxDYcxFkZi
3uWAki2A511PPvA+RdVFILXuqVE0EB6wsY6D+eedl/VFOvs2fEIyGT8hNhOXHwmPN5MGRR6OvZF0
LkiEFYwlBjOUDB652x1iy9rvytL4yhJ4R9izhtt2UeGpRsanxRIrnA/HxT9IIFd+YyKJeQXfIp9Q
YNMjsAsFSMrzwdmsMrkRDiLxLMCbBtjqS1XfktDPMAVPELpFyVt6hOWV6bOrDox/h8z09MYQMB+/
xik5yDOj6jauH3FN8W6WyeobZ8fIH9M2H8b+U1WXsmBToO/Gt6fjWI3xiePp/Nf9+PpcOs4/229S
TIrsqFH/ex50drX96nI57OFMNhEumBqoh3aucztXkkQ4y4HxV4iSKi1P+nE2d4i44DDF0Z60GDt1
7e5XbPnqt0jYkUsQKJivbMsZJPG2p5u3q/eydQObI05xWLLJW9/gTE7fwqHxRuIQVCrnFxHmXQXn
piNQ8fY6dbJpNbwfRlGzprJTPuKfZ64hyvUOaRaB39im/k2ev+ThLI3/HdxiAwTuQtI9aeqzOWoL
FuhsxnsYt/+9IvcEEaGpjYyrVi09gSOZGUCbMffO0hfGZfkix56oAIKyuSpV4Jg6N3emS7kpy+xX
0e4bjE93MkEI/TNDxqTUV/HnLtehfEdXuaCAiAwOL5b8XuypKAJTIRIcsH7Z0GkjFNd6lhPObVNy
XPoaaHnBB0o9AjV/Xb+G1MZdiBVjyYQBse3EHk6Ldd7KhJyZu9+LVtq5V4DxxgGgkfS5s7BF3JzG
paMXZvp6VtcF8DXIyipzsYjh/AfxBwrdJY+wa38liBZbifCeu87Ny1kDwkEw+nZloliwo+RwAiRa
8aLFwOxOExZfxrs4NIBkVXmfDrjFWawCaFVaC8ae+HvXlghEIIHHvRpRvimnMQA73CAm70K9Z0dU
EdYgIyrARxewl7lsm9AFyz+KHoQ1bdl0e6N+kQ+gFI4SZqRnKiz86qyCpHq98bgRhs+Kd5wPVuQ0
oTV1LzGRdYSXweTfjsHdrOJc5uTgcftkg3s6Mn6EM4dmKUCiUnk7gntGwePc8IP4hZjEBi03GpNa
NF887AlCa6Qq3NSr8Fu+Jmql18UlMrMGuoTLsAkfx5ztdg8IPZ1ne1YUS/DSf7M1cs7qmy8EY9fn
185FGcppYJExn70HILMvNYQayf324dDn2NZouTdJMTQiTsxY807VTgWqGJDaZU7vcGk0E7HVhxkp
gVvQwjWGPsmdzP0f+481IDNk6JTn7QYd6Z3dRdksHTi39PHYdEHm8uVWSOjDDe9oAkS6j5UzjIof
Z2JYSB3yGkKbpHAGJ16W6TqpSYiEeGJX31/Q+tgh0vAdoTsdWHatLX0iZuIh41MVtpiqHCKRHkse
4m7QdzwMHAPRU9o8h28a/aWdrkbAAb9D3Hcid7ee59qK+scVkgtPU6J/4RemFnRNdo7ymyRksTHd
H5rPC/sG4ArX9Ami3mmwbNdgZZhJhbPVv4vqeU6755XwrNKYTn5mqrFV5mrIc3YYFxO+IrqiZfnH
TTDjxH85tfZIYqKPLF1yohvVjKl7jdAQ+qSPLyDkq2ySobDTkt3ue+o6c30kQ5MTW3gYeWyPvZYI
9NJ0C00zcy2GXX8dMViu4551TbCDm2ow67OETCLHaZm9YQUus+Z1CDnd5on7qi86RDe+V3Tl9HSI
jGPpz2ayUemThaxD4HFHMhvaikdcQMWaRMJZX6c6ftVkjGViYeqaOsFVO2y+G2gtXwvD5K2PIcEg
lGWJyfC0egc+bKrxsltW1WQO7jIXZ2kJkKFMABHwVXy2YbXxcYORhMglEzIWaEq71GTTQiiKr/5k
Kv8WussRE12lwc91AjKotf6FDo6fX22Gn3mzeEOF/3BL2OdcdtWcRfLB2idSQPC+3pyVj2u3efKp
LNbr2rsVtOFMHYOZq7xN2WNlzmiZc2Rxt1gpBask65F86K7RQqfkq4zsmNtwo1jhtm21+FJdGNDB
SJsV+nmygVXxIv2OpvHdTRrCtXVkhsrwL4F9vEE7FadBLVMcj2LFtQyPLau4uqbCvPLu9dXyZ1ah
PGF5knh4FWn2/DeThDrnKyJ6jwEclfcF9+23nnLrmaxO11oGNgEfpk5RzRp5L1+u6YyeV1d61SL4
lExeIe+fVJ39DtUwTwLLYG+OWGJTmh7HxJjIPFVlqXW/36qKD+QFVEZdBRkU9jQ1+J5+NTim/udY
QEj4GggCuT83Yzd7JkrGpCqN1czwBseY5DfumSg4SnLScysJu2KdLQa2TkJCsejnRPhTsxTv67o1
FmjoCLUKDhqrfkJj7fdUgEAscC50uX5iNgjYPORx4RHOPT2p1jaCMGEagSIumyJXwSIGhzqiNVqd
5RnCddszptRBuqGFE4bsgOrEKl2RkGm0ROpHyBoRwY98DxICJ4jVWSQmpQFq6BzBQaO73dsLpDrU
ETFx4TZaJCsYfvslWq0cmEB3ujHyALdt7wJm21MnNouZyg+oG1ImoXWFelsh3T9ORjXRH1r9FGsy
i9HC7is0VncHvP4IoehngeNxXW1AnVEIW5qi+MwkxtKhQh2k+TnSVGychPVIVPJRWaMjtvxQ0iSi
zFXdzC6YbJfM8JXJY2UC6JiKr4Tb3Rk6uDm2zi/22o2V//TzyRvljQXqiyjZ8gMXsfKSqogbEIgW
qDkKCDIpWMjUExbnfZtDIdnjv1ixWLWcRSPj1P4cTH58zpKJQhMnBlCYzXVwV7YTlqlOJ1nhCo9j
elanKncLlrSvsshfkybAyKT79K3fauQFwTzNj9dwmBAqNjvWU7EH6Ib17ibekLFA0sHL/8eS27LO
OyWL0DE1yol8B5hHMuvI028C0uD4pi5OoYUP6sWi1BG2HGnhahoDcqJ0/WJ828JXoIjBK5RTsg72
j+BQQYLCxDRViVX+KLsPaO7b46hgeItDXuM8M/Ua1JLJP9xVJameXIHbx5HPYwJIHoR+S6eF/dOQ
qovnSeJro7hfCZUlE72MDmaIZMswdlsIx1HEVHPA2CZRPPM/rk4HsL44onG5zqrbWOSKhRm7pmMQ
BNiBpbGtvfisjvM3tcjHA3ssCwv6l4pF94SMrNUXCY9S8EuG+5GUjTAh/E+k1MFM7/CmMfzZ461J
4XX8ifhYvRGPgyYbmcpTe3doZWYHN64+khnOhaK+usDIykDL0rymr8ka4AeyhFNwo1eWiaXxEQFr
KfH6ZTbxAqj6/6gS8reKMccUKpu4g8vZp+OQS4S0j3WS6xYSpbH5/oh8iJbq8gpCYfmdSI/SPtzW
0d9KD0WemxlIXC9sdblY6h653mwvZ7oFcFy+EWtnJAu34u3jcDlLXKyyWrT16aFexe0TjxpThw8V
4SEGIDxnvoJB4Kt5RrBfZ7Ggdeh8xFhlMIDPXcux8GnE10xKI7uyVtDK10CwsG9yFvKPCBn4e6Hk
QTx3zD+CAJS8+B28lM7vzm9K9q8VJs7KrSsVijNm+6/vLO46yFbYYSiyXRROU7cbLb6pbbmu7EYa
e3zg1vzK13xzc+nV/FBjxB9JHXvXYUYU1jhPmkzZj8wFfIKHDOT+PcxBey8db7tOYeDvb6yQ+XX7
U9rWPYeTSnp/CQiNmmb5xU1puJ5wKnIUAVFx6dFheDY2OKA1fRRWo0lBeRB8Eqcxwlc4pi8YTuu8
W/u29BmJIM875JmpT+Z0Z24I90rAf972UD9H9dGzAqiCKL5m5yia5ZEvPC0C+2STd7uVK3uMZksb
AzY0XKdwobGLRusboPwiWDywJ9v+erMgR7VoMBJYFq6TVIBCKu5skykdqYCmiMyV1BpxIUAsxsMS
tN3bWBR2zJFpB/TqA8iI+F0N3EuLuDGMwmcHjd1NOpVJ1VnL99uxqRqzfvlC6nqJKT1Y92fZnkFf
aV8hS5+TrEg17fBPMF/xQyNwc0AW09zwa5h9kYim21M3WB1sIGmQVKyd4ZkvHt5PQqTuQOFsHQXy
bEcdhq5IsttJoyt3BTmmur4bmwYCjRUgUGOiS9KOQaRhHbLoa7dMpCSofYGwP7DqB0JzVBNfgmNN
p7Gp9FN4+QSOzLlvh/8fe47XVdmJeOeUzAc4oP7kPDFRLd67DPYSeLMZUKy86qiImmyzT1iE/jTd
Mi6disFqkzDkZnCS0M/gOefJEfnIVxVMQxuv07zH5hOMnYE7rX6skDnexONeNnKULK8Sh+9BVPDf
lqbrnSz0zLtFAefKyHkrpBr7nDsgvpupm8gIXx2h+Nj2YsgDDL0ffUBtcBI+WY56GKnMxfzkp4/O
4/7WL6RZcsJa/CfkmGz1A2QQkS+jy24ZZ2alzwPqM9vI1E3XU+bbaQWGRnYW0ArjlZLI6bhXMzEu
ns9pm7x21MY9uiS9DOocHl6S1/W4cSnkA7GOCFnhKG5ThI8AA3QwIcaH3iZZ3YoQZ+mytAzcnkYM
nW8GopzPPllrNRZTc+EHiVcBqETRWFVpbgIXImGqgQWIU9U58NUuRHYxXLnvTYiI8oTqwsn2H++F
leyhzzTak4Dh2tl8F1MhRY97KllqsaQ1512H3AV0p+PmCXeLQAX9egDXaVqA6UNxJxuJxJ9u63Mf
1dGFTQ2BrZL9V/RuHN/r9cEbkoFQlSWuyDw0h3AKLIdUsIHZYLJOiY/f5pI5a8MoHoo6D33CRX6Y
HjYmto0MulPvrwJUdKVVNt+/LLrlZBRvoq7ve8neHEmI7OU+TBvxF1oDZKj1w0ggAVYWOoE8ZfnA
3bYSSj+ldOLmwsuBpGe9fzGec2rakEnwhaUMQ8JMu9d25Alk9bDfMxhCSM4gVvgqeDbvxHvenZ8z
u7+s81/m7Z1FJjSFl6QUP8EfSgnjOoL7o3CGwrjhoma+YVD/nbr0n83WHBXSrV4N2zT8Ryd6Z4bM
I4fa00mf0mnZwMhrhZwn/udmE5ne8GgNP6rNw6XphzqIp9pyAJQoABsctUoMPUe+t0Ze7VwWsf0i
dWDi6Qc0ybFf8nbRvXPi9o9JoC5OIUdZVXASZj5majAqoKV2fJ4bJlKAUUkMt1Tt9QqA3G8JJxO3
UBJb01e8uKalsSvhOR1WhUov9au001N8B1NkR3nbFIU5uYxBG4bpkzHhN/ZUUgE5wA1kYHbsbGQt
gjPhrcuBjstBKOxo4BU+JJylJI7wjcjz7+CHw1X3HQx7A0JYvPrbBATpIa0xG5/+Rl7cN2W+KsWF
bh8pQR/TqWuEZEiWvAjMJvM7UgcVUzeoWWQmcqAYEcssvQw6DxyngkiG/vJWGFD05YqeGQwO5PXv
wwOhmSw3w6kX2pidaejtcz8TtVaNIO+MSg4GPUParFbLWbfFgqRXicSBKvFnwtLKtil0SgIK/iOZ
FIIZ32yU7vD1wdS2Qr9JaARrYnGjIBPbdY9WrnznFKBUzpoVP9zZWtHvyOtQLb0SwNJV7eVKeUf+
dSxizPn2GRjx13/zHMp3itZ6CqXLYHmT39Q96tJH/nkDONZOvx8fv6dpwWDUN/Lo3MiXnyjYx1Cy
ZB0r8iQxWpfSWKHrkTWf2Zecz3mG3s1DoiTkYcqFq50Gdvq6DAN7t4ZJi7dDxvHHhirMCsv2lYPK
0s42QsWsEfhJVzUGqoHuG6zwCv0P8zDrKBj8br1tFXchA4XzNWicX5FO6oeA2RepfkVsp1oLeGKv
GRnDdXncGhea7k9jTRoTHB5DwoiixkTjiXk6viwHT3gdtFyowvAKjdBCse2/IE8vonHwpEmN7U4s
iyXmKGH08o9+AlRLMOl2M6xOJk18GKkZ59o2nDCNOUXpMmfuNFtiABJuecX6rnfpWJVOydwdXvPx
Qh6jPnroTwXLJBIu3ixfO69qaXpmTmXEjhEIcspR/yX3/XcBAAfDnig7Sq6gtaDSAYHwnFmnUlEZ
FwdmhoPr9M0i8gckzvlUbEg7iugRZQc3CWin8hKQurzSN4Ct+p1/EHIT1BK8QRwjFvbj6KiyF2rN
Oi9K3pks+KwNVM54Z99WN+svjlUDpmrRfK7oU8Uy7pKb0BHy01zo0GuMc58Wz661JUy9MNrU+04j
lcAfQopzL2Q/YifaIMhNo9vpnGADEYmpoxRic4UaHH1/T9i96YKz/4TcfiIoZUqQssDnlhsbCEP5
VM1DMxjglkDKoa4XsCUe7yVogA+ORqbMREPo3FK14MVRtiV7LXXVJEy1taAeWd3bBJ/6I1ZyMIyg
pTkO4C8nT+rhPo8w0bdWXlOlE1NL0LkCKjO3Q5H0NJHlkRJt0m/YsqSjjxP56Z2FduowpzH2IuQr
Tv/laLV2JdgEFaqed1UF9++WyUBa45TAxCvt4KmEiKLBojhmgPbW9IXsiq0LqeHUYGwYW0S96duT
ivsZhQVCaYpI1ZCMQJifYjR4E8Z60b04aKybFJS+DDfjb+tWGswS3fO48z11QJwFYYdissMDlocV
JAVE+rLD5J+XKgsYTmbOVgec31L+In3CslBQgCbgSF+hNiLIqtCFe8shVIV+HzZerNqCj022ChqB
J8mN8pQq4jKqN8QYVOGPBMehZTJWgCch1izTgk/mfMEfR9vWuZuInS6QHr7QSYIQguz8CYfeNU7m
TuOGbsIzabLCa+afy0/Yqh7CE7hRVfzePqBTK/i+I9eFbTg08jNZNWqiDgoyChPwr8D56ofqEYYU
P1IeiCcX8O7Pe5zpVhV1wTXbyXHjX0A5BOsIX/0iAsipC8/TXKqX0ddHU1mDyEIaNWksPgh+Vfut
e/Q/GY4Fb4Ac/49fVB/mRhLzykOu0ZhZBxS4XEg050fmjNt+H7dG0pY+WpmjENjesTCXIp+/mBwe
PVIVo9y5M4RG0Wehs0gUX1ibABPncOrNIira+WaMdDZ31S+dJPVtOB3T1DjHwjClJgQeK5BaGfp4
xSOtr4LeKtW3QLxYOIfFi44ASfJurRV/tfijsyVTo080JLtFik49oqKEdZuPrBANjGMZG4nHQLaH
8lKgkTtPP+R+F3uRtmMd/8jEPrFY49jpPt/RNCsHT+uJo6VSKy1bcCIZbKx2LLdDKtfJ1A3rh6gO
mahOC6xML2ddJ9t95PC0GsUvCHDCp87chaCvmU8x/L82sJRQxcJheiOOtVRvrgLTHrbUGW8zc/hn
32vM30rGMYtDJCKRMmZnbU+yBtTOxw5NArK1dAKTWRDVEPenm75UdH5RL86NKYZxISFsMFPb+lB8
/WrW5E0abdLcEZ54jH8Hxky30Q+k8xsRqBQMDy048OAsbxOpZ8Zqz1PgvpCUuZqhMnbPGL3Z+ZWK
sckeKjCx2nsuySkVNJBzXf6QvM3AErXNAvvKyCiQP9ji+daXhBQRmNAuSL/SPEkM411ZcCvYf6ur
9Cq2a7Dl9WnRXKEJEwxM+ELHfa2eyPVkfnFoXdjgrhnyZNW/FzmgzPLjOgzryRBa5ghyDWSf9b1i
JcmDi6alRlVpzoIdl3bauPaXweCEIddKkD+XgI7jQJTL40JOIwTEsewo8k7FAVw647e8BsGPdg6t
v7dqF+mXav+03pkV+gxI62LelMgQCx27uFYLuBNpwmA9pOqFuaWEJe0+mcUbbqdt8285sTS0VkFN
FV4fkT/539913kl6amF9cZPuI8fg8b7S+EFy0/40r14c8JMJnmv8u+Vz68wSDOXLAM1TNa+5+Wtw
Mds+K13JanKrgOBY51AM3Pp1ZUblyn/wAyL1lAlCxEv6kaFgBFPBKmB+JobHgK9ccCAFzoHGzrzV
50tDy5hKgGHpf5ouz4xkV1WDPUNDJcw7sRaQe2boWol14vyD1CuhuGKc7tRpstyJ6xDzrQ5SOiV2
nz8I06eC9/kzQTkwoxYxxYRYXm8DILmbGXLpwGMDApbxw1N0jPIMZISAQ0ImjQq0uUJLoTS2WJNS
3ToOlQsO3a6lgpnE+jQTe4hPSamHeakmSQqnEunn+0Rn1NRCX69sR8SS9gwSs4yEiROrlDcw2UW1
lNM+nVb0apW0WPnG489DVaL5seZryLlnoxYuSSoM0Y0GfNdWZcFaFM9VYzPQWQjZ7YJa0ljBHbZO
uK53/e8y8jyNiQ1n4tkqo3Aw5vLSaWxNy7AOUxdTaM7Jz3S7DcW4lBZ9GVHXNIOwv5/oQE+cS+nP
gC34Lsv8/IAwoRyAKVnEMgaCN3n5OvuqG6bwAe8R9lgiHq+ybWkefDrgSG/j0cMhgYijTRaunJsg
DkbfV3dcO4Y6BcKJhebrdrszKbV3VdQUSYEzLFNuw/47W0bA1HE7QdRvrHKh4uce3kfMV1K9V+pz
LS98zmn8GiWM/0yn8aVSat0ZeU8AtjlQc0bWo3GEeaZiVdd2WzVM6OUP8nMhMY66DDQRH64n8mTi
JdwCUbbYgM4nmiZTaUEZ4JGaJNTQL0Da2tIubuC+YmR9T7jcNRVfkUafDffV7i62Zh3HParHtumK
ShylcfQUADkxW7p8qsDGo1lAIeNhIdjrwoV1g8Z1gqiW/oToCbkjwHlNEHdAk2D3ZS/4BUV3HrOh
ICz+tMxTLy9opctnVqG4MmpM0xltj2FpdrTAO6iCij5MwuJRzIqdNfD8HSgP6zHNtCjk/kLIE3rC
9l0kqYbRRJcvg4XC9T8fK+Nyy/e1t4QMMV3vwc+nzVcrOd8+kI622e4vVN/Y+khiKn9v0zO/d5/E
EtLzfapYTm0A0KBmYlGDTGZ0o6XdO39NwnlodzWkaq7SapDwq7VaoA/B1wru9X6sPVa2D4Xjgkw3
hJII/1aLJlTcC2ed3iXx5DFlkpr/n19+zpvDC/p46dgNYgnvtT6a7vTgEoHilese+0+a9JyyOV2O
B9GsqyRj8zHKHNoi2czvRJyT5f2IaPtmC/cAxZTn7j6qQg36yRvUDPxn2OML+DtEhHGnAG+gNWyv
ZqKr5Krs5tqyaM/1r3UhvgbSO744ONdHK7e7V1kw5fVULMxNITowIM7a4FD0pO7sYo/Ba9yPMk22
/jo3I7plGfBf3H8F4xCS8I0TgX5ZHKlQUVYvpcRjVl31toJe76cfFnLX+1Xoq4r1beq/3pkwIlxi
RxONWIRTL8Fyks51y/qQeyhaWKVfW56Uq+iP0PNhU4N9BtX73D2iC/DxgE7Z3qTBvWbOvLoS3ahJ
w02UFg0j2CtixWzzxD7iww8GUM9rh3nNPLtaUj7+YSHCnpNFdnrzqJbxKzBStTm2BFiEGd75vOKe
xh14pzuk6A/FX1Is+j3/7hSXhj6KsRvyK4Od7Ux3XrgnwWzlZmBkjVB9pAMlUmI5EyJDwH39A2+o
4boR2OHDRChK4dUbR/XOh72U4VkFJEDSEapmqB0Mb55EzMGQeJ5dI+vmQ2dPCLqaFneenfWA0d9z
39sl0DtXuxxngu82U2TEtP1Fu4GLyXN/B5ZjTPkCxkAHu1qxkp1wQW3+HcOLXAHy2md8MqBpo9hj
7REmhI24HwTidSMowuNBNuOPwpfCXe+iPJX9usqk2GHSmubKu+G1P0i3An+t5ArDayoi4RCy1Una
lhcx0zKPz6fs3F7jZFZQTDh35cVrZGLNQF8MtW+DLX3mV9FykWOn66dJTKx0e8G1aLs5Cj6AJR96
D/pM93smHjQACJfvtCNpCFMsh2zhhInp1VuAGADLeumQSuCboSucqGGbG2Eo7bSdhXUjfIl7tHc1
140N1vldPnH6Q+/g0cePvXg/8Jmuj2D+7KvRVPH8U2O0bcrs+MMBfGmWO1JKJzomDs/uc3+pkRke
ugLSZs/juZaaY2qk+28mmH62Fzo1sdhFKNhQtNPI50lAktefOCjhwZvaEEXp0ZC5wSAzYCTir4e1
GOteT+6MGy2NcSJ7GZLSnbsRBVDVDXnUmyEQMPfYPqU/9ltdY3OA7sFosa8UgMJW+J2dTrOZv2xV
S6HWAEQns0ZYPUZGNiuWArlwfqnbcPsn1FQqsEGM/Uslmd69wMNt8SCHDq4wA0gVzpQVfaJf5HAU
wsVwooGBBieVahyxqfwzmFPlaUb3jljBnB6FJRAknjtodOgzVCY0aW3A2+sSZMNegfIS92B6ZBBX
1zjROuPBzAo+3jcrz+T8cPOwwbs9dRDk4UFo/GbPTZd4Xu+eSCmLn3slQT/rCCU9ModS9MqkiUJS
HjgZSOVbRO9vgYLTedoEO3woXWWpnUgdAMTbuA4JPtPGXhRMFykS3jdediQVKIbwy5dGf79mEMJN
Rkf9szoZoQzlXuYAjEKAFIq8xg6wi4VFRGX5rGddBxIMUj0DmLu2+4gyxDVFaCkPEFcZBMT2DN77
V1MJoP4IpYc61URu3fVDSOz4xwk/0ybReXOxjCt9XFqWwUIxqr1NJkATF2MOe5gVD/kxilMNxlOg
BHGcGzkte9HRV3V9dkR9mdWeuUJlTwcwvuHnTpj3jhaYCwSzKCsM9O+yBGbm6e57yDrjz+2SbLX2
mia2gfjqxUSxFWPkRUyLDAhlubpuINLr8iW9rfPPpJ5kUa1hsmMNSzyanFY59Z2L5aYuDJrM8Rab
GE2dXSn64DlF0kgjAF89oiTQP2idtAF7Ij17GX2EQABIPHayQwlTBer4Goa9X2TmDU8na+YS6kv6
BKUpNrhOUosurKDMbg++VLwV/f7VFazQX6MByWbfKnyOIa1sn5CdtIo9U8nDclqoc+BUvLq1TzGS
YnY1/9zBA7CFISGekTCQE7XR0XYrXx0IVcs8EWQLvpVhJgiPES12rHlWPtteXIgM0mzFG03R834X
khHCYZS0W1sfiE+uZ/gm2B0HkkOpYDZPMgAuqlg0/ga0qXwdF1E80DjeMJNQnIC18cQq5xYx5TiA
HE09e4ujrnRiC8vjiwMSFSkUry3xqTkgE0AIrnWZkHvpK7kXuAFBdj72Q5Ltk3s77yaowIQJkN7X
3JZ2wdO2xdh8wgnA7TxDMkwS/BpT6LUO3OGxjgOiGuTbogIBqno6E24h09LGqAZGhNr2yzVQSVar
f2pQaXOIjDFGnoarOhjivhw+KUj+mt7Nr4bPLNDtMr2Ft3LcKvtPj9a8Is1eONKDUz7SchrkLmCx
NCEa5dUX9VD9Z1Az3T4l2zS2tbdoUsZcnFhTbNCqnHmopj7cDB+43vUI74aMMHlQjse3tU2CjJXK
QKO4Hb97RMqzDLBUOKAo7X+Xy4MeFeYxjHFs2OsH5cB7Yf6u74wfFTFE+hCwUk3wXNuTMgdhidD7
nOIeRQeIpjHO3ClPfcEynabjzqvudsVQKUdJuLxZwz5hdeorRD6r/vl35oElgW8DSvymvNwGcyQ/
K8461PoTA/sceGyUD8srZbiWq44JzvGPz8+WQcTgxlIKvGj6khuTOtgQXG9xtXVz6E+F/A/dk++W
BM8Bbsy6XClA59dvQO1Xr6ZYQaIQ9LJSuAjraKYKnpOZVk7qiYsh5Hr60U6AQgO7GAQSBbOB79py
BYVbjTk6Tv+ap5xTfc8LtwexJgEXIJj9NqCiEvX0Ggf3ZT0eo/LvT+iYMVFq7oATfEqSuXMox1eJ
Eh50gGNI7NPv+Tsa7RWboqtrcPGVltkbwkETIEHM7awbH4I3JVC5J1yqQsjJLbG29sd0KLdgyqn0
WHad/kfqHOISaMNffMhHiTHpDsFhdp7a1vEcpo/qVu8FLwECoOt+wrXmnfyalo0wmGZYcodAWSLG
5VKducJFzGN8UJFITZB2WfunX5eK/G5facGmCLEFVYv+0OUznUJxUz4jgQlGvBFGeymjkX1u6Mnu
T3Hhb9dNFsQzVprGmZVkGba+QWxvClJopLFnUWyM1aIJHAoApXUwDmxKoNc7irJLzxwhdr1kB6zm
RgOFpb5T5MihpmH3NUT2h1ri8EZD00mRMEm1ITuIEa2emmDQwWrAr08P3Vtoz6Tj8h2+TwCPWjXg
ZcvYgfLBmvaxtGEkoOId8Lb5ZGPGTRXQDXom8hc1s9bRUsMuyGCmCNDHlTuvK84KOa24EPkaRP9z
onEqxUocsUSlyNmX/YC7VIk3yjSvrbxFNW3AEDI1jpTWBTMFDR7ljYENY31mYeFsTjxvQlleFANx
MzplWfLjZFi43SB0Fw7Xviw7hV8Vk4eLXamsW6tMCC/XdkwPlzRZOm6RQPt7wXcgK+O8lcY/54o9
rSFyyNyCSTOtDDIEJX8HGi4z8i47uNVapipeE8bfRZUbyfYcQ90KQY2WGQr9wythh2YBbo2RaTEO
yetxBVIyBlCQN58mMKYmg/0fhCnVK9R4G1tExO6os87FDF5RGKBzyAXbSA1plO9aIXnrwdi9YTr+
BqZEVZBrC1/Xw5R3barF6BGdxwOflDRhc8ng0sIvUEswCiP5HaRHYvwueciV679U37LI2oGNnXxe
VQ9c4KmKeS5wFmgXYSxznkUMVy3vqPua6i1z+AjpoQS5glda8vn/pWqF+QEyA92g1K9AVgbWz7oi
oWMNnD6GqPHkzs9L1JzcVKC8K0epqItFhszbpf1q43WVLtoPaLC+1GnwsXExJbb791TMrcivTwyr
e6Z1LKQkN2J/dbyt9WcQ9Q0aqUVEURwolB/pytsVrvV6X6dhklCTIX2/ZwZBAyBAC8kTrA4oAmzg
m1xGlpF8RtyreYr0npPJXn1Hpw/jTZDlYkQyNNdgJKQE8VXTQ+9AZv8mnr/WF+DmkSvTr6D3mPGP
Sp2ewJbB6l11IdWOw1YyY8QNPtqbhCU46qXbX3nyHgzLHVZ0sb1gQfEBTigIpvN7AFfLrThhJyT4
mAjSMRNgjWwjTqjVP7dO85qhUMPerIDcHZYE+RomUDegLkcWQKC74a3U5Ds7qO0CFPGmGwzhfsbp
pt5HtcijqajFV+6J79M/S2wlp2rjKhkLk7ZFBJxm+nodrLEOuZaEUDoOKDNjMEmu+akno07nsIeU
uDOZopvJDhKDmZRbnrA/vqqVE0ZvSichjf6nhwpSTB57m9t1L17Pphie9lZR9c0kLp648sgz5gXw
SIW+WoeVWUrAYxMaaiV1fo3XQ6pFFq0ale7w8hBkyq/AF0Sg2CQPyJTaGYZoSW+n4n9q6ffDO3Gi
o012fvMaKU05k7+ERau5B1GsIYdmjJS+gtIQL8d21GHe1pI6pA9ImzTpCyP5f7Dq3fong7gsUI0p
72pV3HtY/67gvpRVzgl1OoFXBvtR1xsWm8U/JjIIUR1FNFt6fbKLja1iUCvLo5dWoyH5WIpsilGs
YC4W2/RY5p3iEtCi2sftzkABBVL9WbDQe+ugxL7UPLoa/wf/pmAZqmTL2+BNuT8EP8tBv79HCUaT
pOXeel6nlbP+wSeHTtbcw78t+AmzDcPyWSmBFJGW9T4L5zU3xV9ywEOaAvaN9dSw442xMPAcwGoT
hm7BnoKgNDRUlhWeDANSiMGr11+pPuSYKHK+bUy6W0Jkkx3UZh8mV/gOsWPPS6GjMjbAf27h1tQI
d9m332yhiflGv6tpaU7qyQTJ/Q00XIXf74GzVhuU0fX0AmkXD2C98cLN7uni0z/9+PnRpc3WqsXb
Y4EeqVbd+whmm5njVfYNuz6Rh2RJKnW5NXaWLNFoH9H6QPQGNzL5x8mSPZcIQTdXasEoH1TGTJf5
NBvlpvIh+/bJ4ffuPFd9mSKwl3la3/WF7H71PU4ApVEzXq0gzdlP69rlMwbqjwR2hgnFFqPbrrrG
1qCmHE+N90JAdiBvuM/B9bqRNJoOWnXBGGlt+8wB5bTUPFQd7akfdMLJRY+cTqcZIgAgXuMBfucZ
nSAm4tGOAA0EcAmXPA4H+lnaKyhkaMoQJOuIqFLJTIwhuxDToXaIHYLBDvEQkCEeSjoGVIRXQfy4
GJLGdI/RyyybanTpdj8Zt6dNeuvoh6pCtE6GcpmzAEtAn9E3ArtRvfBOurEW6Xeh+2xKSXYbLBIM
ZEJzyqEhItFMKP2YZLvtuQ/qI5DAn7q2jEAcwVzEpkaIFy7MS1UU8CDzea5P+oVkThHinx0jYYKd
JFitBP3B2+dKupC5kF3F5s4SAZtJfYoLb0uAqi07HSJBSdFxpm/8gfvOeixMv4YAWDQ2xnd9XzNC
sC7V3tXMn9NZ09LGj+hvnHDuh3UlZZe/JQoTu4j/9FKW1bjdsOzC5HW9Y/IO3kifEBabU4R8l1GK
XelrtuahE25KGzYeRtHmJTBS8CGtRnhkjKoycCSCchkWC9qgQR7Ie3A5W2sIOC3mEM79ToTkJE1W
heSOwQf1g8LeQnSzHFZqL/tZ7Liq6C2G6fjRvFivNc0vTWMopSz0KvgD5g+HoSNKPM3o6Gwbe1G1
AwnkQg1omnHGBZP/mFZT5chSibvk9PUzlTQIbKlkgMxPUB1iyVIG74LlE6th7UfW994WktIXvekh
48BsYWqh2W7VgGEtc04j+K/3757DTXoPoHCM5VMImlf8m+T/vXkmYs3ecLDJgW8I80gDC11Z7wHL
QGCaDGyA0KVRhcKVbDG/qSmexQE/UZG21TajO+aZ4E5jvvA8yfkwxNXTAiqAvA/ce4NSLECJ0eUn
YBalitv6L6mq7eVejJ/tzCKyGejcaNfhx7ZODUlswhcIBZ+XYl29CVFde0T5KzeyMZrbijNqPulb
MLWKPmwJerkeosL9iKIY3jfQPoB1kUb3bNNbswxY4i26pt2rwPbfMGZtdK0DRm0MDN07/Ep39h9U
Xhile91Mzwa9IalVR8+u1edE+8ziwp7LDMs6Ezr8yjyr9ILim5VtDIVLKEyAOXUODxDuFm7eJKTX
UN+Y1y0xKWBYRS1S1y5YxzQBTcuUqCyZYXyO5dEsJRLB8ZFWaBfAujWlbrs4qKfGlI8q30zEX2lS
cGhH/OlX0lOdN35U3wJrMe+RYWQqb6w54R+uIsqbrfpvzCkW1P4f0bb6SOA3WCkY1kI8PvR5H4vK
WtPiosopNsx7MyMJJErkpnFXqSwPYnNcyNo405ZfDHLNAsjm95k62shmN6NVHt11hvhSK8CLs5Fm
rbr2f0EuxQe7KUAsP8iLaqAnrjBJ3ea7J/Pkxva7gcY5UtrK9sts1K74Md2TF+CATTDyBEGDstOp
m8awiNDEpfgoVKRyUBN/RlmnMXllIqYQr5gCl0FxHvvBf1zugKWn5mBTjE9L0qxnWxirOKnRQQcU
G1VAu5OvgnzPUNLnXMSfqGlSs6JaRF5itv/kfxPrcN2jv3Py0WpNjKAEpa+2CGCf8DiqGYIxLyA8
p0s3BSrcY+uidDBxdG55Eo3JU1liAYKecqXUbteYLH6e+poKzh6lSuKMx5Z1xM25wNw20vqIDwTx
vG6PdT+qfHeUTT85xukgSuIVTrhMBnxieAsK3BFwj5uYZnBvL7dSA/GdG7+23HLoODxVhY6fMvo2
41TRLIg0eeEuaAIIx0I1lG2BMIpq0avShRyos5zGywbkAqKsdL+XoWoGdR898f8nEr9SvD50hQyI
e5SlbVdTqW2awQq7ccLHMfliLvjRWfxMRNvaa05uQiTcrQXr1NFqKJMSofV7yFA6S9hA3U6F1GHX
YbkzmD+vMPAD7OLSkc8FxJ68rc033rHyxgLshZTLQztjGcqv/s8mbBe4fLBJp+d0BTsepHyUqNIm
+J0lRVbb0O3wRJQQNyTGMvrgOVQGnnOiAc3ZAeJ5MgqwuHhNEYlATLolR0wAtHqBgvg7Rmz+31x5
YFVAWDhx+H31UotagIreZPEqMsKLREO+amGeJzWoMKXNo8b0kkkuAkFMLNq/UJpQOq8tYgKvZfDU
aFG89tTm2J8nnd0tLOrQgA4nf2f1yHpYQq6ezpzt52OtIblIUPkRXoU2xyAp2HrtEboqJ0UlJY/K
HqBnKyuc8wbK5txfSU27jO6cMp+p/5S9WqzWNlvt4RVV2J8r2CEPHMDNvoCocxoxiouYKSM1kweR
PCswXU+7VKhHX8oy4sxIFvJftAMjselLMSB7pkcf5oE0Y7WoHnsll6Pr1s8rLVG/6FI7a3urLU9P
u+IGUw46lLRTHycUETZVIIKY76oRPCQVkyf+LFdDjuEmgz1659qqbp0eHAm7lwBfUa84zskUMLIp
F0hl5nc+Bj1VGsUcfM8APuuvklTxF2PfIYFY6NcnQjulENA8MieM2OaC6w3HVDNTBTOVPVT/e/MW
o46xh+xX2E0LlH38gWwfeu1dSARHrnc2H7+pPejEJB4r82bpghV7Luhcn4FeBEo92OIAzWLli7KA
7W5QDxQ7MpvJIy/JRW4AWD0jGPLY931H5e+eSxf4Tq2l++rdv11RhA5qoNrnoys1tCigPOIQnu6y
7mex+hq1ub1sSUpm6VBvdM2C81L8F24t/GdfEh6pwg777Qj+jrxcmsKsEwl8dU5Yxt69rsRRyUV0
7ON2bbBvnlkRSTBC3/50A29HxRY0QPH7CFvVFkaAMflje23ZsNihQs+yX02jtOaoA5W1PPTydIEe
dAoYDliy6eZ9o3+OCtmv9ag9M2VUx+lX/R6nisP/wUrE7sEG9WZ7oz6sh+p7PSv+j7ICStATmDyQ
H7DVxl/hSkIBSAUTihtWZ9Cv8Yn4DBtUPu9GM+ntSsxXqHL1kPwPlwxp2DyJcWFBjuy4KtlmzYx5
NN+nMIcjJYgI0YhC6RsPIjkqBP0EDTGElcznGPIY1rF6Ijt6RaGFZ10YaIPvBaNsA0fSBmwTfQS3
BUfedyoeira9riIjysVSj9VR0KQ3L6OvPUHByJvEY96gKewRucePtJyx8Oh+SF3kdm9fKYQ3vFis
zsKtexPFVxVP/aTaKPague1pNNEHNuri4JrSV8ks0pqOvfgSqwssyQEBn2f7dplwskebcg5rtnzE
1Qji8461/6NRjljZSuxhXMQrkAZX1J19uv8k2rmas0SFdYNeLA409ZhMMCGV2FqaUupxibUCAvd8
dxFV0DcgbVpqJlVCl3QqNsziKgcjoTGicB6alRMxlj5o+t8ttCvOmpnZnHAHq4s6B0FUyX2Dz2ZE
eH/8ReMbrotwYa0fWvBbtr3/Q/UVePKHF9j3QVeTJoIdsjcWgSXVBANfsgmwOQMUSHWm6+Ojr/uV
6TGRr2rVaMYeVK1nzlWn9XE4mcFnnsOYVgKJqfUuRL51I3ZvMMF5ZxFyOKj/Gc3hhj2u3Lof6inK
kx9px06c0nZM9AW3S2xve4PzoE98yYbHDi9Rgu1QsQ4oHn5pm/RS7aSAySLoTd9bWKl8msOQTVkK
B2rmiLgKBidR//KEHuIOsPUpLjVHCMjtgOeUtNuxQ26udzjToB0C9aFH4j/uD+gJAH64m0z5kKcK
vfkd9oafkuqyTh9NpQ36rOiMr/jyrErLDJAIRIuG/Bo9jxjDH869LjxdSceyO6X8XdKJSg74kJ3j
ij+f80S4tVwHQt+j3lRgzCQBzt46iN6dWONCoP+VhSs9/xNUDhIsp2h3fLgKsDvnpJwo8FH7q1tM
Izxk8cslAIuAsSvMbTSxyHF+ijNal//fUX834eFAW32KtFMSsxBHJfeWQJs4iL1XUKIWH9Kdv9bF
Cea3kue8XwqYlEOfDySiYIGXgkM0KrX1AgfgA1GZzFaRDIFxSpqQkAt5ByuB5PrKIia1TCerZjeE
vVhDh8rSMStGxXfN0qWjvvlq/4a+GwLRzr3CiF4jeRt5UX7jiCqjRsbm6T/HiFbN8gcxRx+ng817
p2ieug5UrrpyQWN4g+Zg7ulfWrCYgpXuDstb+/jic0ypR8LsAaSY+91vcCm3B80fQgzOZe9lCOBc
swxSzN1t13nroQyBD+M6u3rgywXestIgrkqNLHeLn1RFfGE1LIkHI6kdw+kVbPIqmFeTKaimQah7
enLuh726DGeKuSz6mRJ0VjgrAIKVPeYTiOmzxV+RdZoeGBOmuE3YVWaDkA4XCKeTfpA9GMpYaBMf
wjODTj8V5QJ1kYbz0ZsA7mSEA7yCd8ANiqBip2nJLbBWLmxcOUs57qwJlR0rBPdo7cWQb7CxoVwl
a8wa5EsC4Qr0/MJMZ+6mCnBaG9zCvYTCm9c7zdZ54NjmyC4qBFaGsHGnotDnlWwigoW17S091Q7I
0G4QdMa7bVeEUtzcdrIO80OwaBzGNEYZxBxiKEGaYbeoz5UoR5R2IEL0KEltNjdn1pKwLhBHHpJT
sOqxsCOwBOjBtLEPzSLgBaLGuExPBylVplJOynZYG3yIiZOhskTStrcoI6EiNXLSaacKewUBPeuF
KrVxaHrxFvsSGnL8OZC4UsNilwJKOUtFJ3dcarKZCL6FxKA1sjEK6nQsOPUUEtWHYW/UpIWlhtPf
X/hbOqZvcRzVWHf3hvADZX8jeYX+S/88u+SnwGZoxNUfLb94mTMNkDCZU9TX1PfGMm1zh8D5/uOw
ubTX4V+Lvq89LldJPWqutdgSXfl1ccpOzDYVcZ8OnjSrbGTlpIRgH13YDVPyu6Quz8GJaJc83JTD
j3O6hAOan/tASzPVe/JXIrLD1FKvP8U5QP8UUBPNUr7V5ElXxZBKxg7vjGWfJdQl8Lzn/z1MGVjs
DZ793ThF6vJ+bIPE9VR4RPxiT1p4fFtVpjMwP4Uby6xMW65h1TkUwtIwl9frbVkx6d38vdjDlkfC
dUXgBzoc724sA+dp6UCYtTx8Fi5POxpq/C+YJ41WqhT7pYTSbdAncVWvTmNNGnzJbcw/m9P5Hp9K
pI1d/gVTbWv6E/ACMnd4ax8XyVHB6l7LbC1Bh7CQcUNrYZPJxax/UCFFXtPBd3d+r1tYqf9mv3P8
+ChktZvTlmdi7+xQnfNr7hr4O30tAfMd2epJu0UV3jUhnKTmiHfe9bMBYKWZHOMuWQHu6yacvdFQ
vDJVSXPAQbtgmWYqGG0TfgKW09flON/zWVLdBG3EauLsYXx0kcjfjp4H+kaEC+QpyJCU6Z6YV8n2
37WcY7QA4KkdJMoHJnyxvkqDQ+DVfJhKkl8/3J5z7aqlskUqrQNR3dtbcRHat7yMIl/XPCIn6K9a
kBBxFISa/zEtO4Y6WyMb7AZuPr0LRtv3GCPviiVAegAtsqy+y0pn8DmpBh6IEK4S1x1m53pf0cFx
cEeO1uviZPu55r/ruwT8taqSx7nr/NOOvWORgP9ZecvP0T1H8LrbkIrg6whkiCVzSHAmT79H28++
Pj/WDBInBc1v2wL5zgg3MRJDzvZq3IFL/hRoGRW0jlQHtNkb1Gd+kLAs5nxXRnwDnVA17oOIq+ey
+Cwdn36eyqTOCsUJshazkUtpSKnDloVoPGxs1TewGQsmiPpv1qNpLIWYjmel3oVWF0GzcgB8CHbE
t6cm4a9Rk74Yar9f1pwF2Jj1AGv6RUbRaJCwJ9qCZ4rXFYdHhMnVOedMPujwZIlmwHRJbSwiIrs0
t4M/j+Qutd2B2FOykT1p3zeZcn8xK5i6cXk5cL1jheLAno9ZtgG3cLfuF1+SttpiJzIFaZwv8Xb4
w/Cs7tyrgZeSB24yorx3OFEc3v8V9OrHOHzA5UyM3U+pBh0i7h7CbvAx5SwyT2oADreptG1Jf7Ro
YRBuXyNKZWiGUNXg7ecwemIP/+wTdJIb6eGSAAJcOJLdMQZdu1z526DiUlrkegclPwM63a7LpfBv
LROaxwH31eW2X9G1+/nbiOOCF/lWYdLZIdCMBofRPFjdLsV4QPzxB2UgMEfOi7WYWEqLsWJV474I
odAslVSKnug0FnZWOBQjGxIdvb4twvsLwmRfcpsG8QjjMYmAXqvH124oAn+sbFJt2/fNcPTRNxxw
q3b2PROH3P5C5EHmNcyPW4uodbhRMd7Kwkno6HkHSH6BBXDhDYauM4x4AGZtnOSVrz5aBfenEK6W
prGku6Gsb0qEKg+ioIh15aB1iqGxSs/IT2Ewc9V0Zny2fZjVCBu7uqa3vl5fMVHrf+zA5GGojGSz
i4hvfpj5koGvExLad7/BewqjaBXi2WuRjMXa2Tvx01oCCck+WRHJSTlvd7xKXtEV2Swbjyw4umq8
y2AciN1CCFzLTWAc4aCKLA2Y/euHqg1Qa9rJdxQYp7iZ+O9L7UZXhRX3Y2kzeSPp5V4Z8NmMqch5
BCtDs/eg2IQnwI8ORF6pPVdMRk8k0IYtfCuyVehfHDMV5mmMeeSaEyl9u3QxaCFHYlhLstw+0u0d
uBk+gXKXD4pnpV8dNFYw7ev0IFO0BI3PsUC0FVMfBiAGmc9C6cBUy6+NLC5FLHSG5Qxu6CI3QzmZ
7gOrJgoeUmTbqli+fk0glzVW+Rf35CDLKNKVyy6ddGSpx+QWzcKY51i0laeSblX+uO4FaiQuDPRY
3goqY+tZYl/swTVSvAYoWKKxSUMnF6EFgJuDvCQiofpRxsqQQxGiuP6w93atmdCk3BZP9BiyLwFl
vVg+KLQpAes+rywbKXQBWLwcGNiK8c0fRtqpQFuEblkbrxmOedb+PdLnwV0PDr7w0+4STKX1wtPm
Fmvs0V403xrYVVJD6QfFfXooj6I8toHkNOU8jgmF03I5/Hcn/Ll4ykXtp0nH9T5S+FJ9rn2l24DQ
gs1mrgZn46LfBjYD/pLDA/0ZQjcAHPmSv4MxBD4yJH97yLrxdVP92P3ZJ7vtQ0SK5mbkZHVHje2A
Ic+L314J5YYnBVfGpEvRSXyTyVzLQuo1Bu+pUQZfSwzLzaImKaiDvcpPZNQCMENh8cyGg5qdkMsu
Qg9gaMJvxlCAdS4pXN3eAF18TxiKseFXD3i2sQ/h5/vdu6MqRU+xaJNy0T9QJEzWUMhNLz+jCqcl
P15WSgS1vz4+e0InHLOr4XL2ckd5hQl9LWO/dMI+AW3zwUE6djaXTuWku6a+ktL8LKKsKBB7nxHp
wPyC7OhYZbJyHbhaN4zDpyqFLJOEhKPA2zIe0T81atdYT0KFjcOH43J0uiWlgVLc6e8Hs4siLRdf
p/HI9wnaLGfQQ6+1H7PukfOxl5catK+esp7IWJl5jGfWS41jVWnTM1aJI6/zN8MmsyywLxQatEcZ
6JJhb6WP927ExtpyKlkTk0E2dAeUmu1vPR/pRnTxL0q/cw/Wylo4eZ0NOEqdx9O+AHkvt3N2t3q1
IA+6AzAmqB1xubnUG6YCDHk7u7Sp2qkSHFzOgyN8ea4Znjvv3LY10Mx8otRKOKsY1RKbvHb5Z7Jl
fyaLJrDYr7RUNFwis9gheosOvKsd8hlCCJrUUvbUOg3Rghtb+ZiV1VNxSg3waGI0RALPXjWnGik0
cvCUv+7P0nrOgIHzdfV7k9eI+hx+VxOcAQmOKxvIYOAkmuAzOZaLQzkcNeRO2Vyjv0ovbJG1zL+6
ChuWr8CS0BbZd4kJPmtD8CqodHV74EbMdJNK3M5WAzFJHVzYyQgAQpDcKkMwMaSy0o6UZqpOcVVI
ZRSDGeRlFlQSwjSPRzVPr1CA+/0J5/0G9LaJzBoKi8csbcD+Tams/oS5UWDYyVMA7BcKB7yk3VP5
GYwwOph5euyGmTjMdSctArCdlOOd6hgbV5i8lGVEKkQLVB4cEiLao8H86dVuKo0YjWOCmRTxdVkH
csSVUdHpv3hqnqTx12sVjoSzDjNFagtEUjQn6pAps+pSQQIcLKRb63icQah0FfOpsqvEJ1iWn7q7
v+Xr8/rrKJxU4GkOYp6QrZLRMiddXAxRrTsY4b3mhGsos54v7vaRd/uDh3fFb/XcLBWfHmnwy9V2
cnepipYHn1QF1BMh+XU0N54xnAlUouOiY6W91wu6LFbNerhYKg0/aD2iCDgZokMejEh+rJs8wgCA
JxpgMc/sknTDmtP0+cW13xWOg+qYGxSvNNpJRZ41aZfDnotPKZFHK59T38eQRnFEr44lzixZ1fqc
gmqJtwIAIORFFgreFHkCpMdWZ5UFYCX0lyBC1wckFcDI0v1KV1EbDoRyFOp/91oZpnVBSHGgw2aI
2fyLYfAZNbHdFCgVhDkDn7oPXhaSQK3KNzqcEWqApeB4lY8P46HMNruBQ/misbEVoyNtVP/4B30K
xxH+wUmz/jXEis5liGODO51sD3/+9fUOnlT/Z2XbUthcMqcR79M7ET6gswHKkXdrrknUw8vqEgiD
6621XnRq9OoqUOxsYkjQopL2WUcg681TunHXQwFnkEgVVExPfAtrxJf591y/swHYePxMlsfNEgmp
G9Hb2vsazN6xRqa8KSKU4heFllJQwyUJnTscelP5eySUvq9x0NOf1G19VFEdROH9M7A4woUw0xtS
7fCdHpCgpQE8YKZMQKHjT49ZIaL5AZ2rk2cbOBWouQgdNYyjIH1iXTCkHbC0b8hJQBnYW4ByuPUj
DBaAhChkQtgH+mVbuPeOBJR4WDdlen3ItRYismB/5em/1832kUj0Wlxsv9YMmX6U4Ij8Vru5/LDI
p5g4EI+JXyAB4v+4GFYIWc7GqaoHfolKsweLBffqc1wcerKY9kwRtxWSmLP0c3ka1mxtX58DrQHo
u0iuorz+/syry2Rjto7wMTOuP2PGI/709ztDdXMXZglbatM/ykhpvjbJiJ6VV2kgU5cn3joox0HF
loEWIm5Ml5PTfy5yCRgpHstoql+aG41iZpA1/1sNUZQVbCu+598ECqY7YLYh+I/3a8BDAgi1w7FC
lEcXUeHxz0k+cpzyVZQ+2zZKCVduviQT81vfoF/OfU7EftkLqgeWbK7To3jfdCZHg3qAIGik3EpH
4vXTslhgdh/fjdoF4X7qo4nFXN8sXeTD4eDulWiD4vWHeK3ZKBkH92FQF15LYNMlGJnfQpwQc0t4
QTnxz0jwk5IgwlDyH34VSptkcgyXWYwI4ItxWGpFBwDbs3hP/ySViC/5vRWA5uMdyOeZVtJeIQRb
HWZ1FDxJSVHZsD9LkBnf5Vom8AH80Fx7IKsR6EcQa3jEWqv7IfEYMqHVSu2c1Ti6XCf7wXaBhw/N
uO18HeDhPIRfRSeP7svU2gW0bfnFUs+KJ7zPkl5JARUUZvt3Q3MROsbf9jxTihW9Ys79pqG4h6NJ
Kh6l3B84hBAUkMJOh4R3a2XybyN6rg7aEAtVWYAigWGx7FF6wo9YzG+V8RKUD0IiomTQTvQ6UXTY
HJ4/M/SNypTYfUQ+pcir8p1+w2zwfNINDEogXV8WLE6iqcCy/ZcU9KwAEbK49oSuxFwInKAHsJpA
A9bp0uPr2yMtUvpzluH8LeVBNo4tW2lGXGM8GLOCgEHiQ+YZGdWJ65+dExfvdDO/VBY95syJFpNz
RCwpG0o9ft/vsen/JI1OMJlHeU1h8V60Z13uewTSrUEQF1X8DJ4xNPQtbYgxOgi/oMDEFs4Kv+9Z
rfx296HZZw89V/9kf4HD1jKWuCJZmZlJxZfYb0wOj9mVcuTk9UwwMaODkiXrK2OPaH1LfDiexk01
/AQIeypz1avXo/Bsbk1Z0P7AiDRZqfmHr8noco6kMGjqxRafQ+RO1lFP70kfF7mYRFZJv7Ts9yI3
woMU4o0ZbJ7vJsnP3E7TwJF9Od20mTwF1EsRWs2hUgXvlquhIJfCpI0sf9Nr5I79/3djhjH2m4W1
wp8CbCEIlk5D8o8jDy86FrgiOhn5BTO/UOwyV7fG0chnuftsc/fgw+/TNAeNAg9LpUga9jQ4RCrP
zayFYq5jVr6CQrV3uJ3VqGvBbfg/0js0sr6C9W2ohuoEOznYr6YfuruEgaNZ+69Hv1hby2W0yJrk
RHfPSo2ppUzImSUF4yM4io/I8iQPVQz9GmwxtppT/Ggovy21FgzJ4j8xM9FWI07asyoXrcgQEa81
ZCNb8ejsn7WlvRN8f1aNaMty489UTd0L6kgBeT/k4GC4OEvynkQFPa+bZm830kfRq6OFGgjJAghX
M4+/6m91PdxEGctSf4byOEjmgJUnMwQ77CuXwBZPLDirdTe5CHuM7AiS2gvtIauFc41474JtWoMr
32ywYhkAZC9LZPpgYXinKjtVqQsPBPFst6FECQRGRk68FHqPpH8xuAWCASkv/e7193tz2AY5/YVF
dm/waNAacPWLL8nuAWakPd1uxfA57hZmE30mlJkT9Rf3C2sJOlANzVvq1O29KBTVdHTOGzjdbR3d
/VJxZ5texGyTTYmPYoAGU22prXpTMbteOsBe7zbvhDA0VX9Beo0sJ1INxK1hrt474B1Mud1wa6+m
521qpT4b7jjlJ63Kyojri91euDCf4tKKDYkyhDFiaCKxRIwJlbRwkceR8EQWdozqYPLlKPgBgBE9
uAwgBOt9KdIaqATv6FAZkxDPvd86Ic8bUSKFSQdCU4D1z2fkxpyNPPhP2Niwk91Fc5y2dobgZluW
OgXGIPMKs2VoBvN/R1sGCiTvnN3Q9jAwqiWHPD+D4XRJexU72aV087HYY9d2aVWZXJtlrvQjwZuD
mTR2trntY+3ihxb/YReet0ekPexZ/mu1Pdq8UFwtDDVNsBQGhiHztbl3atkwdY/CAQPI4Fs/Vufw
yjFNNAzrEV5Bb2e9bYdttn9v8jcoWD/YYVEQbJkdcD8+M20YlzjToQn1G+rCSaBD5AjxgDPYX0ML
MbA+ByMHh6660/lQmRo1GkxN1uuCrWBQ5nyAxqcxlByPdaJit4OEG7AsCXmRaiwBcvgNGCi31XZU
hE3lri5RBHKProGUILTr/cT9hrjlebUuWsG5SLHkyr09YVGcNS+jdxe4yJ+pPVuLUgjhO39tVEdJ
40efsHOjj72yHFJ6k57NF+5CWsdzsy7zZmNCzrUwMltx8q8j/ObVNLaIBv/uxivrKvBX6BomPJ4a
izbrkDc6sftB258gTUtHBcpg3CBfyEodfl0JOgJDgYbcX25Sc6B82kXnwzsYLPiWmQqozV+jgS6t
bAYC34mV7uUonGtBPA0ocWIr/dDjytSMmloPaud+P9Sa0clypA8Pkeq12hb21cNU3VKYv3LsCbYX
Ay79zRohqXUfk6uta5M81Lk5JxyXIStTCp11mh1qma70VeYpt5ThtIXJjlhfCWriAuDZnZCuJFnt
pSKoGXwS2YERM8ZcFaiux3IYUeyxxiAHcwbqCgTE4/p7tiRg+XhH1B6N0f/u4FJ3QK4j/UVS1Bxw
IRIvQ3TTvnrRba3HV1fBDF2/smoi/GWBeM+SrHDLtiKrKAtU4dQpqTup5bXHMfjRgnV/dWNGVj8I
sZFDdwBlTnSMyMQPBXz2Wy0o8pZ29dQYj6YGepKSP0IxMaHpssPA0d+2geYOvkZjjmxXrxzjgytI
LEFPV+/eV/HZB+8TWGdPm2jJDcRTs1lo6bnwNSxrje4I7iX/GsXBuzWkhbRTDMXQo3vO9PgBtdzX
AyIB9xjOuKV9epqh1IDKJYl3l6koGieYEPg+6YwzK/frX/AqrnZAeGl2FGI7KFlTL6RgOG1Bab/6
CYDir/EladdcViK/CT3zpfzghi73NtBVcljdBNfhTcj6GFK97PPWs+AnX8np5VPy6nPj7bnlgAVh
KmYHCNpy6TJOg6mwKRwIkGjh+JaAsi5Lj802mnIu5cKBC1OzIjOJahFSa5MTEHcQFgaJtM0wQToD
jb1sCp98JMBWzY8Fin2axDqpx9G01P7egsFxnb6HNMo/lUpwzU47Z7BySipxT+wWaIS1BjGrwCm8
gBoZ+Am59GNhL/iE8GNxyoCmzhPRJGkt6oEHwAdBOyXRRiecEvHTI8z1pR34SGNpzQGT6JrY1OhL
C+7NMn5Ttmg0s5X/tNGUhplOUmcYaDKXyn4mzcqdHD5+/hW6XUxfCuXLUSWZP6RIil6OuNNlPyny
PAMmCqxmVR241Tg49RbRwuOswDjDJPHYTtzKlnXH5gEVBM6VJSQRBNK0YKbCWF7BbuEGejuIaIv8
LAWJYkTOk0QTmHC2skpTP603mp1dkQ4onggfG47fghG7pHuQN7Cj5eeuuiqSC9LWsse3Yaq2OLJ2
XZxdA2SNMmEUY1WgJL77A1m88+IJhU2dWh06BwFUvCLJOqVzC+CXePYGybd1awB2PN5eV3X1ClUs
GblyynUYnywOW5+L2aMOyd9xAvtP0TFhuEfEr+7zWGE7Rw+pQSKbxFLIaljqwkW6pV/FrCLm6Rys
lX3QOAWq92H/Fv5VWzTGJRatZx3MxcWrcRAAIIfb60/nJrjWgYOkqWXLtyHXEkYDNstYuD/O5gJy
LMXdDxhFJBOc44KEATWXDOZ5rdDVYV5OHwzqY5fSk6J87FAUhmAJm9xKaUYS1c2WLcFVR6ZpJt5F
+yeV598iMeOmDLIS8RSVM4nutNKPC6o4s7Siaqt3oAZPnSGy231zXB+wbviaqmJoo5iVZzy14LHH
fPGsz5GcvBaxpmeimdzNIeO/jYxGiEDPcRtIy9qPYpR45okdKwH+dDKx5MNXzMamWNGEpk6YMEbK
SORdtikwx68mTh97JZ9X9kxFt3whlYgCjS+r/iEyTvSSxpPVRDJMx4bD0boh2ggDiV/0p+U30eEI
M9qgxS3SIOJPMTOxXiKfZ0l9Rh9mPZ9GC/9fDIM1h0uIFMcMqtGtzZQBD5WA6V9BTGci7Y/WePID
KxhlLxVxj1BzzhJfTbMw7ZEtgob/7lsK4+irFz168n9tUjRCh63sH3cothIdxR4WcJmuEoCBWPps
rDKYoyz7Pr/A8RfOF0V2jGhcdKV8JeOGMp4iV+NQkHt+0NMgEqLnqb2Yl2Qkkc6327NyddOiS1f0
XS/I/a25r0z1v+L0z73V0+t/f0CAdXoI+mm0QU2JMrQoitfMHRSgGMABxVtcMuPNDzPRkH9kmyLa
pGES64nXuPjni0e/zsnkSmG0vW7dASm2UFIZoCakNLxpu/bLODesDv8yg6fagVbzLz6FDU/m08kK
zUxipvX3+77N+G3FUtE+VrJJ3PilmIrBeKA0sWnMgF7Su5Mt9XhzM+lIN69Aj7gHff9IE5AANuqP
BQM7vfgQEXG9VLioUSYt2GLsOdIQecCqS+ewCqQFxROh/5Ee3bvFEfZJsLI2P9yI7zb23vmPM9uG
GayuzLqdU1uErokVvilLVIW38whwdmSV35Owy1ko+B0WKbNJ+emsMbzkPbAQDnzEvpvO3f3aAcvr
VWcDaU4wIR7BVzy7eDruvCNoRHaczwn+uukPJWRvxICZrSp2nm8KeE5P0+PTxkcvXSOLg6QmXJAj
2DfSN6HjGy3oJkOt9mWCdZzbhGpC1HjMrgQtg4M5UQ+u7FWy7orPCp8PK9Fx2y3n3KY8JFlBNbp4
IWwhc9Up3fo1QmH8SpZNweR5GTfnPxd51U+xx6XqbaXtVBYfk95h1zPQrYzN6VNQq+O4uTH/AS+7
Pgf4Yy2+KbRlleok9KitmDA/xUtYiEDjLvfzQZ3QF1qc0nJ408Atu0iP1xBg2RAyaFFC43ZZ4v8H
OKR0P9ndS1716Un3FoC9f1gVkNPoYY+BFzVClUgjdNWjsar9v8aZeLaultC4vS1bje4gMoWJMGMm
zYTU0F3ER2XfzLmHD4tvR2/PL4XmK9b9BzbwAzoLR2RGfntTZQPPumhhNqh0dZKhUOytKQXMi+hr
W+3j+bW2nrgtPmJrCuq8yUaS6YqKBwSTLdj3yBparynJop7qCmEn9yxfPnvkDN5n6c7ad+55hv13
RX/IQ3qDIOk3DPIkbOSIg659Y6w+gCG0URsfqLeYaokjItA9aMKNJEWLSIW+5nWcuWZwPnHM6WVl
CWi7YWI5vEYh+SQKWUO52h+GIFnPWb/7+NHEWeqyKeq5zvVMLU9gggKFFsjZKMs7ic6slqj98/ik
DCQhr9XERPwY0YflXeH49TVKX81Pdx0NNg7hQLIxwErgqBtOqQaqw53TXWkx13jMeG6W4pos8vD6
vNXYUmuFtaOLHRwA+iSFWGDPfcASuuDAaPcfnbpwak7uhuXxgwcUO17IuQSs3hr57JhPz0T/GrkN
tUVIlu2P1Kz4WPsNLQZ4uH/Oh0lOQvrdDrr+HHY5NX4+rbVg//vCjgrHUbxli1l9XV92LHgk4c55
E4KsvTinBb4JLLEDpfKeRMosP8ojCzCwKUkTeFf3lauYp3CrJP+95W3UCM56MEPr6AzGzclnOPIn
tOMRnzIzt4ykzB6McTReAg9dEE6YgKJEYxGCRigIlMO9vsSoKRXvPyqiwJ3pC8W1O2p2D3wt6F4f
yywqyl5p/HUPiXNbxaDfxGW4CNBXtbDfjwGR3VVmwxmIx6MCdiWjvbbd4PRBvLd1FsnAfDOTtPF4
XuLiZjhFyDVmtug2I/m3TgFBGOS+Ox8kXlCnlhqz8FvPZRpM9QHtxgw/jIoZn/4/85rvzSPoZ9Zh
NP4BAbQRfVic95ylVVTIWQumsdeBPIECZwt0FZm5lvfIbOMYOB4VjU/uvY/d4pdbrAhSATYyUWnO
YvrVw1sV/j0g/U5pdCatkDL9wcvRK2/Zxv7Y4y3zINgz4JMcU/pihVUGEihm7h/Blk3w2LmQpxSX
ZFwHNKlPKIjMAK02FmqVpL9XW29Pvu5AnUbAhWIJ6TUL2rbvW+ToUkcjsoo13KaTITuBgpsP5+iW
o+iKTEgSZaby/H/Yny6LIr69cHCIDLpKOBxRR5DnDeyGRvcQkBcZmlyKEn0jV0SS56kCH+eZs+6Y
Mt5pgGhNPmRzryUcOrWAmlVo9ASNvgD7KM8kcpmo/Kmmt4z3MWsCggFEC8uCm0rz4d53ob8xqLt/
h4fJS/AZK0gu23zsBvWhmFtjbfddqIpATlYNdb1hmUR1DxjjuDAJ8eYBXMgRAm8nfhHFSosM1ch2
KYAitz8fZNPmWPlqRDVZF0X3ZupkA43uK716YVuo2KLF+9lzTsH8RCDW8cxxz8mHZXAbyCZBYeH9
jgvAvnSmTFn6lUQM9xe2HIkNoptHwbAOBiz/U8QQ8GyLgcvDdreAnws/Bko6PJFPMmDg9CzeCkoN
0dbWg8zSQoJ5HfxlTfaJG9foUxs2Va14O2G6rJsznr6CZGlFm7fCbY5K1hWyje0sIFnHmH2lkM0x
IUuXIXKxZBxNZzTd1x4SZkboLxxdN8tD9ZiNn668cQOGdRGjZ02pK/5onjzFw2kWaHlCADPWxomu
uusi19m4NEytQbIC1iWm8ulqJwQ4UujQa0P+r8z6FPyWdl13cO/SLz5tfmfwnUPeo1iMBcNZJbkb
U9qRSQCVt4DkFnbmuSRSVztuBLaO+CCS9IT/tma8Kj1ib7z22LLwZJIp81Di15ZHDqF/2hE4Ynuy
/bWFNU+pmau8ZV6GoWCnVGj4Vq6jRrc4cZ83iH3aDHNQ1dxm7DdwZUkNegADj0aXOH2v3ZeZzdTo
0HGfpQ3obFMpQb8lsNP+Lu/h03Bk1jomcmOEniZVdZz20Gb/xE2ISK+QtZyBszUW0mJAAH30q8Ic
xb5SN8bhlnXph3ZTcEfKsISmNXUe5YlFGFYuMji4br8TKWEWyDMmHg2A97sEb6QYjHrF3XHIF4dq
kP0J1IpozFf1D0+bXufl2HDn2H36HZSkUusD0WVykeBl4AqMQg+sWXTcr2QaXUbfiaxPPF8tg4wd
GIw3n2c3qS0rAa1a2wWfhhHMoMbXl/xoH8sE3n/V7dBhjPQk78LRIII4jE9vPksNzZ7gZKcYMDKZ
uaPOP8JxTwHJ7RAc5TLVsj0CUJBbPrYDkxyt3+j7BPV9pLpSeDR3jFIv0B1sBVmxgxDi7f1fmceG
c/syJpsZJXgUQSr07TT3htSBHR6EhhKab6+UxklJR2A+qrpg8IROckQ+++p0EzdbF6xUwSil6hNj
A4nYAfxgVdPrDWw6HFc363PqtuQjtqzJY5Pk3MeO+WogfKfIKxeUB07brBYHkAPZv0+d2yuKwcx7
WAE08bzrV/3mdLl3bEamre0UmtiBUuZwFsMfHA56M5XdkF1I7+twWnEtxGDYvYbcqem6M6+VfBip
22QUhDjvmV76e9ZCixbY3Vd0ZXgBajkP4vuzHB0Ydeu06I83U+P1QBC7fbBWebE8jYTovMDxV2Fs
VudT6GA6yMRwmS9hO1JkdzTlyCCAwwgHpYB9/xuJGSKdt2BGh0O7mWQNI8Y7sRGgnFTfB95ozRs1
37vyYSadUrClkTaWUYxH39jCZqg+t30J5bdZH+r4Aa3Hudo5ND1cVK8CrrwBRK5gkX6+Tu1iwtww
w3iBlaH2Jt9L+7oUqYTd+BAG46Vp2FKudthF/tmzIOHSkF505VXJ/tt7Or9vCchOkycKMvUBDpC7
kOBJ0ioXQaKaSr2iO0jntj0VbTJUmgdcoJavxdr2rIYeIHoBQUxZWg4LxxKF4rY0MYCzKKq5B4SZ
lQrFfRPWrxjA643TZE355+B/mQ0Fy7bk45v8XfCkI1YzKdJ62DK7782tXtAgFhVrjcYwqHiGSbvF
dAc8bubW451Vgmgkode/49GqudYqwebuul9KGvddhuzNmUIhLsAlOaJAuBVJzy8lpzD5LFynyuHq
1aQIFoL9d5PCC3DSEU8o+vEPmoG1K2/nDCbe3oHsm9N/VxME6giHsuaao3XHwbzfTFP1Y1YCegMK
zrmNiFiQzfFBdypzSmvT/LwKJpj5qmA+/bKFmjaT6Bi+Z9qANuKhj7cWpvP9zw6727Of1eojohdL
cDMWKzqJDfu+kzyf0YOq+xqwsIU/6v1GVQ/TS9dv+a3mgL30e/V/k9fkkBW9cm3Z7aQK/lJ47zh2
oVEOX/YMF4MuHsp52IpwZQiKgwTeEDhrxOxhanxOuFTdMoM9aCicwG5n/kcZ+3O/M/92J/KwjOqk
RGsGYYyP1afTaa7ZpBxOaar+MnYNP/Z6bDkkdt2J8jE/WUJBBHp5N5NscsvQ/ziX8XnGoQPhm/hf
TloMjKHbbUoSrEZDgE7sj9GJMsLYMroco4Fty+0bC6NzpfluE591uqbTmVzpC1OXSm2nldSvv8l9
5A3vdIjf26fHvy7Y4UzMmCkJbJU5CX7vOl745BGaY86bkd0vQZt8vstQTgpBOeJ3m2PHY5FtIDKY
nt5CApIQhVdvszg9LAszM0+9GMbVkKWHG5fHQFraTnGsZFPGHMCd7EVO1bJCkxM+eTz83ebKlUeJ
/p5mr6ho3ElvUpVmckzXTMyLPs2dsdnFJV6A1/fgoLCZkDV3TvQGMmguYqWr6ptbWeePeiJ3RD/K
huUI+7f8nv1bajl3I/wwnUY1sryWmHX5Xx8EV9Pox47QHVZFZ31GSJA6vo/ISbEG62eo+mIpDTuA
wBhIjg1ipdMFeFRoyZzLKj8LWRVwei9bSvBxhB12SKL9nxLEfwTF3cYkFElylts+El2wyCCNb3u2
689Z2xobNf0fNkyV81m016EMwWVE+YkwjGIIkqt0kN5FEOytB351+TMEm/+Kd0LbUyuIMNKvKqNQ
hzgzafCPSEDDbY9YKldK1+Ytt7Zqemj25EQf8+s5KRdzN+CvAwzrs3EICgVahzqvHHjfbuFEKqan
9pF5f3SMEZLLUQPCoPKI4zC+H41V5aSEU+VJHfcuiHRwdFy7R53V0tMV8zRY9R4BAn1mc88dxTcW
Y718kChAhfjVhdH+c4O54FS6DBbkZD9E6XmVm0BVFaiQyOqbpKuYG0giCfrVTS2jb91Jry/XeEh1
EtEPgr1Ezuc9o8QCBEYVE6R7AsmVvZzdt3PFcuu2GJfqlsWYI25kbJ49V8xK1cGdLTAClS7SE/i8
zm58MwmLLH/S/KDo/YcjRj8bnrqgv34cp6uAfxA5gDYb9pOtS5E4dME6c8EUqNTZiMk7sL5NQ4e2
Sy1v3ZtOF465jcl0T2B6t9u9HVSVNDgC+yyi/hBn3J8CafVXXwm1wf9csnCCBgQk6TOx0zQPfd7A
WPHxrE7GnC5UQVw1kYgSsBSbhgbjRNPF/LeOYn/nDRmR+L1gzJyT0t5UOC3Ibe7vn9yMF5mwarFA
Sz0CLbJvbof77ay6yhkYJHOoZyQDYN0bJ38tXDXRI/0V6EdoohEYqMhXAxw95dQG/sACaqcx48PZ
BlWc6iaPFyW217ylzSrGtKxNKMjCFg/VvA0emegSxM3cbUVdNm6fp7VhA3Jdl8iA5pg6U/LnqU9C
HKqWTsS90ePOXri7TNc1lXXgLC4ssSnWLFV+nJ/zGDJJLwwyKShvqz7HbA/pilp35EjX5jw9B2g4
GLK9O3ZAAerZk1Qi7IqhX7PKQAMzoVEyljnZRg+oTAVFbDScj7vu6cqVEXzXUExDVkqY+ImVMWZ3
0JskemwE4ZRJE8kA9ezBYcDBWENjbPT0Cw3oFF9hifp7qHJvQnSnKoppEcCOsxzExLlBifQDGb12
3dXZ6pmUe+eWq9srLwVf+Oa0WtpNaXQ9w4ttfC1zJ+DQ0yQJEIGEe6EREGjN1f2Qz2+7IURXihzr
sdNQPJixmHtGlrjrqAp2chIyLPqFguwOFQmI2qKgF//VGjRp6ZpF7Ur6Tr4T/Tm2STvotlRAorxQ
l7DyFteJyVWpgL41sVNEoYnREfMkveqBRTQwomMQ85TcLPbF+klDCH5ge/GnMShWhtWdvw9XlSJS
m5Gjc6VPYSkikqPldkhYnjNPRgpjr7ZCLKTQ95+mxL4+3JlbjZbsPPtx5mGXPrtmH8yRxMmzmley
IBnxc5lX6621+MPoFofy28YLw+Jm9pfWsn0l/oP25Ij1FEW038wVJH18xDJfuPw9NBoZwlAffcOu
wqPsupPCkjUwq1yCNKcHT3lWwZWiF8a/6Ab4myqsFQZPjODCCBhxLDgMrXA1bZWWaFPasSa0oUMx
Sfgkpf7Z/gAcM3FrCTyieiDfjs5Rz8XH7+j6R8wfJLs0h1R4UtJlhFjjcpHOX8M3Da2UdyFjMF4d
m80AuN/38AmxzuIeP+D/1tgtesYf1GO2cWxLQiNM/HbNAxiMNvuARr2vWlbDuQT55Z6cKEyjLrYi
ItB26OqPvj2IEGEQsVn0WXkfnOvSYQ/B0EAtJ+2vPjZ1t8YTr2imkqev++4Q/1c9fdjoQKByUHE0
J2/cN1bg2QwpqGODTUSIFokIjEfcHcnHv4d5PNcwKZKykW1TtBrMz7j8I5IohIGv1I77Y/bJktks
PzIpcVwBKucNXj0pw0p5TH1mELpP4vHu6SGuVdmXWOsjiHqADx97BjoDYizHNxx4N61zUOXVkowi
V/TJ/yCzP7ojnRE5kil4aewF2q88MttG35GfarkqKNk33Lva92M2poB0CjlyWCZDNPkz5+MX53Gc
YI3TtSGOIcoQJHiI/tFz1daxOS68UrEny3IElsmacG/Trb4CfC+VuyioEEmBjRASrBtusNp6bxFw
mxsq00Uqx5z/F5+aRATyxuHrLYpyj4x5p3D4CioXPUQyeuDQa34pgW0QyXatg509pCWoyt9Zva/b
NJCfSrrXR3DpFV71If5hhQ3YcxpeSa8zsE8p7yucyiF3GUrfW1TgM8p7iJw88iLl5xCrUYGXAVzt
fjm4YDmfmd+2yy4Yhd/T1xDGyaGZuBQHUSN1PCz3wkyulrls7g6din46BbK84YiFEIKZE+E8VdCn
Q8vZzzxgJIf5f432IZ+vP2szTR+VoqAcoPp2oqEUlZvIjTKENhaxrOvCzikbQ1qMemMTggcuFaqd
22Lxus3WV1IYJ3XwbbwUDxONST6fWAzOMNix/cYncLw2WzKSlsvX3F2P3odSQgVi+Hq5OpCj/Hfi
2Otx641SxgVxTJv789AM/jinknEfk6qkKPEdeQZ0+/ktfg/4U+v2yLbkdbvlaGwHUSWDkbHnwGF7
Odf5ookiSOcsMiqX5AW4CgYVM0bU64y9YxCky0DGtwmuVkqP4vpSzKOEm7t4nPijFXWV3+hxaVnq
lpqwCyNPGvxTW7b2IOptzXG+3waTF41Q61wkZTEpbiUBkINB+uXEAM49dDZ8wUu+gNo3mEylr5Lh
qeILGwqfiYy3gTIgtL5FVzfO8SCQ+VUrJ09dFrkHoExVCaPjARfMmpukMlA3M9ECZC0h68P2IWtE
fijdeGQHVMWAqrDyVY2K2xsAe3wso4HtfPbcK8ZZro7XnGRtfdpG+/Ui86/QPdqKAbJe22tT7c6x
fahy21QoJPOeDrveRDOprRxLCcoZNFVuW2PwGRtF7jkZvVN8WiOBsBnJQlUICp6DaOKFLB+zMKqN
UvYvIudV0fF79VgYEjk9/1T6UP64lZMKK09jswqNBvXSCAzg0tCE1zqrD5MV1CR3iFl/Mtoh5hfb
gIJlmyZTlea0csiYXkJwY7j7GR4VfHSpEaHJc5wSFVoQCAqkVPQnLUSeot6FGT30G/VTjNdgsUit
bbtD9HtVLKfvuktiB0SWLt2QwWkx/EtlrqrF+uR6yPIvxdk1PthDZxYo8OYxnW3QPhtUBRusD7lQ
PWGXp/6X6h6MIcRO/I8O8fLsB+t/my6q/zka97pDBzg+ldNdwCuA6QB13Lorrb6ppDQgRJpzM02Y
fhoXIX0EzKSFRvHn6FXLapHg47n0rzlf2axvPaP/DwM95DUW8c2w4ITJGEg03TDzNay7B4YGXDs/
AmpIGmegq6ArSl8ppjaTOmXD9t3bJhuhR3Kqg5jx7vArBZiyj6i02l2xv7ciOJX/54bswBFGD5O9
uICzZ6QObupIQXS5GRH6/GwrdBQWXr/Qc+SUcqdvQenEYFPOJmO7GV2GwHrzUTUQHTwOqJf14L2i
dbhAjnoWW7pgdD0Fw4AQrnYa3Ylq7bObbbA2lHP3n82fpCQkAvIPE9fa1j9EICULmh9k+5Lku2iL
qBq9YLsUn6mz2Mo5MSYQaxwDiLl+ChM7Y2IguxRopyj7yHgG0hZ/XMu6dEFi/IKmKNm62HEna6vj
NgxpCmLihDhDZRYe1AUfgEWvnsRNRJ1ZaCJnhTJ7/dx5s/69M7Jh/OIYnJ2j3WAl378QqIE6WQIB
CL9y6L4l4Kp5QY6xEjyv0gD0xgidoTpEj8xtANXFUCYjhcLPYo3MLC2DpyzhJRHCYyEGnbeYnnVy
6QTJlA/ObZSd5AdYg6JDROs7xI265AIUvZX56e6pG+n+t9sRoGFJ4NN9jDEGu1lw6USR289w5UaI
gES2FXmkfeJ9mhpRLq46Daqk3hLvjJR7ERaqG43nAcaNan9nqhg8V8ctmBy28TIjQ5UhkHj+UfYS
+2VYKVV4Mh1EWX7ruZ3NsZk1s4a1Rw/kvrPNAfd7+RnEJCS1E26WcKms31xUWFm76UNtOT+ndP2g
k1T5chvZ3PcDqY0r0p+0Soqu9wgp+7dlbe+om7fKbwT4IiIkPcdyv8CQdmmljAEZuov1tkBdBe7x
JlZ7RpZMe/8ix2rKrWoQ3nZCcawPHW7HzVh0f3vCojL4dK+aYJ+0JGgZ8RzPU6Pou2WSO5ZR9h0B
S552LwKiWiOx5SpdStXx+Lfe/28IjfoCd7eYDSqcHGaR64+KHTeMSpYrS5L6SB0v5LRNvafWOpAU
r1GHd+BnVVsTG+mvqoQkQq38u1rAttxIi9BrmTl6aCBH10d9as5p5OzRL2VDTWI7XQA6whgBIH2i
qH0p/DuzvgRhLrlG6ceRilX+bcp+cqBGz2YXLubvytaxOCCcWRI0sq6Ex4QHK5utjNr5dUIn9xkE
fzXXyAXc5jI4g758/JTq6gu3dHuheBW6/bAXgCmz0hv7ihivCgAIvXj1JBA557ONlBB86YMWA+di
auU9k8IdCfc9n5HyBYzlbEJvSJQZ+xaFyVDO04fcnstMxfs7yXBcrG/TZ+oAVArlBMzvya1/eGJ6
EUVtFUDSKnRafLPR0ulP8Fc7MFabogzWZycoMevJ4VP8WEm2kMWAE6p6ZkWsKf9HsFhga3aC2oAE
rjHb0eolVUbMmQk8IRmRah/zJzcnOiWRJvRmuJgCARpBF4uAz1aV03jgZB+2Q/ZQuP9poXoUtD1n
4z0+tU1dhlqN2sFrENfhw/xPjoZvZSbax7eaXrmviiKW1rR7LIgJxgpix1cPAa3TCQzQJ/IFSx21
0fGH1DSU3bZxQ70jxyMROaCtECCEnjnxcUMa2jszMYf1QDsEU6gEx8L/ZCO3PhYClJjrzM7O6WgP
3dicrF5zUW7MBh4vM6EvHKBNyJ3Jm2sFEB8rDXoXb+jcy4mS2MbZ7NSnj79cQB/7x/0MkAWP9Qi5
zzs4UG4exjZr2pknfA7A2QsvDnmwajQn8qpJmO8Dfj6m6gnyWGfXdT6/kZCkmkeA41Vx1QPABQ9i
GeWqgwr1cRmMWdd64LzjMUr07/p6AFiAAtnNjmi3Rogtl8cLvBZnAgJbXcfFg5Gd2alPK8Wq3/0g
IErJiupi4UVXk09iu/mIrbftcGKQMXlOzYme6For7a1ItP2Q4zkro8bgygbO3aA8J87eUjyJN3H7
kdAgw35QZvUiYweKup2y/yrisOElBfLVqFaIP08z+vwc4n5Gj1sIztF1xu2gFb3n6VmwUfJ8e8Kp
W8EZeVKAfOxF3ZCbPYUEynT3xX5yxqzllRI2pijhb94PfUlst1cUTSh8yiUMupA9/TQ3DtDlWYKM
3iF0tAd560MZBJ5wpWnUZ0GOoA2kXQ1a8l4hV1qQwSzzixi/r2dqA+cepjVjKQDA3Ie0iIfOb/qZ
4iHu2Jc2Xq4c4eWWJ+VicwYS+X+slUfS3uoAXeDWC3XO7iUzjLCp493Pbt0C7oTZspTaVlXOu6dZ
YJU5Ooem3KdjqdDBzbE1ZvEykGVsl1CV+o8TXXak5j7/KrpyCCIbqP6DrtXXuKW1r9D5HJWNih4N
h7LIWwubJ/iHP4QINSl1sPV/WwVzMBmVzy8No40FFNnd6TUuU1mxrAnuKLHazLsNKgTj7+6lXsym
Tm0OFcOe6EoCz41n0GT5tvQgz+2gEofoA/7bGrD84APgHyBHkEfrw9vi2TUiPPxs2LotoubMbK87
BtUFJTntT22EpCmP+6fmDKX5PqfNm4Wujz5KxHqAep0l5GCqh90WROsHxNZe1UBAvCuEV01JuIM6
mmxTToS+v6s+GEAV0JLPpOIk84pHVALhEnQGiC0geXrWMWV2lFaO67O42GCdAdJHtKRT9DdU+cEn
2mBHydr96yCdsi4kH2qqIJfvVVNajsh31QlnwgT+TRAwk6WeXe8k/JBOIl2ZFfHW1ARBVFSrb9J0
sddT1BvZfglsyZ3ofnhtPOotd7N8W9m24QttEkwySvGrjZocR5+/tuHvtOSR2YZ9uJpxyry1CKcL
771j1u4mn+1deswx4g4XXdk1VyPhnEqQcH4GHVcfz1jFe7w0JJl+5VZ7urVP7UFylxBr8d8igiIi
oB7gQoNE+On7WlTHp6jjVDGAIlziijWPDRepP46lQhapGt8v/4cFQSsOdj1gB8pE8EuxCFiwVrCw
tzbWzT1wrshaS+bQYe0UG/UFj0QDUhwtF3x9YEHVZHQzpQtKI1LlEpofNCStKWtol7AvzTunwJsd
5XmSHEIyThJiQ5MfxJP5Yy/33UeAVXiZCdjfY5LclolW/33tFrWfSModOSVm2AQUtjC2RJn3fx3D
yOB84u30i9t+8Y1eOypEWNoLBDQ2v7GaXZRh/0DLDKTzs1UzjyJgP5lqPS5Ac9fq7V/tp/mbED0L
JjlsbhboSbRWD3CV2OaMJdAK1VEwtQqzX437TnUV4yukEsOdni3M/zhF/uSmZTrBZF3o+T6aUf9y
To2kmxqbL7fPbCo7Cc7ZsFI2fuuqPechB3gerYH/C6vd2qkYDqCvBiI5TGJsL/MVBjOZzRipvuMb
9ulLG6PGjqzpzkFT/ClVNYl6u/H85n1AqexT7lm8ET9DOQpLRq15XKAMG92tbUmXCVxb4bOoNIN3
YX8LTv1tpTvj7v5fKCaFglg/5IYmfDYA7iYWzxoeLWuR6AWhf4nWDHab7l6e9WdqxqYgtBw0ugk8
5DmbL7EkAE6Ro903d3uQHTDCuPs8ZPCrGr+2O8U4gNRF27x8b/Mn4gNq7QYwbSyTZ+KeWlaLTUAS
HQjA9k73QJ0aYBxRtFwcxGiDmJyyDiVmFyDkSZL7VK0Q1VMyHeOK3KhKAshcbc1IVSJRt9eCKUJl
BCepZj2gYgqE9QPXqWbuSlNY1mdl+k63X9MK1mCD4tOd9e+pTdCd8zYxJda24F0WToKNXsWmEqkI
8YJAqwWTs5UjUVOk5boAh0IBwRRlc8dw2jJvZk86L3DKyiXN0jj+WdxKWiVEPaVt3KdHSX16WWQj
Vb5SivA9V9pVHuQ8IhAgKb71rafpvtLbBl0ff6hnLRxPYIJuY0U77OrDL+D4+eItFge7CMw7pCQj
yjg/cmQCNa9r4IO0MoZ7lIhBHQ1wayLVz+TwxQ01tR9YjFBnBOm5kdxRunD4bneChzdroWuJT4+a
HoS99hlGqO6FK8AkCZ1HW/DhV6EFhNeDpstofNIExXYXcQgDH9UgTeonM2ummXDHMGdx41PxOuGw
Gj17wxYudRFu+iqlFiEanaxPv3r6KIGXeJSPkjput9OoZ1ZgUKzGY/0dnwTCwtskQimDDgMszX02
xV1FTN1+xWoRs0VzVCM21wyE9zISasw1uAUg58z6bbshVxPKZka9nXJmEed0vlcWINHQElGxR8bT
D4UK8L6PoH5Ku1satmnjugioddumFuXExigWHbILQjKkcHAVWVDVV8mTc3h2l9T/evERTg8kyzPE
ZBtdDiMiTl1DGx+R/+ccAfJylrNwDxCCCvNl5HZEK8tHbt9PR8vooocbJApP5qO/ljNIF7wLq5Rq
5fGGuLfDKBFHqnFIwra2cIrbek1cRtwk79jwg4TZtCLKv805Lhky38wGYQ89wCsCT2eqo1w3Qurs
XVxRso+ryi2qLzUzOXGU+ro9frwetlL7q93yNB5ueH4EzQZoMByYYE/KGMje1/O7JcX1WUY65BXi
k2QSyDWjyMJYPsdtmPOSZ+LMKq3zEZoLYAvGdnSt6Dx5BfAbqmDlnf/V+SMUKpzo5AAwRbv04xkh
w2ceZIdyveYuT7B7Q1TqOH1QtTS+cMPGpolK80qbysOkDeYaHuFywdIxNIzlThAE/m4mKooQ2Iw6
sM0ykS46YQnlskkxZREqk88vYIoYuryjLCI0J/sO2fPa2h0NpURtJFt02uoQikKJHMJG9ysoEGb4
h7O5ULC3kI7SQYQZFmQrFxSPWz6F8+D8IzidxIxXWlOn9BoFf03LpmKoqFZ4vrk8oZjmIZ5eHY12
d+zO0WvzwH0vrRi6Dlsiv0DBrP+myoibxwyz+G9dojAP6I64+O9rR5NLBTIG8xWKvRF+ecNS9FUi
O3JsOIRJFFeiE+8ZhSboTDgWMWqRmAogrKn2QyrJ44V+Rg/7YqmHbV9eFoEu4CP61mM7ojoYS57X
P0mkLXEPYJVoYAe2q84ENjR5ip28zs8oqQDZUFddQcESDqCpcx3QcpKDap5RMJ3pIZbB4lO4blC9
YL4EE+MadztaZl3mtYl4SzDImOlH/piPz1JFl2QRswJesnBlF9FEwu6O1E4pi2lQSjR+zzB2XLba
eDaQA5WMAa56RinFDV/7vha7kzXF3UJUBqN07vrI0JoNeuQiQkz8CWpFQ2J8Zg96dT1o/J9/7lwU
hLX1QuFmyK/tCmShPK/6j6PxCatA5NchrBHhlW2Ev94W2kXj55J0erM9Qonq5/ONUJ7+wAA7Mbmx
YzEFTIGC5kfJSKm349qUYZLWV/RiEOHqXOzGfMt1ASPuzf9HRZWAfJbNUC5129cbuOC2mIzsk0E9
zNZsb8YMYayCkLvhX/Uu2xsCp4xMNClxs2S8VQZ9FWHEFo2fHkqU0657DiODfARhdc6IyE4HOM8Q
rGAa7axeDMn9EiPCgbMaZQznEBb4mkuBZTwFAZSbh7TGTrgWlEdjzuODA0m0eCu53n01F5LzOt/U
4xPzM+yemb/7syvCOd1TIlcJIKFbMRDhXS0kpC7T7qlFGUUKHm3qg3B0wN44rq00z58V1hPw0YQv
qgbT9qoz5BuHae5QVJFY7L1YCZt5qPKGOlBb7CsTYkTceTmyqvgDqfdtVkgXwID0CzloTn7BD0D0
uHqdYmMePNyLsfwfvBipCr2bK0Ctx+YiCUcTunijFu3LeQjn668Un9CnPk6Iea6mxxv6lnG73amf
4Wcq23WgremARaz2pLMWqOhapJBqf9HZP08d0yNkByNsDm6uFB+YQKLa9V/7k/BeJ1iBa8UMCX/b
5bFjzwmEFMuDZu2aYsD0lpHCSLrc2y/ApVmVacDBebub1v4UIQSpUQzSzQPnWvRoYaxeU9WBAmDB
+wttyOnszGq4kBB/v6vQVXOp5r1jW2w9nytLi8orW5E1cHGyCy59JQ+2qJUI4mTULOhi/RHL0bfx
V4rvtRtrK5qWXqEXKfjR+Ax+viJAx3Wq8+PQ9Fu36G6n12/b1uQ9RXQ38cwoxMQ11glaIfpnvOSe
8OKViES59m7U0ZQOXrc4oVtAzrCNWe0yI+3IUSxi7XfKW01oH0RL66EMikf9Q5XfoUn0g6M6BYAV
tR3cuOxYh2Kvg1pKOf0zKhkM52zxqbUyMyq/nWKDt1PbqXzw1ycPMBXBF2Jn7wwJlrHALRLiiA2+
JtrBAE8zpULewo288Vt2Go0E3VdePUk/7HPkzMtnvb7+AdRNUrJKWOOKbUT+BNa0/wQA8PST/45l
6VAPDbudaV+tWHKmZI1tkQnc57ZxStGyjaFKFVxkr9QfJ6urxkhB5OoPkpnqUUkWIo5tYvq7RnM1
dLHZRHyqPsowiKEEtaJnsP5pe/rhsQLGZoPI4pl59OWb6Xw3vqmPwrPzGRzWr96tblVNbuwlhuIC
Vb+wKtkrRSkjZrxJXJAu7b68Bm9hf2nlTv1XqWl/71/Z7vJyHuGtNILI8OyVx7+yccZFOIjC37zY
41ocfD/di/seeJQd/wn3UbSC0d3+3+poLh5cy6yf0yZl1qiUHku9D1pkv944IAqcehDgTD6pihin
CqvjzyOHmZiI7dTZ9tq1PllWMsOjBH9SqsrOKUTL4ClNjlqRLiWc5wLpGhoDy/Wmbwk/6I0RvaYs
z0vJheew0EQyx6J0VHvSzltsvjh3WMAgY0xR14JDzwS4e1zElBghXyOyLSaDgOpg3tOejCpQZcVl
AMrvtkOEYKP6/83SR41VNQ5rAjQoNHsGmWBe8qnaDZFvagqLb4ZcYy7eZCD4tj607Elha5hrLbEo
FyR8V9+GrKP9Z4L1EENmYYfXC80lcInfIURznjF1kLQksGZX6+HZYXw4yRyjitwzukSRfUF5587h
LMgZm5EyiSdzf2owIbKp0HqIt5y5cUZ75sN3ahqCVkIr4ZuGbGRKBF1KHZM39VySo2GmYGVkFy+Q
jbfFgcdRwfd4Wb+xCLaEVdm1mSJ+5gWf3isHsWD5zs5/FJa3a/rzWg6c/ADUDrkPHtBMBRZZQG9F
7iCnUvw6XMFPHSZaPX3L6+zM789ELu6ZJjUmAuvdK/c18vcyx9d7iwKzAGCpCWeSvvfTH0S8bSym
2E1AUgdnhf2UZ8FbOP+/zKEiAAyruuxV2xbcryHBSIexQz86nvR896CImSBDUz/wwPGE2jOZvSae
mtbCxzCwz0a2QJNFvAymnoorsMbnnyzyTZX5YCG72ar2WjBmVInp+H39CoHDxloZjQR8tCVDDs0t
XdSO7IWHcW26Cvvjb+j2QOSAnXhNS2v7OT6UNJW/cE5X5gA4lbYsqSaENgPT0iUNKSDCmwrevkYy
UD8D4oMfInN/JPnH1uIbVz1+EIg3l0smYwrpEZKs9L913o+w+QjjlaIPJsf+7GHtyYiZhvpOUYDD
ibAh0dACxPwYFjcsxDzdCjpXqfV5BzdN6sFAqy7zLPAUQak/jQsnNGqITp76gjir30KT2v3ewSKF
Y6ydp48342LocLcxbo0LE3qCvmdLnt7VIaUsobOaa2l4e2nJzX6hg8D31lFl5DuA2p3Y9kBOUIlS
gOGbsn5TeCqKETZR6Rg2I5zkGx2rhSX5sZfrdnJBNFouLB1FRk5FctK07Xg6JwpCXlWfxeEEAeod
Nqgs3InSusmAgBYHszJV2fwx5MCMuAfMIJTmnSBTgo+Et2g6tfyWKi3G+4LOZ5jzSR74CRhLRDKD
SJ/SZCz6lknvaatLKRaS6I7phYzQzDgkMrpUSYXdHjTZTZS4inZY7RekzYpGlh7VDom5G3veESy8
1z3TICntQHuNsEeH/b8ejBXlgHhwhAV0VnPm+4CxQbnKZ/lxjkurKbK5n0JvzhVEQL4pBDvT7c9u
Dak1JZvIZSaVBM81G5cqCh8QsqHqf4D8ZvcamDlCLx6YoejJph1T+bS/aXZ3GglYVcVmc+th6CwC
E1G0/xXwlmQegiq6rvVnUuPwBDHNoXNXuk3kTfV05FpYyblDFZ7Paqrit7BzGDq+P92p0X+cthiT
a0rEyDFblcshvVPVIKIIokX+gIFfoUYVjbtL7T6Tuo1xFgTEqNqQGn36DFYU4ekwyeHzcEmdznOi
QNEDyXDvx/wlUGulgjnZ7xPTa9OEljyvS5sqkUfHR42RMYgQizM/85g9tJ8IA6jUsDRqBPrGHa9i
L6cLRK6c9Fkxw+qO7kw2Bpqxx/SP9uigDTLXKEFDTn+o5erhasMpcSRW5zs/0ZLmbIqC3QtSSdX8
NeeGtKFFGcUuu2E0xDQjyF9xGFXNCs/4Ge9h4zCceAB2y3TFlmcwvv9cxCrq6LnOyu0+XDQkO5cK
JDL7tBzIVPgzTh/0/+FR5K6bMxe5C1omjQkzFHfXxEBerpSv2yOCcfBULN9yFh5IrmI4y1tQx3jY
W/zda2Q5jGYWaqhn1/ahiP0yv7V0nwHe4KmpWGnEx8eg7BldpYJLyxOoONcUOzLV8nJUhewM3MEZ
BNb2HK1VSRoICai8bIQcLpyYOCi5p/Pr1/x8a0M4/uJx5k+IBBwhN6AMwM2x1gntkCelhwpi6FXa
UtWsdtdgeQ7MTVZXdUMRjGM8RiFcvEfczytnPoDa52JaQB532MHHzZzpBqGPshSQszsOa4qZYhcf
/TsU8kpjBgia8BHMiH7k3PRnktz6oPGVwve/jsLBbHYF12EHCZrpVc4HI9D9HyPgQ7lo1iSAZiIa
WINBR8cFNMYmYUt/9ahd1X0F0J0rO2/ZhtkJfvvNpYlZtrpnMeq4RE3bck5BkWghyg5ADOxtbgRS
di58/7la31TjQl9dawAnQGaXCuvjyYbVoneLgXKq93OHiE+6JL/uPXwk9x7rHnRayEjIV/GAzdro
GZH2hnIM+03dJyjNsIh63Th0lm91Ss3P1UHZhrr7iF/AiRuK1ZNqxfftC85CRZ7xohrscbjWH/bi
FodEEvZqfSsUom7jSgv4lmL+TaFIIZv9jjOLTrGNPH5BLi+7EMJztmhPpYONkwlNHs1ahXcA+wPF
R3xW/oOYVCK97vvyPKpFv5+kZKDn5Uvt8mnv54gtlXVJY2VnEOmaAML9ndcB+2/d5uQhKQz0jDCD
0qELvXpnL0iSqN2mWoU+SImOQPePOICL4qGSI8KlljzkAYiUIXKYCZK7t8JF6RV6Nb4kwkpCDt7R
A//t+CdZJDJ6eFZID4vKDWNzEyPKegVdjiuPTDv8wKkPp0wF0uMwlRbYZkliqOY+ei6p6d8X+aa7
ux0EPssi9IGIRLJ3lm++PgHxWPm1lY97wjWe+sY89hi7O4d/h3BWUbTWfE0S+BHYdAUA6wg2HZUG
/RxgnLWh9fKU//WF1pPKEigIw1y184FDc1XhrdKlIjTcriFOItDx9jR/SL4uJFm+wCE6Cs1amu6J
es4ae88J2PeltmDJlQGnNqTVJ3KbxvyA0PcABN5g12eiqSRNMWHKr8gaM3SCMC7U+5S61uDeffTn
YE2UNNOK2na+JKy6tCEWMJrWhccu5qKWb3lPdaXYYKkz4MqnBpt8zCb54UlAweA3eAEheUcTOYW8
8XkWk73IvPd/28lsMjoeHtNBDZvko10kwYvJIcTJMFhMriw6dxRPX8oFPP/Qn1on3t1UqitunMD+
9irAUCcChgfYFe+QZVOK/bFr1WvhVecZDsXrnzTAlRQJM6hbsggSf1zNs1aeoxuRmXWiCJ1QxxyS
FClw2B2YnZFtma4e4bvNijvpe2Ma9UtrG09ZKdIrKpncvxcx4whF+gnjCTK109YCMXGSQtQkeZRt
0b36wLOVvPhV+6tf8GMjK6neYPfraf+eov4Ls40m4Ty4KQZ++mkwVjgnqhs4SslWM8M3OSv172jh
hgPmAgUwriISfeRX/GKTJ5oTZlyTv4f5+jEJwwMkoezhzTpqaXP7tBdOG6SEtlvFG+KhNpzSYRmX
Ld1tlXHTLWichwRuEHaE4lhoFeHBf6IQYrOwD8iMsiRNcHLe6eyFT9O7405TB/BXjABLo8Tm1TId
3ErJa9LimH3j0JRW98sD44N5FbMkqIwDCY/qD6kCi9b0UFNWC3ae3z2wcQe4FPzrM6FhkPGEr4wF
op7SuoamXDAGacA2h9IMlcXlmnvRFXE+C/PmMNnAPgb8o65+PQmcAXLj/DEwnkGWfCe2uSBidRxU
Z0fUM1vAn95fn8nVlg6IiP1GaPzMPvYLs1mfVE++r7Pi7+A6/JMAcRNLrOBXYZWX597x+Gcg8/CA
FbtcrVmSADaSNs7vguerHimaD4y3O9ESQM3TZgCE0KICn4JFczvh9jjk0JScZ7vuahirHJX3iQ9o
/h83l/5nhEQOxfsTqoWhMwIHJOcP3awHA2We12tCqeKuHTbKS32P/Q1DMnGi8hs9oGdblbj76/Fr
ueO2jCFn2tfkkc00FTF1WQ9RhbHM+mAhg2CIvV0GIQEMBAXzj/8hBETTMREoHZrCQuTXrm9FXLRx
FiFFcfuItwqmH1AyNqlFKM5oaGle56EobLEm8AOhW/dpRHFR5PI20rvmUf8SrQogh7qyUBSRsRAh
Wm01DkkEcft7TiBoLXCFXdbcwk0+Llq/LoD1Eu1C5ZKz5Js24Wfv4Xda25hNmtUJ/ppofSYRY1Nu
UBV0eW5TtEXomYlKd1eHcJOapirgMrUpp/kI91Hl07G6W8CB1k8FbStrS7FfRH9qqwia5rpw7JOz
A7Yt7nBdVMA17jF370tPHhgxcN/KCpzcXg0RqE4JbwtXni1HeFYmENWhCpGlaadAntkN9sIeSIPN
V2d8HzHN44lfR3Glvu4E+VrZJdTpA+oE4YBrY0KadBZ21rH2lKrZMCX0cJRPyfKalwUxnH4iCOhZ
yjufFV1DlcorpeeW388iJwKnvDiCRDOwl81N0NX+gCf50TsxhVzgwh+l02e/VXMmDNMG9yf25rK7
kQjkyywg8XI574Exmz4WSMSol61g/ZJrnI9C0WanbQua9ml46GPcgnQEsdjCgZ0U1vtz2Ggg3jYu
H13ffeZzLHJTkR7tAJz91ymrtUs36g9eDdgnicUJUPrJkwrc88X1v1QLiKNjxdI+LLlGfFD7k96o
Plkr12cpP6cAiS0fQBxBUBRMoRsaGsxegBaGl6qiSLX9HGXQPI1fvj9ZTJmOb6TC7rjb1Kzu0lMQ
O+EBINQwWQexbHIt73VHB1Ysy0pQ14JwJpy/c5ndfdxWxtzc5amKVRrwYbwLYyYRQFocuOpazSdg
/MzNwT49qT0sshKUxkCnwTyRgPMuoeZuXhYfQy8UTi7fmzhD8j50Wk1QffTb88rbI95nNIY3t4YZ
lj2ND0Y9Uv4ekM/e7ruoQTlnGFchljsNw7SgYcSUSU1144B4D9+qnX89l6qtWgL4ptUhN4A5xHUw
WaeXh8FfIsdgTNKCUhEIr7gdaFx9zGugbBBkxQE3+PP/Yr6JfaX/q9ywyWTHmoxbbkmbkIG2zL0a
AYITDX69L3touNUCGwzOVbDnWv1KIdn7YSOPfrMr9fVid0KpdYm4JB/7gbwOziYlrkAlbnTxn7xS
5X0ToN2ET1icRhZ7Wv5LicCFDav4XU1L/Lco51NZ01kkywp2VFAWcCw5Su2CFQt8xcKXW9MsTA3t
CUEmd5off5i0AgElzzdC+to+0VPr/wgBjMRXB+BhulSOyXtrWL6xyvuO2ozpBto+CQjvgwhIw81J
nVJaP6UM9dsoPd9LJJWgkFS1rM9c+GHjWqZ1SiQSoiaeSBMuVaGNcmCZDfs88pjCy7F8gehCGlQq
nciJ9K6ELbdJqt5hdQ0LcfeyowW/sKbNE/Gpe3XJyd49q3So9p6l7o26Du+8YGHYEXhhw5b+zLg8
GBv422uliEZ00TyI0GawR5gwva01SVVgNQ5+VbIr+h4N91qzET0BgimFiRYq9wX3LWhqYWCL9NZF
ApJLZSNc3yRgciAtaod7/gA25oyMybngBtzEGwYt9vbeZgUoFWs58ET4wk77l3nnXPyJGJMOU2xd
DYMRD6iv2PhE2Es1fik4OPcwO9QkiZq4Vuf40u+BbbnSA/VHntjYeWi06B7Vb5jp30oLz819JT5x
tB3cT9UNiFLKrEVoUVeT0Djs5r1fJs+kyd4RgN423r/oEl9bceaj5OleMagTolrJsF846d4ht6v7
DIzhL4PGyHkPCldOwGQHmjCrf3A4fuUZxiB4+MKCGF0LhaJOQAtBMYyD9+3glTlCd/e3zLQ6WJJT
MFNXwKvUfNu0Y7x0vV4w9p1SbtY5OezMvOvHSFrBNWjnN54lbNe8IoVOkEaVlxHlDrSIPJ9I4HMt
oAdTT0Fk15/lHSqpTI7TkfUREY0uh1mm+tXLVNBKZ60U5h7fwTO9fNtXUqFoldOMhHbQ6kprJ5ew
QwZKpoUB6u4UtjZ2ZeVg66TnIpMGU/dRnNmOxROfcQaM4Zb0lcL5ZYMs5erWwotajbhuUl0QTaVB
R9LJKXmQkqczOPNWxdUqDRigFPhIf2/BXmm4h9zNNEn2G/BTvnLeSWIbEHTqjLyWS0+4QH6HMUuZ
9JAo/Q/OTnEJBcH9025HilmS4c3ixYdycOiQqDYF8g0HKdcXx85e90mRJKu79y9YZpp1kDFNYYTX
Wr1yNkPhaykaav9tRlnxkNHx4Te7wg+b5v4TYDlvjE0MhlH97BS0CDW7VuPR+S/NmhLBMjgpf4IT
egd51sHjBryjDRBhcLvm9OdbRP/ENsiqf5u/XbfAoLwA8kQa8yptLvis95cYzGcdTjPmVmbtAfLv
3XjDYr3E8/luIISngPr7w/u06Ozj+4fXLJMrDvkwRnn5LH0uUIX+KU89Yu72NKBAJhQ2qAM0xIYk
n0vMtS5abqzZfYM/MMjQfy4kftmVcuPnA/Ug6ub3EuMPBIC2cBbkWDFHOZhtjE0tGOadSB5K4jmJ
Cqdb45KGq+jG/XIg6++Gx0tkV3bTJxQmOZLk7i48ZGGXNHFC2m0mm/ThGYgn+gD4dMToIIon9dmr
bdAO2ScdB6+2AzUXkLd0NdjGDCy6g/qJjZkeG8hVbX/hD1QeiYP4ENPCsVijaBMjE7TwRDNHW26K
QnnZeMo0lnlDKAmYBCsUAY7V4yHYjchZzSmw3iNYlkvS5hrtwe2IX1ryMq+622IPJ/8CcpZ8NarB
avJ2sl8s/W3esloM0+XL93++uy5z2QGF9mCcSqiIto7yG+6WMDy3yAS4S62d+3F88lji0M+AUxRP
2Nn3bnjRqlG+vI2LtmwR7TS4FQ0Wv/RnH/hPzaVFGIvbF8W4QmgYQooBN04de4HVp1G5IABP9dNv
+PkOm+OuLplOmVK5LwiQcVD4MKQvnQpfE1tpWU4ctHTws71bN+Y+2OFxJ4vGveqpALqYacFNV4Ty
dDnnrSfSpitqJZ2GMLHCRtjL/yVkzWIxbg8r9vByRrlBXNd15eAd3Rm4ozZfkngBtYzpSUO2iIYC
uSGURLkiR8TXPWheod2gTm1j4ZttlvsPz1h3Gq0PVHH4ST/+xPnkOzrH4ccQ3hevXbuW5dA3HUqB
TQa8wp3gIslaJxOAiSpZEnXRajNsCXjLqhoEMe8oDUSTUIvuMJ0z+zh1szrqb9wS0qpzq3DhVcs2
2ZpD0xCuxt1N+PKcHvGqiHM1DYsQOyjADK6PUoJAHAJgftLKav4mpSV1tuPpOxzYfc9BlShLBeuI
f1sV+81n9UAFqOtU7sYLeOghA2dGrj+fbt6fd4nIRKm9CwamKphqdgGGhJ2AKYcgXsMFVP7eeFhT
LCzzWH5wRP4T7qQiLqvtIXzQ9O7KYvU1wqf7QT8OlmTwhKq7JQ483yM6verl1bSAWdad3BpxRan6
3QPALzz+ZuWB7Krxc/8QxH+lnNBsXwyLyEFM+kCcbXAjfbmNEeyP4XvanAhQxagn2bA+mpNo8D8A
Rz7PS4LGYxajIwSE2QIGquviPkDPo6KaXB2DXpAuEpehejksAEgyoY2Q3g5kRXU9LBX7WuVPMMt+
uS3j76oGbYboT5ap8U1eXMNE7apCSFP7uLg4h1B+pkmLRuE1SLIP4SbokZjoSpXlOWAXbsE31T4U
5fL5seNKGsTF7Xqvic19AYYPK/vaGCf2gB/XMlWA0EV7y2V0gtRNPOgWZBE+CgjfUD+RBXKjTxXV
6I0on1yranLkPOGVnbtKt8G0hqEyeHxizWj3MSzMuKtH9pTU9es+FJ+4XBR3/nlm3ic0Dc8eiCjy
NzwtxETSgo/fR7KHC1WeyG3Lfj8iotMxwNAwVPwVf293aGbampPsTN3vXtlhVWhLDHBGyTFMCZof
hDRskrI60UPu9cLk88L+d81j+Zs/G6bCw9x4WbHFIhq9TYjUIqwRKAJMmWgel7TUBkriLuw7i2Rg
VqzGOP7Lc9SJuXkmyqybaZei4sdg4x+LDn+RpVT+ul/HC2Z5ZSICW0t9FLz1TtOuz5TcMyxx4GqU
+Pc4w2ixDwVoTQ4K4q3KNqeMQ2/U8Knyjk1kQ3f7528807Wy7KgFBI91VuAOFO7cIriGuCi88aXK
D4kh2asXgoEfPgB+OFo4W1FOpj+y9pdaoEAiet/XG+3kK5+nT9o52aL3jnBTU2gG82GcNTYL9/qa
k5FSnJFmai578EgV+9kmRZiJrUlgs3LqlG5DzYiAPORlWLiPI58ZsIuwBGKuRO/xWEoVvaMqOpmx
SmyOYbD79qVceiun0WCFnkZwB+OJWWCdvVZumMHUSN81QRYOkb9pB6TeWPSYbamLUwqG5vBUfVMy
jv9rPEwr+KZqlNpXikDarPrYZTog1l1b7y/U8hJ2XQsYPCfQiXjb74eHyHevtm5jHJp2vsjWVO3Z
7c2SSdcNoZAEPj8LdE0NOvTstuTBlL3czgsFIddXicy19XwAfF2oNEeAUZvcXejg0az9kXX54rb3
TiIza96hCGuTjm6uK8hMoiQ3plMxnTHCmkWXg6f7VyTC7oIWMddm9eILggvpvvxDaPWy3Cc5KCGz
86qck58Y+pWj6td9losuFiY+uf7AeNfvXQ1ZJA3agi9ssqsGjB++n0ABkSOvrTVZMh/K92xdAVyh
IQmYXDXPYo3JiCUX8/LuFOvryBdGh31696MKbzWKDD/6OgmM50SW7iIedxBzxbEzjI12dLcapIL+
0Cv0X6MBGe9GRfU3a9sBjMw+haIhN8OY6xbDrUorPzv2w1HrhH8EzSTzKyENti4/JWnWN3yp/tCc
vaZK2EuYuJpCYOf2T8HUttA67pv7sfgiAjLOIxeXclcHwN00wfLcLUu5yrsKdrHiPOGaWH1iykaL
ZeTkJifWa3c98tTjzefuE/fThp3T840t9G+RoyR2eoeECxxrKXSXI6OS1JO3J+JEkn0cgl7ctKni
F/bLj/duosftqe9mbLmu7D9jtVA4rXEpEPHHod8D+D/wswB9FWF9kYLb6kz/hx5ZTdcu9eSn+mfL
OsZTHYrBnemL64TIyv6Y/gtJxEdi8ZS1NJODcwboC/mlZ5MaT0PskEu/Wad2KlvFMspM87t8drDE
dtge9UItJomgLYs+UFzx3j9Wq9SxEzILogGCd/Xjb6vfnazw4gRhEWc25brIIHiKGaZsb2Wdzucd
AvMbGgt24HXyjwnUkX/xOHWMKTPpXWisldlQ+jxxEKEDISr7wVlDBVf34cFYVnybbUv2UpB2LxNl
KchRVjsG4M9P9Lq3fvQzRTBiAs+SKjF5LeqGgGla/n9Mz3b3lGtxKo1MotejYK7VQU6BX/CvZBcW
5BxWr7nYMLN39R7C9K9JLVtbfKnqn13CcKh2lix7JrTGlq4dFsCQMzIkRXD5MCw0PrtSnYQefYOG
o3KgyO0zJw65qxfmgKGYtpb9ozOLK6Xmwprbp5rm7UFbnnTsHsshSuFVHK00wbwwJtlFdtf0or5u
XBt/vjB3X2U0WDVkAFyA+8NqOQ6dR01ErXYc8/EifJO6w7mrCMdQprLYPrJfCaJM/AUrKM35IsR7
JB9NRMDYzePuKwX9RYLGew9y9QcQ55A8QqT0m2PCVVLpVTYtWXQE//lSipkdbGVIWvoHe0EbVtCJ
lwfmX58Iz1p0Ew1DMFurOfjudncpkMMPngpeEzCteGWzp/EQe9SLLJ26NnzjjPl+vp51qCqBvR6I
+S5bMe3U1on7G5NZ2vK7n66Q5Aqv2ikMyAJ/D7pYhnDmae53yrp/IuENU381gtlPxa4qP2T5+Gqp
Spy94zxGSnh5yvSeIehTO7kEMU0d18/zGDB524ZC7Nvk/fUbg9/dUa5MNwTp1rnZxMKkJ8jkTLX1
uk2l48u4SxxtXxYcO9SqrpUSxcZjsQL31jtc1vEYlu+Id7UkgokjEbN2KY99Z8haDr1NeVydEmPO
0i4JGY0aSGNOCI5NPZmMPkg+yCO1dRCzTXUnQgRqr1W3xZEbHz0lZi57XciwMG83UL3Hjytehd6D
mMSpLjFkAs2FF+/0O3pd8wTTyaU3nm3XKgo0dAXlHlFq9pMrYifbMDJyWsQhGsITsOU56b0Mi86C
0v+fKJlVU03y7vx7JePxMlfwYzxfvsPNpyaxOEyed7nmsn8LSxe2Zm2JJOAY+HhfYEGanTAwghpp
6blaxcZr33CjdrOL+AIPiHMF8gdAZTjCdZwdqkHJKRzWOHPmQ55ZcQ1TbNpiYsDYK7/+UITOrQ6A
51AmBpUyRFmRFbcKV5wZqrYL2HQ5QB0u6CQ1syQYpBcvUrILYguDNNCqyDI+awGq7GRe1y8im+Qn
QR501k04/Emq0/X+IKyQTo294ug36/rfM6OECmzvVFJjExOTuCOd7AmLF2sbR7TAa/OoBee1XRiD
/u5EPZABVJsUB5HVfy2tSizMwG78Z0qYgFBUMf3aTKsoztSZPf8vAIjGSXkQYTWfFC2v+v0gWZgP
nAROliAg+92k+WeqkTsWyy65qOlrL6o3xOFapr1XxRgt6msMg35SjUNDiOgU8UWjCy2m+C6y1bZl
g7ipaJ7HHAYvESxw/qmFmYNF/GL7jvgC/SeIHX1e19lWIjlyVPWkJSjzD0uyJjAoB4pQx1SWGtDA
2V1jBtpAE+/ALWzi/rPqPcRVY3V/1VxMZlqE+Y8XdWXazFXgKEUgFLhGb955+zcmpnEIWPq57v7s
p4tCsuEyhe3KQ9+MGotRjRZULseQHLVTRzFZusNcWrV6pSlG6C/Z+W6jCCbNp0McVTwgAh5BZPjX
ikugTvwRWcgbx64XcGn2JBz6MS6lnW/sCQqheuNTs4E/4DErpThx7RKu9jjB8Q2cg1RKyXa2s1Jr
OE+iKe/wKNm35rCSIcxzsbrSU3UpN58WxChoftZidWlFn4H3wneGBbkhk4aNdMp3162bAaVB2DeS
CKmLYUfF3URQHehBqrurdMMApfMCU9gNrd+fBp74/0elFydITf3NZVzm0Ur/nPRfOciL+RIL++Za
MOGGcgUMcVQTZ8q+21z5zeNf7WLgYLPlXzP6vQPMfr/3Ih3PJkjpoQf8r65X1DMk/E8xSFelf0sC
5B6Q/klwzc1MJ5suo3GcaKJAE0ZJmmbUYI1mWpp/kkBer8eRD8oBFdKAZs7UWpaf+D3qjFWSAMdh
sFZk7Ui9BmySwRIosV6kDgoMrlgaLiMzTTFiAJZEg8ZkIr1S+6GnUMHsnuLXpGAzF1+IWyeOtTRV
XkCrgT4tQ3/xzpkh0m22knAALLjHWYGhLl25RJfW/+0GJMCt7v3hhQi5lopmMkdhg3MJDkmNxhqx
1qwpm+hxVgwrVW5v1ntgJDIvygzZzFjJytj41ZtxnikdKr1p0WTGu3+yu0cIRi+GwbqnXDOpiQ+o
U6xht4IAUHLwlCnpNuogk35v02FvMrX7iHttyrElJRRLCmHnEi5Xjx6LzsNh4v+MARQcjV1aB3Px
gEu7lU2kJYTwoTDcy1T6RURpao/DNKPFiaw5UkWTtP/Os5NwJJas53XHhLF+Ms5o9fEfcmjmaxjw
0y9IxVl1wuEfHCBvO5+8kHrj7Zh2wTZBm6YtbtYnexjJ8DRVraN2Vo9oFFAvEZmBnjdioe8r2h9s
b68ksm5FNESzrzfCkTyS32addcdyLN/l6jWuTzdbyP/nosTb7Q/pY855dng6jSVd2tuyqq6YmXNi
je0t+lNbE2t+l2fUiA008bziy+h1Kk+70ftZ7OgT5L+NrfvAnscC1FhrPf5uraq3AtbuaWNsY3Zd
FrsCwPfIR4lqRfdNdUkn0+jScif3EPqAbXgAOKWj6ZOkd4s1dFEZ+wyZYfwqMCCxXDopfXwajUw3
U8pEXTxFCcNI4jWOT/nXoqildZasVmJtymO/fP+7wDYaxRqzjnTxjRUJx8bOBsfapw0qZUG018F/
tjVmnygJjEiQSZOpkcuWG3HtLZKaTYS1zRv5TynJEbFGwjps5ydS3KWg7Dn0hrqWNiobM6bR+efY
C4tXLCAKIUHWdFUbsvXM4qEugTU/4j8KBUmIgWB0ffcQO+RV57kngMHXl7vGuyA9cCxIx9l45ocU
0+1A9wL7m6oRY15Q+huffEZ49+GPF60MfC6K2H6NsQDYHDkrbPv9G5CNx3Tqg2LlirxdqtwgUaSG
npEIHzp91LTO7aoSddjz+0GB1RfWCprawWrWe4vi/ycPrIZLlT+bKHTlhShCBzBnB49p1KcqV0Qs
xfjk8ssPrpf9cd5+t70pSML5PQpAX3XJJVO/zZ7a337/PQkLJgmrFoOmQsIqWzp1TqPlV9PV2Bjg
VhvvqAxct8XzwJjP6die2Bt68jtcrLEvSPK5ALQ1Li+frzpplCEdPoR5XXKjZ14EYIRJIcW0KH6U
mUEub4yugX0r5yPVvJ9kSBXgLkQaTDMHR8EtB/T5M6UTsTe3otULzyd5w7AMeUaPlOyXWXv8b+4j
J8yNkL3wjuYmwpGEZGdDMr5d9WfUhpcVRKLmhgqltR9P+i2+tZ+IderUMPTmreQ37or/LfuLvYuc
kSxs5iQsyIRbjghFHTvRdmloGtvalCShYbrXue1ui2yfhHlf7ORODcf4HGCc7ZGZga0NAcSqjkc4
CmQCoBTj5BOuu72lGuU88xDBtnodcoRxqyUK155qIOgNCgAhEoxQZAQ68kYG0wpPAd4sxtyszRjE
ioRWmpi0gU7TfKhJge7BLhHsO+Gw7K3jDe/2I+KWLdfeeGNlthHfyep/dP2a25y8J3YVlX23sz1b
PCTuhis82SMUKLVvhOM2ccyEKqEkuXbmLLr4EaEVQCwIaBYYyy8EUv+Q5eIGxrBl1S6fQHtznrpm
wDwar1HGYnnLjaVoC6qko7P5VEsiy4BvXf5tmpeNBuD2ynP79v5ZgVt4eeuQjYnX61LGMVYoEFSR
bUG1zyuMbvZC9CAMoC+CnScm54G0jF4c8nc9XFOSkEnV54LtmuP6hWE65XNTy9YGll06DW49EsTW
q3MAKakmGda4lG/YZ8xkpiGHpmTi76NSWSm/3WoqLOMBUiH8F5e/N6N4iO0DlJYeam28EM6pmjlR
fCwOPe2JP63d9lSzpLXcEId9Vjjemcd4Soo8+L/mlzo0Ak6D9AyaSpNw94g92ZFX8ux7XV7zFGFF
Wd+f4jl/9DPa+A1NE9n4+d6fpukrfwrKWa9dnsFxcNFdskBp1l6NcYjBjbP6ZbS1/z1dPc1r6OuK
vWa55mY2sqYZp+FlVGOiqR2jZr+sODoZy6fjbah4V6WUWpFDMgn2+DFs/6EQ2C7Qx+ZxDz7sWMkw
V+a9q3MUH/oPrumODfDY+wCU1mzXNNBnZ5fUb45k0DyNjRP1jTCuLyzDwRh8MSwaIebM3QfwDKio
8PEEU/jaLxWhelm7lLmcWVT52ODAlK88BwOTRbljEeUu3Ow2XTSNrGcSeXlEPefGtW2bicV6bvoO
CxLq/WJnmHSvQ+H9cpD7mAVKqnEnR81gfAt/VSkLCB8AoZ9TzY/xLtYY/4xKuiHhUXYafUDoPRfv
FVxuW62fUVfsS/Ern2KwM1ENnsiLdlWBrR+YnT/yCUJycF297r6zoBVv7cMkEXFFMd0mxTMen5bw
Jisfd/DUF0OGn51Pja5uYEGD8PdvsY9YgDHoKVW/IWDLISBWMsYXmONoHD+WuVaHxXhNrtbYm+tW
gURhhJJ2ZFoDfPvhUiEcVIS2yUw1+9IJF04uzCxXMALSyyNUvKj6G8rhsstYWVT9Z4mvWCFJdXqg
pCD5bfM9AHop3tyBw2E/S0+q21zhenpD5dAZZpkZFcZl6qVsMlAFJZ1srtldRCVp8M/PRHdEaFG5
fW3ImEVEWGHcL+hGW+YZ1MxX/a6ZZ1fEhoAsGR1iihNzCj/mFllh5l7MLc9lwQ11thExJZrBuqVN
hLC/6cYdlPidUIeGsIKeJ71KcNt+Ve6tf6V3UO0dccOOkgnn677UQ8gVkDz/PDvWaMxblpSTDHaj
CcG+CAZrdpaIKvGXlr1lVzztwQPbCiWIHYrn4c1GiiqpJ/voQY4EJ7dx6Ql15W0jwsNFROSnBWL1
thpwvp5mzgLqRQt0F7SymKKtEWLgnrISfvQItZuX225MeQEXasP+j9FkJE9bYfbw8p7/YQU1/wQR
L9cfFMfIC1kmprAix7I/JsX8pOi4VpHhjSXWEqPeB8qKLuDv7XWFS1Y6K9xREG55TqKhRtrw77v7
PaR3b0nwUObKx4zzWjKadsq+PJ4gcj/2eyySGwR4M3l7F5M8zUAwInFvHBfw0+6D75ZO3VDU+SMm
g76r+hwXDc3ectSF2lApYBex/PxZ9Krd3SvWzzTGmrFZYKc+vhIltQ4deRmmAUZDiyu3DeE90mRP
zeW5H6KGCG4sqjYoO99WxhVsoPxhO7Btcov5kO3rQyCRgAUFW2Fb0tnWCjUt4EbJxG8S28AnMWzN
MBWWJGxWePdXHUj7iYtwDYejwzG5bAWgjxKNEzSBbBKQGI5jr8CciVrz825CNRv4J3oudhcAQ07T
/PAldHhb090DGIurf1KZ/Z5VoXEQQJymOArelhaXWzgGWtFHVgpYMTxXiHjW1hkyzdZyrc82AwDf
CNZI6JJH83KCQmVBEk266vHEr8JOSsN7Jl4MYsd65DKKErq2UyvpfquYom7+i6yezS7R3r/pHJMK
LB8BymMsh1YIyq51NUcRwmuyr34OiqTwtjOkMwu5x5BEo0SEV8VnIAHg5iESFMcy+UcPRuln4rNk
1S50fKdnvYSsCXI7Zd9J1/iT4GPPWniHQC/nCMZw9NGP3arVrY/ZsQ+DZU0A9DQLBmR3ZsHnfbtF
BdhZAU/HU1Vf0klNDuWnItme6EGlaOZ18zu4ttlUz1taC1SwvRilrSqcxFN/nbmlKCItP6Sx4Jz6
2/k0hEHIFzULrfI70AbFJi55DzM6WPYfDARG8B5b/8mBHvla2Ca7WFmI4VwlGcXApAqxInZvnVkq
sYT3XY3yLc7kjCHp8C1Y/Yb4ZWmmHCIJScnijpcelMn7+ma2RigfKmw/4buBVCs7aJzhnuMEaRiQ
oBLD2hSPU9TuzraybHhE4McyzoY61HZ4ZMEJ0Zam9/i3XDRXsKUXcAkmv9BuSCvh/8ceDdKaX5+h
ka83bU3Z9hQWJzSgHQSjjMbrOZjkfZECPzoKtdLOOIfVg192/gWhepj6KmxrweR0zfHyxiE68/qX
TBzDVwb0UC6nKIb8f4UM2hrG3fZMG4BmlMI189upioGFqFLNvXoSMEBzeCJR5XrwC+qvq5gYN2CS
pIyyLeeQyC11+PyeyF6Mb8wpbVHJjSI1U5EKlZAKanr/4MvTPSGnXm3dtwLh4EZuYI2l8OoWUXvx
mOcAgupb8GewKQpeD0RUkABeX1WCPYk2zhcsLSeLN0nITMUg43Bl1POGK9kzNuU7+LLpKoErbGQH
ilJBL/FU8RrAASyIxKrdt91oFyqa+4roQp7HZZGsVKjAOXnXY+abIzX3Jg+lpScKM2iiTwJMhNsO
Nv8PsMHG0aBSVe4vOPhEMgwTQhD2uT0EtuiUfd0qKcFTDdquO4YwwE45mm2XScqR/F7QPMgf00fD
HKORXOHEelNM4vuqfKBlU2ag3+reHn5X4GY90PZkgfZ6rJeST1Wm88H95toZE/D17v3Qg8fMZ+WI
7tetVjTUGnVd/mh8z5v7932EPAMQc2c/c2uHl278b9HUEBtHyFfEEjsW4YniPZYJqU6oeW1cWGZU
LgShWtaGP93rcDyZRfwouzGbNM92lb0u/p+yKqRYWgPe2gidIFNHPvhqxMCE+iL//bGUwdlaaWcI
cntJirJb6xeNiwJUXf49200sIeT3ioylVKTiGbCZVeMqfl5ybrv5lOsnMztu0h4eHtI5X5RgfdF6
slfS1aLhRo7w1sAplN36Jz4sXIlrJSS1kfY4V9nng0Ok6g8ExX2ImhhcW7nG+15Z1C9fKFXTzf4d
p9BacOU9TZ+qlZDsOoZlN13D5W0tgv8HAik4ujdJdqTgit/MV6T72f4mXObP7DUUYdFUudWR/zLd
vkEKPFUqbr5ZyfTZ0mdxsjJnUvY9nh0PKs2B+5P30AzFcRj1aWMqwcJat2gZZg5F5eD1jl/sQgW6
HkWakXh6c/6Hx0nAY7cdOrc9g1O3/Qj0lEKbFWMdgCyLulI7xtBdMyUq/WRCMXfQE8muedhMB/0F
LAjylgcFeKn1L5r6ZgdkwCOqHw6XmhfRZRdPMO+WJXQIk6AR9qdiFARlAY4M/zyCjGrJD1UL8fZv
51G5AzWhhoGenbQ746eTbbs18acSB89GfXjt5/jS0+J1Qa8a7nj//4BfeFd6EfMvxXlNOby1RwWd
wWZu0XUeq4tzMJEdfNqp2WV+RmT1XmknMuoXfTkKUV68RNWjUgvQtSZeypHBiwIXE9M/vWOFFZ12
UL3R3WZqL6v3/BzkvCxpqxr+VmGz9eq+UEfxpQUQJXWysv4l7NIxNJ6oXQmV5KO0L49AUWqWd8Dm
yVOYUJ3dgXroSpXyow2G7dZhqSIy6FajFNod3DhqyrrFPWYtVVJrx8yimAaqHbDalpwPKPEHE7MY
B4qF8KFj2ZkSWlLF0qmvH4XTsAW9DDteeJQIkv56NLD6Vqee2I5WlKbgd9+ZWy3XDq24TwOHFjeU
r7pc9fU8T6uKfZ1WHdPjuzTvG/sccOsvq+JUEz2KkTs/b25YYLT98GA63IvY20l1S+IQ31hFDTEn
r7rfmcL1v+ggbj1ROw4P/l1eR3/S7N5PQWeWLAT9Fmi73xACqqntk6JnF7ozhcDquZlR5+M+dt+/
wKOWEqKqsaYnPqGCZkFBuTHSNNCZWFf8zXzpsqfQJJpImGhbviNsa/W1MY5EtonmdJTq/BTnjT+4
XQg0CWi06cAJX2CvsDHuLdIzlOdK7nz8QWJbUsu61ci7cd4tAsyk64aza4K4SpJI3hq+3y6KPiPd
LE+BEhDkF0VLVFXxtVk/JiwK+PXJ6H0SSYCaC2RWrxl0feKovQDDdiEgMGsKtqiOIG93WftuLhdk
8rq7XHOTWft1SqTzvj/K7hUktf7gCX0Fu8MzXutsqwI58OfVtROuBd+MIUfklDH5H2FoKWx2eLqx
rzh1QChvt1DRVBCirF2mQOgI5gmYQjgC0+Eb6S92dB3EbOwLR4nKMZZ1z0B5yhLFCexbnR6MJ5bP
eLJRwjXfoILZR1xJVV86aBSJHbWz7EBwhfxH0o2jAKgrShHb7DHBfKce5TXLLOI9g8dv9Sh6rpAV
YBr74i3/E4CZFvx/0hFVPwYaZ+cEcLJO/h64kYnAHuXLVq1CMiev7izwkznBgXXir1Hjp3I9XDxN
3VFHxdYE8BrYSnVyFgi8lAJgWP9dSFgYpfDVeUopTXfelqKbqbpxWcUe84MzJTlR7sXZROy4fNDH
bF0hoUfzDsOqKnqVC6rqdPT3T8QxOFpCUaRpoUYj+AKQ9CqT7g6c/mBZlsvbdkez9yQi/rSvSVjk
hDe2ROv+NoLEG0Ezs05PVGJitjh+O6qcUVlr+ehHdnkJxekCbUozNPyAHKsghwGNEK0ukE5veUrb
ybpDQc47XzZTDMU0aecdfYKBa1ndJapeS7TpK6GJmpEMHet5I25/j7hKjgmF+B1X/A0e70pmuog0
nrkWPJdrxe91NLYjX5ivjkEbd3d5MmAaxl7o0n0S6Jp23mLXhAfX34nhnnafFO0GFCyXfVCaojO4
5BgebEO1sVmrg+c5yT+RWGOrSmW2RKboLb5Udrq7RQ57V6O92Pee9qEuxXMtylk1m1/RwC3HG37p
/hwhB6YuvptABJ03TG1aNOb+Vd+1dnVzpBgeR/GWV31lsri09m61o1g2Il/tLIcIuV7nBoeVIYtw
Hrq1zh54x7D1a2UGa7MyR8WqYYgDUkhaYrAJqO0cJ1J8a6ve8hVMkP/Hs12iCiphNyoVrhRbFfW7
T5/2rAOM0WbwDxIfuk8bB+NDphM41D869W+HBER0AIFSbLePW4Bu10skHP4lRrvUPc+rXurIsmlU
dlCWfXd2lmuRZGW2w4iJAjQrst0MdSoCaZae5MAiSJJQ/ajrvpG7vuB3oI+lAIEGJWa0dTM2+5DA
RcgNbyVA3t9jItNcG5TxS29Ir3CB7YvlaKT8Ft5SEhoogZqsAyEY2YA0YoM7SRDKSbt7UOuN6kKj
PSprAa8/pIuqk2nHsMMHCIihDx8M0JRXWXzB8UKql47GULdx14XCQt5cO9MOuZNSsMoXyqB8hvH+
oeyIRrlkFJPFzXU4BWFzI4vI4gR6G6lCVDGwveWoLD6SuXJ6PsFZDVE2cVzplFkvp2WFO3kRGNPb
tXG5KtQEYajHsLYHPlS2uvYUmhwZ9vbT6AiWOwiEHMyeO8CsEQMGLIbAn+PNQ/BygxORh5lvGbfh
RYXAkFqWRKRYouYYwJ/KE4zVolYAwL6+MOXgDfiLwybYbhFefI+lklXVKZa9mqvK/PbtyWQNWl95
uSrVlO1XBysIosWHOdpXW1GHZuKlTNSgYYOuoFr4qU05O8EifnaNgHI0wXIDHwy7oIfMC46c1LAA
BOSocjINzf/gdTAwzE3C1ZBSODzt2EEXtHH7LhEuqENe+Cdx3cak442iwaj5ikqq5WVH/lAiw0Me
HiBTQM3/44CDj2xeZ2yDQg7GI8YIWh4V+Eyop1qbDuK7Ql/v9aO5zH4FZ3zInuBfvl+kK6iA6hTM
3ka5wQyYl2GE48Y9X6JM7uXVLdFSv3HeHtVXBmBAoclmEDYuJcfYD0AngWWJ17mZp40c2cdlBzos
qrMltBDQyrauebFN8+NxRw4tIlQKcdTKedwIlU/bnJFLunf0hYvqdB12JGWITJ/nymsNB/NcThUp
etIenSmb2z4XxEDl1fgND5DolCoBKTEKIFhcLQ4tfnNECVIZP1/BUzAKrWeLWHswXdpzeKucBx2O
9nCJNoaGO35pxIZDVVQ7qRyqP3dPsDkKfQ7qHFi6SrWEEDac3qlNY2U2SIwo5AJnadH4RxIGu+Ne
H1HRdnafWdYRfAa6uiopiXMtXP0Hs8DBTMskK6CLsC/rwneGyx+SkBZSTGMlsLhSs24tbhXhD+dU
cqc0KLhYA0z0G8T1aiuN4OXvsP3saE+YTaiKUBOj6gwUJeoNm4A50chAf8+rxsDmgMPwzvMk0Lti
mgmdSKaCsc1Bwj9AykJBGLfE/l2dA9mJWHKgMyzaiClpqzDp6BERyjYZwa2PqEz43S0zbvuYneZm
r94/RP8VC6vIqjLyL/x2G/EFElJ8T04/iBpsf32pVvDmF0tr78hjs+GLjZf5N3Jq+J23SjYLmS3R
8FSATknUL3SAd6KSdLUgEhBsukcPA9IHIOCOyhDpLxiLMfhnhHku6tUWH8aN7Oe5P7Z/oojVnqC3
Q19utUo2g29FAAJ6Z/leOA4zt7fRFLOdNza1+AGpfhkBp5Vx3JEiVMXENWlqHR8BoVhB83NVsPGX
g1wv6LI1dTRvDLmqVBBkE3M1ZB4qxq/XsrEdhdCfsyhoauvRNQe0Gu5wqloAK1Qy3/e+5w72wQxj
MatfrlS5W9v23u43/RqUDRCkAZ7Z1YLqUo2Xx3eCo+VFpLeeFL3vcgHITzGVmuVGI1tCTOBFGxYt
+6vTRoGgRq5QkXUXWo8tqIGaSx4c0LYkO6FUPjF9ZLSv9vbCPWD/bFj/PSktPaL3qx3e7nwhq8ec
jfnGIdvJW1O0H4UhtizI+3Hr7ODL/R9FoWJ4YQydC0vH3ZRrWf9A0Zi9xvL+c/WEcSvF5zPIo55P
TY6Yk3rwW4jwwzNUeVF2ty9VGaE17M3AbGkugQS8awLV1WQ72T4fr6/Rm2Eco+8mfwTdDUxZ4TOt
HBHElmKLIFu0C6HwoDtt9+hkDHpj58JZGeDJXw0tzYDZhXBMrE3RDiCbNeBnYo3G0b2IknCZYlgX
Yl38FptT82EGfRZcNpqvmloxocpat3GWYPFOHr/9zcNAurzwrOtOdfX5jZZnW/Hnagn8CpFc4U2E
2qQDI1w3wxTabG+L1lUfoNhIYUbYscm8qaPvlrtjYRqaJ10wlMeT7hAu7YGNgDpVec4HrPEVCL6D
xoRgRzjNCI2p9OWkeR/nkkWVrEJkm9zWcICg/b3OnEt+U5zTjZqoss27WoJfh7sPXViT0C1tOhgQ
sA+GfkyQKYP/atg/nw4mbu0qXl8UerUUE+TrlM57DzBb8vW7lWbLj0NSBprV88DwZ4qxyeQA1XRn
aqVCF8OdpCM0UxtRaWrAx2B6sZKXrUkB5N8DPAUCJ2sGS2Uxry5DA/IGkXTAlMG4G7xy34WCLZf+
QZIQTiQqz/tAo3MojUXlJ7XkB4k+jT/HzfZ+q6potlm3mrSmkZ2LNS59o8Wo6Ak4eAB2Q8FmkjEZ
q+cb6xlEgg9W8x63SlZRPKzRinUWudaSttZcHzOxgSsyT6m84BpC+uXSAvl6irfbW68YaoaB8pHO
GAW/88bJ4KBlvPy6JQO4FuB4fdz4f4jZ1CN5jFFkhsfkK0Domt+vHp8LtIVeudx19BvD9A83Jk+d
O2g1YGb1U7LNWmHfOC+Q+WQfYzm3Xp65YeqZHD1zH2OEsTCDXasn0T0NBupgdpPGnEuVP2nRhwxT
DgG6FDJ9CD8sYCfrRhxqRB44uWCX04JNXYfdLflOX3D+pAB72Tyw9EX9dtyQdSc1ikXFIp02zNj6
Wj64QWc9gc7J9T42AYpb3YZn+/hj/quQbStJeaiHGUyIe5BnldpWgW8qcIHA+Hyw/lPcE7EAUM3T
HhHjEiJOD0f6+6s3ld77xGx1yHu+tUFtnMSzTLJv/UHT7d6mEudkKXj+3WtFrl13eplrTZTXG/8q
MRat/x4tRfAdgA0zAxhfCykrzZt9dJbz4vK9Rn88TfaiEmBAPBi80xYsl8cwCv+h68OAwbR46sPv
ATHOXZnklB3mYtC1fcbNyTd2RSQZQq9GB4NRZS000TPMSc06RFW2/omTApFi7DMiV+kVlL6SgaHz
Brj6kKX4B7lMc6CNI1ZSG7r5eP7O7Grf2tYwRge6bvp2+ZPoYQ11Kda9m7er2m2Ye39MbbBnnzUq
2yYCMRr/n4WqhNe4sg7tn5H8H0hbOc0uG/35uX9ON4wzehv/BkXKgbQsrnio94zhQv3c2BqlJtCu
j9DOGG9EciQCp2XRmOrpR+I/qQPha0FTnQvb5i9QBQWqljZKhx8EHr0zA7I22B972lWe8l0tVJ64
bpobubi3TGIusvcTwNGBnnJu4VhmMuhQVoy0y+8EhfwTIhY7G4PN6Hd9ERfg7WZIcVbNlFTDQpZ2
8WMliz2no9Unemf8KDrrHBy3Oot8zqicqI/eTLbkM09x7+OboPkty/LsqS4LcejKtrQrpA12DDZC
DZX9z4oDY3GdQQF1ylvaJnHy6o9v+1bHeDicbtUn9MfYd7gLVQ6pGpwwvhhANCh8FqFNG7Aunsb4
vyX+uA+rdtFEme/PqKqemCV3eEeQPe2YdV9ZOAhBdhRvMDUK8sj1ag57nVGNgK4enS+3ytHqWRa5
jrMAY6X8/o9jZ4yTJGaev7Y2JX43Dpva4Lpttpd3CE+iN+yyetP1e+MMjR1jQAwxaAZuPoe8uh9m
a+9u9NFmNUxan0r0DO9jTC2GBMylisCrdp2fn/OTFNQzP70oyGUpKhAGar6KfNvdc+IJgnaLqe0U
82vIfkQuujzShBCKc6WkH4VVN9Hp893nt6/Ha5dAEGW7UYrMMkNV7wWBuPRd04MIqtB66jT+LLPL
oOCDP5koULHGiI47Pul6YOD+2SlLJVjR5u7cUfU8xTwhLuyHuHxOmofX5uYetrsb6+Kbc5fL8Zl8
uvYMLCQNx8nsKtXhsHyd+okjS/O5Rn28VQiciNbROsYrOT0pIXz1v1WQPF7FADOvUhm33ST0Vmh3
jp2F1svnbkr/u+n3qR/xFj8kqXzg0h3sNOZ8K+1BDazzAuNzwxsbdSMbV1p7RTze5i+HiG75a7Qa
UhV0lFXYulY/LY4LrTIPC7c8U7IoK5HXdbaYC7Yar4mAdwYOq56RpELGzmLBzoH0JIT47CXACoLr
YrKvyjwWMEyGtQOB5owEKFCP07g+BQ45OUkP7pAqWgbhIP5P55rOlJ+QvZETuAZh+nZSAgWFBU2s
627IP25FDEQjq3ypM27pc2Kiq9CJkH7nix9HpzsUVe3sUYWinQRE5dAaRdo4VEMwpr21ceqGFdN6
TNaLDW7ihBvbFbAzM4Roz/5DjatlUoFX6sfFeRTVmypoC9TwraPzRY9fdtJuxGgH1pQ2/ozeT9aM
LUGxDYQZw34g3v1j26/Plhd+E0jWEpx4mKLLroJ7G0D/S71HC0uLw3M/G3VoTEkdp0j91crmb2pk
YaIx6u3FzdIx6Hiz2ku7ud2X/CIbxo4Av/0iHs1qe9SfCJ7LZlxdp+OH3u0Xm2CIp8p4Od+FJ0XP
S/RfuYiVwLoyuE6Z4wlN3XPN3nPJzj6JlJzTtCl1lJ3WIKt3HfgBD6CVIgEU+YG2vfa9kAvwvjn8
xwbnEKFkLsqHPN+p103E0gUeviUzg0Dqb03fnDw6+twgld6RO/U9HE7QC4nf4V8VyjSLiGEipUUs
r8x9HRQhNWQej/1sK5if0RrAzg2ZVt5RDDxn6t5qtD/nj9GhmVb9Y6oMGRJprFde6SDOElmGTbns
dUITHpTNC+ZO14GcRMgcK3SOFtQczYJNQmSwz0jTD11zoos4TCpPjoBILzf/EvKV8bKO428lY+1H
wqrWNe2Gq5JhQoEegpngtrtksMwC6Ww54GyZYeYTG4xz6DPzZGW9wdowYwAFwA6/N9Pwp2uo9xjC
Rg3OqUEDFTkkFfl7JCtbpx4++gcQuJttOuEk6mpzDpblQoEozxWcAmdmq7u7IY3/3KucAQxWVr32
cdVfgUaYjP9je4fNNL3guUNCzv9C2UO0U2ohHALiNEwn/cKihqmm8/1gz6cSPvXjsmhe3Y4gQ/Z7
QPwo1ytHZpjXcWQGgcWB6KZZTkPrVvyXRYdRE+Xy7UItnLpge9LHhHTYr7j92tiGD1UNoXvxTbV5
lveQjkFREZyyKEnXYBc79o3BmwoS9Hf5gu9fKgDUKfNFJXpUQFrX/sR0N5youcILAfEZBDDJ8154
KOKUFuDbUI8BP2FNtQcJev4rnCF9eidwzlxKunv0hVPiBRP1HDbZiNFnDNqCiPKbIyG3RbiuULkK
gMIXendETPgzgNO33o8/gSLViTF4IUUCZExRaeqrOrSmGivQshsiRUlbqHM2javkKb93lBzAd6uL
DNBD9BpNdHhVn/x6Eh9G01cWhjWJ6K1e2olz2UOuEyh9nnUSblTdoEQf561SWPnT9mfVRK44Bxcg
OOtzRuSagY3KfeK8uI1IrhIxsz4HUlU8HIyIWxGiWiOhnW3dpDDcht7COrrXyECDOtF7xtvhVu6Z
NTl8fH59eGElY2j16gonWi+y6kZFcREAl+WrHY9TkPexRLGosUXaXtB5/pSYfeiFi7KlS57PnaGe
0PE8F2LyqDbhqjP994OczeZlWJIru0fu6YlbM/kim0PM3cmYb5n64p0ZW/1D+l70Oj+k2D2+ha9T
3aEETACoiV1mFwnLMXflOBb+EQdq6i7I+ySuI7e2f+aAW6gr4Igv93V50mcb1T8krMAScqBDUbYL
8PaZEgHKsHpBw8ZSHSzne6pNVQ7bislB9gVZg5UU0etkFipPcE1RBA2FCkhP9PXAOc2i9sx0LUtk
6cizK7bu5juCTieVZ3Oktaluzufv7NjyZCtppSxeuAixqyv/xPnZxhpD8nn9usX7G8pFp+Ds6jX2
0LfAvxvIQvKq8oht6B4SdwbawSCmWtZhk/uIjOWj5qGmW1N/edZnHkvDR0Ac0RQWnp50Ri+OFIdZ
w+sydye+7m/hS9oywQEJJQ5uKQ1bihhIJodfK3TaWxA3/q9YUVq0dCq5YRaDqMWUbVwooHvCDO7E
KerAJHo3ZxAe/mJxg7Xii7GeWfmlZ2xsWhekdhweHNqvGGaoHHhYtnIk+O5wI/tAAzc9nx82S/0r
bD12XsUSPAC5Hmc35SJWW9H1gt+dulizvy4IhPHJKnyOMr95HR5nlCA/pY0B4te1o+ekIjl52XpS
TajSPzCnY9AbSji/8GI/HdlaQvZuP/+0Yj+SLtmfVsdC5mgwdMwdH2qVSdYdt+lz+mufZkpijbcq
hNylZzvV7oQyVlDz20giIYQi0yYOvZJKx0S7KmeSoQe1ac8/QnjiZurCJ2go61Y3F17Zq9ax8tAg
5/WDTxCQNm8UBlHT3Le66QE7Pvow9AdYA4QZJ8O41xKc086JY6nCRI+ViVprhs9P1eZxCHMEl9bF
hcuycErnxnNpgQCAiH8wZpKs/IAlhvqVgHUa6uVGS8VD8Rkt3CppoRsq0IN36kxLQfKYSzimpUDy
XdEwbFOfdy0NrUFNoy4qiMYhn1Zhg4zbrBTGQhy3wKy6Tn0qNcFZsfS+4IpfQxlcQWyqTAwSt/Hl
8Lv+oGRTV1RYwZ1V6Zy41vE8HP2KgvwF985Ws1+FJA936ojVMpxnxNepYHp1ntkLNiWp4vCv48Y/
ZVqT/tMcpnBUB1XernrAp8YCkBvzqr/l72yVfhGS2jDw61uaQQK/XDR1jTZ7HblaTNP4qwgJleJ4
CB4qXtGmzKaGQGguRteESK5ynm10Gy2frnnfYY8KD+u8fgPlmo7/LuHtfKtzZIuKM7KlLHGEsbH2
4VPGUlJLujmUeQGr4oq0qmXNx78cvl5sDccEDpCo8xYJieqmQ4WrOZ5I9srX1NUEvhVkmGmoSJnj
XEWOovEnmIDEx3FqJIi6TSNDczQHT9vTOOnwaYHX6db+ITqwW0KBpxzZk7R6SjcWJ2Fo3XU6D/d6
iiJI9w8Dix3q2/9qcsx8jy+tk/ycnqDDh38R0Y4pS78ZxWXCbn9iWIY/6bPVZtz+hTc7qolaXvmk
wpdPVJv/u636ZVe60+XSnP5WiXWoCKc23FOLrbuxLefrGGLmvZ+HDHU7bKapozNR52MBz8EA8nAt
09iS/XoZy1TT/LkyAsfo8+ZE+7nEuqwDBPuXWPA2peHOkKlZMAfF10zVknza/8eCw3VUcco0O8rH
dZJW2jKAsD3Gkx41MEBOhBFjaM7+g0U7cKjMCN2qMKUvTKUYXxsnV9159GRSXGsbsDJxllLl1/zC
B9JdFrWKMHNOkFIErIYoCQqI/4/OArv5YNdo22vc56hIRtmj5VR/f7AlH089MqQb85xAofba2MJL
EGYbkFyn9Cw52vS2PhMtFiaHRTotBnd+dRr5ZlqFs8sqo3a1JoYsM8TBi1bEGt+c1DX+1JCV76gL
NJ2Dk209hYTR8DvKmSqKlub+P2NGB1NE6ftRILLlXkLgSzV+dlrFjCXgiySzJpuVMLMeDnuffKIh
rD2mQqwh6OIa5VHc83GK0yueG+EPj0TY4ej1T4ZsnmTuOFavUOw/wRsMP3BKRc1UZ+OtsF3END8W
4+JaWyp1iT7yDoV1DLPa6g9QZ3olC/09ENplYU9MQ7ws3Xp9CHBlyZ88OdxKKS5nYVCEdKSZlg5G
W0pI6Z4txTlONxbicqUthQfl/H4dz132m57+/xwVYosAU4IPaNR/7a+ogrt0g5tXGJ8tkPkYqo+z
7YxIvZ03F4MMn5qMyPwnAJhH6I8d2YaOwTk8Li0TFs7lTX/x0HMyhQROXSELiYAu2YZUQ0HHbNw0
6diLkfJzxH9r/Tx0ao99HpwWFFWGsvqvGyYRco9TdeP/ZOd8E34tdjaqedA+VAkMUpp9+PrhY/VZ
7gldzTfc2SuNbi2AQGbDnAiS2lfv/O7EULIS7JWaH9a3iAIBPozM6MrgbQTmAqOrqg7HWGroVGIv
odBCL777RFHOwIhfos8Ak5gHv5/C45CofCw7H44FySxgfVsjNIbj/pmlImk2x9p/usVQp6mXZfPZ
obOTR4NCZdhJsHNg+ZBI4LAgem8ezzfXBq2tKXmx4pt4ZxoDfQ146pVAGySSiswwn4bx6AfqJcB2
ITkeCPivFOJw2acr0TNuA3qPdEwUxeCD3TPbAu7RqsdYdG4jpP5ZVY8mc/wjji7LEMDNNwpUj04d
kEKYHxLw9IGjKtrrdbiquHOjJkxpdR8hIfgYQLep64YBGmJ1/duo4QfN5yGs8acrcDM8Wem/cAQW
ORfCAEX0R+7XRgY+u6tnC8UxcN7VInQJ2jiXa29RHnkpo21N+QK7M98efwZT7X+Qtxcn+YAosZ2V
CqNaqvQeV8cnwb0Dwjyz4sdXKQEgj8MLAmipSPGC6/AjvzRBFJwiSgHvNjBPDLt4i6vLmsYYlDb4
uvqmsscn1PGB0D/TJHHpPqMQv4gETGD2xgEgROkVWODCLEoSA4KBKKZucCAFk0ZjeppipZ/wuWV3
2njKL9cC8V0dvLHj9xzCTxMHdTwlSWfq9gOFeGDh+P/AwpKi9BmBGNJ+BeU6GfKRzdbE8ZvLUD5l
RRRdeFjv00p9wR435Oq2QV+pb/OPh3hnhWtGjXN5bm/hrQV35xDMBvJYFaPUo0YS+0MQCgDSzR9K
1XgiUg/GPzP1oHo+2GQqt1OnlTe7IH+ELOSmvCjTG6h7BBE0faj4UTX/Bja1J0RlYnMNcLglEPUj
RA39DKV2t3Qjv2RcNrEXqmmcQwmg/SNewHFY+/3LMZJnKufxr5OJSSExkpwUn1W6nerItjAVLVem
dsrDQ/idB+IDbZzrQu2WZfSOGrV+XbyU05VjPZ/xYQAg7Q6F5ItyUCXUKNQgDW1VTOBEShmm76w6
4ibLDguj+pKm/zXzzP5v+Q7UA8lGKsjVt/mw3ad8gum+32hGKqXAAWAiMF4yRk3DoiBq+Ck63K23
NH8IujnbsS/Viq5NU8tA79C1yxYKO1ubiYAZVIvvjWpetJe/Qh6ndIsqIOpoe8m/znfVqi2ltjC/
Aivse9cdssvwfIUbY8/m+vCxg5Uvqll/AKOF0nWscAwt8mGxFwS+mbqj0+P+hGXaU37YrfZ+dw9Y
XVqg5Aib4zt90MIACbTwCgn5A4FAYPQYuHYexOPiQQ9jOjg+gcGY2/qjNYXD+2y06rSGNdqjbZBt
8m4k8MHLmsAH0gyRYejer910l/mIH6l9ccTroxINEZ12KSfMrsDFJFu4G/QR3ImFgeYEvSP1lQlc
cQWf9DgGoaiAPFPb48fw4jRYTCi1ERT+OlMVa6KE3AUfiasAWsPzVR71B/bJwF3H8iPOvjxND4rg
ge4mDuU5Uy0G0q63bjqEdVk5LaYVN9hR4vdqIC2lqJg60PIDghQIbu4L9/RNiCf4jPOcEBTMqSb2
MS7ivkEEXPVdc6iPe3u/yNdcQcF+KDP+9hf9uGY9YNPkJJ3B95/isy5mEIb/goWon2UO71ki5xJ7
uwZR1DZAW3GJbywvmqqbhs/X9E5xzFmsNTswOq2u+LexJ42shVqf8XlyE6M0S6Gng0bk+5KI6HUa
wYLthp/ZCtHQkD5jMT+wCxXcqgxx6Vb7DHSNU76qO8zXHhrEXH27L6KLcLM0+g00kzL8TalXXS2S
aDAETNASjnTZbn/jpP3PfU8Jm3Pso3k261gwH0tzpW8SXhandMrFOMT+vV/cylO/ogBPJ/FJWOxP
Mt91rb/ySedSRVUdN31E7lRLeO6ijWaS72dlcWmrvI00HtZMcs2rDE8CiYCJsDhpaJ3i8EE6M1OS
QS4wxOcz5w8P1RBhGD+x+HTd0OIT/CcFI+TCQQQZAmLJ2HeMj0LvnWGuwiXxhUnEKmagHET+OjrX
D7EApaB9Wqh+XCiYBzfmGWUT4T0CS5O607nnPbINDNoQNwDKXth/a/dH7MqDpwV9WRgtigM48V7M
hr0EsFFVZPycr2jNUbmlu6uRVmUkCRdwazxLNM9I0IsOXoHdj54CTA+VLPoT7GVnvNG9a20P62Yk
yCS/u7oJxNE5Rs9gQTMNsLWIvQJyfI+GGnAb5lJ46e4RgNGNKNea6JoGpM11QNM0NHQDtXdSiTzA
qv2usaSF/nr+JYE4c4hhuIOUK1k2mWqOQmJcoZ3AjjdoelKk/HXXwX9EDqiPwhuXVVw/PyUQaxQY
7OQHfVEdVny8UdOcOX1RzfFfjR8HeMmerOSEOPjm9PsD5S94TJsdxuvAIHLAuboUp89n5bojQMK2
nYoh+LQzwIoFFJ1P0fTQtbsAwy9YoccUiQH+wkeYw530NSIVuCj/0T3B9k3+o4T84dkKMcyz6tTP
zLhG744IjARqKJCehK8Wlhoe9312p7Bg/ld/vtjKIiQXyTsx0HdsDO7JrDiFRZWpIAmfu4MyOa/N
m2p617OoHAO/96I6y2KyOpMPi2wpd92hyT7wskcLpcXc/3MAH6Xf+LYUuMFQVhQ6y9hN+y7HEuMp
B95oUPvWowdOeK8T24mXkhOyHN3GIl70jgNVNPjdIsz55ZwbRUnE1D8ioQ4v6noBnhih5d8kFL7k
QGxK14kf35BCUsCsGN3uAPN3sZLhb9ijxkjnWC0jU56ozNzcJOFIEGbShH6415CqPHWvtssqCFiv
PJ2i3Hz4DqBzczZiixxdofSHcbVFnnN6gBJ+9qbudWfR1p8JTPS4jwURHp1/C2ZXbdhLPGQzEmCu
5OSmSo5Frz5Ulam1MA3ePrZp3y5+y3rEaVmHNsXEPVqTKtxXI+6rWMmUANCtMzMXyRJqF/+qUvQU
dZVQWfn2nkZyKBw3UPmVHs7oVbwmqeKJLmWVXX5J0ztwdSNv1aCp5ANjZWRBlhqhH1gVJ2+88/zx
bPKkMWoFueVlv+nCGJx6+qmuTkdH1yxfG1wNZzRd1aszTloXdThGTkE/txaPsdQzsPXqskqqgJAq
qVB8Z27ivXGk8idziZrKHWe1271By3sbWUVfuMGviXYhgCuz2BOoh1ymdM6vh61LT9HZwBmP2Yzd
g9GpLWte9MzBdRr9kX8uM5RyMaxa2uX6AR5/4Ze1Qw9xmJwxBTbCJMN+C+Bv1iWtOYII/lEsjJNx
mrB85jJEGtUCut8lQlvVKNNwHpNdDKXOvOLeShdAM3Bd8xVh8RNzQhU5q1RKPCtQHLH1OtVS/Qbb
BaO8OsNod7kYN0LSxUiOMjzoLM2RkuinfNNrO2LJfc21XUvYOWg9UqFs01R1WdR1/N705nK5x/Wm
I9FTfb9NrMbUH21znycY03dwoqbRJIGPLZwyg1j2qOcGf71P32bNu305yv3shwrDyinBKI8ddce4
/lI4HFf45KR9vSQ/CQjtW0au799LdYh087j7z7Z3SuXi5UJhNJntYFzj54z5ecJfxv+1/2vebn/z
79ht8COZ8QcLAFRrwxLt+h2Q+Rziw4js/8YzDgVM2BEpdgNl7rNQF+tLHPizF4f5Aba8B0xqMpjq
ewr/dQorXisP9+waQSV5mU1jgtq4G5Qa0rW1F0v7OXtH2jF/W8Q0LX8ukxi99TZGcLtD1JkIHAqv
Sv4K0puuLKmJQiDuRmfW4x2vCcHVNF/ffwiJ1RDh+mYkbI//xoTgdFc+nO3y83CD670uA59G91ld
vNtGWv+Ee4N1U3Qn9HHV7jFsWjV3buLssPN7AL9g9iSnWkQ2m/AI8bzwv+rVwF90/3KhjoMwtzoj
O+gkzRcE+Pd5piJF+U3rKXrGt6L4nxcoP9ZW0uulbbjCC7jq0zNWsU8wxIJl62OWt6YLdrmLX/Se
oIb29EF4wO0cphPc8BcSRsQPYlCqpsH9e84MQu+frOL+Cv7miKa35pxOF3t3lfnwrNhEwkONplxW
A8zt6wgHQxzqWdS0AYHCX1dwE8hlpWBbkQJs3Jm1A0KYBWeSCpbYOooiBloup00aeakl9zkMUCK/
MV5PCBAL5Q2YewxWva0e/PvblmayPwmQo7uYa3FO+WUCmAg441q+Z3opQEI96G4BuWz2gfPaR5n5
oc3LpQtPBJZ1/NKwAZ0IZPi9p6bqYwvebpXsdmnXr5pUaEvUl7lsZFvlK8LpjBVpl9qOq9AkA9Yb
YSeYKt0FAw/Q5Yw0sTPEDCUedNYbbvxPYcP3VRbior/GLU38gwH0rYvh+uKWQ7hZEfPfT8QG7ZW0
MzqMsX3Ito1Ik4BhJyt/+emxy1bAV00hT9lF8CeZI2aY7ve76PqmvigdcrZMUANw5zaqdjIeEG+r
YBNRj/Frfej44mUmpd5CmbVj4YXTrTiwzLs0HLGhPs54fe5IYaGlO5FjHBly/PsIJNOI2JhV3Z8b
vwsqHjpGOlOigo1EYwFfIVVaqC1ImHGYuauY4WLM5VJDI+Ce3rybOezHSKlciz6OBw8z2T5ZFAuJ
3714ShGur+ZszPLIwwxlg5MHTZn+jFNHLrDnUrdjStDZvVX0LXnw8CjcuUIfY6rPxAmKEXZTRBe9
B2xgodW9wSsKjtPtZm8IBz8Cj4/R+tAXI4/f46a1pyKFkll7pv3zw9lb04OlMoCC2UvGJs9TysWD
LHr/Av2m1uTDtHKqAH5qH0RbrnrWLjryoucha2A2yo0N/GgeVsEvjQz29aMn76QL1AhiVy0qfdk5
8iKSRAoNsTw/nIAa+DJkZrJKbvdyMXolVt68Ziiw17RF/IK8G+gROa+JtPbx+dnR7U3yNYdpTd8f
hYWB3FFmGqI/VbES4eSziVcXAFOGTKhugbILcGkfzXkDEOtwokMtLxSLnOlHD/4aTqD9r+hI32XN
7BN4uTuS6609MTwAos/hNjaepWg9KBkpV+yc1INTidngS/zmQm1h4HynAl/TlglvVs9bh6t+HdPM
+nNt5SFtK/IVrBCiMPlaJRXWyZIT/oT8sUab+bVg0Z0tKnffty2mTpYsmyhe5mmby0tD7KfboMIG
veeR6eew1RH6KffsAFcKn27CD0K9P24gDbML6ow0QOLsXLhr0zFc5ZRNbcLyU2w2rOkp5p2+zAuX
0l1UPRA7iXIizM5hmdcnxLfEKvIjd9a/elhd5nGXgoW9Cnq9/qHaXkjjQLzXjqhgu92NGJxidwfK
ii+o5Mz8zgFeyicNIydXoyHUVgjz9HTjwL3IacYnxcRymk882R0iW8DgAVpUJZuhzZxQ/pYWqYBF
I2HKhbm4M+p9G6dbT+PWWDPj4eYOq8OtlfMrgFugPniaoG7IweZEbVI1HbCRSOb/i4ImHjUi7gyY
5bqMPLRpwwG9SSyUbnh9wUFwzw4UTFoIjQYjQWX6IEPwe3P+nFk0Fa5jyMr9o4Mi5Zp9r+WiPjRN
mUvmQAbI/m6mN5FFtFLr0gHxtNCLuDBV8aoVAGSzGFiH871z4SJs0LQbkrjr++8wyMwBSAZwSbb4
n0zqbWZ8R6od2p2BYDHCO/JT3ae0OW9LSHt+F4eVA6tOC3tvxFlTLe/dB8oUZJ7p2fwBnORGUk4l
QCkNaAiwgHo1EP1EbT6giIGtg/3i53PMetnluOv6Bl1v/089ZwTJ7sE5BaSm1uSbef4M9qO8lJol
iDUW+hmp1O4M4T+ZuZv2pS/hHbQ7rolkMW3cTmIBnNiBpZdVzVzWI6O/+4+t03KlJOlaL0//dx5e
7nD74ap+U8YFRkFH0Q7SI3A9wRFIkjYiUrxykqSK2VqHNA6Dn4iHVKvFuqK0mpG6oDbUEkDCwCIM
sTuSIDyX6cSwYvIbzzL5PCz7f+UedbScxQ5/FNn52KCQDb8sxVxqQjr27x1ltVABrn2vzYpuwt3G
qOQO3lm06m/dkFunSR2/WTeeoXmeMBZuMQqsIT0+SrFjB9v42B8sitK6jmLRBqiuUh22o/K72obg
DzctWOPnwF/6ys4z0FjQ9+so/RvxsWBud5eBfAjyfdxkRFAa9nd1uSvKUjtiKMomfPHiBH5Y9pz1
UXD+KzxK2ZvVNWCVjTcgU0qaDQLYslYINa7Mhy9U6bOzuDkd2aS8/yEoVzfepKtY1U96s29XhxC0
j7kwh7TFlZFlcbeeFZY0gVkQdpTHMpvdP/R5Q3EGu7cuFJlth+j9VrazUU3OfS4HIZ7vmy1cpd51
BiJuS0pO6dYmdmFiL6IaVlM5I2eQ1JNWu0OAr7Gzku0WgOMpRSLK0K9A84ed3h7MRt737NVhBe3X
3LVHCoYUDToTNuPh0nSTrX9cHdBeYepEWiA6l+DdraPz8z99dwBgwQIRN5zh/9hH8ZtzHc00x2Al
MUG1G1D7hFb4mAxVSyryJzTF9vl7VQzJCZeOQES13nSchXgoppfw2/rTABMO/imu5ds2ZD1XTFjg
zGNX/amB3b9Q5dBB8w/XTVSBJT3IYkVUiIFFjMqmVfH8ybCZ0EKmF+vJmE+IQlWELkAYDz7MU1Th
dQbiQJPVz6Lf2tWleNhfjgq/cjPGJEfN0neL+AYGOxNJ6Z1YlNbvjXF4pGcjVr4LPCYyxnGTfr83
m3DOYk5dWux5XgNws213V/yca9uaKbMXepJ07e2S8J4CdCN9NHpm4/Ys56Bl15pHIN+APlsI6cqF
W2R/73qSCAThaF8ndx/kOM/n/UngDFvghoh3u2dENtoTC2eKPi94mRMKDKs/9/HeqI/9tjJ7mn8Z
jiM9+WIADhQCuCmwwmltNuk2DBTWqbIHZpzTHplgLsp8SuvYnW42JO4mmATcVFAmuz6lPrdaTrT/
uNxIUsp5NlEtMWWaOIIDgrBi3aU1BHwTzgvRJRkwtaQjSL9XeaqzY8tptLk1pw1h7wLCH48U7JmA
GeC5xuFwKuILUOkONhmboty4YgZu0e9wXk4lbWKh2RqkN1h1TxhsfrAAjMqmHQtXu+X2NeYUEyEV
hOKzQoB6Fq8JRcAxLaqOwE9Ft2WptSGCb+XEMSgZSrh7V33Rh5PI7BouR/zvYhJBAxTvOB8+jvr7
OnIZrXZe6tfU0QzJSKrOBd5sDXUWdfmdoRzmtk9jHgzO+1VIrU+RE7G7jjDJIPznZYI5i+1RVJi2
7p2EihRoZjlsRp+SWiB98H1j+FSifIPocL7cruMAkBdAZxRKiInFga/Uh6E2dZiHsqKTmlMi3xR7
wlZYfMUaTFshUf6PPIonyZBFSBauW0daUCqmx/6zI7VUz6pNZvrqlJMiijmsMH8zaigb4wdSTPIL
3MmIk9Ce/jtMBAbCzG0jaqRJzR9ZVqq3T0qVRuXe57zD0LChIgS3bOv4XD9Q500w/k8DRLhM3GWV
FS5yvMiFY+z794Q+F70bOKOU/mDNuuWUrOAED6WnO0qCoCVuu/CQwzjUF2OYEvIj4A0Gow0lqYQ2
6KFIC1Ty4rel/ryM4jXj1ZUUye/YIZWO9QctXX24smyZ/kK1nu8cgxL7+qZsEuoBNTeygAsJJrtV
ZSnedD3g2zp1ApPw37oCX3MKTM5nsm0/HqDtfW5IP6AH0ggpfccyvROW86m7lQ9FRwEnedhmkbz4
nDx0NsyO0veiD2F4p87viIr2K/84oAtgyqpTcYTJ1iadjVsPC95hw7q0rPgjEHt27VUVbKwIPjps
WqTYaUfBcSvq7U8Nd6TFqKbXny+h+6XH8bjhUsdmidrcSlzDWVy+BXsoXI+U/acAX9C57N6a0HOZ
wAsouNcOI1B7kROL4tlvyeZXityXxbv49xE9ZJPwsUUuQ0FA8qpA7H48SZaM8de/GVqTdmKdIELg
dazE8gZBhpA6LUmeEbdIPh45DbipQrK2gHVZrm2vIoWPtAaODa2spTa//SemFuPI8oScYQHdZWn9
zXN+rpphthJeSAZbNMOpAwbSCvEvsHHu6wpaDsCrYGzXODDCRcCqarzq2w5PTYakoJDTOdeZaT5v
ig8VWcSgdjYOCM4IZf5yDsXyJkY5j5VLzQRsFLMcmIN4NQfFGDf2v/wWDgezlYf4K9CF+ctOXXmq
ssZMNrIzpi5ICD+vGIvdbar2AIDWCz6OcyO11eV/sz9c1CPCji2WidJoGz4RQB173R6GPkgofvCl
VYOXWjuTpcKwOjBl1uwH9KV7T+u8DBhXw+yEcS5JrzSopATt837zWIDK5N2o5zPaMkyLDgp0Tsq1
IfpN5smYZHmQ0RfAw4K1Vpb1oy5o+4iWeITMWdB6lU8FvWnxKOmJXP/DSbAHxiY8IQHjZP2CIueM
DL6iOdOX8TdJXFZKCORJrI4A5gkpBdO8BT8H3TjMmtfazucSRD9j1sdXSa3Hb9run0SY+AyxPfO/
ykz/TOcEDLtt1644sW6U4vZ01TxJwcd1EOQHEzjRyO8IqzYLxe3J+wutr2v1EJkohFhDBw7Vf1Mx
1RTl7pejP+e2HDcL4YIx0l4jPM7ujoO9T/+hUnEjDsDfov4MTST2XctSffKJKmZ/qZww4zVESchR
tzLFgcM50bfucYMXMKLdsW44P2TsE2HWHymlQt61+5WNZpaW105sd00xnCWqsjcHiP3I1mfTftJA
fRIdU8Q8i0iPOM5sks6f61tEkUiO5M+ZWyrUgbpH27aDTccH91mfI/YKy+OjSXC2rENnAihrsz1s
o/31J244GY0X7Uie9BTRaPcP/DtfC1cNYh+XSnJ0eZxB6Yfe+MN7uU4R44W7Q0ofZmFPtFhfDU+/
b8qMUGYbUSAVx6GlSN5dwl2beOjamVOmi9UI4yl2ednXr3qM3wYvLcRZpLSICKBc69JziXEayCDv
VZpB74Ls82WjD/ZQleV0nY1wzMdx2H+prlcaEMcjUnPtmwUyYURXifrJJXGTBCZAlKYinQT4BPLw
QxmXHxq6iHP6O/TrPXB3bBRU+PCUj8j+NaF/xhf2kWYlEUv99ve2PdWQCYsV1N1cn1xRZc7DLgyO
ulWUouV7IxYaZla2ECjW9h4m8PgsytWDBlEd2pY/hOXF4UcQLOdJxRrG9IVy9D13XeQZD/1BFuzr
z/UpjMYJEOt6KNBRFRFv0cC3VkyIvqID/fi3yY6nCrTZyQIzs6pOOtOHbdd5sVWh6rgzlKVsLVX7
kgwmXgXevcthxdrxJuMjCkpsVS/cXNfGuBd8kl2aBP0A8KDardZCnF3XRy9CADyUQz38afKQienx
twERCJyDtuDGBLnr880i6PJdaRNkRrp1JFEhWDpr7Yd1n+Hl3+UX+5by7SdNiKrkSwWfDggJWarM
qaskSRwWzoqiojo4YUTrM3qpx+CgzBGmNxVxgZn/rmhUbVTgaYaDiMvg9Kak1R05yhRtNBK9vNdU
zZoj5vpL1ZweXD+jFW4y5f6SigV3ZhjlNSVxwl4WqNsi8XCNnIvZ3JC1K689xq2+SDjN1VBeZQj+
RD95ZefOTqmz3lD4rIfVnB/HOIaRvcI6JjSEymcj+uvFVCaYJ1ip8XRGKNciklFuksGCE5iXY3QA
r4LpP4lVtgnkD4TuuZBoIOEpsc+U0aDZ84bAEUh4QG729MF5w09USO9Y6SmlWaQK5A2n9Pg+BoVG
UX0F2Eik9f8n30bVj5VOXvdn8ggHq0AVCk1z7RUN0KTog55LGSifFWFzAyl5z9jZPGqvOULFdYjh
J1+NxBfrl3uEK7Cbuqu37iHKMjbicoDI44iho9NFAEqFMHY2vi8mB6j4M8XWVMLSEsO9FJof9pf+
ZY3pM0dLz4lD/5dgrsz3UaiTdK5GrczWXoS9n6MZ+pRNFTEUMTw1DtDa4X4wK1zJPzG1uUcTgMVa
HcaeVhfkxP4d8PDaIn//x81KrawdKIsV4MBZrcOqjZl6+diCQ19f+PerCVjE9e4WgOXMba35IgAO
qwQS+fQXil+N5VNdjrE/qvdsxt/riPO0vaGjMoYwZkL6Vt3dSGMOGDWqoygrfM57t+7lnucirqhu
BHltBLFJ5mRiuwL4JjMt1x1LSnX2xaW04y/+IpnogU0jM4RxOu1tVzIudKSNz6mnw1xxVAE/kP/M
jIR/Y4nJxC7lWljl6zhUhWagTvzmpp80ioCfwMfdBKUwhA6v29N6/QELUAstzFU/hz/1qiDqZZvf
OcsON8ZqHFmfsYVP5Yoph9BmDap0baMoBg9Xo2g57kfG/p/BRw/3qPKvUYlAKezu0T9wIPLUU9Te
wgxh0GQ8dFTceR7bA6wK4BLsN1/gkeYr+jjcfaUdIezPGM8QhKy+X5/WE1b+NQSVEdbcHN10Yd0x
A/mzGJRid/8y1nvsSvfc7/X/oVGFflkw0JLzby3R06Q11wPkXrZY9nzJdfy+sZBtLOhkHzvSKTYJ
WxbyGzvPhAVDQVMHUZ9Ndl4l5Izdhs/XG44xNxIQ6jAzSG0uVGhTOok4T3pTGDvHD+w9UtjObrQ0
TEvA9HMig5sBQGXTIRYrSfWIcTZ5dRC5OQvSTt/1iVVeKp9dqY1pZiCO5PUvz/kOEWzY42aiGUu6
feSuNs+km7tCBZqbrnyV/Qeq+XSInhSJBiiRBo4c8VaBDYIfQJBltjD7we2ZvLwqJXt9wbevPbOV
fUNzP+hpOHeDDnaFV/QtDge1yf6lA5N1ssRdp48Z/2kICOtvIPfBbb5vR6N9f83v9i2Q776N1HCZ
bB9gwz+a8lkNJn2kN7tG97+E7QDoXmct++vFmHu19QbZODE+Ic1nCbO46JGEG+OegGwX8ZUd6y41
wfll9Lq4J0mrFOrxlrD6Pg8aRRyqc3Xuy8i8A4Bey/Vd8T5J0I4EtdJ4cT3XzW2miq84wpqTum6j
kwY+xhibdYLLwrjG2M29kmzHWzSQ3WwDHpuYOMMSty9Gl5bBlKiE+GHlCxLA3odVmfti8Nl/43jf
7khpwMNoK26GZh0V7CcjovFgg92qFCmSqRmz38RUQCnPVzgUtaQbrVraqyOlLf0lrCL/gCHn/CiL
j0tbPxKdybcrIUu64qFoGiC2rZEt+5Z0EM0rnQz2g6Y9DRKexwgzF62tA/3RsyjTWOJr7v6S8FwC
by2TFixkj17teroM4CwLdrv/iujGXlJy7v1mZ+iy/WtI1s4s3vH/DbUcoTZA1Q8JEuRBFFYhF7YY
LSR3fkDSaJSnOhTfbCtP5q7GiyeoNTqEynC3NeGwLXePZ9rztIePxiMK6rtu3HmBWGVpHxbRLLEo
fGtbjS4b1vojtO6lzvQgn8HRkqc7TxjoEmRAczfe1OT8mpRv75IPFqjeL3hQBGQ6z1jWhbUt57nv
zyqHFaaR2lkUhLPmGMdH8W8elNpk7MVkAWcxyXR7tRPzWmztjfS7du/lBJPnVpLG3hbrSLCjAYDa
mtKfoiXWd5gN2XYfMpNRB/20ubtNj6FdlpQh/iVfbtVTt95hkfhFWoYBnJzugnDNZ+vO39mi0BaX
MO9TqLZidNdobajcp7liAbYekf/Ev6O3Y8jlPBe8xtnJVWdsY+WaPd3apH/EVL+BvZMVAW5ujWkd
idwo5oc6a4nqIXUduOz5hUGb1t9KrCJoN4Rva80Ag6tp4AxNZ8Qs9HJAVOpiGYaj446QjUQEeZ4c
uIHesWL0Khy2hQtqDokgWJYcLNZ3gwmDM0OVDgIa1l0ZfBAXU17Cn4X17n2bOxQnGNnUYEcqZKqP
2k+pwAq/78FZlcCJOr0c4NfP2OuQeSyFvoMR99mTv8S3S1rVyMDSzS6ZemDnZzMiEcP4ZELIiRN/
DSHmub3MLeDcjrHrjSmYfH86XE74tMBrn/6OkxZAy/0NYmT+8Tq/ma2ofEpS0n6xuqlEWYedw++A
dy/JWn6v+iSvtPslXYrqpi9o4pOQWIF+PRUL6mp6AP/2O8owo9JQnmhOGfgnKX1a7XIn5jETUp0v
pgSJ3HhNU/SrBCsKCPXI94ZynGN1n45/MPq+kskTa+fEdWJCAo/RFKsZyOiDvRMTanqeS14L2gZk
aZuatFUjzaCZLtBnPj6wL1Zq54tu2/4aQnKYIxdMsDzv80auK4kK+EvE5aQy3hPfR2NGxTS1kdou
YoziysZXVHwpvppKLUX7tCLDT4mgdx8IhS2rB1l+pQFOAT3NQ9PlS9cG1w7twLp++NEPW5hwo9mv
mbql2AcUiymfEdIk1gKpepgRWhY6KM3zEezcKAHLsx/EOMAtP+lkO9SjlWbUt8GU2NdHWXjkNmM7
8jyOyGmrFy3oW0bYJvoBAPo3Km0evAK2Rw0WKvtbEqyR+KXRaMioDEP64XhqS2BvLElcoedAWyyL
WiQZMJ2sqwhVju/fL+8wEao3xupt/xgby+pF2FVWh12mWQ2UwSJTLVuY1N7rEyr7mEVddGqw8o9z
DjUKhxfh4ZjNwpwyiV5H6IgIYbLlDPKF3Gt6khdyME0nQKvkCAu4Q2D4ZJ/MuI4+CbPEWbepLF7W
MFwbjoJICNZWlE7Dfskgd9Gcdl66M9XMhyjCeEg6/ZXvytdyRfR38MoIWm85P0/lDYMcfgUILSbo
YvE9SfRxvqQOh8LlzMa/+TSPyEsgUHkzGxHdUtW3hr2W9/Xrb969SZn7rYa5li2vq4TwOdq0Vc1b
Oct6vGELNb20XICw5UxFl+f0YnFokCaFe+WojxP3h7YKB8LTlwTCqQhSwA2GqpS4mxzbiPDcp71V
onAtoLCbeSnXguwgwP/BXDWRo+bLnpKSd83tLYIf1hTk2itUcjHHDVIumPJ0r2hyKp3eyWUaFzLy
KJMhhFwFz961iXJ7S8VThhxmrCby8SuFkuh0GBUV9PvE8NPdtK1dkF/gV2ngoHioopjJ3KfhlBhz
tLzfSmaiLdi10jvoAj3tR5Rf1WFik7gtfhkpnLQBVlsIY6WsNW08rp7TBLO/TrTXNHN5oBRASKeq
IcwGVd+B622r10JGGe5V+03qOE9NSLlwmJbeVNFnFZvGHk6O3MJXok1yyzrSppwmhoS6t7D0VHeB
DHJQiOsmy8vc4QfHioTCsE7p8p7XiHeFrH/bQecvihGHRsNjJq1LXe8T2E9U5GvKe220X+GRaJ36
mlqipYDYdMYNpEfqDNQ3lLr/2k1UswCASEDSIo+9pKykl1GeYiX6vXxHhh3fzbplY/Dk8Io2d4tQ
T0Efwr93JO3GWTRVW3GSL5LGkSFQX6avralcwicFMVGdFJlQ9mKVJmMYce4kakfUK2miUxT7YQQ5
9sEUF1YbiVlVB865hhcEjA2dZ/Ix/Rprw/nOALtEVRPUhw889ixWyYWMGPvNPi70tZshweUC9rSO
Tn4rLxFNSWldBERUt9thrg2V9Jc6aJOVw1YrZS0R0f5ObndWrgkDUB4UyTwEBjzvzPgSYAIoKR/v
nSFpciTeZrSGLBlZObDOjQlwtAic83ptCmiH/7Sgy2A7TgAPnsCXEGxrcHxs2xuPeamD9Vfm0wrC
Zx18s95kTnRcblCfXfd8b+AlRVvZlO9khk6vjtVKeb94VWASk4Oss2CFT3kxXAsJHgnupC2TfFX+
AoOmcHlXxsquiu+7RxERDMo7A0RUDy906qwZoePf3dE5myVRxAtFDCNU0kTncnlA79h4fVbyQRFc
UL5WpEenoa3aRCyfpPl6yJXJAyxnhU3oKPlWHq+gjzPbhPRI1O5RgestLuv2Mugy8D085mbwjO4R
5tC/mly4ZCdmUts8jhVpvCd2BdFkh0B9qZUthiZBtrQ/eEnQzp0+gdauit9gS3fEMxC8o2s/oV1m
tiD3YFodnaUPwzJWZtlaMTVlzos9KYryS1nbN6pbcnC8yh1jgle/nBKBUddw12h0SNm+T/sMjHAE
Fa5BOaSDH4B745h7RWFEL8iKlrDT1lbqcU47taOqcbECgogL9h5Dp1JvZdrLqSQNnvy1SWt4a45H
9bFnG64PFtdXFKRYnyfi9po46F6LMPhNYB0N0tAddXzrGQF561NTO+ou3fUv8hTs+abL0RECjKM5
oO8yIl9nG9uczNew00exc8l/016jEqcZ/33GywATxmXx8OULZpt/P4Ica8lBjPrXAU8ZikFF6B40
aAwCP9U3DzqGKheZWuVDNLFQPQZnV0c9TZb1beeECdvL+9xBfuHy6MeRk59+aGk7RFvJdE6EugmP
HcchAbx9EgZrRfovv0/0N4xwO+86vCcC5Httnm1rUg7MP1/o9rQhTPmUb3W8cUNNzOmvTAU3yN1b
S0WVCMo1khBLzQ2Mw9sYOhHj/lpKaA5q9OEI4QY5z/qtTWcgaMBLpj/EamN+hipY/5RgcerS0ZIp
+tiMw1hjPwUftSAMmbn22hZNGYUZCMFdyyytR9nUI23NyKEbAJvKVtXMAGY5TjzktLMGY75cVJiX
EtC1+F+P7VUchS7pWKzF7BvXpTXcJJBoFEkJQmaTQDn/2wPlB8UhB0E54rsf0vOAoCnHjh5B74Ft
LNUEVCMDSOMKqQgvb5n2MYWQzYDR2dv/TkksIdLP8wTpi/AnFErj2FpV6WocUqm8UQndxCEqwSCR
slB7JW2jJV0vGCU4jMtffA4cPJUvfq/7HzVkQ3nP/cEXfmkhK889UIsIGDPHs2pUD1OZ0rL1qIH3
LYJaDs7W75x1OhMa3pyIG5kRpoR5267Wa01JucOkiC6udqGdlL6imKUG22MJYCzG3iEZY1CNnnNX
P3zJkPzE2BYtv7D0iT4OHOZ+DVQ3/DRUQ/eUFW9yg2noyEE0KuISnqrdrgu3GeDm6FXE2xEfNYps
8bWUhXYmPtqmaPRXCKt+X1BdYgWMp1hQ62u6TjVy2OsQeE5SiL702EnLgoztRuz3vZ/NFcm8qEkW
XUw+dZAfXxM5B0v0IwvqcuG+vmNd08hNd4EREBuk0lT+oMn0d3rzydVplA1x58KTiLEDWJs84IdR
Tl+vtgvqdafRSf58SzAn6cQ0RyfhGyB5xCfYDgJ+XH2GXgwjw+/rMe8awi4/Ne4fkkPTaHlYQlQD
Zv7TSoaPWR7WjOPYshUJeE1saowzcKZc0knv2LK1/h+x63dn8D8P7pr/oxCu6jWVHgz4UwWKKFFL
biQ2cwYF9YHirqmxxmiWFxFhUaK2Bg7fJmz8LfZpRVK0Tdh541wrWac1hpHiZT6bJlcCaHTjJQsz
kMkvDW+TKqj2tW/U+PierE0HVJjw+ogHK/84Y9wCvRCxSTl3dD0lnoDRvLN6L6G98OGhMlOOpZ3j
a00rq8klKtlEh8wBAINA+TmHoLUhQwW5apP21cj2a8svtYKOPP058h8kkrmlxztBMiy1sO+4Sqd7
7B5S5RovlaDd+/ybCzSv6Lc54xhd2CN++ylGrc/CyJgPqjOx0aLBWMkQICDq0Z2hiMrFhOk4RKyd
T63MWcQAs7PUBqaBX+ORzgAwNBQgA7ONdLtWHdY3xltRrxPew9g+iYZVlI4P8kTbvIkBKH7n53wA
gRUmKxlxz7f/IDmUEf65oBAnFgc0CmfeeqfxKr+Pcxdkzwo89Wgy/9CKAmccIYV0bUprMrBiDQbt
WeOF60/75rVXBIQvP6nOn+SjE7jxfZ5XQGjoRj7jy8nNsJfmzvgq4VV5uQ3QU2ITX6zci13gMgQa
50z1SB6pV2CLy2AD6rXDnyy65UWFSRU+9decFt+3lklAWTUew0sdClLH57DytwUCeL9smHt3x35s
FuQ/9n2XvhrV6THEF8Th3a6+D7Np5i6ZqDqHPmuSre/q3jdsYnLKx/Lq3mLxqN1kPOhuIeqjamzz
j141Itl52wLVgwe+ouzhMvw2jCTQUqhL+xnpJPetE0IXquEBjcdR1gYbiwn+hOOKrlDf675O33K9
HybFIHThCc5I2tlKJ9q+DEloghsPiSwS3Z2Zcy6R1uuvQO+DOFPHUyxUJOzuchHsAtcYouFRvwed
6lFDyXlr9+Ya/lnSG9uj5Qd8RXEa7gkRDZP1wqql77nP+HD6GGdWT8PVACz/XVWfWiYZG2WZ1uFm
OO7tV2kxac/5ehtntvqLebMSlsM2d/n9UmijimMfEgbFe2JOYB+/ILu5iESJXFakAmtk2kyHkxgk
NAK36VA+jdp/xN2/v4JDEjBkSJaDags3jMeam4nnb4p4KlXGxy1TDMgISFBJm7QHxbfMaLnSDlnD
sgT6APABsr4M5vkrnsJW8G1huiD7s257LjWkRqnWr4tdfBmZWk5PJkdPVys7Xo3Yv6gM4LysL+ip
CZ0biI9kZ0KBsj2jM7LduXEvE7BcAnTDmBA2A1DZYMaOrwg4R22u1NsJbcg6A3ch0TD45aiVfZW9
ecN10D6ONIC8I5WXVv1x2NpbX9XV8/SK25eH/B4PJ1FnpQs6JPWr5W4tNwbdsUemiCHFDaJ24hDq
CJn3HvVO/a+NEG9OE+cBS758EUpThIG8BPJRSdKEoI27Ot/3sVonLdfgPw7wJnWf6YDLEbVrvoVU
NB+VaojGYHcCssOqAmiTwyWCWmUJ0uHYfH9LFTT9Yx09Fixqyf3jZN5y4BchjMZUC/7mMAOUMvXs
DztUX37DMf+kJIPSQagXcj3quxquJwlUZi2XslTmyh8hhdPIBIDhLoMhpWPh9WsbiUsgVcDTuNW9
w1c8NqAspZRQx86rOoafe9Bk1EAtx557P3JtY7n39zx6vxM+8U5LfMmNkzuF8ocdXw5jCKHCzxkW
vCTiCJNMkQFrTVh+EO1jxmR/hawoKdnrQCOhGGiqkwsXYGba7bVYLqwLPRjmjeNSpZmYybITVVqj
PWJpB9jlVk6CkFe+OgfDbTauWTtyr5rlXXwMtASUCz43dkRKTC5jVm5b5hfQnvXNIXu8fNQvZjJt
azc/zoSphEO0IovHwk+ICwbDRHQLMGdPu5a/DTudBeklE22ETMUGhTOKK5YdWMtsOWr1vS/zmXZd
WUXputq+23v3Pc6jQPES2j5IEtzbUQvH9afdW1De989rrB920P78m8omRRqjbpjfISFpdVptcrcX
aLet7h55QJTDB0OIcXAOg1IhVjQTTIZwwbD5so4EgyNqKuDO5WqfybnfOi8vobmIT6SsKIUrqVQC
oWPm4zGoXy8b6lSW4rFZ91PLwiZEL6ysF9goHO3AuSGt1OTfA1g5nCUhDy3L+m9nLyGs+F8sZ3JX
LZK7LsTSYZQbLadB57U/AxeGtbhVHxvt7LIer35kSk8MU6RAFRzG2OO6ytvfsG5CEEIJiDAjqLEq
2IVMWCs24UEzdlKEaXUM261qjv8qGrOTuYqDTzXrjENONStAWwiLPpZ35qR/KENnP2Zg97YXDhao
cUK+UJGcnNAss7vyOwiCB+w8uZfG2i27I2Nb+exDRkIYYXSGvHk0nG6d6NpbAkXr2j0zlzKlKWIZ
ExiXJHduoUJDSuMFCKMWV6nEhTDYxIYwrna8VDsF4PD6NZ2ZWp+8kVEzcZM0aUsqLm8jx3BqolHH
Q8t+hjb50RjJMk7BgYWaPKmL+PbAqNIjA1HWANW6gDLEjOSw3a5+76BaTWahsFXApi8KZ++jUsbl
2u+KsC1tJDJ4CMWxv3s6hjbeN/WvIgdO/rIWbl/mdevOJtSvI9jnHlWikR4QhJreaHx62s4l+3PI
B2E9+BrPEsnpbcKBV7qKpI1gbBUqQTVNn+F/33roWCR214TR0P+s8LABj/DDD2ZH06fYrcgBSJMY
ypyC+BvcsRKziwi6nNBpUkMxoUnvgiZvURpxFJKgrcgtfoZRtHlVOLCdCa0bMDRaTGa8Yi6DdB/B
48OgFXcoi13i0j/nEmEbxULxQxW1y46aKsEqEc1WBpsAMDxHBoP+LihYQCo4j+MQY6qX3dUrn+Aq
0Vkv85cteMiX5aTj/ihx6HDoAGw9JPcjrmbUonBrBvclWm0A4y8NHcT+UwZUoMh8TDNkodADEf9q
sPs5vT6D2GgDNguxwPDx5MqHae5ALBQgz1fYL/o1lVKwk0kwEIthszEbIpXbhKYYNXyM4C1JZ1Et
DSiCQtjX+Hck74nbHfVsGkZMTZcyZpFbJZREZ3UcbxzJqEsKt1wUcGWx8lwvxdqqiDHk81pXlaob
z27FTaMujBIaK+/zrAvcLBZoYQ13awY/UGD2gPBadfN/hymmY/+VVgAtwI2UY8tI8AKa/068ZjT+
EHKT8StC3yQql89sVvEXZW7wYIKTmr+jD8hh2Fn0VEDztSTP9wqcd5fZuPmPcPakS49s/6TSJjPW
1ZZiiQivjlahlrzoDSsHK6G0giavgyUhE9dc8T3Bk8cQwVlOSdltNh3o9xmyTFbV6xI2ECMfVKJI
qmYVg0KETc/TFnOZbl4uAe/bGnXThShcWEVxiilqgRyDLYSFB6XQkV3gxcYkBKcqno83+Ytp/Fnl
34/ZGEQTuQWIF5eefdXzjQpXOtN8kOaBZJ2E8LOjExfCOtzRVyuWTgh3b+eYwDzFxWAHTaLZI9FT
R3HOjxY6EMGJQaIPHeVBLI7tJsFTDOvvbToD2zxNlNn5/90qnBhW82xeDgmiDhjxVwjCAVdA2VjF
FBLCrpTi7M9/wq63/Rl/yYDBUzwmkX+OSIvLDC6cMmpSU3KyqXuplEvDiABnV8/4JxvSnBMpiGMq
4EFrGejRyxiXoO8+NqiSr6eXbMInncS/mHyi7didZ4pg+gF9gfqVxfeQhf9oW9a6UN6Anm/1GV3t
QDaFhkhB5mpqKmbsvpEuZuIag103un3B12WIEKK6p0e73vbuMSY3/iLinsiDddoj6s7Qte9hDc5b
vv1PIY3Gw7FYGG2z5WLr+dmnpAFBVp6dxEwujpsbSxBGx13PgSxl8NsYOpoghg4E6ZTgJBZe888A
8uR/qztM3K3mr9x1/BapvcsNTAvSYPSpkHOvuOMFjiOdAOFz9tgjD/+9KStT3MP8f0jD5o37Sfxs
WBChKAdqk1JGWRyziD4wATWwvHNHqhZFACGCoMJLyI5NA4HX8lUnkIK8bGomIKBLpIXJ/aqMW2gC
N3rueXKvAU3wtMEriM3a807Uau8qkjT34fAEGAdow39615jRiSOLiWZkWPYYdVnyQmdXtZj2WRiV
HMnTaHETZxaGmvY7v0Fg6wL8YpPk1kNCuWHLobuRKtGx8Pl/gJtttK2FUyMgBKbjRx3gxYHiX245
PudRswMFh/9MJssgqtXhZ9JbYe5ba4zmrZ3I68jODu/cAe/zL3qsM+Nwcd/i5goaEocOP3M78erS
gPQrQimw1Qa/D6eHlSfO5mASlR5Jt30rnBQ2ZyO0lcTDSf3JoeYNkROSZInWGlpvQoeoCzCgZ3g2
eCAsYGmJH/NHiA4qLmLnOYVUoi9gUBixIH/sW/pzGkonqlOG0UJ0ZLlzadTUTJEvrH0vngmDwSKW
w3he23WhxBuzCUa+Se6HSeB2uXQLLZtZYajuCrJyGhWZ73ERilZogpps2wUiO2wMXllk2iMQuXCD
0/c1wfnu2BrzUIsBn/a2aJ02zkm6CXKaWluHTRLEKKf5KQH5R/Z7UY2/7Q3t8S/VzwNmEsULbQGq
VF/85WCGiB3ww8buHb844tYjEutNjHgecJoIBMqHwb46tp1ewFAZ9A/BLXvlKo/iKQ0np5DSB4Jy
1r0m8ZFp/mho4zwrkla0DXyU5i5lBFO82RXpOgu2X5hU7/yOyVfcviUAownFkYGrzuts/ZoaFv3l
akBYabvWoG8QqGmkQKGKVKlP1Cxwt+oDkjo8YSoBf/Cq2fzqJFEbPcd+TuLFI30EDB0hWeTGLgPj
ALQTZCLgdw8+dY3OmcIkO3uKfbtdrG3YQJZqlBNswLSrGmsjgxJIDs5fuXk6T6o1MUxIda3+VUmp
ajyNhXibR0JBeo0fI6aptKWgRSlikQ0NBpK68OuqZJdDxlhkGApoaImqkApWEVlnpqmMAFSVbRoR
c12G9SRBj3jTnLvFndJl0RTaqA8UlM5kLtHjtab/FVfX8oIgk/CsKCNomRe0PyU9aoUjbzPw3Tfs
ZcvRdtAa+XMSWTBVvPWMOIBTsO2sKZZhxSknev9wzKPUpZab+OnAjDnE3TWMhnZXm05CGNPiyUEh
V1DtdMGaS49ecyxKx9jzgDk1osY7NMgtPO6IaFMMRiVqTISr+QZFi1uIaaSTbyfhO3lZQRVMbznz
bgnBmGG8D4hUTHlVDuGEjbazrstUaCFLn1Bwo8V3SWWQYRZn+LJZGXOpEEtkPLaFWCwV39KHatgk
pDQE5pNWWwogPm8kr10F8ONt/TtjdS/tNOf18vblLOu5EIMkQWUnP7d0k+0Rs4Hb/InXb6EEhZKB
s7ylsVWkYH6zPv3oWxigC5YBe/LehPAWgQ7xn6gEm9yIhl7wyek0ikE1GttQ1cx8t6DpFX2sJ7Mt
X1+ixz3AMDLLNYVCpLBdgPUXEqPWzpjoWLt1GsQRvQJzxGra8Q2UC5Ph7dXra+aP5VkkKhi5u1TJ
GmBsdxSbomznASr4Oti5aDJR0pOCF3Jph3suEYdch3Y0z8/p5Z670j/noQthw16xE6LqMsvt4kdo
gXJMEPfZb3UaqrHuAoUtPuVejZ1adZdKlu+nKrOyUyGpsrFbs13tY7ob/o0ZYbQxu7WPVPCCfaTm
Y+xi0d86RJhGtjEWUhyF09lypIbP0VwupguaHcNoVM1NVmaRgcRfDWjPxKUJS0Nle8iazXbLF76y
NpC4JNDW7Qho0/i4zZ2lO6nc6etik+nApEWIiBD/cnEdTGlcIMD9RKsHb60SBQKExkX04W5RgdeB
dXzh/1cQFPflW2Pf6jaZ9xCyQqds1oX92MAdghF9wsHn8DL8N7XtQyh6gaYKojtCNq5Ft2biw3hZ
R04YeWloHoDHRLnUgnF2rn/dpReZYAl6EbXWGAz3c2zRXlX7FVBPTTWbvWfJDjbPA/E89d/ztKKj
/0qj/kEVmdZjrmAUpmmEqFfx/HQDMwq43F2KuDQNBVgEaaKJUNeBm6jfWx5YSotWAKW+u75gl/iv
DI0xFXg2feHIJGOnyOrGCKcTVvqt36EojmArv0LFqvoIOeR5Gkxa1GLik7BrkMB2n0R4gDogH4Bf
P7Ue+vBf8aqws1Eu7I3j264n40ayu0IkqV+2RE8uInR9dBeffD49BPSGuopcQ8pW+0R0UmOqKuQb
kYnn6+rgIHpb9YW+k/kPxwfMMRipz+pMo6+hGRkVPdLJ/Gz+5mdfZsO6k1IgDJQgajPBNB7+wJpd
ifuDee+BiczhWAqbLYnwpGdUkBOQ+fvWydLY7ZShXeOAo03t6DWEheHrYJE5kzkbuhlm71LbbK14
p9rQZjqvTOG1n4oo5jGBbxB2RZ+KXERvo+st14nT1E9JOn4txKPzLG3fSpWC2XoMPGatkL+rRxCY
aqz4HDsKs6k2PB4IK13EY5rM2HUDtmqfi+nc8dfvmqT/7+dVhnG9aBKZbylJbw1vIN6AbGqKprIV
Dce5BGxsVVYwpibxgBP27kRGerh7/pCv1eUZW+Gbu4mr3+Fh8IO112NmY4G12vP6TERxRcveOPQ3
TEaQijX21g0e8r9DE2nNW5pp+Ga2TwwuBItxZlijCXfIl04r9idbp7aILbRBGsich8/YGJHe8f4Q
QSsCtjXkGCTSWeR8G9rcPcippMiyYtI3/FuevNs2+yvaZAfGe3CLIPr9tRE9auzPjCG5LZtlF4Fo
ATcpVUtPbTVF/e8aAj/ltViqC0V3RtvRsS5u18yRg0sCw/+F0o8OUv5cAxmXNbIC5JNEZvt4+Ssm
kHov2k0oG/phAfxUPb/+Evc4JeOA7xPhVF1fm54FMQN1gJsGetWzZSHhcDIRY35rT67RZnSbkBrX
Q3c+xwJguJsfWUtYNpS2vKotUqD4/sOySDgMFdT0V+XwpEk4zaH02vwOaXyEcW6o+rW5J8v6ylCc
RMVKzzKeQ2SmL/LiE6NsS7yVwUMl8bE2mVkbJATrJgoRl3ps59IsFXEI5+xdUmJAYt2qC13Gu4A9
GShNDrqTmu6rf8+ltJ439on06DtKm4zJTjaIdEZDkc5Aw9ylFiUkWTe/bbEksAAIPx8WagkCU6GN
XaYwqZd/7hwVwMsfP4OafUg45/GIOA6XXfhg8yh2Lfs9s6IKSvPijeno3h+PSfA/yOFPjn4r0fiC
Fk74GqYUYD5gpeTkh6DIB3QcJpvbQl5WXFoB6naYcOKquXxq29Zpl0o+3qEfIMFfFkcV0rhWyrYL
R/Lrbnmx5sOW4XHqezG3EBGuRIBZSNIg/m89WecEtVpoBlKjJ1Oap7WaE9dlE1MGOz6knlSfD7bC
qFjXtPhQu0WNLq6j7DhK5Qlpp5ZaaGuVDtyiHRlNO8y/SDsfX1xnipuTN5lpeX/s9TKH1ukmiucN
vFEmAOPZ6Libjh3dTnnlaTW+6TZ4cmzRRo1Nj8BJMI1ymYRNIn0CjGui3y1o+WTrMUKs7K7YkEKu
HG51Sjf8k4tpQRf5szZNDJ+7yJ0nzFCSHI4DRJBRHnxHK+c3sWvDqPYQZwrV+04/V+1pX9jJOCY+
mVtBt56+OZyF1Hm6EqUBZd6uhedh7EREOcv3TcVBJDsf+U+xk2QhOcR6Y/XVWnKXPJnnCc4eBYuH
TZiqZwFXiLRJ2A4dzxm+NxeMNdEyautkxsvqWOYkxhXXDaWBxt3c2rOo7gpqKXpLSGkiguJnc1tr
eEMsxAsNyt/QSwlJIL8ys2HQMaLVT6uuWJC/ssM+hL/eGz/FjL1vPVoiXykNNtN6AwTEfOi3wtUn
Z0M++buTAypUBxdrJ1KTil5kX9wskT5RDlf+sUTsLiouFbPZzdlD2bnMREkhVG1bK8mBlU59IRFz
lsC3xf5GMyukxn+kR3Zj6ZoGOkTwj+EeFUxH5C2fY1+OZKu3PAtu5eT9Au0sABrkLCfi3fmH5C2F
LX/awclqZPtnqyFeoHITNcdPcZQX5X0zSc+Ots+gmYdPnU8D99PQqIuc5G5L+D7F5OQ9A1+QwUDD
Mc0vLWCANrRz6JzPolOfrfVeVJcgj93inrYlY7VL0lLihVEGrmWcoR8+yv7AhKL7IeSXWKJh+KXX
nhBGCTqY5uqCktyxvVuBPbi8BM8o2UC/nM5GSfteGlUnoOmskJwGKXCQ/rCf1gmoTNIYIHwWsLEG
/paCPsE0renca2TKgufSw1mrUAbZvWqFCVoPTT/0Lgwvo/CtXbNuRLfHV7rsQHIaHy4FlA9jL8+P
P7WlQg3JYv2rS3H8YNBJ3qR6d0E8cq36PC1YipUyPUntcDw22f2hXXN9ehDgpGYsWvB1JwfBxPdj
wqUqtmUSx1CyZXp1dKY68P9f/yT0hV5M/g046cGao4D+4f37UAv7BvHw4ETvEKxbmpePK1q7T4Wr
+qkHrW680nf+d4CHLE2azNt9H7RHpLD2RGDQPPWOG1mPbbKzCq2q1yqW1QyQ1PB96hM9PfNt18am
Q4yXqiGz/6Z8OnZxBcm3Zp0/jiQnpn2lRfvSYuryZtCBOgtUKFHrtyKOKi0PaRbQfYoSlv3lmGsS
GFZ1Qd1uGdtn2zgD8CpzO5QCKCZMmGLoSnMWp6HI7Lw8EAWYPJFpCEEId+dgtATeMbiEmSp5oqSy
tMtqT3THzrt6Jk9HfR+KnmtdQ3+vfMvHbTEpoZ1t+84RhZzQ4zkKIOpyuGaD8RMLQIroM01rl8C1
s1HtAH8NZ/7eI2wh96aYzPgANbc2KC2PVGnFfpZB8lslaqQgTPpLO8GkYg5iym+6TKxSkeRPFWPi
aGaA+vTCvsyiWO90/IrKhE3LoaRgz+Ge1p7JDZ3eEmftA0nJGptmTuLF3QYczCh8WDbM3loAEtUe
FDoUzRkYPGuRhrslv0RQfcyUIgt9LsAa7Kv6bcYwspzvkh+qTFaMX31CK0BD6nlth4M2Lzmdiu17
/bw8oR4pmhkXGExYk+cQk2GEKtgTZXYQdVpoi4O3A9yOymz0LsjuWtLdguJQXCIWAYZsdJhJFo7f
KqCszECEBJMElhZXoCMMC5Vhr/u+PSPgQwd024xnW0kuY9OdHldudUodWCzKD48NNlPJn8Az4nY9
w0diCzDnLcDml7FgwZU7/zhhBKIyTINpyVdVI8V0/W/CbMFg65rmfml52Oebv/dq5w04mYIRKcoW
FJ9y7OVzWE7Ja5GoWStYay7YTGT2uXxMx39JfSGaomYjVNSjnfjMFznXsYTCZrJd/HVaNi2I9alk
tRb6KWaSi5QX3ER1f5x3sZydPs/dhUIuQBhq/XgwP4IjufIzwi0PDmE7YZlmxX0MpQDdxBDz028Z
ujkL8YH44RL3wi7lcwOhUVgyMie9u4c6TG5wIr1r3fG5QtJfm/Iek6bvl9jtYPWvgv3wXdadLkQt
DhyL8xjYGpnUSTdUoG8SbKaJII3WxZGEJL7cN9KxnXvf+0vn/5BIzW/4/U75+G7PpheXusKe+LQO
21r8qJwDWtKJoEdzzww8/xGp4AAJ5tiv36jsUjlaCD2FTax9P2F6Uh3Bm5aMrzbdavCMpNozJ+wb
FEU0vT9CDdd6mjl0kVDCIdBIOjBOnZnkeop7iHEMWzLxeghK2x4V4NQfAez81lcq4QtzTXHM64b4
Qxokoz1BQvelCE5F59/7RCiwPL8KdEFWZE9RUEyvic1lFflNCC8ZiBYzHPwUa4LbXC+4FWLzpDFQ
iYLLQNAF8IEqKnhpj7J3jeaMudRcVgbD48TTFRFp9lhqAg2z8cU1K8KAVI/WYc2v2igbVHj6LuUZ
YX6Kg2XNZ3p/YbdrsBa/YHwlDSJdnw1e7q4RQmZ2jYIcjV1FlOY8ay7MEUdpuQ/LU3fpjXMq+31j
XQxYoHlUeEKhJDnP1zlpP4/x76ONpu2mDDFi6OO0r3wtuCa/A/GgEk8L8mncH8cdv/YxlmHPu9FU
ZBEiLgeBzqmjhxYTgk/NslLRLAJlUTZ47ekpTKesvEekX1anjvyuBD5rcNgp7eaYEa/q9J8OkzQk
Dk9kPIC8csPVzOfmvIpcjcZet3a4/m10zb0s/dmQ0MHrno3V1ZVF1gCTETyy3jVDmo6M65GFoS7s
s3GIWoh73XiyWBKRCdpXOsZbKjc/EjTrfyqHNsOKcEvv/U5DQMNnWNydbhTKvoYOn7Z3pBZqfjtk
C9sgskIAXxARL1aWYqlNn6sfThqn2iFkFpC38x8XlSUd5oJyIiIRtzqjjxReNLFreQedMzLmdvnj
/KvkakCHXy1B8emNV5C+sMjFlK0kfb/GnIm8BL1wAVGNshliPmXY0mAuFygEiH+258a7OzX82mbj
dQtq9CUjS4D9qDRdKCz/xQYwTNdKfbmCwCSE0NENIKrkffbON6Hq6S4ZN9TTq2ju0Ii9Ec/wXh62
mqoJerVIZz/0Tpa8Nl8de0ChHE+RXFK3Ipckd/K3Sy2wbJXBHg+6qT8XDWziM2pcGhSgQ2lVDid2
lJeHUEC+vPG+spA8o1wC4IpTbOU8Ky1aovYi2wUY0W8BTPwuahKo8r3HWMR20iAuQB49L22t7DYi
dKCQH47MBcOVz4Mhl0mbsCrzI8YCRTz4F0rOHprMSNS4/Nsy3Sa1WqJWfqVmQI3Dcug+nP9fZkua
PDxXZZUYzhqcsxaArq2sfE90oqPPdPh/oAbcr7s8SOch3Mg0r5eNruU9TolCioNaR5IYWhx69nEk
7I21GBnfsx/Ptiss5XfsYV1QQB7SNwYbaVGgm8Vra5usbZxuL97XsLo7x1ajB0P1zLQi3CJQY/yX
BcKHUbdRgsV3D3jSSG8oEAqt1uve2nRdCjmxAwKfOb1ho0qhrQZoIl0TQdLQPNso4lGt8gegduR1
j1s1RlvCsNpx+F1nE0W5fBP6RrLYh09bMKxWoLt5as4AK4zTJLfufBKkQJPCNdngIKYFuyuHBlIl
Hh1BxK1bznBqhHzdWV4nNu3K3+wEqYjlCySV+Nhnq7SYl+cJsAo4a7uhzwKfnDinsQDYI+/OQR6l
AbRowLVNQmtfNakCYIsPJ3cFqmKe2EyJV4+ocgtWXOhTqwMAhH4cISrlfkVST/AS9QKImfu11pYK
BtckdNOf5D8cTStwrXexz4kwXlKXcRfSEIrEyvDH8iQLFylG/IAhtBCzjcWJhMIibagj5fRsNZp1
UNvFwSmvHFVaTt7qgdZBTyudQuxKlJ1UTW3EL4vH2O4dJFe99aoIOLHup9VM0ER5gLuKoBh+PxAu
pq9plthmZR5dZNtkYoB6VXX+Lopz8u5CQJMJFeJRucEVm7k2Nx+EHy8F6d3NwEgD19tcEehXUuTT
IFNeV/XHml6eB9sHRilMrRkFQXLtTRUMaZrTCiXg5LsB2CUuDXSBjcesASvD2oSjq/DkKoYwRI6Z
Cfl6P7gQ5QJJd6MtRBQQ5R7oxt3KezE9jxmkZiNFmdh8SCDQOlqP26qTdN/qh0uXYvwGINBy67Gb
JMEObtGrFLw600l72AXm9N76vAxMRZdcXStgjyGM3MS2t/3sTj0/gYvU2KWwSiORwxb+zqptRADq
UScJJ7Jse3BnTYGUWSuXbr9nJMdwc1He9y7uSuteX4leXqI9dwOXhy0QyQD0BhzNkw8qJtXhweHr
zktGlJcye8dlckOJT7Iv5CAnlhMcOrvl47hqSUj9hOvpOWTF2YhcZS8NJoRhxT7u3eRJcPJ1hZTh
vYRruL4wL97QScnwbW82dpH0HSjwnsXishL8tKnkXxw/n9r9uqSfy+2lbjokjIPS5qDzownxskZS
RRw2gtJyHpINz0BA9bAHxalzPZTmhWxrAPqfwiYx4nEptNMYUBWSyCroTCrl3HC6g6a/Lr7QPUVW
57AYojYOo1AjNQL+3Ho/j9nUFyR9H/O6623UEWjTU9XZCvKtgMuvrgG/XCNpvgrjgHCYNSZJmxsh
TVrT0ga/mYQa2CMq0cLNVIfV6aMq8RAcmA+ZtWJWl23QT6nM24VUSvp0JSi7b1zGHV9ng3NlLCZq
izD3SRn6tendIGnLjXW6CNXPZ77UgqymIpXUyFLqqYgtigXoAeiofHiSgup4Pm6hrxk55Y4zD+Bg
4wtO/WHXtPSPmq8YNhYvKwf7Y+39P/kYPtPB+/9kuhVwJ33CPJnhhVRWEV8oh83NgyZsJ09QtFJY
cOqUKL6+pTC22vboZfzIDgFjXebHvrOuMDrtAJPAny6F/kNkaq1IOU6D9Guzd8DgLqMyzdCmd0ca
eKLq+qHBedkptC+8JLGBjHh6kHzObCsS1OQQX+ian9ezoyXWFweiaqtqI0G1uCAMo6tQHHt9J3Bm
1LS5FUEpXMSLj185eoHJbXXLDkX6j9qR9eMetVEMumHyOL0CnldpwqOo0Avn6OK2TNgOpqCutBOD
+VpRtZygLEFSTgsrCcVZC2fqIFfZg23bpCk9r5f+NIX8C9pRQiSVbbwaJIxFej39rkZ6KJUX38wE
wGaDmdyAryk2qVumfZq9qmJeffirRlb3iBhnyFd3W6smkg2LhJPOpo9Es+qRnz3qR9nNrJadCX1B
jgVdf/4GdZI/Q1YlsF4xfPtHP3ljwEeLtlD7rpIzv67bJcZ9kiqHbIMX640c8fTP6Y+uCgXMO9aC
TLP5Du/wWOYWmS6afDCjHtEimc2a5BKlXYwoTWYsstjGZlLSrUEIAg8su4V9boH8TaqTs4WeSBg7
fPvWAog/W2UVByRLKcdWSdH5vlfXQ+l8x+Vf7iQMTDDW/NNSL/66bvAMcPeygkmShTQrriz5xfGe
udh8RHgqZt3BvtilAmJBe6Zyn/Niloyl9CaZGvAGaMAhL/jJqotMAfk6u5onifFn9rcFDN6afxVd
1brWbhjoZqMzW9Ff+cp13UatxInxvl0pu8u2Yy5RUSwJU4yv8GBgZPOyjt+Gy4xydiOGb3FnccS4
0f0qVI2H2SvdR6dr4YF035Up24TCGgglM5pQfzjwolYOLJHUXeTu8UmzaQhcDv/u8BRxIjlpGtTw
5zYb71kdAytFOxBW6D5YQQedGmGsrvXVF95+P7zNkEb2vQHzqoFchgixP2u4wSlXzhgm9j/w0HtC
eUewFhv32LnF4K/cXgfprdNJjmJj3iXUgvI/Qr1CB/+Ssrf7EwP4hH3dGjyTto3kNknUEjmJk3G8
ZYJDE2pXV5xH6gOvc/ilsqtbywtSJAucCsWxbdW3oxDWc/0oUlsuHKhyx4z7N9zRAU+4LbSeuPoV
BMQ6rWpMRCNCqRdRlTykhz6MzlsoqbDQ5/97x8DmlB92jIOyOfj69cf1RgTmjdmpPhzDCX8vRKq4
F9h+luq//5hh8t1Tfbz6ZbeOZAT+mLgbLkPz9cSjro+xRDBrN8umeFGcwNQsV0iNCeOneMLMqwzq
Lgw5lvLZt59xN8Bpy1o/gBBViIjmhKXpaPSFsQXGY/FpdhGtLusNsDRB7UYjqSbArYXl7thUOAG3
dedY+h09ne9+DbfzV6zMh4/wCjbLylm4hA5zYwR8rXi5nq8Iod3mQa6eG6fereER60eW8SvwE4Mm
Sol7ofpmxARxCiu57KxNWGGlDOzXuuyd08xzxx87LS/ZLqAJ1LTx0QV6SiGFNrxp4fFCtYp3BeXd
Bxs1TFzeGXSrNi3ClXxYA6iYQKbDNtW5ikDKArnDpi68xAm+aD1BzC0d8Mi9utSmaXOPh0oY51cs
M90bChhEfZl8ZVDHIkDVvpiuk1UbZ1OysT1idsEOqjs2xyzn5625SuYIdSw4vyO7L1WlFpRBZeC1
fkgqSHY+Gb1whZSrL4ZL3dlbwDbZTr6MUw3lMTk0/BSLnkJAWopEPwqC6KsRW+r0QIlNjPhUCzc1
+bSwKhczRGmv0DxZ7/sHVG0aievIfJlKVxeTCHYyOkixG/5dTjXe7Pk/7Vm0UGKmzHt1QAeNphE8
0w/bShCqN9ZVC7bLu3WehTegH5zy4Flw4raoGWR2GRaAAJ1bjcgLHOU5WG8aP2+KvKXAyrsY6rAP
qZJtuG6bUmUN0l783Ua7xT9JQppBT/ltyE4tPDD8mnwh5y1V6d6mEOf/bpFRLe+UHgDPdq12t81k
AhaXCcYCV/dfoyU6xTR9Gr8ADqNqJq2mwq5i79MRMRRm9S44HrYeqXWL29f2uvWg+F4SD2hwgN+v
VbYws4wP+ZdI0IJ+Hc6R1DLVzJCrE99Ynj4EaRrQMrPvhn+OoTRIBU0Tng9AC4W/T8hyn2zmnMai
k/Li6qbay2tqVaH/cJfg1nI3+gxvSFVCIl54WoW3S5LRnJHR05NMeihQUvYkY6bBOx2tL1g2a+/i
OD8M+qzqMAjkxV+XB+4+Z5ggL9TDhFEp8wr7BiHCL+SWXhPczGSdSW1eWTGDLrZTOFGweyDRTydA
D0boSEBj1CM4nMw+vW2rudBbV1puvkSZv/kSWJxPpO5bVrfQWc0SyheQN/1RQqoAXeQExRu8Lu8l
mrniPZGT3yvTMEaqTQaVEjdL5Bw9IsSozX0ekL6Zpdae+ekhpVAWV476cnbmBQ6hT0pdbT7VWXVu
pMVEq4HIHWW32qtG7qTfwzAvyvmYS8l/KqcC4+PfYZ5xXclhGn64mlHDpiljTwpaJHumqu3ENuaz
JuuPXM4VNY49YRLarnxwdOumTyHN1osE7wJCYSPKPsSOKukQb7244+UIeL2ovswWVnPJFqVmd36S
ES8e9FHwdMODbTMJKpZsLwXzMv9E6ixgRZKeIX7wlUfqg3NGvFSLCwAwPJ3mu+VnzQ0t7x1YqFuD
i3u81Her8KsBczbIQDGE/I6b/6EOncpiiowG9GOZAHQcVB0wuxDj9sNn4geUr93pNQabsBCl1Qwm
XWoQEYt9r1G8GVqLAd1ahn8wWuM19yRpHWjs9SO/BiPw7xOa32WSM00OZHH5xhmc671vs89Cz3PE
UGoE9LI4UnrrAFzmooewl6NS204MCJO/l1DPc430Yl80Bwmrv4mVpvVAj2V/Kcm1mj8lNVx3vuAB
+XZ3r0cwbC4j1ZaQoIesOEookkuHpiST7t9C110/E0UtgXj4PBQX2f6dDnTHsQECa9VvFyTyibXO
4Rkl4hsVvxJU5XKsDrEvYhze37QyCSkTHH+592h/3dckZ/wkphudR7sZ7dQi6vGaiKjgU7tYfxHn
fKBm19kXbZMQ0z3AEBKPXPpS7RdJj5dp2zIO9bqmrGUR/HAZYdap4PA3SWIrtoR4AT5wqqxTpost
RjZoBqXY53Wjg3HkmBP2AfSaCgLlOlzG13dLCx9RUNOQVB2hqXodwQc0eZAtU1oEJqFeDNEKKsK1
lTHFwNrGuPaeWgO+o0SF9kcGr3fSknqIFnW5IFkqvYWGuwpfeXyMwJUJNAaPArVJ0lE7HI99Vyfh
QgrczwsKgPradMN6nMzKD6lD5OkgKr2LXZ6iiCyXvDGtcqchDtJjJPuho/39zAtnAh4L8IPlEY8I
eCofnVfH3CRRrkfmA/OvUCqSSNuGNpNsZcHH6saJHxvr59FKheT+ljqIZX3OqdJ4PlnJUGrDII93
yOpMRLreE57hnQEIM66qxCBFburhMbH1Nc6wiwlUMVAsDfTO6w7u9dNDJlUsddGp+7KwDrhvIpYb
pGZ3VJ1X8fb9QydrbW7/NsyqUW0I7NO+EWOebeQd3RDnfpiH2t0YZl0w04ecG6MH2cj5HjMaLfB8
81RMcKebRTD44mgK/sZ0i1Ny3AeIUXDZLDnEY2g4PbRGfJgd7lExaxndRfNFOP++lyYemGF9UBCl
CaKjzrzJGtCV2dkWLS+P4RpyUVznKjWQ2w5yctaL2yPnjzSsIyawBHdtdilWotayUexuhuiKKLXx
S+9gJMAmdkGFlleFmIpYsmzgpGlnescQO+jKxrdIl/MRBZWQdITHUwA45vDtvNp5EOk87zPeC6+x
e493molYb0eKen3wwKJk9+ndMQP9VqgNSvPMkBVeduz7vhA6qaVFObBuQiAVLTSvsUM+jXPlHubG
nfBx1JQWWP8FC9fjI5LaOoL9mNgm+Eg74OHxadJgSYZo0WQB8bQvHyTn0ulHUsdDNdxYgFa/pKNE
JXIXnDSZfcdZgQa4RtMP7XzKvJSJrbzlI24KV7VD0fbfF0BCSQs69qD2JqxleCHAJKPoHKk6+Ydd
ncU3OY3qRftSlI7PwH2+qCWh34My/hlHYYsDOY22ANTAyRLa0hDU62EFc5FCQiIdTQpHUpr0ak36
XgYjz1QHXil6yMBTFbkBfpHUDO9v8VQrIW8NPlYWqaiqEVKHBdJjtwHuZDrHMxWOZY7vM9rAgHMw
u8GAdto6umSpm603SuKn87YU5t8UVDtt86LgE5VnejDke2unpVs6bGH092PSCTforDZEtFTVxS1a
7wMakV8MkpTObV8pu75qnWiODjRDjucChzm84jouGF5fQLa4DRFPGu2pHayJ3OY1XztqWeUPLooe
7+5Tok7HysfkslrJb72apUejhDoTRSmGy4FDPwP18CpX17txQ9BKE3kU6ZqM7Bk0HtF5Q1tmVlp1
ubLcZdIVj9i0SG0mUUj9uH4/iaRl9pFkmEVohOPu101lz3rsaeCyx2w2q+FDSmfm+cdTVIgCLhFB
Ei7uTqLhq6DK6xbnLSQe6xn4ngYid0Uk236IIVXzmrSUnsL+V6NEbtp3rkLthhmgrtDXhyAloI7m
s9fGHXYA7//5khfFSb1/FlvqNRX0ncePKUZsENsQAuDhIuG6GBeavHCCeGnEzPHEGyKdOHriSQqf
NzKWFC4WnGvkC6W5k4hRt+jFALQC6nCgI3dUQmK/cmBakc9zfrqS0BJV24uBxEpd2EBoAmmU/c5q
IsHjdhrppqfgJbkV0QuinuSkQiphy/EuWF3t1eLv9e7YgXoUCSsUJvHEiO1bndisUJ4P+op/mTe1
jWJvRiYYW7sqqMD8YOd/ihXRONBUU9o2vytOrCq5yyYhqFnBWaiVmUNA8XOCZqV+n6f8Opit8ZNv
m036hvGBmJqEzLD+TA5NA/yzt6WWGLawjhaOFE8hhbPPxfY7MZqnDIRIdnuKNtBW1GVQeNGl325O
BAX5AmCZEPOqANZDLJafZUOtibBIOSwYvyM+6FYzUAmrmAY666JG9gv+RXXcBtk9zCM6zOYbcOTi
SwXgU6gtQ1NSRVKFKdY3Kh+VixXoYPWd7x2wefns4BoYAFMQED73n0beEv5ami3hsUycawyF1B24
a4RGbL780bJ67BAi2KwFkNlp1Vr6Deh+Iuqn6WU/4PzpLo3Citl9FTL8KvdoH3sWq/Gs1vuEtrn0
Wy3csy+h7GSpAnlZESuA5aapd+VzMTMFVO7WDvNLP9iUIgnBAya6BjURCTuAwvS4upsFbRJyVu3n
s24VRZS4bb647Vimog8OC3ua1q7lbMM2ILlGiyaH0BleMvHVRcRsHRc1Pzb9ygCHs+wMGqhb0rxT
OotkQzLVShDGYIeD+7dcUh2/w3WNx5esm06oM389hSfaN1ZwUqnRXRBIZbdeYkDfObiL/xVq75ll
fbzTcrT5kqFaWnEX5xyK+0RfRQZVaAvANMjbc9g5kFR7OfWRM0u8CUSe5gu+LCHj+pe+U70nv7Nl
s5q92mfrJBdmdHA4WkBl3l90L0NrI2asOnj+2r8wQ/F5ulwtyohkCz6SRiJ4wDLispRrW60xR7cT
/8VZyfGbDC+yYkho+NoV6rxzc5sIMEQq0wAWox8zx5iVxZB+klfm1mmCAEoj7RzYM5LvXcnHqdMg
2zakz8m8Eh0qd9A0zcX8XIfP1tJDyI4xFBFFKk974ZN2kuKVDBuNRoblP0QAxsF6cGHeQjLpNB8j
dJjIpxWN7MULUCwnbDHFUnrHOwFJZw8kPWJJGuiGQuKviH9sxG3sgbnI5zBmu+fS8tIP1GCb1TrO
fDiIuTjBx4NKBaSc2djBaBtRDRZ1LgYjCaO3WkhSHqfHW1PYt9uhT6aQ/2UzWZv/4ViTgxFGrskr
zEJ3Hk5bWvKeIIKrerq9o80DJYQqVr9Gl9AvjmHxht1Cz8NzdIljF/K/sAV+B+2rRtlQGYdRfeYZ
TGfQeWk6Bq03Kj7whDK3xxMLRGjzIhtGCj+hBPI5iWv/LXu+T/nqstk0KLS6qQBSdFP84gLb76En
IMRhcak6mbAJS0YPQ9qR3Biie/83p9qr8aq94OXbqLhCPisJvs11uUkTnWuuls9Sx4pUlO62Ozf0
N6HAZFNCO9oSj8Pq0JTxV4JFogu39W6JJdBdBliApII6G2ehLhqab601Fwqsd6e4OYg+3NkH1/nO
wPiNXPzStkN1FB2adKDDX0aQeU8bOTRep0rUDz1RbvSQAWacma0aN/1uC0MQrzNOivVVwtj66k+E
MiQXCtvao5IV20H4LbzWQatKofroWnCBgbtw/ObHeV65pbHXaAdq+WBKL/8h7uQfhtGE66y/Ng4J
X8R1LD5h3RTdJRG+IGjvLXhmN9jiLgLE4QfGJMwQPtkQtxNXaBJ0ogyta6fUDrT7ZRVutoOF6ax0
kQf6Ym1Z6eh/OHl+NrYE03YXbSI1DsE3bHDTM63E4yQz2cZ/woZ76g24Qzuqg8fB9nuSejPy9KLE
Fk2CVAY2M8nx6lpjGhG2FL6J51kNbAeeWTEvA2fH4PBTftdvVYIbF1g3NILDfarN1a7hFRm00CoM
LhKyxHBGLQU8Wy4SMb/TDiwn6Nw6SBFE1ElW7qJFcgXid+U7oOkl5PkHlZUW27XtLxWPiVlnPXGg
Nq89oxvPzN870sdTRaPJ6TWh/SYUQb+kkGOHDvQpeXO57DOGM5yzpNDxWXb1/m98qLWsaxycou1m
fqu3zPsSne/qsIH+tK1PIto3jb/PeXruRWmgQ6c+UsKcohB3USfZCZy63nFqPqvHi2wp26eLZDsT
AmuQHC2D8+c9cNbJqhCJ2hHV+gOwR+QMZIAxJFo4v3ee7CFmPeuKCmjLWS7NIVT/SvqBpghT7Aef
h7nSNmAQE580rSfeJjYrUf/K6mDG9RlmlbqUD2KU3c7/7GUukN/8KH9+egfjgeoSaEYaz3ILrxxp
EeFt1Xp3SgU9ZI1zudibkjNQ+8o578tLfoaX/swqh+WNMOOkMrcruxN4vQBBmd/651yl3mZq9Bs3
6s/5NoAKzxE2UWAkmXUbu3rKOh8SZZjhXRL1HitoMuyufdn8shbzmHC9yVqM6Sy3cHFKYSnbOkla
1qrBU2BDyxCvzhM8i3uTYdnCy4nkIVBuGf3rSPbVkYt+Bx/xd6f+yOrjQGLiVrBUE2mgPhOAdTg9
584YIwEdPKEKUAmPfnNWSutR9Xy9xU10Rpfy0IczWyKg99sb0WO55iFxhWZookhbD8rAEy62+OE8
9itPtDsGMDACpsDBKDc9ZBJ1djhD3pLZ5u75HGoUoTZ22lUM0I3YKy2Vdsh+iKPYARJFOA+JcgIy
86TYDFRm24OT6xMjXkRjpsgwFGW+sKNu7sUsa9RQW8vid1YC2wJmvpL5gK1JL+PvCPB4qvSSVpUl
Qnoc/KFYHKfDU+iYtylZVoXROX5jlGDFF5Ig8jyDiLPu8TXYAYBFfuprXoZoVk1vSAtG2IilNdMA
9sEuwbXss0oWL6JZN9+7qV5eNy5K9lCZ0GIqdXRH0oU5/8i7+EhTx4osW5nD1AM5kk8F7r6kX696
NYXawM6s/hZiTt6kP6VAv7kZfDX94I0hVDN/HB3hx2AxRDAb7NgGWQBN3XfaDkMTLkAGQp5/PsCn
PHne5eRpdYWOzHNKTMfcLlV0/wh17rIOWEFdH92e0bLDlb6LkFtzjsTVpAwFBlhZdWGKFdJCFx+m
UY9cBToBkALAkmEB07wgSjZRtLLV4mjG/6p8eg3xueb/BnrXSO07bz8c6jqGj9RjxJFjYiUnVeI2
IhiJSiDQET/tZOlfcGXqOwWNSJBRHVihFgf5O2k7AgHbFgXVXykkKZbvHcwjbfG2LhB09SBgQ9Si
RgRbKVZgRmqqouot6hBjaX+f9/eNJkUxH7byZP4PKN5zMYEbelyZxsWEQhcqtMnCjmxPuMXbkh7e
2uEsVxE2Qn7GiyNPZiS+1YQUzy+1xNTCS0yYa4vqdDOkJboepa26dCF/cQlvWBz1gMDVyxBVaY/N
4Og5TbRVugYT1gfpdEPXNFVEI+iAMe0AuWXQbqoBXYej622Ri31xJplUB9P6JpQn96/MTIWSQ3V3
z3RGTfa8UVvTl2sXl9ci1TIqFr022yKdl+GaZ5+OVDjhfHLAXNiq79VkFw4BSMuPzdrigZ3hSCb1
eEpuykOeaK32stoc3In0egDmJ9JgstA+prJthTTpyj/opFWNjj99QEvcvclfz7JSZ04GQF6+5hFb
Tua+eRWgK9fud4z9BY7CLwS+elRcY9gAIEav/sKaLXdv1MfVqJ/Gr6VTHNHPA8tus4KJT0A+2+GX
4zN8p5xPH6L3EG/Jig/K2BeF3/+xXawAl0bg7bBlUPh6wmrRm9fglWrD6T4UTEvDmIzl8Eat4OMT
GwHhA9fjmU/Oy0ii6OktMZEy5mEc0p9VFQd74cnVsUnibeh0A4suI+inQYOn59KYFuQhrA42JqB4
WIv2kDSq8e9LDaL+lBugtfJ5qKWhkgRDLNt5VqyUwhNjXDgcdgJUAGlRbL5Gd77ZGAeQH8KVhFB2
2CtxQOxpcAjpkj0HmskzGu3L00Yf4Bh84k9PWx35IE4b8itBhoVcBTQR973ihRyXWlJfqZ502L9k
TYbaCOdq6Mfqd94Ze3LMw0/wSwIYRbUngSIYQJKkr1YDBihoyG0bY60fT16Zbie6mPLJIuI0JkrF
dTFUtVCdE7iG6C7y061Ypj21GlG3e827Fdh3EwpO55IjF5M7uMISIDTIwuy9xBTmWm07q9V4zAMJ
hzLUQVR/XkbQ4WzrEEDAbmLJwZnj0hMBWQY+uQ5L82A164sfqGzi1oKITa3lAbtrUbxVT9ZTkWoY
kjWBR5Lb0pXucwNZ13omtwc5DPadGBKHQnovDp2noTnS48TJmRaBr8lGf27at5y+iXWDFUc5osYD
CB7AUsU5Z69ioQFJQjrh+pfp7L+w9IXviFyRchrO4LdVQd9d9MEMR+RDx/KrizuDpr5zYKSNMLqF
JDYT2g377YD+6ZUy4vcqGJMzUc9RR8SzRCyGRM6dU0y294skiuXJfSgJm67MnndQZqagatH3Otcv
I3VM4Qc0CngVEGbjdxRmXHT4no+7vW9yqZY4UDo/Bz/m8Ybcxvik7HOx/NJo6WsaarYgDwJrveFn
1BASwsb9TyI34WfBP8p5YyngvBOxK81BBvlb5i3cgi/8kobQcJNkuxdw5ZJO4DhDwubJn4TtaXDS
bBsnjQRIfSVjRRU1jL8Hh+r/5a/NXelascdNhUYRQRjpUryWmB0mv63a6NHW2QjWOICo0lrv99rw
l2ngiDxEBjYn2D9YZkJia77F//F7YF6RxnpvsyEMnIsKOYUXsR+Fvo6hWmTRKZb+ebRMuVcpQTtU
qpH3XLCir3JBorV3ZMueMMBw2nyzUmhaNQeGxkRPgLQDA6Tk7K+SmbTKh2ZQcGCy4MGATfvU0cqz
gzBz/lpUUC4a+F4OYnibiJEJopdETI6Sx+Ncuodj6J4/PAe34Gi5bWoNm46qjDbmyZ3dnvT5cEbg
GpQLsqt9ishvXzbtKBM8+xYDmvdd2LfqtO8rsHEme7AR+l9xn3LeILWTXPEstOvxqVMvI8CCECfO
CO7VM69XH2E+vvtTQ5AjL1pYvJUMUOGyi43gfQNUM082SY04bVnV/qq52VoRdmWS2KGmkOaklDuV
BX4Nhl+cUZz/8YSfNAgaXrSgcnhrcmpZFtd+7tUNM40qeDyyaNy4mB3UYiCinWxk0eqQ/vbmfiV0
Gyz9y6Lh7ZGgx6xe3sAqOp6kgci/Reaealzk6ovKFySs4G0xOZvF80grhEyGS7jBmNaVn6zZClOa
hePAsMTITM6wxiog6qM/tg5L8Tyza+y4jCF1nYARzv9+IS8iGluGYra06Wxgrkxx4S+AMDEaNs64
BH2vZMpUxqy5P9emZvSm0g9BqVz5hwrUJ+Mm3mi5/wdBkK1HU+1J8Vh39tQktuTKCgs54ldGPfpl
jEpGTgiXqURPXexr2qdJvE/88cBNDnXVlg41jGR5oimavZZZ8dGtlLk0mSi2F+MeYewrJ1lPyScK
tCja4KKc09wH/K23wiX0YPgj/WFD4p696Rtgas71O5Jnm60pE6NSN+okc5ZXUefmcksAU0BSkVQM
TZ9VPH3RJ7QOhueiGhd+fKjv2Rx/ioY6mcUN8UVFyfrjhcsxzHX33H4obwagwuNbzUKVgKvtxLHn
G037riBM9hcHBu4EYswsm599DNVUNN7LWd0U2my4fJsu36jn9RqAVl1tCxCifORP8yOlFH6LlynO
KTqo2GlmaJNADGcycdVMk2yISGImEzy5UtSsODPP3CoYrU1zxyV3ZJLp5nP1XBR/22QtfdONCQRw
0bX6lW6WE8n1rZTVjZfOO6U7hgdUjUTytGjiC9TIOQp6P8EnaEIPljjpaaytdTP/YyMhcRwhIiPo
QTxYodgtrYeYWxS6DjHeOctcGrd/rW4tfqWdLGuf1hJ+PAnUQ2qRU0SeufnYd+FOCeWAi1N3KAIb
e8xTrlKSkbFHYra47KGtdUcBi6+vi94/q4DXSGLkplnsfCju3slsXcJRSWcWrKMddt6P3j49nWlQ
flwvol3+gshhx088i2wJuZ3BcNe6CFh55puuLDmXDouti0dpZ2OYifQqbBPYm6eFsIN75DrEwDfP
AKS10Ep029aS7Lb2yDOo1ka1703uui/vkqA70/MhZLEj4ullGjSFKr9cxx8HjSRxjDLdWyaDnJ+W
xY3FZxSTvSyJk/P4mMu1rSqmucWUAKdqYu74L1UoCL8F0E07T1wRpnzvtUeinsVixkrioBcGE4eI
4+csIWMcPfqSBjibjy790XZ5h+pJH8VWtmcZ0VKbp6WwHS6vuGxRZvUWRX7kdbJZmVP5SxSjQslt
arcEcoYbK+CAN4YX+QkYX3d0giuTOcJNv+zLHlbPCH3d4dg1zt4YJJ0lj3xDxasjzuJRnClREI1j
4imRWtYTaGpeY8Zz8Xyo73gFsxpWkoslUO3AtbHJ5xc6/b73Cq7mfFHdEFYo+efneAIdnMCIM44a
wYTwRkBEJHocT1HIeVl/ws6xSIp3vlcV4JdsPIG80no7VbZey6J2gNsj12hf2L0EEtcLeKKnmHEo
JgECT3gm3qYjjB5mx39W+0cQGzsj/0HXKm4/8D6PR/aclfE8jbGI3rHrV+/Lz3N1FFn+O0o93vlJ
p8xoii+fn12xshgUhaVC9HvQ7fLXwwQezwHwzxUm6TW4xHYKm+ZVDJl67BzipDlQxVFzkt0yRCB1
gAd7ThObFB1DjE+tn8MYRRwd4Vvn5a+u1+PxV2gIAHlbz8gI+w+w1mFgFpoICG3SN9KlXYx0PUNc
1My4NmKGMwAdOmZwmX+QJck9ZeR5RCGJWrhdko3bR0XgfG/Be8f1sQk/4oxcwnCqSz7RCqtaHELQ
AttzmgPfKaC1N4rj90veGV6xR9MJo9CgHuYTYbsG3F4HmgCokqlXq1FKfcnCSzOVFtmKj9Swm1ms
QWvCZ3WPB0stH6sQxnxtUY2qKfzwUXF8SeWe6P8kHkaPYJd4pfsHgbBDuo+md3eUOPO8T7d8VdPS
+6ib1VpVcKeC4C7RqQ4GeuKS/1ML/0cN3WByCOXb32lPvqVAmShlUmhBJPsx3HXN4OSEbCVzHTXc
9X8HStpz8RzpFN2rU55B2GEPWNZ2U4ZQeIK5ENtQlv0ID8Zr2+wth4+inl6kATHPpHcmu6yYl0u6
tm9HUFUKGzx/aKixnGUaj1vfDh+eTbGgrkFaFsM7ojGUtaF1VJsM1XDNJxxbZ0zcwNl0oT6Bc49X
1mf4K3dQtmnO9wtCQGD/IdmfmeUbY3dzKehiyI6rcZJArGbgmFrRKsqS1bq7s0TTdbBVv4jB4OcJ
ncuiugJrlL/RfsIONmIc2Giapt8jkWRaEKwoEqnyL7Z33E7/PHe5knQwLILbw3hk3KydjdcYdLrf
SVCVM3ZQt8q+cP+HhUYWz5j7sZNF/bwa5zVcJknGy5sCQPUd0Ni+pdipKbGFUnH24xk/SHz+cbtr
j2/7PQHC4+GCrvVRizlrj2x8j5FeqjwjQVMdYXD8d5Gy6Dvd0rh+8BJDY7UwzxvRfaOnhbHE+Pa9
q+gGIMSiGbb4mlWM6VQ3B6SusQGfYu6n1J++gQcJ3lt9x80NSRQWXjbQskb204yr6Zq8KSgchVjk
Q0P0nr0piAirKkMe0gjmoZTdVbB5zj/P4lezrWlO1gM14kWTb5s4niufKSlmTdN8TzhlSFGPIrc7
l0lDKQRY62pa494N+i9g/Zp/RER86mb2aTqtSjXrt6Pgqfz2F5cYsWnttlLhBcLf34WRyy5fGANJ
z2r1zH7tw6AB16MqpBug3tDOdWcqcQASJGd64Ajv6oiKRUqucCxmLPrkLSI6YpzaDxpFQXCWGqHy
SsxoX/6XRVx6EkZ8FenV33BvmdFP67hk/c4yBc+Z1l8PKfRncaZEBKhff8e9hVmAFUXxyxl647Pk
Ps6fgZf6IFYVMV4RVJz70TDFgUyzb2P5X4YiWxveJjSvswqJdVql3kPuAkuQAPoDVj3Na6kDEMuF
w/0FimnWPA2S3uyeF+WunlR+8CPhlXj5bPh20mNM3Ee+In3hnKrldRqbSJZlgekRtTv6Y8Nz4Rr7
3ppNjIrOBiOmbwtxVem/oxvgLm1NFM/wA8mRKDIdDspUK2r2C9ntT7sBhQGHc3goNRU/ZbkrpeGs
AxIhCPyqW022/TZP79FyE929G59YYBPV2AetTQ2/GAnST9mHHsIcLZF8LQctJF7a5gZ6dVenn+1U
jmy4Zy/1Qit0t0dSeivTdtKxc0CKu/kWSTBVgFCzBdLZull3N+7h+js7+2Kn2+Fhc/K3IApTUXKc
9HA1fiRtp8BtJvfjy38WORrRRJdKRi3fMvD1cokhYbPKKOmEZklHF1EIeJlLneQpgzxS7tzqZW/N
lmWtfZszj1qB69t4PCh38uzSeZhq2Z8kELCf5TvzmC5cK9CfnhjyFAmUp6LOFzOsL3hNqzVSemBV
TqmVU4WBIW7AfTvi7PNUp2UC1UT5FBmaAT5di+hOPB2+wMaQLHzsfFgmaLoyru2Ye+cTyVzLW5bt
/tq750VTcfHFq6yJbxfFIF2ZzbXTGOHeudBqH+FcmqrzEPlLhmpQ/q01iGFCYtheMcP+T0lxwcDm
qIQ7RZZ4/wEZs/Aw0chnSxaBpee7tPupeQ7SPwoNXBcbW6K7/8qF76KwjjxjeC8C2WxI8oZP8tv6
VSR+IVvZ1Xwdcgp5BfvK8A/D/blqIe8Kn54rehsS3hvXSqDnzW8BJZDKhHzJ8X+8Dk36fqVh2J2j
VnGrZRiBxpOQkIBPKbJrHRXKYljjbiNTJczqSUXQKhqipAe5GfSSbuB26p67WzsHR/fJAGkxJPuw
o8gaA67IhZo7fbdxe02oGi9KBq9+ZjCDHDr0griuH/LjpxYac+7V8gS056hopSSL4L3V6bdpPYdO
MMWHVUQ/hQy/IwA3zNWxjhGjeQ4PU5UHLSPID/bAgDBlIq0hqKFbTKBBbpCEfdFnO9mIXCCZoh4D
i2+e02EKvtvdMVLGO0ScYyfGrGBV6zwdt1mAq+aHFPbIUPNuODfYQQH0w3QU1ZGffBtvg9xv+tHF
mI7rLwHNndPgXF3dAhBZuy90vtCJva43dW0GTsvMiAWKpEm+Nf1R8sLCrDvLFn8kKnZR7tTlrNQS
fp2nSfZYoZFQZeK9pzYelymhk84G4SRk5G4TOqOKWyys7nEEnqMFGziM8IdGGWWj8OWGAj3b9RDQ
qkfNNmzBvlrSQw1eD9JCHyZoYxbtaF1mg/gsQ71Lxa2BQr6IHq2Oq/YfTnf1yra2uOZ0bu1bVmSG
NoTc1iP/Jh+g3tzeC0fUStYQWrIFaUgi6vzKG65Gd3CbiC9zU20bZGjm6uBZf4czLzDjcVAUMN0L
Z24rmGObTude9EoFrlfO3eZEvYs/p8ELrJvuVFnNU5w3os7RXDduiTt4Lq6UYWsmTNYqq6OoHz9P
oYpSckczNlmsNhgihP0XAapuZTnKkkzGQq987sQEspzYbxpFBDkgnKipmeSEeiY9V+RHWUB3Sa/9
vj2VynFOq9q6qtwhjJSLam8kcd5YZDxg5cohzZykQI+Y1l6KU0CL06NlQxw3x58OBuAu/tXgqyD0
fsUdblET860+AqVsGVLph8VUbIDY9iOzR/yfrO2QTHoYwIfcl/zIDA9PelwKhqUj5Jpr9T3uRSll
XA4PcJDDw9MA5fhVbSIOuuDyi4oGn63fRQqpwUZ5+lDUzemNsQWobcctvd78TZNEe+RCPAILZMhv
f6pIn+C2ivGOhlIVZtneedNh/P15nRzPqbKMnceyQZP8UXNEKqOvltDPHjLom39ghTLLwBPIMG1w
OnFP1o9xjKp+Dx1JHraHDKqehfEwuHh6L79p1NcdIfJnTNti2eLHYcrMrmSprfryn1F/zL4pLqZc
ew8RHVSvlzHY7hn6yLIRwxpsppr3Z3y1J7qr7Qf6VkoFYuPLrSziDcB9tNeDn4OST+sjkhDhhnxu
TnkGSnhujUuHR+RuBElPCQ5bI4yqEJjashRQrkKZz2ImOniy4Bmc/5POHQDr19fNcM/JbvzNrSqJ
LJ2umXVJG436NT/0JwFe8nrVK2P77NNk5Vh7pNokmBRJ1Lv2xf+NTP/ZooVEH4e3MWqE+BqjRzDo
YFlCZEfN7pKal+KKPuC2+UJSHV1mkY10EpX9xDjftuEM+J/uCFWNwt7WFRx8doK9G1sA1rSfauZ8
FuzaCtaPQwTODMUGQE3qXwsxhroFSRdgN3k+cv0wQgIGO33ah3HX8InzblhzjOn+7eIMUnzm7r4I
8e7To3lik8ZfTTYwtVz7fq3icIePCxsYVKe3/yFueepQK8d6Zx3loPrIrIPGOawv3uGKFYH+5NLc
PIXXb0bWbCogPIA6pM1w/wjwlLK9xoZCAAWI1PuRC1WngX/yOAiZmZFaI8RTI2pUBwSaSs5D1e5y
jeepupuDuEjwr7mouWxzHqkiCw3nad2tTbdLx7pfLyiuOSROfEl5DogaKIsqUuf3YTyf1RSO+TIk
B/FVYknfOUyd2PsqqMf5fFx07DSCoFU3bTiZgcN722b74sOH6IVIvEx1x/nvH7hlp1gfId2GMBQ0
+0Ggul2vMzDu+kGYRXuQl3tGwF4GrdXWXZ4tUam7v6IaNQbOumA2sclNFDX9NQqT6BvOGIY2ZLuV
pJqq3loEIKlcTM1Pi0OFBclSy7axL69HhqPt0ylQtFR49A0ES7aHycQbwpBhg99GqS4tnOWPCZvb
0suudsXXDw+O/GWDS2yBxWIVxsu9BPX2pwPTL3RnXd9t5aCY90137Eeq/zX5/ZL58lUTfXp1gLIR
FzTscr+Djv+5F0XV4hCDSBPOLvSIcQ7xwgLrWha6ArTtfs9kCJYjE6dMJCJJu7FvqpozScMd+49+
kOSrPBmxgB9xoiQVeU/K+YYB9fJOQ1iQZZEAnUxkmD2XbuNJ8MGXAhUfcVMEeOLOBpnh3dv4pOZh
k5SsK8kaJTYDOIkIhfaouAebHOSS0tpAsGuuc+qhkhDhMdYiyvstJOeNML62RXqh5E6+IdIwNLj8
eGRQHlV7EgBH2mfWA/yUF/SO8nm6nGuw0fsGgjfzIifCgybgtHBUfl+wIXyA4Z/inRSFrcR2ay3F
TotRaasjCm+7HL3P6/lUzUzZfhioZvNh/Ih4LONVG6JKMKMiGQVcGYValVehVI0QNZ58VTIEa9Ko
G9MdeMHAyNi/UQxXXhLcaMiR91lePYvoG/645hKUZ4MUIMJeR3Xn1FX1m0rJo0B1qbrkPk8k/ZUO
jVEblJi4YUVQbHrAeixCZ/WqpQB8t5yIAiWJdJbjJ81YmqnCyYytdk3afrAznYSa2GSe6WhPZ+P3
7ccjxfKbFH706zI2hcnP38b/l/r7c1vgx/uJEr1seL5Jjk2FjNJ8knyrxo9ViefSXSjPD0+4uxjx
YZ9Tm75hH9QzfU/jXhS/NZ/3zjTAmnvq7cIpvmnhgUEU8timiKiQrUJqupQ1NP3mFKlLXPj8AsFd
Xesdd9JN3CazQfKLk9f3td/sec2A0L3/hhGt6GxCwYYpRLkGDcUZYWgyhoSZLcyODErIjIaeGl3w
vijQ+aFkP1G8mfigQrBmjUAOIanfWiRGtdBLHE1QLpGf3Eynsemng5iSHeBDNEYb2GZPCCjJK8kq
EBDH0RWbM72lTOOnqyGKsxhf1A42cis1VMYHyvvptJo4sea9jAb0DG3ewdEpNuctHFYqg6d40IfB
UvXvOCUz/ZyOgTdcvYf3Ihdx5QVq/yhq/w8seTzJo+wG85U8NrKy4+GxRQmyxKcbg79bAVCdRO6V
ckXwXCOhDWZ8ZIFCI/SmDMzC+2SvGf9pkaOJPDERDu2218qndQvAxxLsFKX20std6SL+cniEkrNl
neEeCgIbObg/zBXWVL/k2Dqw57/81uzZzNinjd3KjDMIbrGVzzneTjj+WqN1y5U2djUuIUXghTpp
Akte0g9oVRHecN7scT7ZChbXynvCSABBPxu2PSCmxNPFY8CPul16TIG6y0VtmiadIaL9X8zFf+k9
n4wJzN3duePIpTsp1xdauFzcLwOyRvYbzbWk3P9w/vyYalnJMOktG1y3z4wwtqGuk7WinTOMQyim
rArTq2J9f212RgcuRh7CYJN7EdAvzXHUZ5/Ht4Hc4hQO1sHJac35AmsQIt3iqzFcs0r1Kfqh74NS
8jMzYqXd16we7sPmU2j6Y/H/cdmFeN9OHtgZ9Ecq8ZVKxpwtFnSI1AvNctLKgA+qJ8AGBhTZSngm
t+TSjdvo2QmtGWhxwaQOlJ52l+hi2iSwUqdKlyYZcvJjQ0Mea+8/SDbyo337T0Eeww4Barx0Thy9
i1NcWbRmtEVZ7f3vxVi2UEw6oBV7J89bkiP9LFPfeTwBC2UxLl3DPCNCfgzF2IhZDsEapLdKzm6J
tSwVut4JfInwmhbzOfC5mmEjGaaQMPtznbsPKO040AbCh1HuBXYorL+kTMNv4UwlUcvN3gmiUMIO
gTpAyuH1cgYshZUibGKPq7n1szD87Mug9jiNA0MyNhQ/wDCUxJWG/jrK10HDPXmXTbmg3R+emLEp
CzL37aGw7PDwIS7XBZhDLV4W10r0xZD3bf4Eoc/scfrSdLzVmKgOQ++zbq49YpHjF2W7U7HhCsbM
Q6ZHiWxCu2LpBU9ON6OeITgq6/CkBOIYYhpcWprgpUAjJuTAMbZAL1hH1EXnyQk905ZRKRjQG8B+
fhxZDtB21D4FmmWatogW98PLtHmKGdP4HcjBB5vKMQW75AZX5uG7GwmXnthYlvybm5JkA9Lynvht
c48WQfCwm3cFc+l/DsAfoV7heyLt7gPD2Jn4BFrMrffDEquDUtoDqsgGnxUjmXc91IavrTTPR5k9
ZlaVI/CNtPJMeKXaar6JOT+3hNU01OVYbl04DAON7yyAJH32NKnL7PryzzU3Lslicf39TJh+fMeP
S0MMUKPJr8OsD78y3yFiWgVQJKpZof/17Qxl56xgkXhgKWg11KWhXdKl7uYHvCredC0/aW0c+6MG
NJZk/wA834pdiqO7s1Iy+VvVEbABcfZDecPEspzfkoY/g55CI6Be+kqwCc/JK10V68xhsycvNu+D
ubGUkPMCywtXy/HgIlARXFd8A9RoRuoeUpulibWMU3jcj6m5IyuNYPQsXNN5JrYcq7SajBVz0EeR
qN9gft72ekeJvsatHUehWxJgnpHV/vhamOnQ7L0m1QMKiA/Wkp1zXykCBHao2vWgZCLaD0uoDN7Y
QSrXO9W8+hvzJPrjGQ1E1XiKluJxec4xrHK8rKK3n7EAFHvvz+Ej17TICz1uBh+NvCWIcj4K4Zd8
4DTW+8I7PTL7wfUm7YHEEwBvmNkQS9dDFI4GUTzOzUPEsYwAz/HZ+WuGHon5soXo37CuPAv7rg72
JGiP87QyOR8sAlvrqX1IdMNzjgqMZ77iU9wmyHkjsd93PZoxdtju9ybmRn0cVWtNF8ij655q7Tnx
Z5eq2JmYOdmTrBlNDnnfZuoAC/4NGlmgQUuNNMVZ8XzwEEhFM6IkZhVTlrSnFUOscpa87jvdYeJU
0XIGQ/iDd5vyrVSGd0LjwLyTyJClnxpljqWJx3YR+kR1anaZzslH2CuyFY8oMUFJHzMz5LC/8bZw
VBAQuKIzhgMKsT5FWC9TS/VP3/z0WWWWkI0YFH0yH/azz57kJ9xf0w3N+K2HZtpiiU93nvgf7g9a
x9p+6Reo8Jm9h8ZP4XxoYwMfzL/PGj0UmRZL/91ivtuB5zpFJt2iSI5aZpux4SJouyRyGES1gf8+
SbYqrFBOFvzbD5cqr53Y8vSaIqaP3fMK14sgqEi72YM98sENrc2S3qAgDieWqkBl1QG41SjlH/2n
0Zz5XHwNyXYcatJY8sumCjiUkJpgZnUFN00et0bTlr4w+QqzkHknW55rH5IBftWunybdSAPItNj0
sjRXCiMnqnKKdexZq88oH0MQ4ZTBfK2VBpY3sBAVjqL0lbTc2ScNzzZ4VwILy2jL65zjC7s/iBdG
aOy9Mlx9uiKtMduDHFk9W/AcDBHVxXOlGMyKNlC8UlEoDa/QZYl+GH+ePg9W2pOTMVm8JXNnGaMV
Eem/HO7Z6vNiJ5Oldo40m9q3VNTAkwRFQT6nnpAl/QMjXEPUDumUchFXIQU4RNl2umHHZwYlQdR4
sj7044u580SK+/mV0/3lS247uQ674+kG5+POvWkmi+9u/H+OcSFRTKciCrt5TeGhwSI1RSg8kGXG
M56uOg/6iHp57SPoGkbCs2x07XejcCegLyBB2QiN136aGXtUtQFT2ie1UPgsTgZoDGZE4RZiBzVA
6Zg6Jo+37pbO1+jFQZr2gTXogP6g7h24M6kgm14ju3iBXivh/Fw0zH5MJPB40Ecz0DUUPKDZkNh5
R7E8p//DDZr7oeOpzQAwOyFxz8WkJSZWxfE++HPWQ3wuVPGOcUYWaifXotquHRsheIrZT3eTP8R+
u09s5Y+pqbSTXwJKtnwr0eOZjSuY+JqdHyqNKFAJ8Hv1Yn+TyVxEfXvYzKVtPee4FU6ePixw5GBR
IEdMBh/Ncxinj527TWskTdsLoAe/TJFCtwlGaq1DR7SLZLMk4hEpek+EqxT4uyOV4GjN+FbqLgFj
sQ25GBf6KmmDEDoUWmVT+dmEf4rjs1fMa8xCfdpGF2Pm9ZFe/BaOQTxrbVQe1SSm5pkdmXfIsJC7
rrhZ1gcgFrryuOJUKZpYvC1g6DfpUunQn6HtoYm3yj7/h3erAdsWmv90+hNTnfJk2K4dcTQb9FIN
1JEAh0Sx7kl5Ku8/XZ/Le2yZ8/+KTyTgE2KjbNs805coDWVsZ76+MVBN9xUNldyUsBvVJNtF4TtE
42G0J2/UWXFpwdwgLRgEEd0trvQAOZbTkJDTWjWrk8vvd1dSUCQltf1x+P+4zeCYkRjhJFahhRmH
ESaOaSEDHMVvpArPrX8Wf3PAuxyumf/iRU1XdrIW913GppwATngcIb2gwiSpKtXnJPeowDc5PnON
J3Uc/+fXE3Qom2TLooNfP0E3kyJrVdNg5FnSrV14FOcl+9U8gmN2A1uRZRZQQ+EaF5XmvOAIkJXV
DhMVNiqquLFzuxyrPSJAV+Aw45BSkvAZobsGMP61hGkyQGiwSoDoedPU0i1Vi1/y7PS4tx9DFalh
WCud/b9Yxv4RT2YOiwiTV2rU+j15wt9Vk+oRh7ffizBNDFrXvJXSC57m+NWjrekr9mLgruilagNp
OPbMPbcsNdv1pW3v2fXmTAW4ks01TuDAvK1ZGG5N/iULfuRiiUD0v02hzwVn+xnCDRiTt3nclFJ/
bbx0+pLMCF326/lX7yQGOG4Rx6+4OSway/J0CTWYAB5Vl8j5zeuE5lxDMXG1TWqY0wZAMIUr/Ag3
Vv2wSUsEBss9dwMzF2b1yC4iPNSQHz/nI3Bnw8m0M2fIjfVaTg9U9g7FSVFaX3UKxBCliwddT6zI
OqWHOJuh7e2AKQRaroUdJP8QgpcebDIcWA/MFjMNjSS1hdAbaX49Es3XzOft8NGn0cWMf81WSUkk
Wl9h5cbXbKCPVUMA2m7AcWiHjbiKCOn1+Jwjj1y33cAtJ/3hDm7eH6z0Gvb8J7kco8vspNODWQ/f
P2ZWVH5LbuLSzMxx6FbJqAdEnOnkQm2PgTUv8rDNxJPCZdsVD1jZl55vcMN7sPvXpH/vbDF6oE1m
dWXmZTtk8UoGTeAdQt5TZ+R/JZN1GYcEM3n1AJisG+nZ97r95dNQjCz5uqYjo8zu0rd4aT6mPj4Z
Q+RhK+33p3/7QuqJqGq/NQuw3U5yJ0gcKEwHeoER6H601UipeD4MO1TtYnLESPWuwn+c5R0/hI5v
yp7yLEL2ZRUlv30c1+LnRkbQaiOZE/uZOgRQt6OctcYX2+idXwFTpR9Yh6BaWl///COiKafRv6Y/
boJHi6a++APsEpNmZijEyoIbzGacRSu9nlnTplTm+0ZHtjM3E+xy9xNDWobaMC2loIplexRRtBAv
4QVex08w4uWRYjzxwrZOYISUdZ8+dVEwVFmASeP2IGungvMg1M2NjolzR1xNUkCpZIZ/iWapRmx4
re+ngjlGFOdy+Pm1zKBZzLfJuvcn1rRcaJX59ykE8N79tybPyXsExXcusTUZZte6fbKUXhx9LSFZ
RBmgGEboIIGTjF4TkScPYsERzrDul4DUYYMy5gUZ57X4H9dpg541b8oqdiohb+rCslG7UDQNF5B5
iu1jVbdpwEvNzzOGx/l2omdxF65lKmhlXJYddFqZHpbzxb7Om+C0kA5yaz2LRUzeIA/LRziyrMbk
/WmbimIFPgFPHlCBII8SorUI+pfEgcepUWffVRvjCyAXNXJoVLY0Xrx0QVeCX88hrVGha/t+T2y1
uDpyTMkMe+Qu4S7WXeXjNlWJFKyS0tx06kBz1E+awksTnCo9TnCKva6u3LdZoim1gsYNaKvOa8qX
hHvi03MV54cbU9AVhDocXb8f7C95BltAK4v52FN9yE0WDI9oKrVhe0nYQNXN+ijrYsUuk4mJH/wS
JnyuabHBKmIVxnWj47Atdek/6ITSMvo3gdG46CasTKHDLK7aQkdPyX6chPB0lWlLo6NLLNAjuLnQ
+a62TbDD+MlcwjKMTSsW5YmFP4TPvbr3y6FsmO7pHs9SnzHo1Dv8jUzK5ks2QIf6GL04wfin7lfZ
Ti3zO3M1CCpPbAX/oCuvKYDlfd3FF00agCz+RnXdgpP72d2Ej84BWecjqp6fR5yVfMcPyHv7KCrA
2Lsf68w/pr8lXoeiDCp1k4p6cjc6MvNTVPvWt0hxPnqHTRCJjalPC8Slo69eOboMih6dPSE3wLKq
+5QStfieLHe9abPpui96U1qAmfrrak4A5vimiVyXypWIPNkASqbJOtNN1X0556UHIH1ZbCynVP5C
2rCLoefeX3dItcCtQsCEvcEeaSpjMMFa+U7huggIgvwf9ho2qlvGHNpj72QVqa1kFiqXLSoyiebi
ZVYkoyjvqvh8zgmjv5Ww2BOYehL7dqE7S8Dgh0mso8YaEmGu+3jLCp5tYCCpF9Rva1kkt5kN5UzE
ZKVdrYZ+u987BurVZB2Jzb89J08qFmCliodoYSnJl6Mjdc1aSHy5TDGL2DUnG6dU5o6G6hfO9Iok
CFPDSqj8x1qtmPCyg6AHjX3+kF8OVLJeZOg89Q3G5JiKlSM3FKXxKwuxR2FK49sC/oYlwPd2HdoD
JCuXXpoIFTwIIQNq702mBKHi4N3Q/IUy8uab5g+ze2Al3rvOyrXoLzGjvS7h8z+rSzTSN+c95c4x
321dseVxlvLcc9xdRWYiSfnb9xlNufZdNbQxuECEUdsn7LW5BxGmaoTJh8j90csNYwQ1aTjsVhdK
4Pu8+U/oDew97GuxuJFXW/FmkBY2ddTRNq3NXch7Ijy0ZExQ2uOC9LhRJdcPABc7CbAFQznMZ8Sz
zWvnQQZVegGvh0sFif4x+rkZYf3DGy6VqC0eC7+vnKKGBjwO9AjwuQanysh9ogTuKvG7wTbeUsHM
emFZb7dODKSi4PxlECzNybr8K/XrvtCg7gyMIuxbXkVmJbpwVnKmDM+P652y8NH4HtLneK6Vijdc
6arV1FQMod/H1HBaM8H0YEgz/yBmv6X7E/X0N4ikSioMQtcljFsopuvy0xL+PeNm7w7rLW7S1Bq8
XoMZc6aZzMgyPy6Et3RiUwIQ9es12UlYwcFibD2jom2IFJ7dYNos+s6axmSkQleoZ7yf4o1nszIf
jwt1BsHsbv13sK3a0lv/9HgpbSU84FgXr6kAP8un1VjsDWPQQ+xrtbNXZ0gY9AJIzwWI+V7BQlOt
toda5t1EsIDs4YgyZlhKeowITMBZulaZrkaRj5DF/oHW+9tzoyR8lT8mGDVLA+lB1pZv4QrnYZ7R
iBTFTKDg4sNZ69TJ/1QhPZ8sEv+nKsM+l1FFrNkCKh0DIDYbwo/XDAYfSKvTOx8D30ZS/LE1ZD40
hAPaa4ehp1+kzzSRzVxDw1KWOCVGCr4vBlNQY3x8PEPGXPSbxsRBZzD2xUu70TlSpSzDzqxGJLBl
5hbnggrj2xhbQYwVm624UlFeBeoCHLGiR10f/Se7kw8lhgc9hu7Vejauw62kmsUqYGkp/0oHmDTV
Nm+50vVrFpvRDYoEzmcNr6Lt7SUIb3BPT60ySe3kysIA0BkUtXEDMclbU5IcyKLE1P1HZ7f5BWEH
6d5hjautum9aTHoMfuOCxurXBbjp5b6n0UCzhLNN1KjlMGla0G9vls4BB1nQS2LI0Br/kl0/0V/N
8YfQIXHPw1RQGI0+Tm3e+5Va+fG4i6DI+DySWgaWmD6pLsNuvRonjSL+M7OcZAcjaNSZgwYEerrw
0MUPLXOCA1Qi7Em5vVe8i6vqaBosXzHHrqIEyqTiJE6XuwKx+Mf5KjKmjYTFqSSSqoMDzXdbC3Vw
mP+kZ1P1O/Axh2nWbvEaG0kzH56p9Umry4Bz+MAFYmPqgUsFGsviB9JBqkG46BpNJKETp5QmXpZ3
kRw4EuPrc1krmHcdAbdTX+wBgx/Y9q+/wxC2d3BagVo27zNF6LXkMMLutmandBfMO1UxwP2oBTwi
RpJZb/oo9FOuRUD2CQl3hIhv3EQ+4yE9OPj29fImYhVrVyMVz1WBBZrKsXbHN9L4ND6Zx6u0nmB4
xNh7sHvlj8s9DrYvO0oqE5jkVpqdlMB4bL5aoVew04H63P3ddbhA4cptvbpCCKGpopyiQPM5NYLN
s3qbw6mQsOjphdSXI5XMPSfFQBXZfjBextg/v8HWg/AchtAgiJoVVT3IlWttPImtORYMOIuWuVyz
7QnO3CBkR5j/QTrlvxQv1sUKAjfGeYIW3J8Fs25qlLdpTPr0dwIW9KDH22X/do90RQyioMNLsB7c
5Vd5WiPUorm3tsG+3hckEqcaLtZSny0gcbDrV+qdb9KULv/k5lvuh5tc5qAAMeHhdZrxgYjsQCZQ
L2+XIosCgrLD8gt7YLgH11YcDaztuXjAidMcrfsvHVNrZLEoo0ehvxeGGQ2KTSFmc9VCXbxQbEno
hoMdQsIjwGcC/vim4+hDTnC+uKBq6uiOWeBDwiLYzI9MWoNk2VXqaaWNC78hJm9iQ+d04gI9iNIt
pZCGMelMETRvEpb+URX9wfH5XMFps5xhV7Yx2gbShizMwK1Gjd7uFivPF85t3EKZfgVii5y6mc7v
S2/BcptrPtKqGLD56b7ATjzMunU7NBUda8qRUTS8k3kT5T6PCx0ts/tOxtgiRfyaEXh3QBIU6nfX
uJgYKKROc1q054sJOjOhr6XO9KRMT+Lp/yl4egj55sjf1+el11joArkpqNz1sfD6BjzRjzUXDUM1
7GIYmJvZYSPbj4qpwm4jOzLMG5s74l7UXEta4OUOkPZsf1bbZF+H97pARndhCtNu70Gs2Hz3XTDb
Cpf9Gc3SBYPsjn5iRjk2ebZDLnBuHoE0uUVetQh9gZ3yTV95+xUkxappD+F/ZCoN9PfKTocA8Zax
fiOfyRNeL3KqI/jAl4888bNfi2a5GyeqdIYvmxRXRYPAEGFzNPB1E6Qw2T42pZ4qvQNBH23ZZWf0
ZVRZww+90dPyOmM/70XVG/UPvp5zU+ETSXJNFPC2T6gZKOdXezC9PBAB7YBSiUay1+wFoZb0J3vz
F4Y3R1jET52S6Az1je6THAMgiuJTjcs2XoFqhkhnFj70+tqsC/uPm0nmFVb4/sy1DZ5FBjIBtnrh
2bWcz278oyB8Jytg+UphkNkMuI+EL/Pxff+t6jlz+9HuG3Q/Wb1N7rifL5WUcxKWn+Qf27REcY4k
CczLFyyRlkLJvfl5y+UaiW91qaQHP1B3Hd9Kt08IETRvU3KvoczdWwjFlxav/geHCkXIyrSkU1MC
VxZKoHC4tmMNdcOLodabMWlZN5yU2EptK4oqGfH29ChCySR+F8mNHjqhO9H1uRgfH0mIYzwwAXgH
XcRA/zg2QTbHngsiHkVToUvtA5SyoR3Sea2zNHNQeEzjz187iLw5ZIqhGrL9aSJPbzP1zN7hCA94
8mEpl9suEx9VnlLo2f/G3QtT1fRlSm7KZXaeMowrX2VKZDOV3Tbl14QAlwCPfsP5900e84t5aaGe
ZPeOZEw4ubYjezYnz01renkWz8gGKDeZDGS9Ykl5/T8rq1iTrkyQF0kTQ1t9XrOpBMjNxDrJBPuL
mAwL/IldcB0qGZN0ZStHPdminWtnvP2Cy4PVPrIz7XvnQyP7DP9pktZCCDm3GtSf381anlyQO3rJ
aor8ep0Q1AQCU/hfkSIKaZ7k+gckmKBXVI3UUo9bK2pSHS1ylAYsi/D/u/v58ZZHtv73ORWbA3sE
EDkkEB2r7OyRwC8vCvrGx4vELfcG26Lavj6FoAgWMqcWuf5sjslvlLCkt6zjaMxEe0Bv/I0oXYsA
9v1/VdcbY1fKMv/LYp4E02LxPCWVjMv1JqLF8uXEUu4s/6UntpucMqwUs/QRId/aoyzbEqbwd8jG
oM+ug0/UksTGOZLG9Q0OHffLz54ufcyS7aB786Swh9WIZHWExLuvZSeHlLWqV/KS9t4VKkT+7NaQ
sDv6qlnIPglcGiBhdFB8HBVNJVTXe3yIyy1KPb5jaiB5xqQPouZpvKnT3b9syHF3qEBRUvFctS6q
N1mwXXW7UQUsmy/qVnczPXr2iS/Skjv9F73VCdeCCYhk+TSY0KlyKsGdLLdQ6vHbdyPUmvQ8Y2/i
W5zij8s1luDO66zDkymhxVM8ktHZ11QZeK41gkIaY20V+0Bg91GfgAHR471CkxSy/nAjYltiZABz
yinRkcb8P+FYk6sqmZN9oQf6tjybJDrf+mSVFoSVr8l4Q0eLAqymXyYHJdTCraRQdPnfTcK1oHkv
oFWreq7e8dzfezTv36jh0n5++zxOJKCH442x57ZZcqqNRlRPL7MKWSc9jOpG52WcbgiuDArs61fB
sLvhnCbc6s+EkJ0a2+h3JyIdy3KNJo70hHbHnwGv/v1drCbL2kN1QYBccjq/ZduAHW4tsYaqMaGF
XUBY3yCm9p+9j3ONzsEGhgQyIKHGSXLbYpitEvhYYwFk1Y/NfIvlZ82Dhe6r9wG1+29xZPA0nnDY
qCCsDeTmENdvRz1ONRapcJfb6NBJKVmttNSNij70SjD2Z2eEQSNiOSfC0sZY23zM9AgMFCqH4rzq
4BWt9yYkxE+Wha2B1wQRCWgh7YT8RY6N2nSBH92vJNSQBIAmYCfPLBXpR6wiJPUVbCjfd0XcJOTf
oiE1TJencrx2xOX6xdumUEmRdHeKsT7L0gCnOpIlwf1OMABzS6iKxpx1lGREYI2Ir3Qrk29dMi2D
CknQ/jRZB6RHEjUZDiiVgeq2LkVSc3bCM2+P4xSPC8SKUWckDwg+39KbLBJh0pQZ3x8IE94wxQ7w
tntR5orPTqF9eygHvvobGDxUroN+/Pw5uLZdP7OUxuN+bdTQsLEr9FMrE1B48HjKyWWryOPhEmL0
uoClHqFKO+vrr7Aq3EWL1tiwz0RaaX90q9+gK5+Ev5Hqy8AHZxKC0VUERuo3idFzqwcD8+YiC8cz
U6Ft1BsR8YTD/lNVlrac0S0d5heErS69zOnYYUiuwA9hMFlbslsZTacBVsDXD0CQDmlTVhuZZM3R
AcGDQr9c2oIIc1iJYLh9c8FOz38hr1DxwiG7KhRxdutSkCiu0NWpI6fTOKk2sF+Fu4Zt+YYx9/+a
PA4n2Q9tu+PJAKUxBLttJVKF1CiJYtI6Ud++WEMKCiupK4TCsQFPkTh18t42R1m4hUycJnm3+kW1
2NSA4mO49PRZ5ao8K9wRcYmjk/7E+bbzMfLZg47u+xKJbt39Y4x2delIWELHuGR0ja9yibkDVngS
DoNoVJxvDBX03uPYXkyqvaUJzcNAvS+gWp0gderHpsNGu5g+vx4uY1UGcVTWhEPviYabAiFJTObP
5mMsNRDYnZQZIOF8DfIKlM7Fsq0i9nNMfZVqcXHub1JUi3hu4GHH/8cjZCEsyckVyqk7hijNl5pf
OwewDlusqb/Z9DIgz3f00sFR/O84EgW5FTNqR+MT/ZYdPWCnXSax7G6qbdRW4gzJe92NHGcjtsxg
rqxzwtbIZ6nAyqyPA5TviGzDnrWmvg0fJJePNaoNFGZ7x0X+GV1J+3GhLUf13cmMqFVuQblLVsif
P0Vn0b50iN0Y8IcT4z/JrFH1Lzf2DUARUhnsrgtJipPgRr7iVTPqWVhfyP23t9mce47C3G5N2t80
hPj02qj790YRxpufOZv/RLOcSSPvsmR6zmE0lsIKNfBVznzBLLJ/k3DLpOeNuTJLY8RzprxPqTS8
u30pGB9B1Xd4nQfem6ZxUvuJFIgicHiVNgeIx/ef3v9bRKUvw5NobGEGtjgfOwNXPl1nVo17gQAz
9f37DIX/N71x2sEGLLcEWgmutB6OFr5Bf6otfb0p2DQZ3W5nJ1PGXeV1fcscnls5hhGoqx7+Vcu/
eQ+8ZdbkOo/j4hjv9C9yCNwhT95IuyrLXlZB0ELTIqNmiFPCAnBSTfLbBZ2XB7WmwOmVuHyR1Ztq
JWNHtszJ9mCDmzDZ8W9qbUiSsggqPAAwVhD3vulLExqJ8KcK0faGjtrsn/jao1KrgB70TbtksW1d
A4viV/q9FCp8TeQqLybV+OFTxH7ekhvxXtfJ0jfG6bi4n226JZRcuaX0etixB/hrwmVgtVp+dz/n
N2pvRdaepnR+Ddn04WGlK+5tw8tDcsuqlCpv3ZCqFbzr9m0MHi+X70NfQqlTSt8prrBWaFyOE+23
b3jwaNGnNcmW5fRk06fcMe0RmV8sAoBa2KFoU5fymtpZw9UpZi06K07i7A1TADgQJ38lBX+Ynxxr
ce/h8ciHs3Rr0uFB4zoYbwsnHBJ2jLYIplFfmKI5vVTBJLog+SG8dnFrwR6uB+7nrihIxQrdq1oZ
5cL3vKi6yIyK01l9x28gWAfFvqZPZMHqBj5sfA68tOhpzniNz8g41U+sizP5Nd/qwXtAwDhhIsEf
VbB1GT+Gs91FcyaTN8fJO3DqFWFxXU7tB15u2mgljZeGq2CVU/apyovX/zdiJXpUL5Pir22ZVcJX
6bHOEk1ScfFUhnK849hubHI/6KrVK5P53Z7QEJleTbHRog1nzXa2/4PIWteCJMbRyUiOw3tpugHq
Y6fwhVOwIDajjmcurVSCM+3a6kg6tcauBPc4Y8I8G66oZd5oV8aAaQ0MmjwfmuzNXPrO6aU3UO0E
wR5sZ0xGfR/oaFgT6v2TM6lR67ilu+xF7vYZelcIkFnPHdWMiqQEa+sP1bphVkGL+JoSchjg9Aiy
Eop7vX1z3cie0R5HYQennH4A9BovMf5sJp6qiL+Vgfq/D+8lT1qkQL4T3bol+Rmx4uokRHlzG4nl
afheS6ZhxV8FW2TjJSDiBzJ3kzr8+MmoskZzDCO6SDTPKE7nV8y7jI+pCZ7Oc0nBYNqSC/vMgb8C
mo8jxOhpFNOYaEjanXrHf3RF0fKigSFD1N4LtqNhrdz+H+PToQc/V96Z0Aq1qUyGjoamMLxrNZLM
tjryvkPSTKGYTbhlzxBfxKbfKp/Ighj8zfRWgxPhBUGQenDjDW9UJCYje7/2W/dzETxdtAJy2r2R
fp6V2V5V4eli5Oxq7Pb/NXuTASYv0VezK2TiodnMzfZ0omxPZIb49T25FgBcxo1aToxnUG5a1bPz
H5o6l+qIrZeJPYxvhxOgL8egpei6/NiP7Gc6ep906mMxEm72k1Hibav7GUCjFE/y2ENr330GVdo9
nzqK1DytOdhdip/ilbabL3cd0Ol0L8RSHaScS7SS+0O0h1NcPGkDNjpqSq+OS0HgJrzFCz+LrdT/
C1r817+89rKgm1QfQeUYyGAI1VSSlh5Ep4Uz8c5efgFW65F2zOOunXP2rQRS/q2FW5K4fzmZ5o26
GSVhMzLXVeShK2JXFpRG42HaHRq9vsH7FqlbpkEINmZvVEnLe2mjd+8bCJhzaLuUkEF38eO+mqx5
Tehd3W0O8ESiZh7IzSQYIqHj+qyoqKUfuNv71T80JDGUBEgcWXdGcAu7cLPFM9wul255tI2pOhol
6dViwaAdDo3ro3XrxscIZN7LU88g1Uc7zxIB7lx8CsKmgI/+y3VbPKi7P+apZBDnSgcGa24ttPhH
X7p9SPDAcIkizdnOa+z3FjfyV5oW700C6+MTQHGvvqnCyio4hpvl6wbvV4DcX9AVj6IaViXNg7ss
yfYR3F7fqAmvrrhHQXjsJt8rPcetuQ1rY5jdqzOtf3dZMklaQH0NskzORRRoqWYrycL4o4+aSrSp
VbkN9zOShtvdD4sesoxv8dO1Jk80KGmesyoeM0t4mc+dhj1hP7rEsHIjRX2k3WZWagzUb9erkd8y
sbOEOGK3RADeI7kzJ7ojQjHp/Wx4T4dAhTggqa0nGArVO5LNc3ATSWQP0An/AeLxcn6U1Nj7Hbwp
nZYnxF4hYmYPb4864hdQd8h9fK2PIUj69ueixx8smWXSIIo3F03+e1rE9sCxwqUNHZ98EyVQCFcx
STMNYqFGBEutjK8mzE0KOgb+jQLyzKlC9oIukimm6cP3dXRsQ32MUAd7+55BvukWEwnu0zEZHOTD
8UjYf+GTN4Y7cOTsn9rrt7ylVO6AuaqAfctNc82jPPCQu5n1JjqPqG2lfhX2SVXlcz5rMyQMx0GM
GIA0EmElwzcZe5PDHxLEf7gnfie9ZRiH8pD2GNX77WiX+KZHDpX39+BPLklgy/knk8IrvwXmMQn2
TzqVY3XgEduNw9Gq87QIb3KwXsi1vFJ8V1yPlLuaMAdhAOp9zZx68Oz+aLV77TWuRqI9bxqiv4tX
kcWQH4X7Cn8xN5R/Ku1C0siDYTIhfH0SkJQiiiY3lLEY6tPVt5uOK7wuuGlP5rLnfSMskg1u6Z7b
6JirNfTEp1OvCRERR7jdQ/q0Tri98MgaDfzxe99vfIz4UmNInUqnQTxcHmdeyHiBYagfvRW9nhbo
St6lluEvRdmso5Ir1vfMa6m0Nk8Iw6pRgG7rODTfOSeg/qWoser5sNaO3d9nncbbuleV6gcXqPLr
+ewW7AcWrHSFlvlttzo1GmtMnmJaS6hqOgwvw+3fyJTT9wGHhM593aiF7mGRlH/UcAifLUPRFcnW
4mW7LDQdQimHR88N2A7CEgrVR92sBhqmXpAsEuxh0oa2/ghMZCrAWtUVq/sg+C1dmAgxxXDC5cg6
2clHonL+DbBNZNBFhylAHgUvvuWQ4giuOdp6lsGWfkE4AlQCBjPdfdFYyBW+uO/GfgIjDsx515bd
z26Ys7QR6F4uQIXtO6GNKqS5kzH5i1lyvOJjrw4oZJJu2uT9bXQoXs5oCdc/yOVxMhwuwdBlvhg+
p6qbOXc+3HYSfDx4DkNZoukS93wQ6I/NIfQhoxgwvrOUSlkZPcHtokJ7vZFt5N3g0BeMM0sJRePY
4GNPlLdBq7VeisBSkSQCHl7sAvumI9brwGK19lHBQamjJu6B2VoY4S6G2jKD00l/LvAp6MELbw1K
GfUUGBMUCy5g+VxfzLD/yYAn24vjjiz1WUI+l4OSByhNigRoifhNQXXLankXItM+4EUKnvVz7/0s
82l6yRhhxYxzhSnc5PZVGw7HSfWZ+Z4KgnPYYtgtwVSS2kByQCjYiLKfzrdOsBKtbvnhf2B+geDh
RmjW5io/ppL2y3FPxz+zxpumxIWlBJ2OyW2m7ceSUyo33U8zwTQVDpf3QVCvyEs6P8FYsl/W9GWW
1WWzX3EeinAYv9rWartEF2w4+gqTw6zlsFkqMeBcoBOh6bFfKjR+XbqJLp4zYw0aJRc6YlpW/F3Z
fr0mZ7FxQa88sri1N5024KUxBdlk2cYq5rLHWwNIdjmUiZq1XjZxLAZl1mqHwPbd6LZswTUuB38y
0gzpsA5IuzatAjF3ugCLpzfrwEvZawIf/QP2Pj+tfcf+fLRzfXHfdIlOmhb1y6MRE4qyVXr9/jpu
YZej2cwsnd2i0lRAsQnvwsYiWFbKE2tZ8Z/iMbQX+ulPJ7eGWDUzqRRihl0c0FZd3NbWb5DwJWZm
y7g9lZMvWKDTp+X2gtiXGSVhTCrResz/+RG42VrQ9I2AXAmJBOXbEGGkxJ3/oPA+b9HIpf/RTDSK
Pscg7a4jq+TwPJHOi3X5SMIWrBF7dd04COaf22wN0qPXuO21uevhSF+047lRFKLqbah3OtQDm1g3
ygU29oPPIv3SK+fMNvpB6uVVcet7wbR3QEjSyy0e8C4DQfN+YsbLerScMIOUKOqFYUqjFE1Wz3zk
AZktKpHa51t80xoEGAgOm+Lr61nya9xkEUBc1XjFsgIi1Ng0HmMY/n1+0j60uEYRkLfPZcmrax5t
Bq7EfN1samO91qnwZmaCW38XAz2A1cZtecJin/6XFPSFxYn1udkT+cegkb4eJc6gilklMT5faiR+
STR+yS+qvWwV3ze7WZ3CAD6SfvDfKD3A6PwGWxS56hCwnk+J/U/vD17Knm0fstnqsBiH+1B8eA08
GbKllVoRmKjG0nsByMFl+xYTwnvjEgLVJo5zY+CnnPuf/40ivnJXbW9c4hbhycEfYsMgYaPBKScS
BUtQS4a+CyVOeSFLqMCMsIrM1jJYNKGcgsNF9FBK6VHchtLR6+8foSRQ9sOpErDNIULLemYzNHSY
qhPbv3CgNXts2yckJjiQu67oUD4qQzlBgLuQVCiDf8VR1qoGdV1m3ucD4EUu22eyXb4zn1oHyT6K
yIiwdzyjQuBewQfHwP7aaZqOyfrq3H5EFw1ShLJTEhMzJ1uzv2abrQ+NlrVwokJryWh4hKB446bT
29LtQ+1BU1/UaafONg6RoMJeGRQuQNcVU7cuyR5F155CXcTmalweYPuB1i7zEy1CSL5ac08o7lAn
ISLgeqOkMzlophlZ4p+o5vUHyUWkGamjtVInBx7fZExBMBw0MwwZZ0ypJnB5rfpJ2sqHWS2YoJUs
0KUy8vQTOaL7tSkyNwEyXyNaeryemRPEHI9N5H4k2oaffbJS9G6YX/sYT/lA9QZiPgsRAmPo+U9W
+YmpfjQ9pLqsvoyUnuiDg4A4lrs+1eJpmIFJgT0VSz4bAbuX/A4e+QFp9jycUOsiwGZZst2DL2po
wRA0FQ0Gw30XlHQIrALFhho6vaxtJbuqjU9ZsMnGodxacZW2sRFpZ6rMhwYTXdYpSMfihLGHAvpF
xemNCOBBddozL+7rCvG7YJUzeuO9ho5mHTiw8apJDoXkMCiHkX8IH8UPOOcXMjQ5bwhXxNRkC6Ha
7s3FrvqQBYV21achhCK7fe6OFxEsZrPFkqxj8DLtSsnUHPJQvQi84KMCFz4EcTFrmb4UX/DO2aE8
mDBIjX/uBvPAjf6X/N/eyFX+/TVJj0xq9dfLDb4edlUCY/0QWlaI0LEgMLy2f0SPeOQ5PxAvofsK
oeg256R5RDcuOswY/e/m66fNtMh0zSur1tNGUiNyh5UVPnNUbxOrOwGEHV4x4YWSRa+6Xsyu+pU+
0+4+BOZvbnsd1S0NYwVAaNcUSvNrxzUj86oxX/jx07FQHToxF5bUOVQrOE5QUOqXB7WcD80CUYou
OcC4Y1y3j4PR+o1jT4Ohowhc97Qgp7dEwDmoT7UNWT8iSUZ7YRmwZjZrM8450k0yqV/hNXOrwGK+
zP0GH74vRu0VTDg/fcq+isiATMka64ifmTkfB380khWSf+G/LZcSrdp1dtX6tXaH2Baz92UAGWY1
HjREZLKLUaHN0umtMtpRF7I1/421fOzTy5vyNNkCSdGzpIhu2IYgNjU2Xda7wDU8Uc+2OyndSKs8
6TCd+OEAyHChGdG1a+JrcaAGqZ5sLSZsO+bGi+xTvnO0P4MdYJQiU4A1YxF5HHSSOTXL5eYKM9GZ
FoJP4IseUhsteGZWpMJxsv/1OZq87a2b8Bv4FJjNz4c0RvhKJBhXAiwrMyNk6qbBzmQSO5b8EzXK
XsVGXRIUsur/xUS2uF9F9NTHEkTkpvnouvzgCN0QJoL5Nlf1KXrGOX8HSDJrxMGzRoWq/VLQKE1n
qoYDw1TN8y56xHujvLVYrm7Xov4hDgNRph6b4KpFVRK1ZXpQJskGCVxXqF7d0t8x2+U7MpyqByFU
Bc/mslzMAhKAIaWdVTOEXn8gkqgaCVSyOIadmgOb0VwICWkCFTgtm2AcqKzcQOJNXDADktjRk/cS
jc1nuJ3HbbxwvUwwFj9crbpr1JJHtAKFuWMuSQKZ8d2GTZ4MIjKDYhiYh5H51nxsD4mWjqeEOeBQ
ubZfR4T5LBCVK5gWohog2YvhPFYrcRo6Ihq1sLNaRzKXyotLehH1fn1LjRl8jCOhXwTqRPsK1kdR
l7l1MLNRZWIKog40V9oVjHN7nkdEd0IIKfXgtdzv8n/Za4/rXXo/b8WNfvww6k/gptssrBz0jyWR
ZERgI8J0eBZCrQ30qI4BcpxOQW7ReJ7V67b1grBREimyZLrctlzMM+yum65uoN6I3jgDwemedTp1
3FhytW6fLjL/JHBP8Juf4HbuchC81hJeQvYVfQ9EeCL+/J++11Jwu6WkmeTAVyNmhWY9lAC9EYdy
+xg3dNG+no0HzLBr3tCQ+n3ZFGgIdM8ECz2libKgwa2liXYgZa4+22SWspfuj33ljR2zK7i7itM8
UkHXFhK2eywinmsrG95UUeQ1eZAtQPImNiD7MyLpP7DxO5fXfMVPzqdqqthV4hfUroyhEFEk5rfS
eFNQ6sR19MO+t1REypmK1czdkY4x87+m/lUC8eyvPC19mywgQeSEmFSVVb3RRzb4H8EXLJCJgCf6
VnkkFHV33sOZyt31vJAjjl1vIesoM8srfOz+xPjiQ2pBjpbqdQmTsBWHq0wKFtf/ESKTTy1QWDKt
od79rRinvfQC0Jtd1I+uMLPvbTp7wWp7IV0K7fSuyegFONy4duGAdZn1P/rjV6JH/KAu439iwbUm
G0Qs+CaqAkB/+pGjBkLkpzBXupQCpspuEZklzBzzcTMUvzJLup4yuIfBU0qiPMa7lXqGhaPi3iWb
5O3CtvrZohg17DZqudCVfqKdRyITAQz3priBQ390U7DqN4SRuAXTxjX6OyWxl7DNNGUnT+vbHNRw
2a2uTxzXW2trHdF0I1S1fuSULAyb10F85OJrm3UAthQ1RaOSAcB/Tdv0QPo44VyR/AFFBuemI7PP
BdOQaXQHQvDkckTJuAnTtefzXteHOCRoCtWCZKBIoRfFuYMJiyYtu/G86oEPoP66B5OtQ70GsQAp
bNQhXCAxMNH6oIMIsuZ6kk9b1srLJ90z4ZiSb8+D3jKtTYpB82d/27PwSujwPDzFAE+9vQp9dnjL
tBuKpW+QMquJl4AewD3kzPzaagKJA+A/Qvl8UPjPE7kMcOE8j9GvZ+CbGPEdKXLM29Tt9IcQikkp
84QtJHgz2PPtSzFIDee5iDePADBDm0pfPnCn1faqS2QGG/NwfA5se4C+KXLZN9tEIchnvPWlGqZZ
chBaqwjpt+rdRk9lMPESCdqL4oJFk8eDyAwIic0364Qqe7/b8shhbg2RdU1CW2Emhi5QZxJOfsfA
6h37PS0F8h/l1eREzTL+Tq0XPMmf6dyULiyX7bbG2D3oa8bUBLTB+c8PAMWfWOaCwA5+mmNWouKP
nwzj7PJ8Kt5PCw9ASGZWOlYICoNf21qbqocqj8SIte6TbYTokigJeNYwJZBy+i72M2yxUqkphvX/
fo/O9i1UumNz22RuDElFiM1Vvra3cjmnYZbxH00WDRggj3fn7CQW8D7ER6FeoF5udZ+JHRCvPNSL
NgXLR2/ASr3vIRYWALEdq/u+iZdJc4dHqQUp99CBXtVQCNIpxeZoP54FySTE8SM10ehrMuE2xZDv
JY/v5htXM/nNKXjLCrVA+d1CnjqB64KqR26tVzeJMmc2zmYYl/IbToLEd4XdZLcgRKDCNj97UC1s
87CEnxbSloJF2SBarYOI0+yLeNN5wJ+itljPh/C29U6UCVndtCsE85G+il0IZ2SzRZ+U22zL/NEv
kf/rDuIM97p/Pk+c9zAY+BuoUE38Ma7haZ4r+8WmCldPg0ADbV20GJpVkbWVAlX0xXl1pwcqvozx
TcFVFCu4tu+N6AdDXZZlw2k+Y7k2ZNND2qYn5q1EdVraXsUOei7TWk+QxBDEiWeYlQZu+6WQStyE
XjczDHKkO97xoAip8D4pzHIZStsyJDhcQCaaxi+h+tqlPo2kW7aK2jzkVYLDzJ6vZjmatgLjucYR
linnbOSj9BbPT9jgDPRpnvoh4gsg3PQ/4qEPLk5FZA3VYZrwnHIVgJUQ12AH/gmM8kgtNe1t40uM
Gn3QxnNntFroSvgQ+EG/xSuYItKSDxqjDpVRs1liCrOjhr/3vNtt9BIuHFPvr3O12H4wWLe3aSE0
/Mz/2DZ29XsUiW7dmiqNf42+5tSb8ERC6S2VSl1wl4/CvulVSpSzSWJWng6bG3YlZ1lF4cPvgm26
P6sPiPpaMkpg9onTy8CrESUn9UK/MulcU/dBxsaVt0bDtFOIzgOqwEaBon+ScubR2oYV4+3iUSPd
fxo9D2PeEZ+Fz09r9YlNZkoGcvGjsc8mUbWycmKJQlbdQymrdUGKSiKXN6qn/QDfQ1yAyW14EL1e
hNrKJwxTQGBZDnzS69b/K4c+00QQI7OXeeWJeNHsyk7ZupKl2LdEpc4KRbFBZYgJzt7Bhad3+A+N
Fd0UXEgkZO585FyrRFVfx61Cpp0OvsXVloUw1egcwXkze13vpC3YILBHB1X8+Cenb9ZA31T6rMu4
C1d9KHdbvlcYGYFjWx9QsgHZwlmXBmy6CN/W+Ni/yuNg/W7KCXs1CJHoXjl3l+8mAaPjKL+P891G
HIE8ZW1iwxl3cownu2q+aO+L1LlRsMwnsjDPQnqwqnZsrTIX/OzhfLIBg81wUalGLliaXfo13gUQ
DMNNS7mwwQdMvXnQLzO6n6GXKfEB0mczqfp3Scfmp0HQwlSm/91q315DFsVGUH7pSHosTLTBvaGk
WW6lExmDIQCogrbvc9097y1BAOmvBiVVhjBhcwSfLXSQ9ocq+OQgzERd6w15zY3Pdoz9GdUkszjQ
bAy8lCqLoyOFBw2EJy3KQquT0KqRC64mcohqb2zFKDrb/5pvgwt/+sBQYQbAaIX1BF3BUCYB//0b
6oml+XfBy/Izryx8mITM9osN7Q7pVJpfZq/8Yj2CRO+qreml+aXdk4auAWd0qxfMosbibzhn/XUN
eA/rENLYrRv3KiNGuKxSHWltBK/9OZzIg649kDXR+v7e/JI71SJqhmVHVt+JIFXYU4tXDdIUXb0X
AG07ZfXz1u26hXU/gUFgx0UTKB+PkCxK7FP6qCV38Eh/q43EaX+2Jwl9zj8t6ZTbr+gC2Hl8OHbY
Dhzw70MwQVynPgGbixBBA8yUrCBXFy2xJdGpj4GRHLxUqEfqjKAiTMyI/j6yPN1k+zSEAZcqK51y
DRdHUmo/Pytlqcxt/j1FwHpqlJ0ckcZ/cowNcp80ST30hi0Vvk9Oq3bC/MbUa1d562NdP2v+oghZ
6DLpjX4eFHgZ0CmaZ8teRF2XESU3noUVom9eGGJlxKgbNDgKJgjUNFkQ7wPZDZwClt3sgyWtzbRH
AUpJHn6CRSNNdgrBlzMR9BCJXEzCxhUUEUJf76qtzlC0QXtC6EcRWpOVeO72sazlg6cdyJlIFtu5
HL3S7qtbd3OKkzoXncgbyEvk3Vzp/jzCl3a+HP0QzxU7E0SCAg/4x8+AeoEyvd7lj892+cdRxZTT
lgNX2oZmEmVsa+f3C7h2Z59J4y6ht6sEAsIaiQj+35wk7xHzA8mrcEquuRU+TX1PoTNwfYFtiDnx
vGRwAajpqPD5ZStHKVnhfakm87ww+eUQ52oXcXmTZgJP4GiNmWStoEEvfmdqfSsQCOYmt9jBDYF8
2GFmFKy1PJKNyF1TF6MGfrrsQq8/Q1BORAZBT+/eriNs357dhojNYD1itfDEvyfTQxbqxyy+ocM7
0MYbB3cIGx8VAx+uYSivTYDiOgDcKv4LLWxhkIzmf6V8litgKAgeAIzwO7O0W4zANpWKSHxLy5G+
PJkSQpe6Yuoxj+OFIyEAViX/aJY/2MT4O+daXKQA09/xqOHbd0KAJWSyHHyumN4zotSVs9l+pAFF
9ntiwrVWAIEfc7/6HZjicVZ0vVNTTEko0jZHzOgwGa2+eXz7k7KRGaEGDHC3HjaHWbXnNzNNlmOw
e+3f7LcBN6QI/l084Q4deiGTbSkzFfDe+hHyEntfc0XRG4W8MgKU1cLPNp+M+74s57VGdxLPlf+Z
8jSj9Uq1a9xu5hCEtQeSP+828CUHw4K/erInLO5OFSDCVl6Kb+bUyXU6tZeX7kLyOMN+3cS+LXjP
BY9e9R8AFi0GEiyNykXjSMOEmmko+d27nNQXTBAEnnFXJ6znHutqr8fKHHa6d7HykPvNgpw30k6S
LMtYPsAiHb551FtK4nAkE4lWAiPN0F+5MOXZAeacxhH2HLeANDIDSmPUn9nthDpF6SIVLHvlmvok
HV4PZfUQEBTkofqpD+m2kXww1unZAnv1ZFMS6TK49wKbpsGHlcEOznHfm145IrbjNdgpEcFzGagg
gv1/u66LeYFahu88ZSywXBM++5R0SKab1adShr0NirXLljEelBtvgW2Ox2YM2Z9+KO2dwMSv9h6Y
ZNovgaCsgCO3XXaR+yf2aePZk2lWduwTLwtAg5TalSKjlx5HcnwNfHh4qNpF5yUxqVTSNLgmPZEj
P+upNIOIxWvcjfc0iroEaxLVWI5Mx5sUl/fM63u/jXI+ntMczJQtdS1N8iwAQ0yjtRhmBP3cfcLC
hvFIw1F80qcbb1pBF9TP6H0Uv8h66hxRkDnf/nc3UPUER9o65jR1WfqDEvNCkzVQnLuUwTxP7vfV
2TH6LxutF3YsP+O3vSy1Q8durmmo1Eqmx1IYUlIZVF/EGV4vumk+BU2Za197SNRSlYY/S8I1qew0
c5BNjPcs/dxz4TB1X0hvHV6fN83fi7kT+xxlEjSWb0uXSl0Jcu2p/HLNfZcvghZzi0vmZfCgKzlD
InbevRV7tIZRQS3Gv/oVm+zN/XYGejM9lAsJ5OGqne+GbCNbQ4cSdy0fvblsMCcQ61/TvC26yglB
Gp45AhHDBOB+qeqAiyM0qhtRhltNUOXSJRsrgxytDaAy9yvAi8vkZqYQO8SvvEwB8dDRCWtEu8zm
BrTenssLmtsaZMqd1IJBWR4PDpOI2jFm6uREA85NdcqinUmEcLEmi0hNNqdfF2h5W9+efGiMuLQn
xVrlqnRd+hsX/WwU+qNjtKSXLuXG1WV7JTmrLSlC7W4LbBFrJTOyDHh+GBcyE9aCHDovpQbEq2qY
gXv25gyaKQPY/YNp7m+rFOKPr3Eb/qvP8NNFfkyvFqn5DWRu0RWKP8xm/Hr8zAJ8696McFeL3yMr
bz8ZXaL9bkyXoKjgiThIwQsQGuOZYxH2Q6cBba2PBaXU0B/i/T3iXq4YJYHLugk09x8o0bzcOFM/
ZMxBt4ZiZqRH+ei1nCxauRxcH/0x32eFnKbjhMs0U3G4MkZGpmUCb55aqL5WW7D4wdyhJpAl4k1I
Exyc4jqu+/ZRLT7it7YyoHHzFeNT/+iY30ruJARW8ggqkaJ6+LrfpLF/8IxqvdOyxwOD6NT17rRW
gqRe2Xmv7DZQwG3E4G+SK/69CV7oi8Sso2Q2PKNfnQSNJ5FpgwxgwBBTr9gWMOz8hvn2CtwA8URv
ybiG31LysN4CW3s6silTCcPk4FaD9GCn/RKKR6COu1I38IMhWACkz5XdwgTkSE4oL7mD3QCqbA3q
6Oxf+pzk9Y7lpwkBIxSLrnllepbDO2EcWd48quibfC+cYYqzXLW3qsieWGdMUnf9SW9mI8u4NYEa
48fjYoUhxny5/0IfNGO4EiGOtyIw/N0qLbTMxQA/5+v3XB5nrQqLlseBd5jNfHKfkFazEePNB2aD
goJAm6/t+F0Z8EXvmy9lDR/CPZrq3ql7PISzQV9Mg9CtBprO2ssFLIrZnqbM8/OeG+fim/jKjgZ2
HMiOF6B+MhgGKH8+OStYGPBPxsqJWHTuCPsts60K8WgDh+KkQUYcg518/geDdGOY7H5LQcmZ0mVr
eGUwWjyM+7CUy2Dov3/JED6gH/zKdQY3FiFDOYFPrvi3Vqm6ff74pjhaLZ6qMV0aMDvPJJic9fsr
YXS02YAWUOZ/Y8Bf+X4EekcEkX4nGsZAs1O4VviKQ20FVnoC1IoZLqPf4EIdUlVK6fh/hCf5dMG3
zOOk3tZZU6qeJMbbUOHKDWl6nLnNs9fM1Z+VR/2UCQoQ2SIsV6+rzgejuT27I+3GVjLW18mGL/Px
pjtytwMFtAMKCloZzjbQZrnlNDI0Ra+aebUS4c4EBy9I2vySzvCtR1/efwhzHnAu05ILsYJbMyEL
XbSSLX2Bi87Ffi+sSZFgLaWc22kFT91MwObin4DfGsRzfC5mZ2OZ7iGIZCyRObKVeGByvU3FKomB
9dmziGxv1ODGETIClusbTE0crYEpdd1Lc2fTHumNV+C4mGxT+eaRBCAAk0mmgV3fZdNvpm8lKpyQ
EfdksqT5n44t1V/0KS0vxp/Tg5o6PRGARYEpWqKoNJ9BIsP0HNvSyVoi6yNfWkUlgMGMW/S7AVzw
YpUMmbcm/anu0d9Y8z/CGYRkQB8QF98BLKQT/RAD6GyD2KDiyGirwRK/PT3e+yxRVRju8Ts3TSWP
sTJ9Q8hOYz2Q6kfI1mTJA7pbCC8Jj3rSp97V8iLKONU9lkVWxWIXxtjIX4UwMs2Ujx3lcc0ahfKT
4c/dYBXYj/H0iLWzDw6jz51U+7iFA1Hfqo08G+yNm6oKgl20oDzn+H0uQz0MXvtXRf3YckWFGPt+
JsbPI90xf04LcroweE9Jv5j2tTx5DRqiu2uao69CeUfPhSEEqsOcfcEhHDj1/zEr5vmytcOkMa+y
ARl68wHhZIm15gtm9mHuTRicImgWyUkFhCncJiBt47MNrWCAUc3eA1gK9k0lz9LZFoAV607RGzvT
vu4UG/t5H9huAghtrfjkMKU7gvp+NRlafspNFnklHm5xgS4jCBACrufQ2PFlywrkZYVR2DLnWu4O
FJ2eAk+L5EN2VjSHv84kWCPFCwmj7kZs1sTkjKl/B3WEl72dSSDRwOYWH4Ra43s71e0rxNq7GHzi
tJ9ZsVXwPkBuQRnasZcVKXVLWaMLpsAtWJILIY7CoZGU/yWANhlf1XsgSF/N5lYbvXANg2I+2xn3
MCqFGt+EbhZlsIPs+FXZI1SwYzoSVy8rqE1Mr17Epacmt3zMy8w6YPwv/VUzBKwI0BnNVMTxzAxu
NzA+PheyxwFT9Mllje9Ws1H8XqKB0xtYZBRK1HT8+7EOsYm74EJMi9LkuKqOsy5APMqviV3Fpr5P
0fnXMTZdmAMV9UxvgrVCaRyXkU1L8cgvU7BkA40G9+s7hHHfl+dvdMzHTtoNkFZ9hPiqF7wDVSL0
yLXZkm9Z9Osa0h7qIqWv1F/N/JMLyen2WnkjQaTNz61bWhwOVGn+e6ixuSL8UVDanP2oLce7VzO5
1tow4QWLq0yZeDd9E4P3e75bBdxccsJfYFX2CfyzAFDvCntZ6bph3/NT4uCBWWR+nru5yOFARoZf
WalZbX4/za6VrAv8WYorex+yGtdT7rlpfMWmBlH0Y9u8TpTX0H90jVr2L4mbevlchDeQF6koX7Fv
8/6gNcdlQt3B9Qa5w3PDw0mWu4y1ik0/1yVE74hjn6UOstoQGe5LXkrYnxaEITNtpFdxr4Xbx+5d
Zav3xv9uERExJJuClJ4/YqQvb+JdDH0zGKE283VVbSLhgXdFvFND0IG5EhJKBtLuhk5fcMxDJuaD
6I3GK3w+e929wGLmvZLnHhrENJlmmm0MbJ5dzonPXW7Qp7H2HiM5DKI9FerqzT8zEY4oKkYzwd1L
FssRNvBFdZ9CSzp6xxqmeDHTO8FDD7l6b10hTWQiLiehCCQPnLGYjETPhgGiFxUcO7BevUR36nRR
l03yA2EjrdPpA/I6hLeoWxtBuNasLNBIdaSsdVfuHE5axAl4a2KR7f2gpMh/8LxkxtKiYsVOB/tc
YE1TbbGvIRtj3oMAEenNwJHe2p2xpFA9XVP0w6c8NDjVXd+x2xy9s/pjRRvvIqOoEGhqPBIT5Z8c
2acr4vQEMpsIAiGGaZRWGjq6HQD/qsvFxoo8aKkBblNFylUe83XZAQgBbX0wj/hsgPqGmwDDwkYl
TTwggCoPdeg6RCwuOSDik49O9I8eNWMUHzEpC618xXWtvIvAFHIGLcKSfgLj94edGpcamfMcvMc9
YJlR0EIjFvjiQI1WFxruo+h1xk2vdZDmxr2IuN98aTCPxU2+PcWpJIbi3dGSc0xhPugvqMTCMtAd
Q0SHd7HQEdjGzmaqajqo+vei4J1PtxBHvvTUcYeCgoP2LZSmGWNVYixzzFluzUiBdJsIsEx7yRl2
X+PyIp3rdCXcPhOhZLLpbBcEZG428IuUzROA7JIZ/7f5S2udkcXqHA81+36mA83EoSU+yIoy1gAh
3nZzrdys19seSHlM8cZ4Sg/K0aC3BpdIA7j6s9f1TcN7ORyaUbA0kOBjjjVCr5+OWsBYQj4Mnbvo
SjK/HZk29TuY9zKlIjGtB3AWNzWXL7V2gsg32+bsHUYyS3ZtiKMsFXDYCnsZf71q5hlJoBc4lrTm
Jg5R0iRszASRfLuxWTRJllrfOE67w3A06YmW10RwpMDNnxYeTE2BbR4NiLYwJx7hTEOriBZtzocu
TVgEa/Zpy26BjjLQUxERakbn8U2S0siqUeM0IxXguSNLSfjWiIMlIME5qXboICpfdrd+goBw2Vak
ZhPDTuD3muXu+CvEvb8T6VoV3pgnjwCgETlZEaLB5UT9nSXm5Ap+VouZuL1f2w4DgMwcN/Zjd539
OzAf7J5tlCC6i+b6FTqFwx5OCwzMvQmhFKmukxachz179UoEXY+5xr8Mv6ph9Wv02wq8uZkZFJue
vDPvgFn4kFOeKD0oq7/34I6USwkOx3Xlzwafe6lABvrtUv9HZHV0+/SyQPdk/Pzfe721sCQMGpOa
2LNUHaHuTC88FFuJk7UarMC8iVgqVNKdEBtgKE8uNGw+2ZKGpOKbUJRlWGrjgdckJwGUMBwYwzm2
8K9fbLqKYq61BSFo9n4rbumb0L2jdHHUQNAJ9CCi47uxEEJY4qAgCPA8Fzb2G6jjGIcQPzycvhhP
Hdn7Nh4pFiEAYk87UOsC96IidAZYAMT4vFmfrDw1yxoA6UEn8EK5XF9b6AN2qZMtacUDciZiJIFh
MkXA7HkMyXbKn/vzJvWltT3gCKmNciXrWCZjWhZxK3x5ep09WbkGDZaj8Q3q3c5qjYkkVPSA7hQd
/bOkNTERVQm9hyckHHaUmCxM1pGW5oqy8z96ybVNDkDTo+ygYWAioFaFiYIMs8ALM8MWb/d84P2B
YHnkNdKXRrwkUKqZfOKQfY02utbDj3tnW5PoID8eXthTzNk5EKhq2ww3bRttfUyN8oA2cj7JjMcL
jzIPCH+QbHUqG2iCxRBiwx4DrTtZhubZ8QPfE54eb3Mg0yTcoQRpJEdtuC12uOvOM+RRPHzzXDGh
ggXlUOkDn1ncXLWYCDW8a8m7gQYnbVPtwNG7xMHjS9HdAxu/CE1UQx9Er2cXHg/Nq9y7o38osHrM
CrFuyH5UnMb7AwnlUsFXUDe2sanisw/LLSt9sOPofXxP2a5aRONhh6sICDA645tKXOuHAFsi84oj
kWYzhdfCO8w2U/vfBw5MOzdOV4KJbtbwBg8aDAuH2wxfDJWuMselY1YZGoUVTpZpNNR2xmiWEFI6
dn9xIeKBzAj2NRG5zhy6tcQbiyOmrg445dafbiVawdOlrUZ4gbv1kBMimpYcEZyEM4wVHOoCm782
MsBk+7bCRCWm/j7FnAdHsjqG/osljBWbJsKqT/3Vojiet79vcZXVfDr5LEHDAJ0QLAv3ahbrXxds
xX7jdw1lFqukrCWrpLwj+/uqdbCr7NHtinLtkMkh1ioqOqSJziR8o2eYjJhYWLZDuIAUoKZRsIQ+
dH5p2X90KuFF21UwLeHMvQ/hnfH7bfqK2t8nf8kyiQ3iQvHnr+cZuQ0V62gETTbmabT/PERjLNVV
QADVwXgDas8soDJzyEqkxdLZjBnyV4bTpU/pLq8CHIjcTTm5WAGAmIvIfOvj4edktgb7asyN5qgX
S+iT5d9Z8qJDf/ptX4Q0HT7IOdjeaDOzNPonZC+xgIEzMRbP0kjd1yLCzPiJlitgHcLswIHDw8Yq
0vjF6khumQnc1EmvdYZKtACM2iN4NV4fgNunzY2dXqh+738+Znnd7gIeAHV8zRO9mRh2vgZQ4KjW
I3HYRMPu1wu6jvG7gfL/jL/iUs0QkiyPDr28fz/z4WbICNf5/vKAAL0KRyEOQnwxcxRyE/9mtTDr
NmGdn/tZQ50mdM1Q8Y+lXWOAvq1kko0FxNfsPBuS4/2q/3ETKOzo8c5x8ogQ/uKcd0ewI1k00+AG
+yMCJKiBBkK1mjOdNmlm2Ei5Y7d3x92Ypqg7a7WlgREiE2vmu9vLigs73n42aCQfgSVGQ/+fx01s
OVVAnDvH60PIOtb5BC5+VKVujRHl2JTS5IOdTGpDGX9No6WCtJKXqaVfKSfls4eHBgeTYQUvfit3
2V6XcfEp1rMrKkHsNPcZbfrad1Uhd2J8udLJG7ySsLFBjzRXkcHzj4N1o1qAtiE8pE3F0kIgRH7x
1VxqHPamEOmCr/mfvuV/32Ezioeny5venCYmZqrkAt0nFHOGnOee9IOTPV95IrNNq5MSQZeR+MIe
bUIkOvNyb5in47oIoJDNCJg7LuHG8YhQvmFHoDNsr7ovB52dlFtrrMi1T72VfhFFCQ1gsXwoj44D
QVo1Uouzmu0MaFYhzQ8Yw+CG3rI0oEHPggYG0D4SAiHFtHBLN6XNP0LTrWziEEhePg13rG0vArCf
T3KYW5sAGny9ee0hctri2CQpq5579ZPuSiJNQdovogyFdQN/RdiYIfB5BRrGUW77mouyH8Nqtb0/
5RFzWJzLbx+uZ0fEPA/JrO+yR4hUWQ2wqfNqN9j5tw98tTMfoYxrSNZayH7cdvQxCa4U4a/9UoS+
cZBAkqWrcqNer1rhz4wkYfhWQDpiGlfsEA5cE2SIKg3fXDY1CKWIv4RSY4yyA0nzswXqMDG+2L6p
6UCKLpJhQY1AfHA/v8oSW6mRyUy5cgYjLOODWDsccpsHHKxwBDTQGjePboqQOscY9Rk+THgqS/6c
ou+nZbIil2PsEoLn5hKf1qTs0UEkeNVidZIAZ1RYb+Kc0TN3NWEH2nDxFx382wyuWNqurV5EW4YS
dxQEQoh8+p7GudGS08zG5kW7bhxEsSqPQ5JGJueKs9ZVpsLQ4RqdUKa5Gj0BmKBeri83He+ABiYM
zCyFG/FOGhhf4tjQB+hUyDWgwRgtW4rB//SwgBN63lsQJMvH1r3AitpFlCKLB7Vmn3Vmr9kKxBHf
m1SlBf8UsAjM2UHjOFuHahojRm6QrzlPZfO5xqBFzDU1fdcQkwKJ5n5n8dzRKFgnXcPCR0EnaFMR
XH2hOsLEUpUlyYWgEES8/lKlxFMyV1po79d9+U6mg7gCd1tcrcpzgQrPC5kKd1z0Ff9uiwaV5lnU
NO8kEJaMChCZCPGXLZTJDreaMfkxaKINj2stIMchh0AGXW7gwRfEKIgDB3zSiu1coUez/V0QBbTQ
rAQ/DJH3q9y1lbILlYFn6WHKmKb2MBWsbPuLkX2D0KaYSFoJJy7EKw5cWqENUREG6HhJ+OQZ86Gc
n7CPTHa0oKl3LMZxTfZiB/avcitJKK+caGV9ACW5EeJrqn/QCCL0kNvz4DwpYmchb1UsI2pwDj8H
zPKfXR5yLt1WBvwkvHsZvI3swovi4vru0fj4/f9RJ3y/IhcwYv6+D8WUZpFca8d3KcCu57G9s1Ou
36YwAth/Vkhw0f6v80sh3r26N/9DdFvllUGda8XsQFi3XwnCF9ouTI9DI7s6u8tN0jUEzbqAPzqM
evClr7lLsXbV1BMfMzalWNDM7hnXUD/c0McSUuLcquOQG+xsaA2/quuhXLwexdKKNnIRB7WkAVZA
WOXLn78jKdWJSSawkpl3BarZbC+D/7w4Qte/XZ161Xtz8ONokAgBX6ikD/CUzA7T7csJ81GNheKX
Tdj86sitmI8dpymLDUvzkp2oCpy85PsCWsfKYkthIxpFUQs+z3UYhxbOlnEqgzmBOJZRmuF58sVd
SVt/JxEcRJ82sv/KhKkGFRA6+A/TSUD1SgqNoC7izuujo8E4xDymqE1WZyL2di+6Ps9cetvU+JaT
k7a2bZlaK1wkoZZp7iv5E8x/a8O0/lw8DDdpWN2PxcN7UNejG125++SA7hFrr51ToPKZO4zozaNH
aqfZxdTNMfclkxIsWFkd9ZNz0JjkFYczj9i9NmyOwti/xJuf7XZmwb+nF6B8KZ9B2puVWPUxD6Ct
MD0ieTGmLdhgh1EmzGiknZPUMfzsuzQmXDio5Y7/VRQw0AZPiWrq9pNHi934bklJX01F0GBtYkJE
zetmOgr8L5Sf9q3bj9rXWLLr5deBB520CT/1TaLck1cStZX7/kXlEBSxQsP7dUMf+y4e2k5xtP44
yoWrIOC8oNGK6kVb6awcSY11uBLt3b1D9rmLiH8Jd+Ya63HJ2GFTpPIITbD9oZ8TGjgM+N1aoyfM
wQSJ47l3gFkBO+TG6OAYrCeLq/AjP8vsnoTvgAR+XKlEYewlvk3JM/8Ez8oRb/VFKuH6FNkzRpwZ
dJBauNNMEKtvQJDAotsQ3P0g2xvCn/R/ZnGYTY3oIbgk0NrKFTJDGoiC3D7c0oa3LMbNx4QmHboh
Fkj2xTSpft0+HNitmbkTjfKPiDVdZx+hELJ3tEwuC5K+IMSVgP6JDc4ND/dmC74Mi/qUUayGtJ4n
3rjKauYgAcYNPFShO9Fe/Wv1FqGvrw21PHCFYfwNPYqIP3cuxAWTn3J+lvcGvYKkvKI1FhiS2u3D
gBhFj7w6e1l9fZVJhd7X4RavJ+21LFLFSZsmdRMWKLuHbwX0J1yl2Xzc+UIGhbULYaOxng5Gf+Bd
59oBxlBwMB77lkOsZBWOYDVNR01F8537Dfjvc8QZEKYfR9P4ZWQlhkAdZMIXWftPstHjhNis4DSx
zvmTxBxYv/2pUU//Hsm5GcR+D7YIUAApxpFlQ3wOyWECssf3YOWLOrPPCge+6Ks2e9dPGvcEtlWz
DAROxP1ASsWPrLBG2qGHBF/JhB1Tu4eHp0dqYtiArkEdrwsYQIyXTz2N3Hy1q32oqjqry6nbtzL3
CNiAbICd4ITg7izvvMpaL0ctKiJd1j5OxFOpCjX8g8KFUP2hNm9SlyFSdNjeABs8wGJhotVAXemY
yMYrg8SVQRUzluoIB/ULfApTHJ4M4imMSz1QJeJhD7oNSLbBmJ8YyevV505zLGIO4B+B0WHJrWIn
gKGdaiVShXYtBYWlWlXFZqkIWCEmFHQxm7ym2I01WKFGNcGeNyayjitz9lwE3jVcQv6Tko0mSOsp
bPUADyE1ebUPl6uuuL53u0LkTOMPjcbkKQ8ZuWXd3ffDHSkAwqLnrv5a387NfKXGywJpaUst0dCU
rDYA1UkXJVnGaeVTSqRCOzZgKbOt9AIaEJ3C6oU7g8gar4iNkpdKG+PCuYAMbNM6c7SI6woF3RIo
po9pHHQAxSxB4FIhsqJO4hS7S0TwLcYprdpnhnhnXeBnlOhjUHpPVdTZ4kmCeLVpVgQmYy1Ad4pV
yjhDxi88oTtFWJAmzThW5tIFSgw3MIbvkJNWB4/XYS7LelLvqDkVX5sRYFCEWyAzoEHBe5mPikAY
6AJnSB/I3cCPK0+Z+l5q7swW5BrXz1+smhYrravu3I96kx6aYmhBiqzVDMR6Vz37BMt66MszorEL
80jn9mM0jNgDfbC9dIKfmA7GbPqtrdJE6CYxfptfQKdrs11GPCZ99/ELpYmzmIJznExmPHlS5/bf
kLjujp0yArOkxmF857esUQgavsZL48L9gkSrLhwnYbXJKnRwUJaHM7k6tCS0Gg8boCWZznZXCIva
k2jJxIH/LfFw1y2RzSGLapj5fBZ93xq6by4rtT2KjeRDowvtNZX/QCMsdS4XU79Ah2JsJDAE3/8W
tfdasc1dmONQIgm2ilsm8OiNWONGmxcamnz2jDdZmbVtfl+uoCE4ItaIhWAmuIlrc2TNhRWTlqYN
9hX1/uvh7+a2mTKp2ZZeX2v0OWAyGWLEqVm+XinGA0STh5ehgwBUDAVEsg2iMx8biHzS2c0XzLkt
4JALZDv/nA4QcdO6t79uk7ERqSusTJi6Viaaa6RwYeY6wu2GXBY39JhI2iy3Frn9RUJcandtZtWC
wSw4mnMs3K85G/X244ec8JRt8kBs0fjY7bSOuOhLRiNfvwS78JfLZ8XPrs+1Oap+9QRpQJTBjM99
HubV2HuhvOBH4xOekdgA1MfFcOysWO1MwgkEyxJtMaq0seeuVE2qJCmqSvx0JjFkGsYgxFPezzWl
9+ahBLU+WwGBd9KW0FeIvnb2Zlue/NiXsjH3Qe4JzOHC4JFsALhX9yedOnd9rlFIBaNeHHvXrv4K
ZzwCuHYIkR+4BzmNVaXTonhKwdRbhMB2nMOQ7aWMgSQ/VSQM/7MMNljPQzhQv3xqU5fNhm8kiorL
cEv4rY/VBiBWGmIQ5yA05A9/k4C8smvh78gHevndFGvrEX6vf0GPikWJca8JxlZtqbgXW9kIXdg1
Lu2yos6vbhIFq96XArKUrQ5xZYqzIse92zEkSTpA7ViolQdlYtBgvZMO5FaKC1mGlSvpVH8Emcv/
BkA64MKB9FBCYm5/TDDXIZCZQBsvUDmlrAhpVW+vJS0vHKJXOci/tGPlfq8gaBRMMxpJwGqAmdws
k8PT6o5uMZW1c2SvoW/p5RA2wWoPAzQIqalhrDqJ51rdtYPTqntsXF59vnB9hiHtcof/BU7xWFPM
JFyKwngnh+jhA+UevRnOQpB5qAVgnxkLJyF5eMIYlSlAs9ZXNq1LygTUjrqJqY570aNIUDUcQKD6
zCSeGFVibjFKz67l47f1b+BFjKgDrqt1CKmhNls1ZhVq2TBNsxGhDUAZpWzlXNb5AsULlmN25XTI
GDd401f0kTFXUYC7uvQT+biCgWIrsHg6nVoTn9wC+je9YCsOuLUFymyRcXfrWBSLDalJZ2pIzkIk
Wvl0LRA74waOa1fmWosGcJox+dYfxKjwxUQB/MI6URTLvSOnURw3qiAr3J1Y4AsCLZ2xAtUtFfzX
31iTQuObmPQJVNVahBeNGj1oiA3UyAZzGifo5AGBreHR1hPXplpJwu2Jyo0D9GYDScGWSHcg82Y+
q+baJzV+4XVVUSTYTe6uz/hvAE34bNly+x5TVF4Cpgn1GlamrjWQnUc6amrygNy4nOTnnRrbbX4E
B4w5f482o0XqB3yZUDx7aafLEilHQ3xXRsrCE9jld2gOI4QtXgp4rFBSn7anANolR1MHGSXGD1FY
oGMDrse1aBaKWnFNdGozrWGYytSrJfO0ScglYlnt1Xd1qGJQv557b936ZL4NxyMar/fguvl/Ruii
UUBFA+c0higUiA7qdfwMNP3MMj6ZfPqrXO1d7ioahLEH36Ry1k67juHDDqNZKDHrsaxwz0cBVTY2
ULTnJ/4ZaeJUCgXhpX+5EqDzmjYGiIrK0bx0R/LOhWn331E59Gj5H2dbMT6m/wUHvqT4qaDkXqUO
ELykqHnnlmPNY9ANaYqvz+YIg6Bqrx7CqDJL54fGKRVMTnwMO69s2ftEESll7AdSelJNu1Tf4UWT
FkmFL1Kl4GH5DXLviHu2IjMSV/BSS9JHV4Nq4eTuF1/ADj97lXLHo0HKmui97AED+2TvGHHj0qg0
azh9sQwjuXLE1D056RJyb1UzTNfMyPgA7OCoCj9q1TRT2R4me9dfvsH+USTclubisD/sweQ0X50+
ysa9DnSN+SEXVn/YG7fLYzfvvyn9K/3nL2MmpvAz2IL05uQkd+MZQ/pdxwutHi8jLwX7SHwoVsP2
Eiql/urRojrmBUmMejgE0ZBLXOkG8QBlZVna35GPQsFIRywoiSDPMRjuGKUkjgl6FPR53Fqlm9Gc
IjMhBKgPDAJfrf0Lc4hAyG9rIMp8izNvtTipVwsr1GCeyvWyAJ00u9KJIADpah4ILVxey4umIhyk
3A22Zgw0dxIf9cK3XvKoEBt+NntFohjfFq0RWOotH9fe98SEmbowAHeECthZdFdfbIa2m2z2k0o4
c3HnEf8/RPWWWlWGrmnUWcY0hz0k/6b4r+Xh72yw31/MlEG+OYyhchjqmf6kQu3egGQky9ehi6E3
w8es//k5jIBsIjBYrO8w/gJZSnyth+jeQuJAZR+eI4qJDbU3ThgAUeP9ELG0CKE57ezP0IhMHpNN
rUQzzSfR7IQFUOOkr8JzffIBM/KLSrs4d8of6V5/F+5KqV29gS/DUPfXEPlgMILi5AO0+faT8Mln
G4GxbsI+ltLtButlu6kFteQ+Nx5zxe4ga903q+GIRRauawzB7FQj78Q7eGvVjl6nVPg/+dPbVXmD
7/csd81nbCxjEcdze8fBta7+uU9ywom7pIUn8+EzjeHJwH5XmPUT4GcS9LMOih/v5gDU2UGOzHVU
zwrwyEKXl1AYAiFP+u+iBFtT5miilwzjjg3i1nrdKe3zOG53JdbRjl1TNmoZnYwKJ5QKhI3QWV37
tWWYibgtId2PlIuvXuUXnWhdrRj04EmcT3QwtnKZwLtjrw/7qvz4gizL3UffQKobWxO1fpJpXjO9
Cj/apEephnF6ywYJyTtdQl3KO3bOdjd0wYoHcLfGuciYg7g0G76wJzJFJWZliRHNHz3nij9zqyaZ
D+d7Z+G0Wb4fzISpozaOIrcJfEtKIURdHtoN3YF2gpHxleECjB7dbxMDBPSvAaZxp92yVoG6CaHR
syIu8fg1tewE4OjOsm9FBgXwpMhOYCVO9Y2ZYVzd6cE45S5aFRhOBjOzdOiMv7kDja/l0WqgbuF6
FXh+4B+wkdj49WDL8L6LFsJ62nl+b1uBrN1vdcaTHVruQh+REYESBDw/+Risug9bDvAjqAQBMLca
RXipO1azap1MzpJRLa5K8aAUW197YzK6lN8ks7U/hb2ojDmUL0KrRM/AB6SQdlMsZRqLacC57ji1
kZIziTzkLzZ41+ZuJVzacemz4KPXFA+H2rQrfJhlexWmFSuwyTFIPrwWJvo3vQPMO6A7aBE4VkE4
SrNgWEC2TqQp8MHSawX77obY3R39xz7o9/JlvBQej4qSbehw7SpWhvw2KK5XHh6zadtQZbqZy/19
antpu3vFmlSyKJOkI5GYiX/lumQzmt3EPTzJZMfzX1PC5/jc/Eij8bQ9J49vqCdwap8w+F7GupZm
E3XfaTcdZD3bf2GfQBAQ3xQn6VK/q1xPTvNYS10yCVuapQVCs1wcg2E6V+Tre3BaC2590AJAQKiy
OlitMXzDxTldG0HaUH+PK3VcE9r+SOtI4LP0XhLrRQNgpjvs4eLssNNkc132N/qHTPK5nXdt61rK
x36+4r5KhqOlbusYIn5Brb+kKVmNxPg+oWFHeQo5ceU/qqQtx6QHa9A/UgjEXbx9D9jKd7u3TViA
8MMTUzjkcCEXbYCWW5lQJEL5ST714v3Q4FdXjDePODPwyAHNfqbxOKxzeB3PRRpMuseyF3n0w6hq
LbMLO3u3Gu1uPsGiOY53lx8NFniU2hWXomJBUWjb/g+LX4EgdRBBgGAdXcWuqMrBwqIO/Zcxx5zh
LtwnJNervhaHTbXzumog3N5l6LVOvuKuOXsWGiKCB4KPNGhZFFpmsbzhsTB21C6gmNOByA79slT9
zaOg+WG5S4Fy2I6wXaJtv8Stx89ngirAkJ6Q4Hyp8W5moapaEhj6Qmi1MPWq76WNSCV09+WAZ5Ie
Qh1hyMQ/A7xOrmwIlaaXweI3InSE2lIR98eeaWQQF2waHYt/QhxASmjiQ8y5YGD8FsFcByI1eHCt
enPI3n8TB8lm9FNcT9lckNDArLWia1lCe77wyPeigZWpB5BDtCGSVXK9I27fx12Hx6xSnJgATORL
ekwpNX806gpSMva6RhPl3BQm2LjgkJbFOgpzWBlLnDwORB06bQCwRX01YnNpicrfiM77weEebQMn
1rmiuME9zQzKozcmTS/sgxZkw1hC9tpCmg3uMpq4Qlf7+9k3dPgQOknenbCMYLaFu0syYDj1pw8I
yTx6gSrmSUr5Fq+9awjwWZ3Z9LXlT8N10NPt7gKQ9ELzqha/B9CL/Ng5YRoDhkWJbO0CYH6aTff7
SLueQeeH52SqOpbcy9aketGHguavPmqibb/nTV2jKJVm/xf3kvtPHh+fqBDbbzlOnxnXSIAgoFhJ
YX3/0YHUUK+dsgTXFVYhZ3iwICVmTdTFLNna5YhjU2p8yRXxlnac6O2tcxqLCVng2rY7xE4uBniJ
gzdkxvyj5kZqPsVFgtQXauxUvvgdeUN+lkeTuJIRenNyvxJB/hkDfduVjUSlPzQfITMgxZ1NnlN6
e+Vk9v0HI+vjSYI2Ggx/mqQHFeufmX66ie7LTxRN+Kv+q3GPqP87RTBZKSOAJE9UR/4Asu18vTft
XqQE0zndP5+2ZZPjdMigl/FwhDcYlJ40CbZRZ6va2NPtVgkyDFhUJ3bCa2/5r+pQCmjXPb0WV54N
aYva/9470b46d2aitTnnhclnz/1RmilMkrT18oo9ewfCxC5iSlQ8q6/jIlg6xq1A1mcoyrdroAF+
nO52WGUuCJ/eTIJnnOSOhb9rsjS0yfy1+TOtdUgtzlog9HpAqxHSeQKiGGxs3Zt/Hxp6lrhP4X2h
xdafFxIjkBrjM3rnHq/1UGWqFK5CWV1l2P0BBBzuwAZap0w71f7o+Mq5+KMajqHl+VnPLkUqTD0E
R34TCYBgU9R16ahARPay9pPvVqGsIjbL0RVo820/lnDCVEiFVq2/fsivjXauwl9oOoOn6M664ghj
bJuFbahajNSejZrELvNzj8ZmrWOQgq5NO4wWpHDH7FYnkivVMjg/UpOlFLHqlA43fwJuVQ9NfSSN
OFcIdu2TbHuwsozSwlJZKoe0om6dtWp+AlN2Jij+69zxqyESK1aKXcfmnOmR3x2mg5zJBMPGFgss
cQbIjTp2bA+er5Z33mqD6hGq24WOdRTTrI5HnMKdkAHNOuuD/x3IeXjUVsPQLn67w+V0aTG452RK
4ubu/PLI8b+kvir2575CEceLwZlxLOulxwdCSkck5IqKOM5/QOEvLYWFxGDASyAaqAvyRjPps69K
6BGjkr0eUsmPQf+/PoQsZcJmTtKxp+KD5ZaoeqN823TdO9Wv3luED2aS9IACEdrvr9xcjTzK36we
/cs3uhspG3LWvpVGbRJPoiMepdR+wzLkvJnUDKgx/QuAaO2NkVuVPs5uj4EEzrOu0UjqnBEEVwmG
lFRBk4Q9oqdJYqJfWMtSNajDseZ3dfWRhK29Wa9Ch0acTySo5kAeymjr8OY5GCdVtIEySxTy84ML
FuiLTgPSrp6d7QM7SFBIMMDgubk5Nxf9aDYhKFODmLLKmp9wrH/f1uZGfruyDatFZ4k2IOnWviox
5m6gXXBDzxEYPYQ5Uk8+Fr05bR9IXlSN7Li3QNxKzH6RY15PrNDIF4nx9g9VOwrECHvsV/94TCFZ
HrN21Eujz3iQhO9dqwPk2CdUG0Wv2uDlXmhthrk1LomT/KUbtExVYJVMt4WkTF4+mmNwicmOvXba
xsmwRRbZhSD/6NWxh5Ze+ZU+RBPJF2eIvP+B480SSh6FJ97o/f7UdF2EFyBnMy6AB2XT8Cc8a/1l
IRLp2qfG2zZPl/Kaf1pkZytqKI3nVKHtlbqX1ihKsHDvHbNdF4negyla6JlXflPXuGasnFbeK1Sd
uk+Us6QJHeF5DgTqejdZyvzRbag3xjCLSGhxZqa4Yz3PGbt012lq0rBeCFbQQRPwkJCIulvwO4R/
IY2kwUfj3WpGu/6NfxU5kn8ixG5PTYtj8Ktq8/3QITA9H81byxk7CI5CjNJeHO110N6MjsS6Lorh
/irMph9r83MGOd3gB6Vece3zFAwXUHRuGhhohQleXdA1c+Qq5NssGoI7TLQtOIKS8yJiAbxKicGh
93s9m/nMUdEu2eHJ2QmfLNle1I/7u8C+x82+i+v7ooWGnbGO516KAY6AVb2+bpcI+JJPtEFHrbCg
rBsDiKKFQ+jiccpphG5ddmOWBXqEMih5IxTwvsk/rRe4GeEBOh5LJ9IeB4KWiJkKNF4yrvTO4svu
QqnO9lei0ve0zwEPq//bpYeaWbp/MoFp94ShgHKm4ALWUmK376D22f3IM21SoNRj0GjeRITJ1DcM
LTkiFDnMiHvU0XZRO6kLnV7jJuY/SMDBfW1SCvGzPgNwRWLrSyi/xniVhKwe5jROfATsklDxR8S/
3yoRtR+J3TAGYABacGTHj0uML28wZ/GABoVqoqF9NsTq1H7thbU+Tp2EAQkSxknT4drszNTH23Fp
O8KQo46XQEtHwyOGTTi2eOqcvWSftUbWlsS9bTL6S7UUJ3h1dLDxxTuN8UdTBoLrddUTQ0+3Q0v8
CbjOVZT7Cf2M9kEDgxDweDwUL2E3EHBtsMbGZhM2t4FMgKTD9mmwp663Inw9EGOgql7PsFfSQa+3
m2O7JuMQcZFrjab8a85RpTSE6NxjIrUAK7CkCt9+zqg2KtA/ipHDO/4apewPZDY+YzF03eSfjtmr
fQblos/H6aNmvZazjg8k+trQKUT407qYnmsn53xYbYtY6mS3amZtIaErbDHc4dsWoiB03MVjuNVN
rLLrFGuDQP+oP6LHUFNHBpoQeWhgENfDTa50aZ5zNFGSPpZzKTm+KpOoOYYPED6LUh/MA+JVOY77
8xVsE5UxBDIzsj4+uOB1PtVxjx1NRiKwvav56AinYUv2si6OSmFyxJDKPdPx/0QFRsLAE5tY7cba
65gtk6WtH82fiw69cfkBfmZttrzhgiaRrlDxrEexW6XLnXMSBaqQaNOsUkHvDN/roLBBEAD/Rdry
DTqnf/3YJb9coKqVivpShfrLeVSkP7Nozb1PcZCyrj99niHcNyTt0rV80cyvcuzKkke1lZj/ELjl
5QfbLBs91fyi9AS1YqBxyNyZbSAneErJ9lFC4W2EQa6Qd64LR2L/9pA/xPfGtcAJxF5gN2zOia2i
RXJjxGfKhW1PLe7K0dbSrXrkbrbaGD9VInNHeNOWw9vTM+CNT5RYtTTM8KCbSCzEaFOw62WW/TTs
QU8MpHe0h6dBfnjAeslNpccoLiyqZj5K/5ivTgYmz2eF8ks4X7FPvwVYdeep6GcudR473U9lTDwI
kIChtNcV7/xuvSUhB1KFsam/fJcNauEOpeQNQzWiWc8kJIUYvOcDwYinD+Pxyypfg76yauFzxoSH
ePH1HmQn7YZk0/0rLgYLx5AIVxpx1cwK1XzbJjzwWcFjrfaYTX3STz54Ub65z8jg1F077M37IzoK
2hK36uJ+0uRoPqKsUnkEhP4fiDqiAkOzsGYrndDPKCeS5goeqHv8aPk/rWaFXuf4pNl3ZrB5qlTM
4B1gZ0dfCgXblZHqaVsR93s7fwEe/+ABZ53AucCQS2vhWuJmEd3Qv/eErXlKeDTUWmkocCrXHLWt
yWyxX99jheRx7EN+CbUZ0zdzZyLWhyuOgDSIUPQC+HRsfsszJFHSLw0PNHa4MraoHc5HHGJ46Q/M
qReeAM+EdSzjZadGNx3hW4Oal9TLtfoTFzDE1NDYqPGW7dqac7poJHrKkmX2SCdqZ4BjVYU7J9FC
JLI/sT3wjGA6yvY0Sj3xim2aLsIWDK6izjguL7U9HBjEoSITNIjKKW8MgsD6ewVvIjPDJ5ePdOAQ
tSLeva2vzgkiHE1H2Mi1NvjrV8OoSBKmIniQI4fw36W0r4amhxs6ZgJu6h+y2VarMnsqCc7zx7A2
7wTnSRC/kv1r6dnDXNNDXoRmFWaZUHuopdMh0LRNTD+K5AXoD0Qbox3HHwmgqVXDtSgS744E4l9X
U2fi/5UOecxN7mkjBMuV8WqYk1gUl+qTbI/TY/iFsLbsouSEfH/X6MN45D4/HUZN3bqEiMbFMmj2
dm6sO9Tb7mOVSjE8wMtCdYOmjwGitoDTb2/dnZ52gi4Fa1uSU02U5hEKh7RSFOg7tw3qveocvAqr
OfluOO/yoMleKl/N6SCFmg0KadicwgtpePTpQybW7SdO1VyH0rWncZmQIpMBfW4/fN6HISApGQ38
ENylPMFDMx5fHMS1lg4QtfU4MiQlOz3N9HsGyAI1Ac+WIuf6p/6qRD25HocScnU/dTQgU918vdJp
koBpd3tLE4+/NGGSYmVIO+6CO2mc6tgSX82WvZ3vnobRhOj+6xnpl42jWHIJrWB6G6dX1Cl7ZVYB
497F5H6hAE8qStVxDqfqiv8oDbngx2JAxmPiS48MzvP3Jf7/zqqshl+SP46diFYFezKUFX3Qg3LM
QxP69FePaXQN/GMEz+GYbeq9sLqaLEMfVG9adTxFgMHwFAMPCCuXHss/ONKyKN/Mdp4zFIG6AWlf
ynLxqhtX33oPDwEbjkP6WyAbA2i4gbnkJBJylo9Fa2knjdgEpGhbu7IzFZxvU6QMZ4h4Eui9ZTCF
YaKB2+BkNW8sNdOdrZM4y+38Uunndsn2KHPDnVrS+E98JO6bG61ZSz5ROT74+kz4D4viM/Cumvdr
5o2sWmXS8+gKVubf76ktRo3qdOKUgdQGQNL/WP1ZibxzLCHblpqHB5hsvFtk4pcb0rTCMWUDfge2
NhCAXOh29U7dawQa6mlUMD3ASD+XJJnBbNYybkCYzeZwONWNHg2qXP4kj/SKcbkEunsOf+oYmj0E
9CFNwV6/A9l8NS/1KR9R9l27hRhADA+Jmreo4jBPlU1gcbIWfbpJ8KfN+ODo3JY94cD5r8gJ67h1
yzhuEa4OIBHpMQwGXLGzYFdFJqmPfna/FTXpEUBn5gktq5D1WDIKcNrT/xUXY+KNlNKNVzMU2w4V
0KPZbYtayIufuOW5+Z7l3JT7v3l+0h6YFeo7mCgmrtFOq4w4iyjouCdPH7ZH//NWbI7+TX74YVNT
zGRBKepNpAtJif52AMHb/RmIp8Q40K8+AicM9RAa1bcFqCwnykmQ0DBpCDU/Jtns/Xerf7il5f5K
iKiQuzwy00A7fhKWUDUJNtxtEHGSNhHSFm4BDAdpV/fqGEJOTkNZ8LM7TxjovkjZ/0XyKktHPKm9
EcJ78ENGRg5CRj3a4NGE89g2YUOyWbJuZ6Evj2fiqePjTj7/K9slL1ElAb1F6f1JtaW/RZPspPzB
LMLrK0ymPcEikY3/TN+7LNoI3CeXFETCluy1MPAF2fGxpHkPmCyiXSZkmTc4/Ulp8WmyYJVDqQ3j
D2zIkZlkUtd9QCnGABIqy6Kk2v7B4kYf0jF1oudRtxS/gd66d+is2S1YmAmFHJReQbrK4Gpmbe8B
fim5DXJ+uD57f4ZzJxD+yhlWENte8nXp5ovK1Z0LxcaWtHXgnqCn1QZSAQHn5q9C3UggqU7xq/5F
sI4aUrK3UE4XD6zgQWabndhLwDr4vjGsPBDTIjDbKiRlxBgpkWAP6k7ciSBB2ovdWmqRLeN6Y/Eo
CA5vVPSQQAVfopdF4Bclu6ebM20YB6K8hyapNzNgvCtpvnx0tV6Oat0AXulmrL4qsieNcinRhNl/
9k1JCNlIgMLWPS5Becf9EI4F3aGOt+l2T/Vwpr56drRP8EDLUzfpZPvRClr+Ba1/jKuoiOU4K4V0
wPkX+UDxh4NmjNFyB4GdjkkK4HmyYunr7k+CUf5h2hwHRmJ5DDa0uooMyDROs2RZ1et1cx02megQ
RKHH6S6SEHLPk0n/l0vBa1H/9npwxmuuNVyNIjNuCA7uXpNImTZtSGzsFD9/eRF4bwGLjQNOIhyz
j6vwi1FlslVxPJPc/ps8hCVQUZUsw+82OKQpXV5/bEgf7fxvNGMr20XwNOL9SCGOFzesxZdwYjcO
rLyZKsH+AuvZoEK8Fq2rHbGN5hcFKTYfbUapoVkO77/sEM6IE/2DaVmtWVOanUxAESUBRM5J0Zt4
CIJ4iujtkk5YlybTgtNdenQEi6bWwBKs/PKyh9nhEhmKzHuCF11D6TLKNtPlp83fK34//Cn4NR3Z
cJ16cn8//9+TTrylwOzUYzcfRSgcyuomZnH+GIyLp5OLihpwXrUr4cdNgVH9cPr83Iw/+S0Jw7WP
YmrMGarWbhennSELgkfV8eRN9LFr3ZjGVhwqSLqDh+pr8GQc67MuozP1ekXKBv1LenHIKt/M2gp2
TEpwTR7FEUDwpvtLD1XaVZ0ihM7+YUiYrbRwZkHFpHPpejO6wsMQXcsfkx36WzMWxpaqcKf+Xpgk
5mwy9t7CS0gXcs1yVtMbbo0o7kkgqwo7TGE0+o1NZclQ/Bwhx1tNLABLTHV1kwLvXSuKe7Nzz1sY
CQNJSh9bGsccCcNPQdxkzGArnDITG4RTd8GqFKc3N/E4nWCndHPmQWU23t0Wfk2A3oMYKUs9hTva
0eGAORSmiD8EUmnsUQwVMjIvGuzvQ/MS46eF+RKC5zJU663wItbZFnZ5p8Z2ZOvO2eAtBO/c59je
oDe61hFqY+PNug0trp1abVGTsMHBQJoKWKJ6PyxFv9HKWFklXl8FuxRrAXR2z5ED75LGPHWkHYJ4
4w+kTY9uNfPQmsTU9KcCne9Yq9LeHIOWxWOlP8NRONhilr75oQWpuyejXpEonfoYq7N06+D1+JDo
ljiZQmItt1CqxuSyNnJ2uKdWZP1NgczsGuTn10OzWQEQr5QxVqs5vDqM6wEsMgDyaWYPbMP2dTOK
Zva+y9ZWgTHNynpnb1cIhZVSbFhEVLaja+2Wl6OzsdfPYADydP+0MLTtsBh81LuZbZ8o2u9zUHph
DYgstex/fGzDIZjuR/C5qHitxf9sg0ktwUN7R8ZwYot7Ls9swUvmpqHY4Q+soqfitbtaO55abPqS
Db7wFlmm7lGgSQUKXho26oTe93Y/nsT0bIAI+iSTxrwzEfer6wuYcG3ngyYDilhxstfMFE+Tjr/m
xZadYa+spIkE3mG7WZG78iAxmpwNQXV4jN3F+VD/DjqJ61QCgOn7MzCdpNEjefcE8ZpnPZaWQgtB
E8KFUrd1ferLY1LWBago3ZxgObK37TEj3iNBhE0RN0JUDhsXG2Ih8bklRtDZNEzF098s+sVbBJ75
SwpGKUx3q1PHt+MMECQLjQS0kg9hp5xqAjVHZ0rUqBI4Q16snBga6cVNRalBqC4WyEWzkgY8wu2U
A0DyBhky5AqkLSZKELpkMWQDvn79c5TTjNxkbNTLUj/N4bm/p1IrNLBoaKdHj4o2e+QpFPybPbHg
bpOdxHUM1a5hYn9tnzAKrnBpfTKxTGw7orqpgQt+lPeyRD/6xnfWlofrksSzrbbfZRtUFCSBRfpT
9DT9ocmmWHnC6do1xeFNF3Rf2mS48wdK0Z7okrNbUs0EHiY8SWXhESYKflyGyI7PuMeo1j3FTyWc
fQCo8nNUDOh1F3dUugiDIN39OfWbqZsFE4iqC7h53BjHtGFOY4Kx2P1SGDlWRKwaVLDewN5iU6QQ
KR9UEoGZSO/G8ABA3TEna/nVxizlyvWULWq4zJthTy8xCzq2wDNpeGEOoU5Uh3/JTGcgiRsjyAmA
8fZbw0QdHjzaEzW4rw10N43PWKGN/azrjeJibN/3C5h4XosnsOyJbW+I1uAqZlO2MvEV4tahHbeh
PagtCiwBDspMMIkNzrQoaLePj990K8PVHRJ15kGlFZYg9jbY69+mcAozIMDbQUUt7MkTt37cXNk1
sjeB5dmB75hiWGuBOcsJift6mJqSZEGldSQ2bsSCMvvHwO0KkpsFTq0rCZLzQM7au/FbcoNWEVXH
OUg8B3xCbf7UEJ7NlLe7qASNs4Zd/99Qz5vKzklTqukpaZlmL1YVNCoRI34mQZHQlJn6MQFaX64w
YuALLJBWjYlJ9mFTC88BjpAnxO1LMM+MQohFQ5AfHH+8BlCZzIv0HcKQB8A4oHsRJV1l4aQ9IZTc
iFbuRekJFuACmQmPHvdLOtTZ8il2hDkeCMZsuhmceXcSNcnoaVpYorSEXTLtTnRvoIbl2l7fILli
wpeeayRbf+vQn3/CScYzOaVcv9w84b5oVQIjindndTD1YgheYyfjUwbmPfYSSDQjW4kc+FAEZZ7S
OVTZwfUQgJr19fri9DfkZBxPymkY3oAQKNz1VAeGEb2pWjhPzcH74+Gr0jrmeCl9N/ONJwa72Obm
GHcoueMsJi7vLSPHfguT1miX2kGORKuGrGgDc8Y0BPd9d2rkPCBqiM8Um2W3TdvINIpWRaXWjog7
sOCWD1QlSRK5VkrbCngOrOCsg0z8nfK9407VMFv4joUrUTrFBMsq4vOCv4FcTIFZU9DEOC0gfdRv
9WnrvwCeZgApM5oTbNPNEDOJIhcJEJ5ap4bnNNo0Ai87fC77AMosSQfUfUm7KgCKdstgrgdXbcHD
oyTLmpMy4Hl4Ockf/9Ii+WksUj9i4FdGhKEAda8kePQs+iVH3B4nkEvXbw7FdUi1ZuJpoi/1n26O
VITRQFzjkp8j0HLOKQcK7Omz7jAEAD68/sUvNb3kV0QGW+WK90QLYFwiArS4djqEeONSJBqyi2Qg
tNv3yan+LoRj9blnAA9znJjtROjlHAzK1xI7L0UMlZHQz37hgGyMT4RfIpqazZ+6JkABBUU6NcYT
uI6eqdkmK3Y2GZOAJJRtZUft7+k+67PscVIyXRj+vgjCdatUzyGnbuu0Y405tsdZqqecytS2t+Gr
tZmbRCrWU6tehIqxyERtqVPiiZqvaaye2ge1rZbBqxsgUd27h6X4BM+o5T/gpJAjMAKMwbLdTJsI
CWq3KlQBKM9C8dLo99WLy4hOoKgkRdM8Obf2PiY6wLVx04Dgai9nC5sLM2D9D3sz+LtfW44/gCV8
8IyL5hM8nCpiMJXRgJZTLor2u0LGO1tMYey1Fw3UKKIwpj4Q4UX+vK/QtzLXJSrCPxBs9dPFWEQo
bVfJMxZ3o3NMghG/P1+9Pj8HbMNehDnLoaEvBG5m95OKgMRga0TeyZihJtKSPKQzYBy+C+cpeTQe
P+jg7YeWu6GLJaD7hr3G3I8rB1axaFRXj4OCzVdEvCsEkzwcf9uZzxn0snWh5KGCtZ0WbnMMUd4a
WXnq5HMT1/vu6M1uJMh4Q0QGMsg6ReagICXTcDRaid9pPOeZapEfhyUDOWLPvhrMzl09GeTXIE/7
ieP67LlmiuSHzp6p5vCytgZTle7nWs/lWr5YtNxmoLUiEZ8RE9gu7Yh6d1Zx+1lq06TYaYZh5yiZ
fU7GCb2oeJu5sNEi39U+goFm9KR/6BfFsR0DgnqS1Ysnp4yy2/ffP2fiDXIvh+lUeGLBp6yc44jp
jBQaiUc0vDIJghBb1G82gd8EpEM9gRgYu627QVG/Ynnp7Y6yE+IbTy5HzqMOVfdOibWHWqmq/q/r
QW2YkvOC6WafFJ0+HbSL09pgF80L0MPHDyUyqEfYKS5Ob9PJGEifOyj3DFOyHvzZIuYoCUXrrmhC
kuykRFVPE//VW66LX5r3KWq6J5/V0BFlTmfFIuf/4Cbk22NbQM8IkapMNt5kWuxaL0c6tUJjvadj
uX3Sxg//TlwqyZouUW+ZZY8T1GL66TvMY+uxYFqD4zVoT6DOkPyNV1Mva5gxlbpgZACOt9NqQ58v
sBCqfPkqEmI/pRvxHEDaO/XUSye+DAw0zqaXhYz/rkZJWcOzfpYfva6OoHUX+Mb5XmQd7ejFCgPO
Yw42zhOJ2XQu8vFkiUcUEwWzznrMtqCbBTzY22VQMUFJp0muCbPFjReCIyKP3S6jwkI31rHUVGEU
L1PgX6VD4dCzW/h9O/UX5rgIM+bqdN25JWTz1jbT82MHgomVpTugOnJyyFuAlgfqkjKEwUp8/NaO
6sYYfuUHUtP5LiGJ/wo2R4Cu0grU1NS0wkbs+d7J40JzWiALIKRAweFcLFWzczogxUT3XIKruxrb
u61qXWghonYT3+1LT+Hf61xgFVXAhn/LsMyy+h/R1YasTtKntPZTWzEp3ttwDcn9uFjF+tU44iSe
LE1D+mGNrPGvZZwGBHaqeguJT7EP8UlD1qgEG+Dq4uinv72064ZyrGdskL/vn7hIVS5cBW0efwbf
Z5w3h3jnAaEDs/PF7zjVwJNl4l1+u953t1y/sNJQ+d9/zjRbZu9mMkNK0C9+gRQiobNieAsR6Ged
0nqx2Z+0uaZYSZ6CMWmkUhQRfJdIWADqKzDEDRQkF6WZY8weudgQXhMpTPQXpMWJnvs1GBkkGKNu
qAAYIqIKlKUidZkyKF8uRUng/fz8rGqBxPJmXDFG5T2OSXPZ3xC3qY3rZxmaplbbShGYrHUYP8ao
ukr12nP8zL8q1Nn7KdmPUEgpnzYCde56qiJEgE3YomPGNwwKbfvWTfdrid7jlpYoa5ZDt2ImhBew
EcAy+PboqWLU8lbVFtb7gbhu2+yqtkItVBzlvB9U/f9sVhosWjIA///yiV0axN8YoE9uegYIkIpP
Onfzz4NAUgGDAPkwoWM9b/Hg3qKhlLFuitvJhYGLcbaYNs5WjjYJe3zh/P1ImHKM6bRU+XQ9m5/8
s907mvyhG7E5IEvC94g7+6ibMNCG05bivE84JzLb62xVrtfLnffxWi80YOnVMj15XJK2Dl9+FHlD
mn0+Q+noS0Nm9P/fP7MgcyRhH7pupLkPA8C6gjNPA+cv9ce3Vv0r4eFnAyM8g41VbSmB57CISrlz
VGvQCeoX5I2BVlCEewHk8SstyTdjTJguaSusegFHt6sJMG90pp9NkxcMCpSzi8dfBwFJ1+lXn1/V
+9XhUAsBIQJq/F3SxqL8QAE+ZttypBtdJx6eQJnp94N+mM4gF0VoaEALAhhsHU3FMkFJKdiAemip
uhTbXVfDS0HlzXidrpEKfrS5ZtWde76Ll09FoWib+Qh/yOOmdwt0Ym4hN9BL3kn+1N5cA8IEp4q4
RSiK9mVLwviB9KONVOxVMH4fMX5TW0AHfh651ha3Pt4pm8n5vmE22hJ0k1o0mtxx7cSvCtV1jUZB
HkpeU/uj1y/o2XHnxrvkKukTGyOtw807HQ36cBqTwnnHxAdo7VebaJVbur9VPFhwZBFywZ9gVrd2
dJe4nAciWIkio6QItu3J84y+k4dnJwpOvmwaiBn5Rl6Hz/T5ZQzv/lkI1kHrxFb85rQhLDIU4fK9
UFbMNBXV6Ee3v0UGuSnv4GNJ6g5wDu1tx8neQqbYG87ZlCI2Tr7NL0kkn01j+LgQtTlzWe5XlZ+N
Syy75gfJvInewU1e2oN0HyOtXTFnz5aYT00PgPlcUAwucyl56FEhYvZAmmTD90IdDcMK3w3uk4/3
GEgpMkO3GIzafUn4TF2mSZTWm41oHR6JlQRcGqoim6n+T9Er5TZk0drwFmOWh0AGzNxeP2yOf86W
iYErkmmHZVhfoXBYezAvawUh3g1Ts5WWijYM7Bq4P1Ty15ZO+rsWiLIrbVVTMdzEHANSgXV0j8S0
A4xffVl057T4HQlYG5AiTbbaDAvJUgtOeTFTulm1ajrklfQwDw6OzrKCkWr4ugy1LQd2KvWGPDLh
snXNbdHydXlu+Vc8QhJ4UrC1Iuwz34+7oFWziklI4pxxA8j9xTdOkPlzApDm0H59cvIsVPESCYnc
d1C1gQ9fynObbgE7bC7bju83WfrdeHbImjou3nSnTJ4FcneCuoc9W7caX0J2eHAzGgXNgBYOOIXH
nWqA3sYScT4LMjTbmYaAiKTNTUWYavgrFmi/eNgThUr4YltAn+nF4bxdGbfD8SXdQQ/mRfGc+ezA
2b+eA99ILrvqBFVUMth383iIuEx3B2SgCxBOb6/Y5hSDyv6o50IxUXpioxU5SOrqgwLDSK8hzlt5
N3oKCon+zUvQ1M9rgW1J6/ZNmD2/BZFAhM/yjGmFCtu2PrFOuiI894ZSSBZNfisRlE0JNmJjLWpn
hzwXq0dxgCxUWQuBCruh8KdDg0jbNGAE3p5nckaojLPO/Ww0Wa/GB/vzHTf7zjoThYOQpVKFuNYI
aznUqpBaqdmbqlNe8vQ6dA8tI9h0eYy54RqhLqPAYNvs4PpNkAaNIvDF4z0LkcgFi6h4WV9Y0mbx
xbH9fzBq0vBRB74RJajp1mT03RIu2yYa/4KKFQup5EY3njOEI7hwQoGG3qBETrumGLS/aH83mY2M
UEDGSdnb4L7/wVyKb5MFLtIs9RntqjtPUyUemyq2p5si+sNsK7pc56FQ8oZYprdpJ6u4erYkCVJX
iSBnnupNh00afQWOsvFb4FGIvXWuQCpbeVbhp4BU1zaAd57BVwJLHWVhU8lCEKtTynWDvTcAI3YA
/7SYq8vJKmprDW8XkwK8Gw6oFQQ4lf0cTmINbeHN5NHYxoy7F5ePgqiRREx3JP+Yq54a31pORIrz
1o8PgPdp1gXz4qqbnKooCuihcVg5XLh09y+URDoKIUJkSs+5XeadspUO9siEUfXgtV6Meecp5pHp
bpra4lytVZXDLwWUsNx0wPJ+DJa6/EunayUc03FhTKtOce/obfxlJzb0/+q1NbPQyjwrXPfrZWZU
tPmQ32aJyA+ebAizIKeeEm2VdEsT5+7SZ5S5brVgJoFdPUF4ZvH3PQ+PrbYpI7q17sQHYbk0wqI/
8AjVd1wyDp7HbVO2V3BhCl6aGW9gAKvIdj/s1kIb0DwxhloOd4K9j4lEOLQD+/4G/5HjQf3jvZVP
ls58JGOLWoFIvCKwp5N5U8YQhJDwrPFbXZmFGjYyBHoeCp77YfWxI4C+LQ83Gv8xgM7cFLQUouKl
XeqXXkDreyVrn/P2SDAkouyFy3evO5OVk5T8EQCFtESG5W0OQPv6HYp8hu50UbQIy99PnzBFcCCU
iFFl616r7x4C1RTx+Ia2XIKtZyxaQomPJ8VL2/SzDRHbHY4PkKf3C3At85+zs17RfpB/fg4r/xer
B/JIJ0fvEulvJmYgEphB8XCy+cBfqKuVgCZSYVT4SpALZmf4jSo06DbEhkhDgvSnF9QFZJzKM16+
b/GNZ/ijE8Ddm28M3SVs5Es+ZPcdEmS0bAi3R3prpGDuoq1QawbsAHC3ZSzwj9uTlI3BaQQu8w+A
j9TNNpx7vt6vYTyh39fcddDFLb7OEdSVeVX4Uss3heZkH3EXrDLNIZV74GKcnOdrEGp1gyArSg2y
s4HvRqI5g5Y5BKHubzP+qn9gCcQUH3+I25HpBHbwjmuCFt8DZqJs3RInVhatjimmGr3ORkGyYPgr
i3VifwqvwQN7K4UvJQaGehuN0We3ewfPLhyjQY59x0tx8p0amp/FFvtHLaOGVXznqwyiuIOHD/La
QyMGE1m1dnRWTVUeUE8cvmOX+B3ffGWZEDUnFY2okxVjI3vlfSPq1kdmAzihBokGreR/aApbD4Z5
EsuGi8+gFgKynHN2JPV8GnK+FC18cPBPj85STcidMs6kVD3UP8ULYIJ4aEZhXUkpLHH0P71fzFVV
mnGpVbrciCAYdpN2nYeG1ThW9uGRSuAJ2NpUX1NzxVkG6spoMwndkCZgo3G9qLzkmnUzKCX90Y4D
VmWFuV1/dWyeiUrNEhvqGvXaLtvaimEvBAOsJYBnTLdmvPe4pI7IlBe/oy35nqZqj/S1VHI4hvZ2
7GJ1D1MCm7/xmfW1fODUkhZGnHVA5SWieqo2m3+foFJuwqnNYtJYYXBg4J7rb3sEc+RqP1xbmsZI
9MbnQb5wA9AUfaLdZ7jR5W5cKCvTWOK9pCtT8vBNdenvsqXrNpAvfd9fg52dpqp11HRtFCVt1gGM
hpTVvt9WDM/jB7Udd/kQEfarOeuuAIP6Z7SlSYUBdDJuS/tBXplZF5oyQuhabeQ2aWieGY1DNMzD
j367yc0KlPp79fRlRR5qIMUEtP73ZBfjqFHFTCs0qohtu+rb1wzE1fE9kq1NpvxO3iFMk5xT/ULe
XpegOh5cy9pUHTkN6ajbQkioB1et9MDShj9C+kflAS6+x9pCDbzZLGGWJaZw32wtcdtdDfYtD22j
E5M+pIv1cdjHSmi9WJgZlBrEt+5VmSWQ6Q4pjxzISbt7pdYfdKK+ed3NJjVVnmt8kQepG6IwGsT4
HmFbq+N3QLKqkzexL1ldMh3qnNfE26aF3JXmmoF3MkgvREiJKnQGyrdVhlS6APLfuA/L2GzV+Mag
tU6Ev7QNmXgXg3mzAnE4x6Jgu/mJDv8LimKuZvkSy1+q3wq+z8qePGsKfRS26dD/nhxRorDTLQkx
y2h+UFY5fQNx2Z1aJ8ZMDxsAZ245g4/7HhGyIwOSoB9YMdJfopyxK6q0OU5RvUw+o6CBvjFpwLHn
Y/pzOSvqAY62oxyzbqct3HqvPuz/XKRstGBwcUXKajc1saUCNG2s3XcY94Zm/OnQ8d/IgWG+hWr0
hRYD7wnsSrltZbGoizh1/OmVg1q+KTPJE/ySeCSV7yBOB1aYaV4S+2oQgHuFJuAgMH5LDKWyyJ2S
mWpUdAI01Nk5OcrUxUNLCQbNFPZUDRFSXPEAnurEp1ckrFr1Z+JfrsjDgoNQkKBH/wDLnQdF8tmP
8CauoykmKlaay9IgkFh88lBWVZpQ0u5im6jgpfRq2QzZEaOxCNEU8tpvHnyFPM6WFBabRxeXk0Ab
6ErupAcUX8ZkDnazRe5OHZH3X97XyL+HgcaHd7QQAblue/RYfw1GPbW2Onw0L/2uE/1g7RFZRM66
ntebW2Rq7DvZ6c+FACCmlL+R60Dd5VYIRdale8JXckqki2UVY3NDfz+iFiiED9/nND8TYVK0ODkz
XprSRj1YwheeBqrWpSASgftWwIXitdlBrIgzi0eHFFx0+5evsMi/rkwsdnb1aSJDGUfYIU7EZJpI
/3oZjTvS9e2HJmqXiEmOSTVMkL5mv3L+eodyg6mBgnmCyX521flFhgl53OR2xwMAMAfk19AW0j6y
rSZAgKgMpXWq5qA2WqC+yFOuW+s7wF7zhID2srro6WtqdtF2tQciJc3MhyPBaBzyNSquGkdv352b
OvvPi2K3QYqqfbCvs337kMNkJj/jOKq6kM0LHREg+IMxuXZ5xdv5nE+E/tD0g1yy5gFDsoGC2rD5
AH/Nmt2IUWRbcm1jhQ5QaR8ywKUIHBk92dE9kN2AvRAGEx9nWGKW/lKTiA8A86Ngzy6qwlJGT4vW
ZAe5/oGNsUX+XsKfv8iOXJLqcSvWNo6lLuO6GO4HnlazgZRXjFr/Vmr9RV3PCqnJy0NTbO4ClJF8
QkjV/w7yIZeuJbxuiXMsEZldn4kAJGYDDb45Rq4T/0eSMxSdMbVRFhu60bbcHtqDlpNjHbXLECTx
oHUwBokcIPT7TVSMhwZSPLA68xTYjFSQesoGcm1Nf9R7vTPsun61f9nxALxhQt1gDhJLAFtvK11B
1AjnVjoQYYgYq9yxpwDJ9o/hbsR/wgIe2jHgiwikmL0rWnbiMRjp4jGpji08T1BL8wrHPynbZlGA
7j98seYtedLzAJNtnoDOZBTKjkyaTpd54Eh5wy1oFslVBcTYnCW70PAAQG74mZ2pmlVlTml6byKA
iWCbfFCySlVk2c64xCbeZmygQc9ZXXvyHVcIU2xU+WPfAgVOWEQpeOMHHHyomNqN6m1cvSKReEhW
XjOZMssKe6hEuUa7yOORM+84FI3Akz6F+7GoJCWQV+AlPgfM8jsueEnj+VTf+7DnqUnSLNkAtbaK
FApV1/TF44QPRMzWtVqTNCXEjLtNjMeqGCCdRX6ISRu4xsOGu9MVbfoHa0Ajb0YJTLNRl4WRBctI
8hvu+Xu5Wodw4EPXhdPJJmoFydgrJwk3kNKMsycjhBQXcWoC6jF2tLF2/tDegm7MtCaSuL1pRk9h
a1hFAD8JTI6koLFo+DqixnjkfEopan+vchxWSiKiVXmmYZxHP/ptSWev0MRAE4GkJubkPnwRJeTw
aVUaoirgxf1197TL4HU9Db5trQNB85edoOsk8t5h9ddeY/WSYFZfSa94Z1lzAps1b5PKHi7w22Ll
qcg7d8GMTfKDdSK1giSa8eQ55JpLNN5tOWeOzxE2OiU40SSQlZJGe26znicr0T/TZQf4PKNZG4nN
yDUOXOW9RIn7VU7Gli5U1/8dMV1pF2ZqYr9at3xJUngUnYbC22H+Veh3i4xBDeNnXxnB7wx4/cEk
ebUNNcvpC+HcIsPB31NX85edsCNRxwYHJqUok1nnQxifkZPgUcY1l8KuaOZOACF8dS2MRX5OJTuF
22POS8Dh/1RIpn90nKFvW/YVuFUDsz+Wn/GHLWT0TyaYzXNY/+txk3SKnFeWJqH0vWSlBOC7GCb5
m9+iudCaQsHEZ6g/Kv/s2auHqUZhpaDpM/CJ0UDY/rA7Gu3Xdvgj3DeIZyc2a8N9zDK5QZLIleLw
SrbqcKQIzFI9NYKzj3VHUX4+mLt0A9xqtG4I83z8w/1Vl1UhIkv9bB8VTSSPvk3VdLCyHWedNk4h
9dvHKMgmKBOmOEr7zAXgLkQcS/Hwvh82dmJjlSrt9e4A3kRVtbtpPRnU8gMIJrifO51To1Ivtq5p
LcLrtsnLxhbeAUqHKLXbrxmkSdpTGR/W4UepsJGX+JjbVyK8ggXmpNs6Bsl8hehHstExe9ZTOA7o
McY6xOiLBH91IYV344K3se98JPkgve2jUYoX84cNeFTiNsqet2d3Teg7A+jYMkt1C6IxjXQibVCl
nQFBDNrXBBh356/IDlovX2iNfnvS3jfIOXAQhQMvCsPjJEN+/ybopjfowi/cliIasZK5W/DQjUWr
iGQ8qeSEXcGmSGuPp9gHfh9iwYWpbbOb9pz2KvmkFYCGEoFrsKaiE56hCWUkfPCiqz+4AxgLtH3i
w9P8BMKhEiyzi1sMp77Us4ekuO5gtRXFgmgtVWtjFZSyg/JL5UonRaKWhMwwklXAtaKJiPeCol3q
nHjlpNu5l9LzFKAfcgYYfWkY+ZU9ZSNmJt+iIoFIZQzvcr9kz88wMnCn3bAyJ/GwTo/ptaQ1i5C1
o1UrvNx5LPE/W0I5XYov2ryavC9fF1g5Nd4iC7XqjfZuyX6kC3be/RitBqRJTDcba0w3NOnH84vZ
T9jTCZRcUhrCtJO37YokdIWMG1j3Tv5gCsRTCY3swdezBx7NF5smDDPIgEMuRTlv5GtL6eVHHKR4
A1x5rPg8Ikq0byrPYJfBYgyS5t4nuCvNUApi/tqEkgoqELjo8U75nkkprvn94Ey6yHtgr5JKGJMm
JMrVEKvOC7279OBa0MEBKX0e3/l32pwj5PtbNlyPi05/bDerWNeKJwLq4pWpYs7TUypmnkSMGiII
PyRHtvstADpXo2yTychLragQ+zfT3OXESEEHgm40E3IXF2xjSgyXCxeKndV5qEeJQkGmj8bBfHpW
lwA4lGwpadeECWpmNiXvrPznBgDTGCp19hc8fgIjVcIUlCPfTvwBpkFqY+25NNZm9nWxPh4XH2dO
IO/D5ov37L4z530+lH5LgALobzmvM8evgZeAP1R1J0/kvArPXUXsB6CtLa+SOLJQyoeDrZ0m6Fm+
yZHnO0FaqvqfLZNTrBt1eLKa+9Cq168a+NL7IJEHgkQ6gWLZApq4F0iV97YgsLDbbKZjpwjC80qQ
TXeV7ExvBfJg0Z8pyDOGNWGVCi5202UQMat+9NSf6dO5MeVwFcKkx2pttbVN6rAyCLpJ5lGWFNPR
Js56PHemvasyF6PLWdPZe2brjDikwGDUtmderWv3iAtgP75QJPBPfYhL7kVaj5YQyJU/GoJRMsee
1XmJ+AawT2ezjo6qLKMJxCz2BK7UStt5dh/VFH5UYMHKZqod0NQR2oK6d5KChbh+RkX0ltdEf9y0
rlzINLeOJO4++shVYeL17y3jRWnFkVO5ujdnLp0wIOgGS0iG2/+JNOg7EJfAfJuCTzYbZwwBE51z
Q83DLx9NHFIGFVNVlrmBisuMc6LpTZryRMQkber4wN2qVSBtGdtR/r+fyci0xgqYgKnru5UfpO5S
P/SjFHRqiqXhXf4S5QHWN2ZEsbKJV0Tc+T3vn7hNxzIq1QjcNiW+pgFdP+l+Xa6p42tuNJ1BUJwt
QTsJaNDAvJI2NstAosw7duyP923LarN3RzXa2Ebk6TbjyUPBA4yALUafJjXRCr9eq/QiTNzskqqH
cJOd0PL26MD5oPpiOL8feLmdzbFIQGnanPq9Q7UpBEAbnaNygoleHator5Vs3zlLnxOhV+iUn2G1
hAgyjt/s9xmLpc4qFn+KFVvQLd6wCUIoCosyHI8mhaB7fiSTZaXsszoUrsJ5RNO7XuxIVDjARypr
ZEc2WIrTNxqM6OD+zasEMVMaspblhSAA9m+Ip1CiQpdR7l1P8AsmbvkFMMKHg8wUPvZUkLfIKAJY
XZjE2KaBQ+m/pjZPbl3Ghc+pNyib0ft0Ve656gzzA2+1kvm45+sjtguJ9+TAHl52CikBTNUXR2Ky
hMGA0vqi8cvm9zEVYwO4veMFcK53J1+8YnZVBGbLXhnFp58X+sq1R9awxwH3wAcro8nRLi7iSRTd
puDTXyhbp/AW1Aqh8hxNE6SFoP6uZBe3Bw2r1x7wZXUfji5wB81m+eYM1jD+KHKaE7gsIWaLYiDy
hiczyhkDXwuz4XUFNIR4nDcCohPNgOY+7oy6p8Hm9sOvKSXJWJg/6GL3dBBFB20bTz4zoUli1o+R
MXNJTyL22XmIuRjSqhFp47N0yK5cCPdwRMOkAjT7aS5kmtR1KqAuUVUPfRyX5MMjJ+fxlezIyaD6
VtF20kNBCFqBKiUS06jUvJEDCHN5Jn8XFS16kS7N2ybqYhTE2tZSflXsq2xiDakAyU01CN5DZycR
lPZ/G2/oYYgWCH+QRcLECLmhc4uLJZ2J9avibLE9m3A4W08wblSi5w1V6OEXwTF2VPs5/dwjT34D
sWIHCxymZ71PVlysSQLMSHX91UNywFxkltD/CQDEcKUZK20Pfdcps/+am0+Sk5bgQBlZGeIme17j
zseInic9ZWp59gogJzPBoh02RixyLJqrw27bROp1ahEwnTngLtcxlJYCWiHQn2YyTCNoDx9wk3fN
n8dfCOH0DAICs4pQWgWcMpVx1+3envwxKEpnQ/nioB0DchtDV8caO4nLCZ42asQXVzj/dR7hN5Th
JnCoxt7fVhZWhPdtrstlYycB3UCTtSrW19BkNS/cnWHWTdDwzR4uk8eqwNphCJDw5a8VAMahS+9U
wPwut/4JuyUDsqB72CjJRKvOOR8oRSQhytykqgZmSGKvj99zSr6U2sQYhSbm8h272AViJ50+OtL3
2b4et3XPNBb05NhxaVG84zWN83IqxIA4fMnkId9Fk37G8GaYHNeBkS4Fza8AKV4zpXsBS+rG2lUY
fsDTNEesiuscaXQb3u3l9Q9mgAQbWebot4RrE8FmF+df3OaJJ/jFTu7UEd4aV2sfzVYTDSBvc4bk
1HiFNwNRn9UaYwN50rCb12jR1fWX35OloE2RuImsGxhHYUmMWB9XalDb/JCtAqOZfGnuycti5ckQ
f2c8ejR8n2HPMmYZbLpO3wqS+qGueypEMNqErpa3wIXKOVQ1WGh2HcK4KWaCYfb8IZpkBwVyMbRT
Jgdqp5GQxqS3V/SK8y+oaiEjGPzABejonZ9ZFPRqxyA8SMFaQHnor+o9DfLvwuYWrE8lZcG4yYHZ
zAUjAkCb9RH7EmtIbtXcRncos/fwfGs7V0NnT5+w8UPRzeuciMBxYc/Osez/EdqfFxaWMvcr/35v
0jposDJtXYKyvoW/6RI4KwZMTjTN5/DQ+pp213c0f0aQf7rPf3cRZs/JBxl5Yfoe4wXjl48jV0SH
tTsrUQ4CDBBuDovEbLBfSSVIO74mrmI0cbtNW1Nbb6NQg7x1/NRlm4Fnen2huNkzqEG6+kpKwMTD
KM61YOY6POexEBE0DG1SV7USrgDDNa/ZJ5SZ6/68dpl0n2ueXWoJGYv+HL/J7RGCDIKbBpXd6kxx
gQdlBRhIaswNr1+ADDEwFhG8CpYmy2zAfgw6EMyZ1pyHIprqmbL1P5fEOHzLU7FAaiAQYw1HJNyU
H2qMkySbdJ0qOxwIwyvtZq9JNlOWRtZVq4c/uE3B0DbNCTr4N/Ei3b5hUd7yTEE/61GoFe/4lm+9
pPpU3vns0BpO0JQEaA1fh3w+r9oM2u/PT698tkxyK53qXi6o4Cgk4uJSprAyqM8JG8UPQxN9/+/b
vF5NIYomzqylwpFnAjWTCkEL+BH2Rw9kCX34sPlevJgtnFhw3onzUWFpvthdO4vm0HelDHj04XCW
mGsj9K5ja8icUz6LwK1LnoejhR8bwQtNqBKWjtD2VyT1QwmxLrf207jeMLb1a71hh4bLOMrZWeA5
S6BYnStuUXwDFa8f2yytJHxJIPCYgQXMHPrxfSFghVQPz7ottz6PfP/CleBnqfbhJynNTaSO0ZfX
nVDQR3NfmjCF+hFDaTu/kckiSLfY5qmzOKCcfhi+luEuMYRZ6kBTNHor/uACZdXFp7mer4WlJPlA
oRDIpnM1958UUfSyJt/L9cDNTPx5AzqcTADdoeCGLQ+PSYeOJHS0IDJISkLInYlF8A5wkfkY4dw8
FThGZGM8NoceXXvEN2aLireu0edEST84bzkWyLnjkwxYgI2SLrq6wIylbkQhFkv7wA5/lCdPwSdq
z0z+gqvjfdZyRWyhOMfBq2K9XONoG+DTx4Qu+fWEPqkd3PFs6jKwYB6XZN0sMeU7ng1JYkL13T6G
ZQgT+/8+SXCjpgg+zuA0zef/khTIROONT2tU1BqJdFRmLIp7QE9yS/UCI/MgsTA7QVns1qoGgKlI
FmTquoaUH5EX7m87thesGtvK7tL48pdyprPMFn9kkZgl9WN5qqWeg1AMQdGayGhMXFyV3fZf+mVH
HqJoc/rlyq1QNwMUJCJBCkPC7ZMCd79uNOhxPjjNReCBlOcy7hi2pI16TOuy6H+DyDT9222IYlCP
lPVuOyF1BLy9IvsiyjVoMbxUalhk0BCjPVQ5w+bG1ThnUhQ2KCus+gl2RA/L0gQQZe2p0g+pFqz+
CDApq4o2xkYmizIfgZHnLHbOs993DU7Mj7fWg+6WB+9bqKbdG+PXvf+cF6KxdHrcalFdKBM9+wo5
/2CucZQNs+HFXqlXfDMiAuISg1qyxGHq1y9g3boTGzqROJ+jRcBsfrSN+diK1FColI7rq5lp5LDs
GQho1bPY68+CW9SXnXvgBEk2T2y/AwbxZ62hFvw0t2nsQFlEWj44d2dEwNYn499Ejs1WtjOE2Pvb
SRc4XqOWO9MNOjPtQOB7SoP/myIlSRi68i5dSZsjj9u6TDI7nSucCaGXo64ep62jtxJIZ83RNdPP
CXxz0Q1fSQ1y/7ljM92BUaUJVa7I06MlcuGnaPs9rDfRkAqHKDEnyWPIXc4P9F44WH0/JTzGeAWT
Ka7gY4ILgKGmUdNB6eYEjWStrqLj0djdDp2TPoaArMjgtwJHWKARX97g/JQvA+o2s6tSBbGCcwMA
Zu/0CYvZYcuMu0UBstqg42pJ4+bX3PYvxU54yflrFmgEoyRbECIZiY2GsdOV/D3s5Cwi1TxQd/4E
sr3X9WlFlQVsf/f0pgeSLg14akqhfkfT55MPTjEXQ4UfV9Zo7WjW7P2fw84pJ+gh1TK5j8xNiCrA
fPjGhAMadoSKnIjj1O16Yfv2DNkN7gcakTJ6FjhWJFudSJ8axvRBbcmGrAERFcyFlOjUlRvZJFTg
xROq+glR08i6/AZOiypAZsbjSg/YpX0SeU4eIODZeM9bFqJ5w7lNjfjSKzLy7RTSxbpsi/ArQqBM
2CLNegR834C3cMM/7XxWnA5DIDoQu4cMJO5Xlj2fXMpHDowAGASJtsD7Bt49rfCtNUwEDA5AG4A3
az+7viJLhM8xdvM/KpzlWlyaaFqpQIiLLmd3uVQPT8UcH1NEtDaB3rVJcsQDG7FrxzJhN41W55sp
EQb1rmMUJXe5G7/7dJoUnbIL9zgLlOoMf2VmfkO2ewD+5Ds4a+2zp3xQV6vMyBjBPALJ++yissnk
Uk0i9moD11oXA/jM/25hEbuywBLkw60YeeSBOvi4iFEk6bxL1TUFD+aIQvJqSirDSkx6TXfbnRwM
jYlHZjn7gzW+UmRYXjDBAcWcr5pvZHcT8b8F3kIodJIePQZunH9gBmvgLP2Lhe3+LdMYm04znJc8
57AK5jYuqF/S1ZzCRJLdZk4xPgQOSSRPDdHMpzVv2clQb79e/7VN5e3FHJzMi2lEIPJ2zP1skK5Q
XqU8sm5CX2hFjFEsHXfFt16LtQNsaCIkFwUpkyfSeFit6B+bY/fipo3AsezpPXx6+9J/2DTYiK/z
+4BfcMPUETJJMn9AfwakszoyAQbI5LE6fATwU7p0cG2+uY0Uecqt4u+kssP7n2lRvMFS5xq9gRlB
t/XvjgUD5Wzv2Auhw7b2gGhShKS5Lh0m4An5h4EJbGyt1MW5aWp1hczJVVoS7bX1juHDhryXaufN
Fa7Z0ngJNRZ75C0pDe7BHyRaMfeE0Mr+NQdCZNK2MAAprhAenYaTqSsEKmLBcTUZxcsFAahl6L1/
T6Y1oNdrgs+29QJI4d2U42mSKUvKiYLND6yCm6pyiPQ9VQvNkVwt+vYnJp5+TTKLJQGe6+LE5aHu
ISLodZSojEE0LAQS0hGZyvOJcZOa+EBUY+K41KbOSpwjIm1zW914LH8wj6N97L9sFkHTKNG2Z1CN
Jdkl+USxaXkasndX/UAG/R8UV0d5d3weOroqJmMd2xupZGfnuWcm7wNnOdWe9AJA/1ZIPpgNv0MC
zbjFv6PPAgoSdL7UEBUZraQMALNCbOZ3AJaTq8mAR6QEX+mu/SaL9U7NgMjbnchqKOnnhKpr0/FB
lKAWt+8hWlE1Sb6kVxDGqxmfqZfcSzMi4fhS0+3FvMZRL07SBFiWNbmWVB+ODSfNXNy6zo2lfGxV
oQ/nGrZjsvDpCgHsAYXaCBJls/DLFstome5LkMKP1+Shz6VAF86r7J+oHRVQiaKIJIlvGYWK66Lu
qaPoEthKAeIKblymaiMjvhQIAamGggSCTDC1RLB0hQGHdYCttkv74KmuT4Qz3cTVCEz/6REbX2tq
oM2wFwINUegFBiwwfrf02Vjdflobz+FudYZrzhMlq9x6IQ9m6eWeXQyhw5E+t/AMCJ5JMe+mHpbx
xV7Dte2QX1Jx3SySU08bUF0xjZkKXAIN2y4USN2aC9KbqRgJs+zzrHlaxw5u2XqPp7w+ix+Cnt4T
gRaW/+Zypsh9zXGkRmhwuGZqWDUCrpz0QbFDxy7bQZVDuQjkhfReW9oE7X69pT9ehxp/ApRU4Y+a
qHDGM7ubnlmFc67AH81vSj12yy/wGHvyIMykyWW1K5Ux612VcrMKlfpHeTm1tiBrxqOxSybsQ6uI
G/ZTzMI+aPEXt7HyoMK95obp8QP6AELvkI0AALjovda34we28Oc/67TNZ1cUAnuNmlEGizd4XeXR
FJJDE+reEftvLRFDWRmNARbxN7lR5sNKEsdOkts9wqyMC/MkQX5wQBBMWMK3ZAgYXY+5M1nzwby6
Nt7KzN1YBCJLbSWACLbfE67I3heQJ3/hbnrYXhJrAJ33z73bFd0g8cYAx6VSrwGMoTVKrTwckmKd
plcuVDeAHOEeGeM6PuR5RUIQMlsU1qD+8H9FbimjsYEklVVIlXzB8QoNml9linPqCSYHjmslU/S+
/o4mqjhPq3o0Iqom3gd0/++VkN9we3Yn+4K4um+9jGzjCHI7TNKhI9n/JSnKBBTU3f+n3BhyHUYU
+g7OJHLpMZAxQ9rDjA4UI/To+VvlerzGRkNXHuw7gMDQsKZ0N0odYGcd/HrkqXiDo5eBE4vcDhRb
JF1Oiht+qBOL9L1QJIq/ZhP0RcD8ObX1ZpDbktb5sGRG5oOFtS9dBqFpLNA9xrHTLXB6C3aabLhW
yAMeJ19iKFG7wfnFxxXahYx3SXIepgpY8coWwXgl9btiZjZ96Gdns0P5K1Yl33eEb9loh8RWGZ5l
xUzkl9TqWj7fsYNHv9YaZQrsJqYtQ4CVOuUTh8PCdD5ctonyf8rKxfwKhLnpG9vgTSdrlvBdD67L
QnUONxxVs4M6E/sngcrJISs5kQRwRS+Y0Jlekts63kVC45wcb9fogG1oc+mZ8yzNby7L0ax4srQk
fO7GNErbrtw8hR+McbViWLOm70CWd35sxeRK8z4YwVeEvhL6Zdx4Ht/5Ca2WH59inwkes60s8eaB
MSzyRz7v27vRw81PYBbSzqLgVZIYGw5Ks86zPP1fECzUvDu6fLfPGE/Q3EBFTWdjAsQSGUNh3xvs
P5NzjjsVaWh2wiVjJN1131HGVI/ySUTpUEnTjOanR5RIyC+vlCQs2TM6C/x44B3ISsU4CR7xTKiv
4prS9ub0aKjF1V3wqvzkLUfBEBfH9jF1+jKdQOuNcY7svbJydkVY+fkwp3pmXwdjo5/yvooGLmeT
IytWu2FizMOB5J6DqhOnt3gWJPYdID3EpC/WXLigX1ykXoJdGKI6so1pXRe6qzB0sBx701EObIuL
w/ocBjmRVlHdUpfoJJGWmEVd1vUMBZHuTmGNBcEI8A5XfGpeqfnBkRmnnDID2+h49fW9KvFFYxap
Y1T9c64fLwOlxKOvN5ujk4W0WPHPeiMn//LkzgmRP7PoRlkXfOJBRvCpA+omSlOt0qc1iinNAK1M
2kbbmAB07xScaCBJ7oSUDLOldPa/+aVSZsvcmJXZu3+WdZ3H5SP0yDyqn2vH+ZRO7fZcdkn2MZdF
YE7nSbKwVSetPaTJFddRUrmk27XShASv+9affwe+CANKYCyL3Cf7xPIfVxMyAoobkNGsUVpYYiwv
NO5vjVkzblDY48R8GrkOdZeFXAhDtzch0VYB2girjmc5U3hO3xyARcDitzYGGZpzFJUXqk4Xd9oB
3w+yYdpiCh20qFZEAsbGzaXgo7eNERQDb265bs8UbiWAyJo2XuZnuMh+hGL0IUVa3+T1A6/ZeH5X
KAsmprZObp+DbuTiiBPcXChQ8NvGPcPom6ZoTFV8dl78EtuUwuAp9muic/LF8QeGaRK0JrBBqzrz
TUdAb67z4FjgX4frz+DQL1vMVRhwG0+LERxgTv3BxOcJDmQh1FWaWfOfTNQ8Z67gc5XKKtdagoT/
hDoNdkq7+Ke4P8NdBAQHntAOS6+oRy5qkZPXO4CXIeFDitJfpBx1OHfDHHazcq9HlXxbQ9IA/hgM
VhyB2HRLeWgD/daOrEHAAt2z81vvFEdo3BXP+Y3qsmY3fhdUeApmXpCod9koYP93p/MrMXktQbyO
UobK0y2VwFgWSVqo4IvqWWi2AAsmsB3hIHxnSpsTwKltF5EnKpGNDDur1hMFQruS0RUNfKA1jT78
1XKX510AcnLMpG/GIh4KrXkmaCaiL+FMOccdMU900LlxVnfwNIARPvo7ogYMEu/hVSuycYvfTx+g
DXBe/apLgdvhBunCY98RfLA9Y+ft0R+5PBSLCaUyAj2q00dHAWujeajrYhK6uCYVS+bBMSe3hMb+
/i2HLrHSbOzu5OW+4e3mGm5bUbvEq6RrVM7QPnjbVPrN/9anzo2J6xhgcsY/gqvC/LcglF3L4mDJ
qdit4u69tqeEUhFZb99q2dDeYl6vaiFNG9EkRhH6n8TxSvWJ+0QwoSkKlnJ2Qu7h91Gi6PNxsiEA
lsUQs9nfJMhiP2wu4WEYDlfmbO3YTTpgksCYhtAGVCYT+wvO+iSFR2g5ORBjgmofUddahgx9X1Hu
LlnRVzCxzNX1jxm7iSUWQd/c3wQt7kX4Dvrfm7OUBfxejzJGj9Zp0emh7Yxfvzy0WZncHprR4nuw
k2S6WFDxkpV/uwdc/2Y5WVUVoiQbJkHWwTv3zXWyCLDL2BDWSz2oejtfLYIG9yb918uhA+k2LYGM
0+wn7t7sCLXtWOLgjBZAL1engM7/B/J9C7ZGXFEAIOEmJAFNJgTI3qYkLq8UgRojc/VLEwEa7w4z
BW+7m94tQ01866i7Q+Oxyqois3LYQijd5MvPa/kHOqa4jFe1+S5X6V+kJIqnQuClYcDw7PJQW3Rx
b1kP9EAyz3xzBj8SLxtyXqbHqNXQ7nFgJ/caoMy9UhfAtatImpf2rOJQgWdEZptdjHL91e0Ni22k
nt/R5+4AhleKX6LhGfsSidBoriTJ1PeyXFUE9/yb51RwMoQg2fiE1ajZ2VgBX72i8xBuXo4cOYhD
o3ljyO2AQYWej15wcLxqI8kAfjlKhxulTnzhzvWcxQGs/odYSpHVPP2/1NfRyLnPscMy7R+iSOc3
nkJNBppyoPABgA97pWoTd6oAidLCzFMzvXCWsKxcBhx01VV+XckXdJfezdoBID3NLCrmdRjIsU+B
rU5U6bFFE1B3XN0xXBrdT6yENE2U+JfIwRXZ/sk5VPs1e23c7b06zwos+XawRBfvxkoEfU2LrLc+
Y3KRGsRCNfLzcBg0Yx5j4Ve+LS/clMsI8qwo5QiIP4F2Q6lqQ1YMXHlighYXMnhjdb0ke0eijXqk
JxOPkylt1zUO90iDk6KUctLEx9Pbi47ZkzBFdfUkJ+WwRwnyQzqBqW1aCJFbcGgzF7BqYnnYqXS+
ghyaiPzEdKgDgkJ4bxE4q0TZdwxU7wGcCrUOWQCp3SW5S8ojnPsICAEaUCYVfwSKkC0N0Qy9oiKI
TeqwHx05Nd8P/YBM7VmSvcwjzgfJrD/YaUQPneO8Jjw9AAoJZKTpSp/jMgQHYdabY6a6/2Mn6zGu
YqxtYryHpwdB/t8XpKu2b+m1UlgOMagj5sVYVKPTXf4NFDEoOwupRAbVddAMaOofIscBUshC5ppX
Bv0AyCGVDdsBA81A+iOs3M9pOcxnn8FhGi2VXfoc1uIwhvCFj3208Spqg6BQhZtpJUvYMMD7l/kE
rsviPFvU9vTf9ZMoqvBkmkw1TQbP7kqDiP202b5jdu6xPYfEohQpU8W/tPRSJQnum/lnFGyIROKy
O99lwF1ZX8CKbqvfiZwORBnQyKYq4CCI0JqkmDp51NsPTeiQ8MJC7mfmd6M58o6MPrHcNeCiA+/K
LBp6bpnObdQkotUF+84ZGYIpgdPmkDDn8p17O+1uQRwoVtpqpkkuxXzsYlJAUYa/uqwS3uTN4SyG
vYMGfAhXeCWcfUrJ7wBjpmzjBRpLxlDKf/EaXWVzMGBODIRA66Jpdvb2JEAR+H4D7QwBKvCkax4R
yRd9xJm/HFMLcA5RmNwA0iHH7sEPoHvw2W08x8gnt55vOA3yWZAAY91wns9eHBJTsu8SSWoJjAzT
H0zT3G6khDdZrlnJkLkbJZM00R+iD+gjqMCthMpE/DD7/ntEiGkByxE65e4XuTxOM8fRjmlQCc9Z
uyKj56gydol759g2wRQCIQf/aWCW+wrb0To27pevLMEX8t2u6YPQUIgNnhhFpZzzoIkzFtVlPXR+
kS3QLv9WkAkZsT0DTEeVfbx/zUQv2AZhujqDBmkM30rsREVIyn/8ZeOCNiBqc7juY8VXnjHiJaI3
41Q5+frf31SC2aBWo3rh/tJGaVLfKLBMnUrygBp1DsG9UAPBVI5ty689ZKN2ffKDtdXdOHgJsvGY
Z+mDA/MsKBi3mA7mMAIrpVP26c0HjbcyWbm5TwOI+tj0jG0xTGeMAIUedDUnBEjjyeuIKu+B/Xqq
V4Gtx/iYkI4EnRP/v2oy15AbZeaSbFZDFn2YsGqUE8boJ14Z7igsdmZ3g72kAP5UErmAGLa1w60W
qclnubD1wbVypJIHXw8yM8XcSjMqrU+c7/d1Mb/LZOmwdHlkZj0HLjXLA2l8KgnHH6nP2qpSKFQS
nK0N7LlqzlJswQh0fjllk10ZwCxojq1z+HPv3KcvAvnwFtiuMF2MH9QcaZdnNtY3SHzNHbxE/GCO
r72Ev0pa77xzcjnbKRmymjI+4UwlHq0lqh5Lf60/J2Xx+bn5RAoF8ClOKhlUczH60FV2JdQ7g1x+
4wqa2kd2TtWj9MnQP8pBd6xTWoU/hExXkDE9+BpMwJ5HJfkSdkp2rC39I2iJk9CNNAkgf1sdEEg5
OUslT5iGfENsWIHLyRun4bd3PqpXagocdqApJkiIuz8X5xCo5v62oyOwYeekLLMI3bL2zGWjFGi5
pxHhJ/WpjP9Ywq517aYhhEidhK1zfQ7QJUQRe41VfaK2RDa9goP2ZBrOY3cXGO/8cIQy+9y5okoT
axjkHIvzMcc0F2inYUrDaRxkycZiJ3ILi/U34o22M4186SCDj9yiYPnWcRksDt1e0oNdXIstbXxt
PyNuQQRr8Ikuq4TkHB+gAgV5ZHtvR8arKWoljNoDKL4t815e0FkRrtOseUBaJa683VfderFe18ep
PjxaTD2nVNa2V1VANv5mMAQt/chbzgewjHfIZUePH34sSA8m7dG52vMg8LLDIt1HzCt90HG7KyLl
6yZhSKi8uenM/bz0sJvcAyTV3a9gEFj7UrGtcI/tGFzUZVWfVo02sy/c/8I4vD4KYKKxVZ4sbcTA
48vs9RNm3FYoiHqWfhWxEE0NgxE7t2hsmYjBCCIKhHjV8ys3MNtZa4klAzA7a3914veiU0qty2Nh
jEv1fnwLREFvC2s4hnq6yOJG+FpfqzWyeyrnMQLZO5RKqdxQ61ifDAtmBj4IQ0I4hR2aS4mhLmBz
1rDCjhjsNTG//4hheK2RNZsfufgUOzdiToEh3myEJKipQpKbLi+fLwvN+c8YRgFz5w4EPKpO2DUH
jUF2/bSWC7VtWfIENs38MIt7/NvTVdXbLuk7zXiXDEUv2m9/7svzIaco+VJ0p8cHAJEO8rqcp3xN
BmtmmbE4Z2SK/Hw4U/S7AIg6sGKk8FchwQvrOO0lgLc3uafcwMFR8muYyuWgDw/7gFtUKpfmlWCu
fByU09T1eMPMBHYvDQHNQxFV4LBLKteQ5PL2HP++Cvwbql5On15hrC7zxZTeMxnT5Bke3LkUdIVN
vOZr0KcN2N7+t3SvzHMjPd4n+4ZPHRHvMvPi9OD/TFyGe8nZyyfU3SSNEzbUjFfvrTJVi4iRpOWA
SfLPjm/A40xy9dLIVmcdOYyds4jx9KHT7hFrMjXCshQsS16s5K4UgqnPyjiEmAwDpBTJ4/5e5Z7E
iAgYxjLDuMcqcdSHbobjJilANBGgtLJXANZ5H1ioOfbl9UcjKso4I8qZGx2j5F+ug+gG75naQUkJ
dPSWm9Q0O2k3sRcJU5kvgh6HSg14sVTjgfjhyNKxhThOb38JlpryYPEIEdiaKk+1Mns8znv8WA0G
8EgU5BlHxAyqW9rEQP06NfTx9OESm7vFjiFGL5kHPxWSukjfSichUK+32yszUZdTrlWx9WiJxPt5
xZ/Io/NrXFEBFL3n8IZmbgqH9UiV/gEClQXXgK1m6tWZtAG4/+7vuaGUdph+yC+97RLey5vGohPp
g9ufoRKq0nUbJ07PciuKZ9dgzN4JGjqN2Ze7Ly4MCfsahLsKqauuDzmYUNc/qtCA5jjDJlznVWLB
ZPXyIsAvY5+ui5dNbWvF++ymNHOHx/wkRYRi2pXCwMStwFEr4HloFCkeuxZqi4Cv+/a13Zk5ep7Q
LKiidYxj2FZf9L9PBh+3SCmdUobtb1rxvk9ls6o5VSUVTWmi/dAB8kUMdy4aXllzXoEvyX+Xk5Xb
NWI9WNl2bn9gNg1iRl+fXwQAGRlpNMb/5Ntb68uASTGXcde3ajgEID+ksixBRYcVNhjr9WxEETR8
5tlF++R8xxRPd+ELSUIrE8uRgBCLhLg/GLoSLt75d546Hosohw0fKB/YSLibvHR4abxynCA0J0XI
ydGvC/fYOq69kNmSa/nGvQ67g8LcA72Puz9QFO9+bFDF2FbSq1KSogibsoxcnQaS5beAtcE9SjBk
Ks39vRnxWpX5AyENaYvzz/ZMXxk75k1m8TlP191oKjLsa/WngXuEp4OUoZHgc/KiJG1WQDOho9/m
iKFeA2g4cJC0AluIT2RDG/MTsg2MAaWjAQ8SLhTmhyKBPG1LFBIwKgmoLTcBSwzbgbPqWx4J3eZp
o7+A/UDEFuP40CeoLt9gnbvadVb14Btdg9xm2LNrcgKVSTkfJzoZfv2vtH85W7eFT+h/DMe91y7n
9p6UEL4uWfKUMyTex6KWHyE8XEfxxzpZB1AyByf4eqvhr7pcdE3EIOtMEFdsQS/SzLzU7z+zYY8m
vl25nL5igYeBEZDhUYSf9Jy1bZxP9Adz0A672Rz8AvU/P4OsnqUx10EDd7/W0It1qyTKMhPBoLoy
WE8HY+Cz/2ie5nyUdpFf46MoRLZoiPjB6ef9zUvUI+5+EeyUuRd9b+2ovZFaClX+yDaWwAwtxCBE
G5/vIgR+7zVydypi7wZl9malr38WJgM55vzGWZWU4uZ345qu8hkzD/coLi7ZX1mQ9tHIh5+d+bnx
y3VjNnecdnv5qp1RENtMYnn6OIep1ZDL+MAWAGA0JNQXjYwgJGyrDSfseDs3zYXQu3PlmTHq/R21
j0kKnyt7+KS4Bp3xS8Y2sHZnGlQM2QT2hwtVN30B1Bh1Z4EcasHPSeo3OOQiN6B2hMK++Fei7zRm
Ye6Ry2y8vzaCu1WHVOKRuYs8ZShwDzlq/ZL0H3dzSaPmwG0qxcKtFd0NgaMZEmDSsPdEzmXgTKj+
pf3ErKPeMemaFy607SC6jz6vieV/qoEcaXChn4mHbMwi/7g2G7g3rP817WB6Ja98aOIgIuRBfctD
1ObDDHz57O3JwwFB72/gBQPiagBAiMZgvFHFdEr7YWs4PRMWqN1IDgKG/uf9wFc9x8/HQxMJkrAi
1zXQIsNRrLqwMn9CDHhYVrhEUe1HrbNqU84UDT2J4/icYbrxGQ4bCWrRaW0mfsXJ2rx5Lxcb299u
1VrKMdgU+0JZXtq6lfO4vkYALXNTzBJTUHrNDv3B/elZx7/NX26etRA2lohs3KutuCY7iRbeke0d
keSdLZZRsAau0mWaFDOMpAHZO2o3T1nbVHuNWbXktOfrRSEn4RKMX3u2r7vHL86GRYShxdqKWLl8
DSVA2DveyIoTqEGDYWjsxsv26HsME2s/RzW+mD1zpulMiy5kDyoysKBYZ4ZqoLkOrdUA9qimKeJl
ciJTOxkVhY5t57PmKFFxuRjNZE6A7MUdoNWhi38HaSzQLshAnJH00gJGl5zbI0nBxjW28RH9Pnu2
dYxVW096zwd1lZG2P10OiEp511pwTN3WnWIRsxCCm1fNl8z63mRO+/VtAhyRNKqhGlMm1JKfWd4O
1xmW6WgCxbn516Car84omJwAxiZ7Hc9gbCDgcqhivqGeI4XAwxc/5uWE4dvhoeh/gyl3Syp0kCsl
a9gZtisVARwop3rT8Hp27ZIvif3xraPtPtYgezQufpDWY5C6DU2EFo+Lt0A9EDsZy1pkWV34ag5A
MYcnz4BiXbHQohhL4gbN0r4zVI5mjhA/5UCW00CoCSfg6xewCNEj+RCZC1g85LsVH+2sP6GIdn7H
CV1XM8pRewzMkJlAwn+kjJZ4nXDGvEq5UwT6LzEtXSAD234xNai783Au4M/OSQSAHBPQV0QLKicH
Y8tvKlImwKq+ZgONfZ4LG5zDRNhPAZSQWcWjloKwbFU61TtZYMgdBhSCWlQNJ2d7Zoawbml7HF1t
HcrpJ+6XPVY3q30CEs9IGOENHe08SOKw9iYGUMgXls1qycwbnFR3v4K3xj4ev6IwriIQ8GM1OxY8
09JYbi9UPJKu1r0uL3X6qRTx1IG71ZtTANTuyHttDsvXlQYMcPnlvsoWVHI4v8cfuJSY95xenRkR
1r8J+Q9L31O83piiVZ8GCg/Uoo326bKtuXmLR2U5QBNQK78A+WP1xqZjiP35IFn6H753SmJu7Xe6
ac0ps48mD5dJPI64jaVlfe90DaanxA8i5uc2/Jc299Dj9/46UZnwDWNQy0UoJIhxJbsUbOEdiM2x
aEqtvxh8zIBAfDPcT1NGz2+7Qqbx98SbX2Hj6HItfR2UotVAQk9AjpHmmyaq7sXDELJ+ZvkKw4k1
FjCHBEBaCUcPlxZR2IpNA0xdOakLkyrsZjhC9cyXOymV1pYjmzehuEXMw0NP4k5JK30ThKx3jWjz
qPNI13XcyQXR5Sye+eGVDamyw2FqEr4tYjK1+8XOTFouUhi3SDxDBTqguAkonMmMJC33Q6SY/+oJ
qYNUestUAuMEg4ry8p3BZHg+5w/7QuMYKzVQej8Sw5ReEiVvNJcJfDz+2JGx4mwIRiN7WS/a89RQ
D2obQQ7083nrZu6yboQsJeHlyEf55WVwp6VxMKM/qIFYQulgUGjtQ9e3C8Os16syGn9VSty/v09+
gBwdBR6d32SG9P2BN+ebG4WrmT0ZGSRr+33obmJDV3tguLuh4LdxPa4OWvQr49SLVSPvW29X97Ms
Xt+TCTjnZsBvRa0WinmwBICwYDwGX2c6PyNfGVfUU3uuAO3wOijDy6p5YhChZTEhpqb3EslfGq4g
yn93bCPaj2oR7jhWFyAk+TafI4yocGU+bKUhRwUXlk/t7QP1b0o7ErY3BOx9Dm1qZx44owNU2ays
vkDICxnfaHRlfpD5qMDT/7dstlR+CWIWK99R842Zze5lqYb/OHl5xUWFSf7z5cubXY37nD+GMWhI
DWIWgKB1qbXl5bKt8IiLZGEx1miNxqTJhOHp0td9CxUPRFhA1Uk/Sn9HWMrBPcFDXN/MWgue8237
rf811AVGxlyC506+WEgAXj6OiNuj8jUd2GuuB7xWrhIdImje/g5wmdowu23BoYD+nDYtvtLR1voT
nUMpWXdZBEsm6tl4kCmQ/UldkIcQfz/0AYsy6+Y9b2i2Xpj7CnQUEMObSFuaJXZr5i7gmnZnk0mg
qhBZMt528hzQkN8xQ+KvFdcfsgfS6BkRWeO8suCG/ZWquWUWJjp4vmC0mYNSR1OMj3iPy631x8wD
2HL89Kj5oawdF2TJmN4kAGXDILPBiM5kjLLbuhpBC17eMvDkSfWeNtbu2n+d4cxgP1akBrNHyePN
0jY1SXzrp/gmtNJVgKpZqYFjsMqc2gqhqGr819vWX215uLOYcQ2SU0kijv3I5M9QLRZLuioR76qb
U955VzP4oiHW/6UMZO+Y8aEEhAbP5g5kLO+KPrXfGfq/B99WLIW8AJrx3rtWQhvN0x37/f4QgQAt
JvvaR+sNwlQutEF7woEUP+oWxJG1evlOEciGPBbU2sXAiJjr3V1JEfTm2mqTgDdGIfmxx0+7TLxg
zCwjIEI92qFtgTfp8uH3vtnYDTY+JqFuX2kQZkH3tFl7pzR8Vw9o7Q3WQ0L9f3ewD6gvff8W+HIE
l3p8Piv1BzGXzsdUgnbo+ynkCMuDGtqBUpWyG37eSLCkzHbPmgtvlnHKNfGdRLfFqk3SM84Ql67F
1equ0mHboVa4UYFzZ7QwJZumN4472HUN+6uV7Ou7JeM+ASSiyKsiumJa79CnMZEWlyXmuNjtFBHb
/BpfF7eTkBlt82pqtHBeg+szS+VhziYCWgdVuJvj9iaUWxoC2F+OJopk770xFcLoWaz1Z3Kbt6/r
4shtqTjOGbj146KgqUJokj0TG67nUvyiq35sUXz0H5CEZaB26CSJd5Q3o3QPyu3DwV9dtwFu48dR
z4CeoESgIyAtcBID6EP1XajA5RgZZu4OpUQDjMYGHNQ1pJ5g19YD6lvW0xR8EdgKDAo9/xsCLaIJ
LTeesyQB/jGoKf8R8cKRfDtQ4u5xf+GChFC0AQFmXSe7TOW8emC0DHbPSWH4CftppbbGwqQr1Por
fkYhrnS3Prn8+VUF1Rh7WrS5Sl74aYzIemQ/Uq+S9ERnqm6e8Oxp6Rl4A11JA8MlmQAX4aAcAqqE
BogEMEOrT+qPbWKZHybiwjDoloQ4blZtuGR2FJXtJ4pmugtYwg7jmSyVIQj4isGRDSGHH+IQp+KS
Nk+RdF6tBIBrjLsvZjwCCtRZ4HJQzwxL0z8Yvy4WNB8nNI69gv6YiGTVkXvlsPyhnuCOl8joo2k9
pKNzzcTxHxdqqOibjenzfYdLU5tbrVikQYqu5Tg/s/s2dSl20088oaKXQVUe6u575dspSRYvz0La
9IK/q+xyYBh8KhcfESmEE4vOCNxrdFWXPsEnk8navLXdPfl65lDH9ZWtHSVAqHR2i5e3PFCcRsCb
jnaYgZOwocqxNg4cwhLn7sMiJJA3kp7SjxnFajDG9k1Y89YhQorf7NROtYbjmzW6LU3EljnAovLi
Cujnl5lNCl0/g/+dUvtuZbWqyIhX1lYvh8+sh4Vxj3NfU3/BzkPbyoU9yGsU6IPDIKpbvU/sVVEp
zgmUv/CE97+Zd4WEB5bAnDm1wcBe9gaLMVOqhD1QowsH/ODRxYQjtbfsQ/uKAecFxB8pPdlklov1
Ep10cKuP48wxNutxfE/QUv4G6+V6oi9kNCjI50pyTSF7eVTLQ28pnq9WgK+R1HQRX6E3dvfagutt
+A+7yKHVK0ABpgIJYsuVVb0rLyA0KP1wBE86/Z+oake8ZavFROe+xHrRY8zE9rtS9X9DufU+BLiI
KNPTDgCFBhPlpQ0gE0cDNTnc1StLBbury+fmfsS2I5QVmHST5fkS4CtDZAHC87M28XnzFmR8eSaW
W/HSu8mdW2SMqraLgAcV4wsABAtFWFdMJp709U0OBbyM4lVya8DaF9UUlOWnCMDTdtMj4hMnv3eV
tVkkIuyJSzIv941U22C3WBXgD2rxSeO4DNzMkQicJ0NOIekwY16Bl8SjrJ99e1+6DxT0jdKDL1KT
FtYAk1+ez8gH00EwQ+tCADqRNmRk8r4+sQGZSFvBZDjzC3YyrMFFvMqdcbnmITl4oCB3gnNFiEke
ywDJh+eOOMB5DUylN48P0LlDu+6FkBxiE6m+fRS32r8va/eQO2A7UkLxCxTSmvtWcXjHOj1sTzA6
Y4MOxXfXHbzyzfC12FqjAUJly8+lxx46h+yOxiIe3TeQA7g8xY32aBb7qglgkwGRJwvcXAYEuy/R
T6EiWPqpHaP5kcqUGN5yAwW/PsXfgzwKAFQVkfDzl/ZL9ZdKL5jJ4WWNRE4YxBLEMuvgoTfoGubC
h8x3dE7s2nYorM5I1SGFXOboHMLWKYrPWbYn//4G8Qqql2BcMjcrZyUhS5wSdwoeulnSfTngFe30
y1Denx3kdzVTPoj7q/cqiTIhwf6ayarNZoSKX+VPCn9qr72PrwKKaNWqdbR4TP8CTVIhk4zXfq/l
9cmf8lG3NWtnM1zUUcHoAdTQpeSzrGMHClSG3M2znPzHqjf2wav+U54shs4fKSLVULSIB13+Dytl
YrBpzXRA+0uziZS0DiQ5qGN+QTR7rNy0MhkJfEMDOKCZIgs3QeK0lJGtYgIkkzRyI7xUigfgLVsl
3mpuFJ6E4ShxZ8P5X4vn1haN/7qzTFnmQ5SoSZgqc+xX3bAAO/jcMXUKs+aQK2JgbfQBknAe7s5s
nmrjzB+g3csrmnKcE+2BhybIMeleBaI0g8TJtCQqEWRFu2gMThnyRV2CwHsN2GfFEsczH30g53w9
ydR8jVc9f566R5q384gOjJckqMKjueDXKBCXhWTz4UYHpSdcCHb1akYMN0QYR5nGyXgpI/1EEk+o
cS/AwbSHxyUfwkpUTDPJFdrlgznlqKVPjPxfGlJ+UZoNbZSi+l1fGWnpwsGKNoEcVtM0l8V7huRd
QoYr7q0v2xhzygS4/0U++5FRTVg/ZjUaGSV2kgJfqfBwdwfRmu6bB6qLwUxDQKBG1CF5lemCdtc5
KE5ue38gMb1GJBgtbJjyTlE0s/MFNJbMrmZYbSD6eG7LFvOgM9if3U/Kh4u2hiv0JA1/g+JySdrQ
qHKDAxWVQCYiC3mne1oicyvhBsvqZbnMtZVUK5wJDlOR2l6+GEFa1UBfuWd1YJmjNFw+ltDyXxEM
XxNnL29zqd+A/bpkx/PB6a7huw1PM9vX4qQcj9PvYhbW582XO5GgFp+7x5Y5zy964Lbmi/Nr6Yw7
rdwSn3T6+s25iC0lfSJTBfjAdem6WEl7ek3wKbR6+ALTPndbBKhFTBi8YWj1hK+nCh+7VY/KQbLu
47p5v5P+vGbIiaVh9fgLPhYjGx0ga1NEVh5ad3q1ehYIIHsaFU5xv2YSPihSkeO/0OAfHy1nQP4+
rcgtXXGmGs+ZcpOdcKYUrdsG/cajJfKLCQUiFlX+6ZNuXXwlV0cBxjUHKLYcK34eLAofLUVXVCev
rBHD81qJQzKZLjJT2koiZNCuCa/0PjR2SxY2LndtACGSPltGnS4V2UmvNbsSNexoKsFeNMZbfIM2
bzo/Uo3ee8N+NdtQsyWZghANE/+AGj0oSuhyTbCQgPE/cIH2Ulbv8X47jSiGWoDL8XY+NYB6oNg4
vmnIsUPYCSk3ys0tofDmLuSe8nut6DVpksN2KJ11bEjrt4jCPV++2f6WZNF/8POLE5/wCQTEBsMg
wrGBqO5aZFI5zTcVmjc+A8u40Q02R2xBXSRFXPWCYO6UmY9SEJOLWIeCu6qzQ5mZ+yo0xjPL9X3Z
fvWmMTOQ7hmOuCovcuVwzU8AIWWAqXTBgyR75zPD9dcw3pVJEOfO3Es8wZXTTZi076fmdj1S2QZb
mQ+XjuL9BReROJX8rE97E+5YiAr97UbeauuQVwpWqZ0pF++usuy02kkHGT+Ff4yZm0zhfg/ktgzj
ZfFfiS6p20lf3v2pIjF7tMZF8+7zakJO0+oyLVO3n5SK3TdICZOhtlwBYz6sY3fE/fMCeM0s/WHj
WGWAADwgJaZUx30sbJlDjmwAwtRQPldo1AdrGJlfwyYL+TaAq6w8FYDvvwAbushYJfovQglgXyHf
GPUoqHkRxT7LXsQOdxHYfnB/GjwaVFT1vXEpL53Fpp0o7zf9wUdyDMBbwgjggg/HMmhY8c97sfC/
7Rr7CYtZzyIj5uAUwVt/Fr+Uxz13t3MReUkCisz6Hq5i1yiyN40ptjUB2eGHmVAFtO6TS+lWBsQi
q+Dy1GmHo4kcDhc0czi7uJ0u/Gn39PA7bnPwLbBnIwMH6MjX7xTfegddjQtHz55G3rfAN4ZCZNvg
pSW0F+4BE8QpwrhawFXSsz16J/uCgRgR76OwN/J1g+HMYogIz0DFlYpKm+p5Ov54XRoszt9gokSD
YBUGP+gMLn1opwO4vj68kclk9y7ILIH3IfAvpsGztTSjvtjcXglGO9ySnJr3NxBe7ZyNJ6TE6nLS
Xni7XaUFzp6nPM+uemrAhJBNBUcOHUGBqVuEwXQIYBb1chbbOHkUsHeQKiQeLdB67r5UARVDc0fm
oglFUw95mrfYv7AsWAVOvZtTLOjCKN0x10R2rVWV1NOJmutexK1EyNnH55w+qe1UyDQbxCnOosaj
Qa+UaGGvrWBHsYFfx0x+FRUDmYVhl8yysTk8qYHseHvPI3rpRUaVizsbUHP5h70b7v1T3e8DhyYH
OkQRm44lfLiqxXaYMgH+0yKKuZ1YPYvGioMlevejAdAHrMSF506fazsjCAzNpe1Y0tDdPMVpD+1S
eoH8QxHunabKgy8Wt53jqLyKr/xaiZZRsyWfno8gv07ir09JUuu9xpVXHkxdKwZUFPYP8BdWN1j8
+jxZeyZelHgW4wARjYE6D/NaNguoV0n1qCgpfg1bGnwOoej/X0vFqP/3KRTdHzSoQDsOkk7y8uDI
k45oK7t73J2e8oE0S4gFQn1VCaVhVN6Nz+Gq57ZnbLBOXmtsYznB8YZwF8PjtJiiHGMCU+tTEGBb
10vo9AbITadf5mIA+TIZelbtz9K6HuFI8scG2xzLMU/huWzTDYu5KpWPgIAKmwis/w9OrAIvRvHk
q920cR/pLUaqyoFppDPyphYtc4C7cczfa21pm+oWvj06Xamf9t+1SaQ6rDVU5vCPPSUvUrbbfvrF
gvA3K4uxrCrdDX8UU85fo+CJ07qcBYrv18eJ/09loabzyjrSKpkAexEk9VxswSL8vemzr5IsXwq1
72ImoAC6ejSyan4oZ67MMIvoem1kNGKfJ8CwRIqfs+Un6Ura1+wMH7s95fvHlVSA0ERo3XMRNmK1
Qj+xeHwBLxsf7ItpRQGX/kHhCl5QZAQKROC6FNno2NMSHOnQZFyNtIhm2RujGJAFVkxIqfEcl0s/
xMTjoKEu8mL3JA8CnQhgotg5anFKQqrgFeYkouOBQOz82WnKXFCWWPqG/WmYQCXSFerZraFh8TQL
smANfHn47Hw2cSQ89HAcZqVm+nZg9dQN0V8067um82EcTNCDp6G5QnKjp0s/pzNGQ0cPomOvZlD3
DDXrdEEuXDDSNgKxDfLeU/EZ5auT93L/KLJa2ZgLndP/hNXjcYD+BCmbc7JCTH27QIvhSXBlP1LN
Xw4g8VilIAWuoSzvjuO6WL6zK8tWaomTMvl/re07saqg+u1vo2mXH8aDJINJHcS6IrTmGzKnyRl1
6x6AXQfiU/v2fBmWb11RusSqYFhuL1866lNr9c85M3Tx5dSQeei4EWg99SyzLINao1WzZEzYjcfh
2Q0LuAVrRCavcPKrnwsWOamoSS2JH3kaHhHPt/xG3MnSXtJKbNsZoHGtHLOaVNT3gxaq0BLYjCqV
ZShdkWrBa8eI8F3ghNqDZtlnEecdQc0yqpMClPMgzmTmEzS408fe5GUkbPho6IUCP+b6CDKNHZMg
T09CEcCTWEjpSVzbGomJOk0eV5YGczdHsWLzawdUekHylxk3JAyrKyw3Fm7pFhOTTAva+5F9Y5cB
ACj7ulTk9SMzAm7eDfzRABbcbjFxgCr2y3B7B6cdjvJHhjE965OJDeZMaq0WkDKyb+Cx2XEZpPXo
6IK27sfP2IP7+HTx7oI9PTBrUZPULiWD0xeHjfiPXQOJSKfLmCwsQwLSSJAMNtYz4PPX0hbJDzVt
EWmDzrveXWA+c2T1vkK32oerzACqiOcPHzJN3QB3gehR+Ky3EDGmlYs/hIFhJXOPkU5+P9vXsiiW
hx/QcjpC/VGnk884ktyXwQT5NTqRNFahp7uEs0dWzqEGIFPZXqSuXOtJdRm77BKgOHzQ7sSY6+7M
0DBNa9HAK2m4H+G4hXmL9hCnJmrSo0nAV6HFgE1BwUI2d4dKmHdPL4Ia3ykTmKZ9PZ9WhGKmAv1r
g+AKHeAyn72D/E8E7LvIAqi7TLXriR9z94SdCGBg1SIDPH1Znn2GvxhIfnI8/OwwCkF7Th3Aq9FK
rFfijMIBkiBh6rtYzg6WYAvwyKNDm7DJM/eaihI5fyzEDTNYjR0pXWz1VJ67kiXkEEkeI4Ip9Rdt
ED5FhtB19Nyb8YiI3svwGrPxW0gbGBxaOG/g0E9MZ3QL90uyl/w/BWmtJ1heZEjuG4tbkKWl0it9
SRy5CleiV4OgtmSp1ts9m0cEkMkbKcRZLHq8aeKEBV/Pv2aaemXhHeYHEyBrSNKIZN/WlxjDOtPL
Ihq5zT6efkO815xXJ1ZwB8hjVcpr2QVNAeHwiDg79P2Sg6KhuDv3iKtwl2GbxKx9MK4/aVYYe8t3
LsGwubA+V/w2d1TJu2Y9itm6U1yg+pZ42elBOe+fArQvpb6mGzw0iXteFJIIJmguQf81Ax2vHTNS
WyMSNWH8Vw/lpCrXJSFk+2Cf9H0kfxh2ZVSM2/qcu1oECxRzdT2Y6hDv2Ayc3d9MJW92Tx+xWjms
0olDywq+boowo/sviqA5ThZ7pQsihO8WKkyI6qheXrt/vHR7oUdjSjHdUZ0UCKCaHLToDr4d1Lqd
hbeEYI0UtudtDmcaof6Y4gt0BJZev8BGN3FiRkKEV02qBRNbDbNQ7tqe5Rqa7pM6liLcX9qAR9et
QPhzh3m43x+KwtAp87cvd8jKh6M7k0ayV/SP+vNFzN3Het6ozMQggPNYl343IM/De1amLI/OcqEO
eTpUNWtiRRnPNHwXZ72lDXl7PQ26g73IRfQHKegUUdbG5TRhgzpckyMzpLO/qbTYt2U/aSXVcvTV
YoxmcRKkZ5JMsRQw2rFviZwmPE6bdesPoS7A2T+PvMTW4uUG98sbrbzE34zPadIZCZd/nyRVuWlM
MMH8alRKzxO4wamehnI+rjcpl+OyZHI936M/bvUiiTGIkxlVj3Ufu1B0kzJRmdHWO4mTPzs7ARfv
A6Rq7WM2KtjO05IZY3uKRaU/x+S19W/vvxH+T7Zx47seSVfSKQ3PWl4ucpqHoEl7o4hYKnBE+wYQ
eFQeSEQIQkiMbA02Y0B0REDeX4zgYPoRDh0utHc1PdEDcsApTwyPk8DBJnX19eFnn+9PbAdEPUi1
I72uMDfLqSIj12XFKFABVW7W6fZu1H6cFrrsdUDqxvZyuIaIxPh7dLBGbJsUbRovhKABRKuFE63F
nFzy2Ro+dhSPQ8X9HbQEemrtYmEn+LDE+Mo1N2kxll3hbqvppdSsmUC3eBbAHuh8EliH/hO6vQv1
u/tROh/yjMMof29v/fqBu/RTyyMYfZTXkobKz0c8Ydmpj0GzI3W7acnVmahfhGm++IsZtntoR+Qh
/s2SIUeEmuHzkPJXwNh00fFHO2uRUpRuH1BRFxTazlAs8Zuuqq1q6j7eWVqwQLEN0lRNzuKNdXAT
eASIbIIr2WJs0Thl9JAd1iosufIfkYLx0JbYF36bKcP7coAYT/wEGKOM3OyhV6hPMbwxz6S6kos2
uhukL4IaILhFBjci+cR009Hddbqul8rMCuZcukeX8TgWK1nZVYwUud7w+W3ojVGEdoTbqPh6pIn8
VAJb9Mx8J7MvGQaxITP8HIgZyd3XKivlM9u5txbASLUURhhxA0tSwztpGit/U2N4YcgiuNrD3gu3
WE9T+rdYEcM4HjREceeP42lcLyj/Spzkb0F3ku7cByZ99lhX1Oh9Bc4Toji2Q6GoGnNi8PDv90sZ
fFoHkkUMV+UPXoWgcSTv2X+m8Raiy6Zjp0Nsz30pC6zAGmYC1u4wrgyx/livuvj6sTxp0mHIhqm4
1XG9Uv8QgF5ihttp4pxPZhyYf2lICX93w/9yMbMvHaoWty/gdL81nDhx28FBLjeS0VupkWYiala2
8lqnYF86N9YP3ZF0glTikTwjjoIRGyZER6XhMYlmTs1vCqEKjbPNiC88MnF9mS11/8WHJBtYvwu9
feQ4xzjAX7Jm13VxLYWeL/BspGTbSxxwfa6lmJjOMXlrDF3UUmmEWzb63BswbXwlm7cdKz1HsMeA
7JTvRaJZ+0obArYaxHkySsB5IeoLbiTO37RiC8kBD4K5SJpMJFQRFwJL3FQ+p1lLlGw8e9gmY6fD
PKl2H6hdusH8fBCXOfdvvxQnm1UwgfNgTsDC8MYxTR+zV6xRcYgMQhFrRo2XmEtFm0NgvSK5hO+Z
fspfUDfuHRgo/L+F+SFkxqlyfolInAUcnJY4z2J/QgASwVDArf+GhKOVzhuOAJyN0xS2zs8QTfsm
Qz5J0zQrF8BLNpYmZIIoKFAHHSg6MkhYscIk9seTeqYMO/UhiqGseBjTIJPTZ3st91uEXodoeCuf
QvyFaS0zjiRxM8JlCiB4ShhPb/ax55+gLJN+cSSRTWhatpF+PzR3Vj8Q5Dg9MKg4g+L+efn+wZ3E
9wTWPMVXwxSqfsNRnczjZkIaBQQYGSggKIYWpTbABq5qTRAlWzsF32HfOZHoWwXTWgbjrRPVyNbH
VnV6Y4ksYCqTxnOVkcJi4B2A3PzgsBKcTOg1zKlkQJCC6VznW5K+jH5kropIgV7/6SToWAgs4+EL
GG4UM3imorTPtNoWpIuOgBX1qNRq6QJEHYa0gz7KOK54mUKs3mJ52ThQJD/2+r8Kg5HgSjolhKDw
hucly5IKQc3b5jN7/zRhOyTo7uhgMqQfT5XkjZJHt8srICUKgLJYvk7FsOf+0IamlAinuZln5WkH
F9aFPIuQvv362uvSLSp+uPnI7yOPVYyIFsEZg3Ev9xpbuFifL99yh4bI0dZ4qeRRoYCbJCd3z99z
bogHRDtMnSPUFnNIGbp443glAIHcxPsQ3Z5UWvM82+QEqR5c9ij36gOhjKgyjFYDi7TEE6evOvzR
IM/DVMecpSkNsHug3JfOHu1fKwE6aE5kmx25uQkhrLBZeAYAf3UD/7E5r5h1uXZykcCqhqZt9Hbj
zd2GWyJBECM4MhcBXPHBof/olXqeyIXzRdW4yQYOxB+i3wZFaMy15yksBaWD4qJURJbm/U3l0Nke
/OF/JKtUnkYgCPouJjoVw0ELRnoRkvLnoH3nUR5OC+Ju7kNXOsboNFbSzy1Cws+G96/Bs5LYX85n
lV34zFzsD6FrCEU0XOvyVoKvvyePjJKXz2udFumyulm4ZcZStwMZy8ukL3LC268NepVnScDcCF6K
d8SSPgLS2VDyKQOco4Thw8AhK70kKJfILF8KQvTDLx7zRHzokjVD7tdQFQ5VYwRZX9Ktzr1Tly+y
8+xnBKggaA32nfzAKW3ZYn0sCn534gdPyPx2DALC3e8+eoO1kxdVOyyImkICw/O8H0SwEMMY4iVG
mvBTnbev+JqLxtVu4W6suKkj2BTtXYdzdmfCnvwKKtkZpPMupYyh7mMCXb8hUpMr012k4NIyjzPQ
3SJ1ryBCe81AN2ieYJOhYL2pfhEsEuEtcIaJ01bfn/cMBRJwPoKw2xTUBYqoJjCpxEazHdmObeuP
ALG53mKMUkjDjyVxsGa0WgaXUzgxTiJ/uLRF0R87CTOGmAK6RfyzsQ0uwOUrU68wyUS8Df9iwhO+
alMWOerLzOjH0X1BtFIo28qSoDCMpKPbKbRdccVENfTawvyq1Ae8B+qlwuJPJhr5eyzXpp+LFXH9
aaI3RZSPv2rYcJGXJc3FrFnRQv0KcoqEyTU7x1pfoWpLnvHz43jcsuppby5LUauXlvqAWQMPk2L0
+X8+/pQUtSvAN9wXbARgGAT1FXeI/aWPdDkLUnUBeO29wLTKn7cr9Vd2f56HUveRKmeRVcm4nUW2
Bs802OHnNhtQDdlThdAZBSDqqTTYJ8Ts/Pck982K8i4k+clOkRHU7gVBftRgfepq0JpObThZElyR
A2BsrsQR4BgiaqRw/3/KmTwTMvCGkqJ3ArkFkOJz9wVHhFrlckmk/6M+1U2YaQhBd6n7ROXGcFy9
fmAfh+SR326y5xkFs4SNwaUkudHlY1583r05gmPmwLUTcntrg+UJMmld+UortsIY1ddmHAc3Akrn
wX/SCwe3SAEceXUrfthUyagw7A3E7L5JgAKw+bIln8nyoEcWjMFLwL4Iuy8hFTgGG/ZkwvPc1n2h
0ei5D9myqy4pPh2S7baxOS5N5Ks6If47Bc8V+y926e9lV8m/HdEZPa9KHsSMBo3ByeLtrspjtRlJ
+sJTyZPru51YeOlGBIU1H8jiHqUz6oXdsfht//NwpxuiHuzTvEO/uCHAWyfDmKr3a7xgxZZ2BE5R
AjdsUGCR2GQHCXOo6awv0oXMBKLnckfnniac6AAP6nd8EMSiODHbdJJa70TuJvpkKYWLQaX+/QCI
fWS7NZ3XwPhJsPJ7092Yr/PFjYYQn7vT74WEQaeN6SrOw+uOwOm0k9pFr3vNV6jxHAXa0grbohu8
BG7xd1jri9pwpoGiiG6AogIZD7UhlXp2mNoGe6LrkOUqE9hEM0QplY/IoDxNbU7grEQLIB3Ef3QX
zD++zN2kCioLkLKv7mmaYwaP9b5m47SphXy+szZsIxasKX20vU/HhhtHX6ngDn2Mui73sKf5if10
y//k3EjhkpE3Cuwla/ZcpqbXl/jGke8VXYHFCZqTd/qie/D0UmMIaGarGcjV5J8JyjLcyHdWJfUK
MUcQx90mleoF8RwK04j3PIcfu3DQ8Iji/lfVAKZmrmd4SaFXlezqq+v8qTjD3CQPSlNzkghv8FrX
F2Xp3XmhnFbyeErzQ4SLYwr8LnQHWnHj7srTe5UbhgfReGIalfXVXd32OUf7B0pOveHBBrmr6GBA
x5n3qDJUjI69sb4cMajiT7vNuNKKbEsIOQXnJ6hbrnULIEtWggue1oux2czZsv1+B4hZXCyodwmM
BgfBnmw5e6/4sNkAig8BNM+rUzm/uN4AYyvX9h7NJ4XT6Zmpw7wDYD4ZMAdxtESCSiUgv6oezar8
Na7WnGmEAiUyOLUO4iaNabkx5mPwPQoEEFrx/QWIQwVlax5B5tWARKi39edgnbec4A4m/IxFQU2d
hw8a2BmrtVizwsK2vcjOV8YNMF5JuxZAhUsxR98YrIjde0xrSubqHxQNIBEosqKYuboHtGWUDown
JiV3UqC25PX5JcHT8DgR81WSrbvDnUlt2/rXoWcIEA7b6VhRr6WX2p0SvuTroF9ubmRWEkuKvYDu
FXGgQuhK9DJneG58DrA2eCGXE53u/UM0m25QcLbgZwhYuS93CW0yY9HpajRBdFx6qVRMmY8qd0Vj
mUSU5Fjybg45ymPDjBiemszYuaeGyjTNbQFDe3RyYjLFxi3+kbIQaDtRIghHqPauTeiCjA4khS41
mZ0uPHX14oMgV2JMccYUvUIlQmJOuokhI5aNrWk/At3eMrZDUOC9dc6u4lxEHHPGh/Q4bJXWYwCB
lLoHqfcGji9tV1YDum7LVrlM8ga2AueM+oMx556hINgMyRDIYKpdF5jPVrvsatBYVy5qUaprip/h
zb+aSLF3L3f5OLgpEBIxRdrKBMaTM1jKvWAvvPH6SsQS09zCxHrfy7wlRhEwySKqP51SAbxlSf22
3/pqlm4JhmKWqQhG6e+COCGYwMJVBmWO62z5n3w/WR+9Fcxil/Vifw2wDhffydiLEwF4qBZ0nQaf
YGT1hVwjyEqKMse2+28WOGRU6LAVukhYfYhNU/Q9AzcRcsOS3qYygLdEeE2QxupXy29vLOBA7HuF
5YM2hvMlEV3u09OJWheSE4kjD8wJrDQlEZ5nClMM51mxIRtDR0RRs1Z2r0kBTIWpsYGzUNfQO95E
gCOBa+50dcGyFAHvT8MqEhW4mzguj7Vwf6d7RaHD6Zb6fspg6YrSFJs9Pl21JL5dBplf1/UlOghW
9C8Gc/r2ZBLMnGwroXRGKABiJC1qptOfz67UcdITygYVEQm1OKrfvYLqZO+7/fjUtWm0TPHwF6g/
Csfvx2WJ9Sv5SLZwMOrdATiOQQmxaASNMkuIOa85DgoXqHxUd2v5DiwODcYrheM78Is5L0HfFLQ7
sseHjQG8GkhabV1FOVQmm04D9IKrtnw237LJptfJPsjEJ8QEltA8OZKiVp0H/vQaqyICK0y9W5nM
o43Uw5fpU9nCQj584ECwtxKVcbf55VyrtNWsb5ZMPx6UIZctKEhUSMo4bUaxoBszDzdciwEo61ZR
ibQVTs53//h/7xfWYMTHorbJaQIseiUvvbQkTKOt+/FKeiLEgZD2oiYEJRT0v2jnRPddY49XcsOS
8Gyg8JuMk6iM/JzTu/jEtbekiLUFG7UOiWcjq2+Ng2W7WYsDDqhpQNCWho0YIeU+FdAyUPTjpxcq
Rqgv6MG7tDbtCvLlHMF/YftoGYL0OGkOXW/j+kfRFzCda9j68bh+9vd+TjCw1mKlHPiQsCnlb99x
wZCeaNoPbdFz7S7WTZQvig8iunqO/+GF87wE8m4UZmigBVYmlvcgxcNQv3i9c+srTtTW29wCo2fL
GfSvExSkIhz8mnBEYrk85SrQ6XjADWC3vhu9wJv5afQNQNY919tnIq96CAPQ06uZ54R48FY+1Y2C
uJCPHU8xlLmSi1n4SRA0o0Y1wKLWHWL0Kd7QiBP8JZ+y8x4Xn+p2lLFlmA5LKKr1K7i420x0RHXA
Mg9I7hM4oXlllmVkW933Gnu+bR2VbkAap6AoSOCVO/dJy2cWuCu9AP1y750Us3jgcpXe4HrPWmED
UytLhyJpO9uAA9VnInyU8a2aS0gQECXpukm4dV0L8z5fRqs2pBHTWZQcobXX5AAV0NwoAjeT2X3U
yiyRlpzehVtkKMTSLojM/a5lJ8IYd5ZOdMWYUzCexwsTPADrSh+GabKYpJyinZ7vliF/zOK7SBTf
QcW4ahNwi/G2ckzxrcVaRAjUUpVXYk48ODWR3hs2VGQTbF3XimtuPVL+iADtyCdF6PPqabM9/w2N
LzIiWlPIyiBvQNJ0PYc2BqRdLEl3d4blDX9/RVKdUdaXSoOkCyY9bVMNXbrdIxxS/oNjW/qRNJmV
uqs5dUIw010tzvPjhZxgMpxAzLYw25MRyyQeMyYcrVIPmnh9GuuXc4ZzgUtMkUQzULD7Ws7ey2Cg
xZflYK/eK7wBMez2aqEQEDHrvvWxWRZFsiepm9oTcORyaWOZUf5LMLBdRMCMs9bsMI9sbvYiIlH0
DWLKImHbpwKMxaoo2F7UVy43XOLSRsvpaiMwI1HKCxYQtZLt+j/3NFleUoWlCUXMRlpRlrJgAZ+n
B6aTrDCiNmPPkhYQ8lO3ECN4iRGTdjS0T0iEUyzW/oZ4pyszFLoOm39/15+5G8LIj1EMdtqZ6n55
+keHi0inyCRqm0x581XJPhax25wBTeQ7sePL5F+NAhNjyNmzA14lS4mtzy2O/8xM/7kO2LHuH+Fw
+q16Cpt5S6FaA6UTIQqjynAG9EGnq0OPO3WmEjUxv0cZzmSEXylS8WSqrPTuJK2wFm0YUABCjtSR
WDzYohNe0GTwMBqYoeoawQrTnVMWWV0f2gHvrVfbC1XaQxgg5Y/q07vY4Z//45Sxdb1l+SFp2Qzp
GAzp18xC85PcsG4w47VBpV8i306unRou1Ha7vEiWh2MUf+GZSn1wETBliHFrQNFHIr4OAr/qmwxS
o5WQANEpXvQ3bq4uC6/0eQ2pMBpGEWu8SJ9CwU3vcHaJP9Uu7sLaY9vt4bchZMRVuQm5O+NZRo+n
dY6rkZSguoJO08tVcLQcoGaAElu5z4CVTlKkZuuCPcQPi9eQozK8TrRSk8bMUDzt3n9edCItyIVn
CnY06IxqAFY1VLACTEgD34Y0kKmACiwXla6MC2aCXqRX3r05Gi9SjbiSnss6mkQ/2qJGlGBRmM53
4JWuLv1aff+UTr6971vCDPaPNqVgyUhoGnkU5J8iMRskAAFkr71IYAGU6yhGVB0q5pIwGXdx0qqb
Hf0KgUocLkqX+a7OoVMKHiwEk118NIAeXjOb668gBylSutELbxUL04FFhkj440hC2kvxbzsm5Iw3
ifSlnc6Rps8onuusek6X86Lpagy5ZyntHR0s9KJftDxRig0wY0e9F8IbPHhz4l2/AiOaxDezg222
jt9Sv4i7UvISXv1yCva9ELig9PiSu5tTRwBE2vlYmsTbckOsJDHjcoI5qHNHNKn1q2l+Ul6vLbrG
jYWfhg6KOgvyJtPg9elTdKPP5+vOZkpzfTjCF0gCY83CgynCDh2hh2U62CXmsL2pPf6BYH1xvChb
op9LRHuZgJACaoApPAdbukwuP/xF016G0Hu3mDKJ6AgEzDbPI+v29trb5qoIquNM0wfIDPiAPNs+
W+DscxpAHZDXn0QpTMo5KpqNWxTA1rpT5O1+KGc15RnQepcegpq4qSBNCPVceH2PXU9S3hrJ8m0F
tbUh1TxLpD2hSbzLGxFuMw7LEYbOX0g8ep5GQB4BnYM8jILRoNwCOJP5wLBdJBfykWNlHxHXGem6
RfnEPXOn4GfmTNmrKN5kTGKY90Iqhn67HdrA60CSp7+7PB3uNbgu45/jORFWeUXilR4ra7/riUbC
0Vv0q1g9MVKjGj7oSDGjiyjRbscHGO39IIot/dgd956YdAfOgjCVow6FsHn93xzSXQjRle8ZvZIp
LCP53xx3HwyXIXjt6WfYqDYn/f+vmULqqZ/40787ZuuM0vCdAPkS0zbZMRnfiVx8Nh7+FYtWZoZ9
1lXO10gCUIpMmIVmo2dkzSjQ3Y/Xb59GOt6L4QEfmZnqiOehpQDJJ2AgeY81gz7PWuhNhfU1A9Nt
6nRvySmITWmpmblCYemMHqgNcA+7YGyVANzevYv/E37Vt6GWH76pkD5POXMRdxbl6vDqN2osjaVx
pWZr8Vgip4dtwqPKWQfpFIAGfSCB182hy9Gv2VswJPhhR+zj54P+qLSy1hv90j9u8W3OvmV4ah07
3P5Fc1L4vAZDxgJLZGIeog3HXCXwWjAmVgspGAwgJsZopasyh2gY2u4SISdWW9LdWiqmvDj94o7B
//Fs0TS2Y8X67nO5P66z3eNIpU1W4p1Qln+hg1VpKUbx85z6Q2dtwRv4SYsztvC4gEVYMqou/Rlb
VpHjw1bNSF6O0D9FT3y6ZFDqOGjf2FmT9tetxTHLeJSoFQXcvQMg0cqSKk/nqNmiGZ55AUFv1Ecj
SfnW+y9wsLFCc/E4EuL6VlGQuxhYmofILPz5qH5m7zU00rNHLm6X3jhwg83KiwqMYOLIq2w5zOUJ
JiKfd4gBqX/6k0JWYtF+DtPWMc/SG75XfaC35cSC4ZEBulUCEtn04MQzrJtZEAEVaKMcA4yrdrEE
NmHFLO9OVIKlnGjRze9oExWjMy5LYwDqGFmeUnGNQtQ2cQbqKdIKfWhG1ThXW9juf/NfqmJMN961
FXTMU1XXeJdifFEglLFq+INUsSVooOvP0x5saqGwW9UZOyx/oefKscDJCDDiPpalGv1MehGa3NOm
RSSa/fTR71oQC6GSboKkyVUylmdLqdVWdUp4W8ZXojlXgtQIPFAzjA5zX+tPnB4GC8knwZmlPuWA
mCAfpYB80DqnpZGdAX1mBT8vpi8WfJggaLB8ZJ/niwe6lFpoojJF0mlk0iFNCciVw+dGyhqtJRHt
tpnnDfSqIQ4Qs8/sphnDBo+gTAtGk5A/tqmWAgTzwtbVb0k45d20mHtcOKpTJg3NcMdF/gtG8Jng
go+OTDIQe+hKXSFemZW0WBzA8q3GnyDaUZBK90PTWvi4qHgsJNv1KUHYdSFLaEuy1rgQl/m1rAQC
M53j7bhVDjBdF0wPSvv9F72CzExaqR0gpDQxI9fbUqWAzwOeh0+z1atMUdNV6pp0EfFdqxp3HtJr
+0gUJC0JH+rcXiIIxHE/+HmK+pAyhxd1yrjkqSg2dWVjIexzQ92iDRJ+tQWAhouRvKwl3AGmPsIm
JHbM7PPYtM+5V+IQW1WePSnHKHLW431kODSDdgDPADR7W7SRKq0u3rDlIrJaCmTuTTukaWbRVQZP
iEOA4mWdPCZRKAEyfOc6CcGm2OkboWIp/ZAG1N2ZDE1uWnOUnDjLiOFAk3gGcjhbasahRoWHNjYu
lQgA/DblBladXBvk61Z6CywRDKK0SDEpUV3K59SodcvTIlDVCLvhz5KdmT9Y3qOi8doL9xdiXniY
r1k8OOMRk7hr2vNUvnMXg139qBzRLj22LDIXtFN9xVsrFAwftbFa+lABtWeI6AAbuQa5FAnRcXfs
XT9WsL+LfyBVnxTw0pdkaWGdNrRXyMR8PpHdy9JSYXYvnfR1dArc4VCq8QupfMIGbtwA8iyu71jx
YTisVFO+YRpAndmF9wLi0Wr0y3jZIFwMElogcIku+HjQMUOihfv+yrNkcVKBC6o+RnDgkVALq0KR
XDpokg/JwtJYUyWT5ustoVqWOEWDC3yVZSphRAKQ57Rlw50dcdCWv/TUh4Xqv0OthpGzuFyiS1EJ
l3VMf9GvjAHGdn3bfpWIT86TvGd5Bdn9joHXkuQZETf3Fyw3PBWS8VesxcIVY9cfDIMfWrpYuqqi
25w+7uS0B9fqx15RNseG23ZnPpDiwiClKLNTcIkiErHo6V1KzqbO/SZls6OQf6enUR8BYLVj9dFA
SP/sjmP1lrRAfcRm+WzNRg0uQWxMGA/1dawtCmEVJg+kTMOqYsjdxITsx44+tUE2ruisWmLmWPUQ
YElx1mxe/rhrt4UnejE2naqsoTiG07+LndsWt88pXM5GYTb1BIvljC1jjK3elh6SULnhb8WtHcSs
cQqUgk0U6pIOIWrjhPHa4ffbUFGflEIWHEtNba4OVdB+BjMb3nJj+Jnl/0reBSBC+Ny9dpAAmlWA
h27GUAvnAvC6sG764bd4V5vStDI7gK0FzDw1PjR0Xybr1Iu2S/p//Zac+QsuWl55vPcU+QUTBzVA
2sy75Cl6K8kHE5hZXXDOHDF8JeKA6+4LqpfcxSnftaU6/ZrfrrsJTwMWLIFTqKXblMylTIatwL5B
bzsnS3EU6a0mu/c6Que9ZxGWqF4yOGMspYXI197g6AUv/78GsbtK3PBB9x6dpGcaFRFmKLg2hv3g
8VBt/XEd93wSeiIhVt59YLcdXO8Ry5sItRjGjs5Hcsdt3vkNbtR+ZbvnGqxAJ3tee4E7kqmgBEap
O67SzuneWY/jwOkdkUXqlz7Vmj+2TQBIVjOJTmMcl6xpxzs0Wpquqbci0NNl8Xc31L+l9H94SG5V
gja2pD6eqW9ROo2xUGxbjvWdUcAoVOA8lCzhdkGGuguFGl1lp25sgxGdP61yXJGXM94tTPebHXFk
zAU3ovZ/p/xywCbb8G/6vX37940+JsHkpGGdmEU/8rTumIigR7KtMyVpgYovMaglaiojZBVCB8jP
2HAz7JxTKeTldexkqgbxriuj3SwC4JizZKA28yEroLlFQiBhLkuETwUGJVQPD+jQKN4qbn2ZBOqV
Mcfb65vDvpRJON8Sg2hndsHRADYUZtScMNgy1EOlk8cXo8xU3krC+q6ReDcbRbt7/NDpT/6IRs6q
IDWsl8S+MhYP1DBwmUzQ4/KO5VyysQ1+u+i02lySQm0RAvD83ClieoHsKc/Utn/JZfzoMpj+F51+
L3VgMuzeAvuU6rm4pgDNYIxs3CcPB9a2QxtzOofSoIqTiN8AzzDbb15kESdN1QKN3z2O2bsuQrmq
OVsj5M3bvqL5BRPAfqFd9tBs0wTniKR93pEIKgC9QZx+nCHhD7A11SO+l8Td830TPbm6aBV7kB8i
BmJSoNw9K5d3ruuYRgxEz6A0SgkgbHUQB0Lg7A6ICbyD0y6D7mkuKTul9jQGjuR20gP4zC5Yh3Ub
M1bcHu5CrPqW90gxI8GWJ8vCXoAzP0twzQEx+oUNiF5FUlxW99Tvuz+c4Ok/BtcxmrHO0py8AWVO
4j/A56Q8M+ATYLCrQ4lk3MIrriC6xbTYB/smQh+QFf+MCa2AA9HkAK7K2to2T2PsI97hFHRFBFnQ
+FApTas2xHlGFNPSiffsgkEM2efsG+E1DsWHSwfzkjkQoJZTT0TzZ0+JsQOj/Wv9TE5QzZbWu2WJ
0qDKi1H0Lx/kFoGvrWRNLpv9aP0yMPzYi7PtHhw3QfTTPrbfX59k4m3QULtWjou+hNgSYTQ5Xomo
uYTVuukGxB8+qv0BNsCudDaPygyQsD6OZsupqYUnotRLVFKTg0gWpGz6XA/cBFQoOk+O33tiuG+D
hwEPtLb1jP2g4Y6ss3rBTd3JkrrcQNdzAo5t40Nd5T18rJlqeZ56/YIUcEs2fW8q1evud3MFMdot
EToJf17QffFlSYoT1DiImxqwfY3wZPnKbl8AhRdFGgpI3djDBL+t3RhOKr9dqejOrRXKzkO8V22S
3gEe6GAeyzhEoEY/qKbWYuXjpIVAk0tg32LsGecrSuCsPM8fEV37X249dbDSf8pxqU9+CZU+xhLg
knb2XJHLr5uMEBJx7+bjVn9c3kPrlH+b7eFPr/yEFi3n1iDSLHHovBxN7PYh++QxhQlNgWD560Ii
+F6cNzfwhpL7ATT5v27/cbL6Ag64Kh0yKB0Ou/EQT5+VL1z1citHPtQ3GqW+30szb9VOMj62c53T
T10Ij2HLyO91GRdQB7ITtZa8vgH9rFUj9vWAvH5O6Vo4bK2dZ/nZNqT+WouIJfAZkCh9QCoH765N
haNAlg/vE4mz8OASlfaIfNqFX5dC4WecbTB+t7hpM957moBkgts/rKdgBDDPFadcxkfD287ug8lb
Ti5MVenERDnEP577oilKlsieuRxfxxDq1rmERvRxrmVvcGTBMpzBXXBwbonBgRMCJhFn46NL/5MF
SxGv7HaZRBG3y69n+53pkcq2fhfsGmDcib3cCYanRg1/zYkYVkiEs0Ab3UlK5lFbTH10vd4uCQpH
F/A0OqBIgKl/IqzjoJFyF672SBQUxONLu4ytf6Q8eWQHV/r1sFKje2flD56cKfRNmRdezrfMXxzn
ZSEdA9XTJtzCSYCyi7RxxYqP71XefzrbC/HipInVTA6YOPQZ5cl9lOroryUmDiHWlE+zQlCtTxqx
/lTjj6Yjc2A5qfvjlLFE9ok+a5wl5hS5nEF5lPxm9+slHYD3temN+MUhsf5IriEGAjKFlpOFbluE
xfKVpdDJCvWPprG4klZqdxt+RbY/kXSf1ivWPfBbbwGSFsfPOF6lIFU77qSYMDk0U4wAb1MO+h7M
0j9TnRi/CXIANDRdmm8iyXoRpHBVmXxSIg3+DWT/bUH3Ni3KVxL8BvtTLwOGgGb9ZVP/vEydZ9PQ
Dp4+Elbe+toUA35Z1ejUTcW1lmFtWv6pFrUlQECJTS/WK2QAJloMS6xHkWT5k9UJiwtIKTc0+ueO
zAh+ETtihr1rsyKMS4M/Bda1/cawy0/005OlvIRR67USDtOuJID8PMmA0WYo+PE30KqFJ8SlfuBb
/ffyhKpF/Cran3OUz59H5fjZSmsALLQVqZrRNCwj1lkgR5Avr+AQr1oVwmevtSUC9yz6fsas3KEk
cJXlBEmjsRzJYFOfbBSIvqGMRP6Xpm6jXQGK1wfcTOeYspKv2RJrh3X8BulGz/qtaUvvlQis3nr2
ggdo+UYdsTKlmyBkkrA615SWNfl+vPWTCvhuFiC3IgMI/BBI3QCwonKN9szoshmTwv2YEJPyDxDV
WLE0Dr6z5XLZ1F++JrMcbLNSk5TxEI3s/xq/MCzwzTOM2lKQlJJ6+vxOQCIyJCp3yM85BBzm2PY8
0Wc5Jjt3Rcjz1JhBl3vMmhPBA5PA48TeYH3GqMsEoI7b9wcjjCY2dsGXmvqhVbllfnAdrPRcwHPk
TZi9HK+jdNcNPCalVoSADn8fkGhon1CR2S99YKUsUe3nL/YvAdOp7oRkAhyP2qdaFDQAL1AQ4QDD
lQiQVNuWdQoXOK7w0t2Q22jKbQmXp8xJy+c0kufX9SpOgBvuOgqy0h/SG+tTWjcgPVnJAKtt2Uvk
op0ahKEg+89r+9d0RMBMTvf/1IQ9oGS5T84SUMrQ3kaBIvylT8BZuZncZ/GxRJNqjMgEwTyR91uM
3X6yGVRTQTM5dpvRbZpOggwVhdcIyBWRuLPsf8PiGyPW3oiIbA/4+8xi3YCCOrk4JfwKTzKGhwRZ
8gO9NjVMsbkQ7dSlBwrPOf7+XkQlq89DztyPPGVBhqYjtFsZyltahcuxhBAJClw5CRQHaZxBP3Zt
PIBj/pwCkBiuzuColJ0uFm40pIjRJ2632TDCToyXRxWZA9TkbLMVulqTvvCUIIeNrgJ9/TUMc569
LZJAf3BLLMLWtS6K12beZ+wAKzBp+JBNE6VxjZlzQ6j6JwWU20eb60o9mfmI7sP1/3uKPxT7Z6xT
bW2gPwEE/WdK/RewWv7o19cKLeaBvGzzeqbe588AinhtUuAfnQflXG3MKaCE9zh5EeK/JThCduwc
iQ9QIpO3OMEfCaaIq90dmghhQc9/8o/Q+hoYdh1tCBlu3/K0iyqmmwDXEVqzAguCkIArMBHcot9a
FlqUxuiiXBCsfYtTmddvASHhL1Zi5QGDVZzD8Y/f9wKoD2TRrb8vOMFexWIvu6f27Hudrvlm+a8z
V+9zV1YH64IpnTBQIL5Qy0GbTpR8hms4T8rMq6B96zE9tbaataKkDYbiWRTmD4SOD6YPZwja2AL+
A8PIIpwcuRQ+gw3HScj6Z1dabFvZI1c0E+5vdkxcY4blqBkbTiS5VtRyuwZHTD5gbruE+l1gOvWx
wGz7nlyVseRejJFR0zNyETvJ6sOwcuCVOBq4f8cMED4fMZa/4kY2mhAxa5kO+MfGDj2yD3AnVOsg
HULIIJrLY6f+FOn/kf95/WYIvHxYnz72rqUw318RAsQvPIKkxOAQGcRTWdfPOuGQPzoXw1GdMm2E
TIrgICw0YLnxlwjssfB/bqbqd1u8M1TX1at0igmKob7uM8l66XwaiWFlavD8mTDUrWxBmKWDhgFO
+BpxyKc9RWiJ4Z5KqOikU5G7+5kfz7q7HjErxmrRJqT9+taU6SI/Ev4NFVLmt4TsTsqrTbLCdMrQ
ZP/pFJU+ZA7+5WLzNynqcBktgPYe0d8xkbg1putex6ziOTlzYxLEkzAHgcOjrXHY3s0dimhY+VCu
vJB99H/j6yQMDtxq+7ILfKv4EvtWYKBb2bPP3u2yzlWjY9eeWjVKyJE/GLsE98SY8ZNWV95Y4wM8
uGVkwqVB/iVXnhBSyAMfzPLefIJG0863F9LHhSUJbwv3hCu7B/Cdl4I52AfZVkfubsNJccCHzdYB
Ad6k9Sieu8j9XNNs6Ozl289YhE6eNL8SyieO0vECO/HilBp6BqJTNC7FjM0qO0xldQ6Omcm+XImg
rlLBEJ7qqZOY7/e3tPv7OxCnKw0i3mzJcPY6l/2qyVPRUjfTU+uUkolOiq/4uyQkzArnflKNkUip
v+tWB9tyy3Wx+wnxLhXdYe7Dk0dvklJCnff/0bTDTVZ/WXiX1oIfSjrFKUL/fknPynLVwmF55l5w
B3pr5CEWW1q6Ac2loCxRRwmfm2BBwsjNmCff70RpM/q/R78QNYi3gsde62ULT7bUl2mtVB91SiPu
L2RoDk5q659HFMEGZIP0fOZou/KS21Xw/7A87NRavTRN7SsfN4VAz4NgqkfR50PftfvZ12D0lHT1
dElsJRzvU6x5aCWuOXYe3G4KTwlkVk4nHuG89zoVArh38X7uaiT6+rwNnWFiMeJzm80prCvf27Lf
3Huot7ymIngtu4nhhBAwlwVQ6PpJeCSZlAFeqo2vrAs/u2O8qJ9qfR9df78JjW/duJJZLm00n49z
VldrVj7JRvciN9y1G9OmQznxO+tGSB+uBF/WzZKxWCfFVIEbTQwkB2tqnQHOb5epUQ4T03LrbjL9
rdI+yAXLmoQwqwwU8V7P1ri4ivW529uAm6LL3ve3IIvMH55oah9+bcW45Aunmyrwo+a9ADw3y6Px
jxZJw0SY9GQ/8+dPuZtC2rrEuu9OMhDvmCUjtfm8anLiI9TVpoO1EMZneuJCJhV/+iSqcImY68w3
0saRdRr27HlB7mVbpdmwA2VhNDLBMZT9161Asamf7m8IOfU3A3ksI7J+ZQWDVyaDJd2BeUTjweh0
ZzfHBEGRrLtZIisKh9iUrO+1/l3hmh8r48IeyMov/jrkpHaF+ybejvZj4Xy64MwuQnyQwzrHH9cM
OZUaKheh1Pb9TElLcBsYxsNajUywiyro4tY9H+x42SlBj77ogGugg0DkLD3/AiYy4eO7qppc2eix
U4OjXoXI9nimLzzJFA2O1csoGz8mbmwVbHL35pJwaXyjT4f9svGq9G39Sbl+ldt4qRPPTWvCpOeQ
2Ad+KWKJ8xkAha3rRwTVLeJnweB0Ea/vwScd1UKLOFhEBAQiwSimFw6JkQS3uiv8SA1+37Dk5IzH
3twdwBkrsglC2nAEum2FQNNl74h45yqK/o1UtsH8w2UMJWWnfovLaLdL+JoZF40Zs47zGKXtkje2
xEU1eS/o5nvT3OwUwXcOKm/UbgjP0Vd+cMSXhWmxxTGOILdzKptJvpflk4UCCz3MEzaEnB7rACHp
GbAiNISUJJdaJrWGt1l8Kr/fswANMCVZbdQ5otORWREz0ny31kBX8ac/5EYKLc+58XUdz4J4W+mj
8cYk7DzxQrzdqwVs97dwveitT1JlJkum9wG3vJpxlfQLJzijsKgEgDE4PT2a/boI1+VXiQCky66y
qvCJ9jR7OQH3SUX6Om43xiaFJS0EiuZlCx+WAJqQ6aO4UhA5BRgSLPKYV3nZTE3KQcRQGugL5FJU
hyfwxM4gRIYXfJ7xshgQkLXU4UL/jrFVRWVyf61RdfKIZ4EJivYRv/342Z8S468jkwbj070m/dGI
I/5ZZJJxpa5tXfXpxFa8DbUbyHnjiv2cuYesQOHbT78dbf2/xDbuoHX7VFRPk6tO2IBAMMBGTrWb
gYXrTjfEsMOEjcktGP+KD7l8wJVsx9qhnXM4LVT/2xBhDNJOJ5jSC5DS08mLyxPJ88+MRF9AxAdl
kvUFCwMNAOkRh9JU0hE3CkMgxfXh8X17AvpXVDnP5TiIhAjkcnGoME+DO97QLm+CZDhpMbcr7ewW
4SQ28iyX5rk5TKlmJuYXoILPNy5UYvY84wIcEjFZeFftH61z4k0jXSYPQFa6XZpifdqRkCWBTMaG
uVlkTGjmo1usftP04J2sVzq7YkS0H7sIJhnoy1rtJdoW1xqTnXLM9ge08baQXQB7tTv8pdxtoPRM
Vw4jC4rp76fLaY+qlbjMwP2a+ifCjrFyJmPKEAnabrHX76leE6nc/je4HwoAekTsWlb1oqAQQIlf
cppBhWiOnhGwMJhK6yTwkCOHT7txHx89NkO2baaXXCKJ+ErUfGOVu7m9n6H6ycsUDQ3xA32uKrAG
npk7LLKu9JyCO7x+IMzz6xzqHT6I6KNgHfkSyOl44fkWJaKtNCh24qNcYlYCNhKZP46XCXTD1UFO
lDpmH4SURc3WFnlHRVx9G294iVZlcxGjJwZiupuh4V7SNfJ1Brda/IS3aUKmzskNDejDXUqun5/s
QUhaFAzJibS47xOqvEak4E3Pc5NWFT3MBSMEpaDBoX/sknD/EEn6LsWI5kBV2i/5eP9wSjtx3dv9
VEIB3b2kwIUE6xNjWgA7M3IEibdZXlHvyir54ssoIZH28g79sl2PcjuSuGXLvSiR+oj/rpeZxjNS
8dPqEZO6Cvi+A3A5QsBZ6/6V2LDJvz95gZRs344fsz2U+b7uL6FPsVHz9mKIgQluyS0mpL+rkyH7
hgqBvJtQEIHOzXmq9T361ue75uxSWtGeel3uG2W0IEVW5BpnRaLdNKW0Mb2JqZgDWzajPh9n3GJE
djFqOJyK2SrrXp7BhHeOipCMmdfNkRPivhfkYcJYc5bBTT1hIMogHfbh97PphzhTDfazkV7CD85f
PxCnD6GnVVXOcFzv3lnay/3g+CQGpIQKXx8jaRe4dKjYmDD4GonXXlThh1nG6SIhUtnyoq36gzAM
iVGj8KSxJwYhVrB6nX0JoFH0PtQVByKjbvYVjNEYqdnmhHuRgmqDz+6ajVwAsds9VcbhlA2qzNnO
obqX6qNj/tnTJGTNiGesOAALKScCIvSHEEYjhm6IXZSQOOzCzcVOBVbrvsyPjBGGqslajB7+5ksI
Zr64/eVE05tALQ3KbqBZ50s8k/nVB34mFBfqIeNCouLHJDiE4EOZS+bInwCh4kNPzmLN87L3ZjeV
QxFefiFYxbJ25NgXMgNgIyqhNsATWKNrY+cQmBDKiUT+XQlYe+sc+0HiYsVusMwUb4Z0vT38mWHS
6Snd3M6VSFL0VAW4DdxgjcyNL9v7V7FWk71oGMPZy/Jf2yaiIaDH4A0QIP/7bJ/uH9cHtek17M7D
eA/m+Pa/vo59uLHwm7oietwvxuOJM+0vhvxGWXQaZL4tRjIWz7vlmwd3rBLEf3ugf731mMGr8RRp
qv3N+S0/qs0JyUK36B7xUdtOhKNOricxbmqsfBBOW5v4MUhzB/h+I5uVgFTE+Ri9KeeayZiIqrzD
UTZI9TwGZ2okEjNnxxyvUtxHDMVh8YMQImpkU5T2Rfqvlh/rC8ydsCURIVDevbK2lsKlVVKJFq03
YyXByuBKe3H7ERqw9/hOvwzIWcYazzZsBNqkL7iX0vIDZbEDaj+/678aTlYbs2UOdVprbbXnvh8x
1DxoY35F0gAQ4aAcM/xH5EFFWi5A7E2tq/JoM947Ax1hPT4bqaZTRBAbQJJqrrflOnzyAjtr7Q6H
8jaTpEiC/tbh8zB/k9Zji5mFi1g/xgl6wQ4CbwhXKr3tGKhJGpAq5grUY7SRS+UrVedjODlX03bk
efHY7pfH2yfcHd+ICJicWO2ktdwh8A/U1RIAdUR8yMdaermXJV9vOpolc7E+Ybcg5LNJUTXv9B5q
nw563mll2Ohjg/JAHngEhMhxBy2OT+vjWroAz1uexxaIvjIPM5qxt3JyEDT3NHQS/QjQtdNAb6fB
LGKTWM/TI5vL7rlchz0N82we46aEVufh/hntky/AQETLshy949k+kCnK/T+xiWfHneznPaYAxMZc
USRU/MMpxddqoCY3oL5f3Lhk35Qr4rB+mqDGmOz+PcQgZ94R9d+HqORxevyY9CfRWQGHxWegwuhg
OQhSpT2eeBjacicP7X2Xzp1KQJSNbytG1lBYJHFwEHLlNkj5n8oAha1fliw+TYjWCmLt15xjf+55
nUGQtLHuKO+t4jXJUASkBl+QNf54Ss5mnmPp723RTi8ZTwAeiymcdVi5xo2ERHhxcKoP+iJmVP97
AJzPcCote4Ph7+J6+CIeQrTeW1xbQrlg9L+I3BMJpY+OJJet0XFcIcXF+Cxlfywjz32z1toYJ4f0
pTKD8siWn4FB2GAyzOBFoa1HTzHAhiy3fW8dVyAgc8B/yEGGZnJmwGy4fVqaGsD1YGCWcM5J1QEZ
XeuWGDUmYg0V2HQcSObzsqrNdCNuVo8tpwo6ZkpVY2SnYtA70GI1oW88yu4XazIrtol/QBPLppat
p9uw5uIfVETsl6x+44QwDMLi3PiZnpFoVbO4hFz7xpxzBDg8MROsjaAQYoVdH+ZN+ICjqFTaMV6h
rCr9h8UAZIFqeVpqTuAIORlGrahd+0Avnm0rE1fT/lo5+QB8JvMLl9+EzUamfQMprwX1xLuzgGxi
dl3G9YyB2ZM0YGS0ZxplJ9Lchjc2+ZbeoSexy+fFsEib5tJgkiVAgltGxp8YhoQmSP5MHEBcdn2g
B6Xosy1MdUh21Z08hQRUT9hPxjf4MbehVSEgS1saZpxoXse3YGnwtZ6HFw5qfDXVvXQSiIuDUxcE
Q9bTQyLyjCfJg34Muj/OV/Pw0lj07ew0AhnQx8txIxvVhCv1xKu3GqF+ADkwbwhiF3DSV8JpJCX2
a0xmaZ4+ci2/EOBbFaf/84vBQQ9bsZ6fJ9xtEwzW4MRvY6AeJ2KqI4tnl1rj7Rg34LGkqTat1SGv
UMLq2aKL5vPK07CENPOIOdQJIEb+5E18I2ZiTIFQnfXukf9YNLyf5x9wIZ6rY04sh+wtQ9JBOF7v
G+nTUyM1UR3ulDaA8OfrC4KWtgmyAuQ3/rctZjorjhn9HTX83Ve1f2jVeGG6Oo5KMOSAdrjrCfX4
GpnsYUKbbm2SxIEPoFAoB1SpYHONAdDNcdMntQi9/+qEpldCqvyRkPBhVqaU/NkQXBoKk6zVURD6
+acQP7DrB4nJNXXhEpLPaU1cR4nNe+KgzBgiATtCqTPwawYwSctfCxIPpSZ9DJnq8IsmPo4LMLz+
VjGX61yjgyrrU48WNMjTt97w+EPtaeSqEEjiibLooPrXg9QmJHVlk+SwcjA1qmFI/6xGo95NnC8m
8A5q4iNHkQAqZCMlxhCgCY1+M0LYuNGF7Ccy8R+toJgeISxZWuK1HnfKLEBR/bwI06BgG/yklCoA
1eHy0T1YX6MakpTT2lmK5QpyowYE4BsC5zQEu0OH2/dDI/6aTorTmE3o2pwmwLn2a+qe+JsNxr/h
F25ZUXyaif+XIDkC0By1jIHptnq6LkGk359aQCpNM8RG2zjUZxpnQexFqiOkG4LWf61LsrEIzkuz
YWnNYSE9jy/WBm0jT4LKghBpvDqjX1P5qiBb+vx/WiqksiP08kw3uPBYs435fEAkeho/OuDIRgEo
IR3GMILuHAkwKfU6W6CrnviZ31RVQA7CoCCiY0UJgKF4O+jrC2/vrnbc+iV0FmF7OmmS3hVkDRL3
R2SBgdQuUYpyXqNBX4G6u19GlQWcBUYCJsWthZEOTJ24Sil/fEihIgg20wxSSAOZOFzCIzdLNeWu
UQeuwwdtzQHkMFfgD7BTMyGdgMryrbBRAEfEsmM9siHlXADyntY7y26bA1z1GljJhCatRWQ+joM3
vVT/O67NtwnlK38iCKRlJf7VWuUtpmW4yBfT9qnVrReFZW4lwakS+8VPN5ajI6/zaihkIvpsOG2d
iByIIgdPOEz4EkDzNdDSurazbMmrJUjQuCzhmftOfbISFxnU0nRn0zuHvTOkHZ/TLWYgjAHlZEmX
TVi2QdD4Y9mlFGagBu0PYR2i/2qybplM0YA/jEQzCbK9p1yP7Z+VXR+EdAEbjW2GJSqj+vGUDx9W
jNnOR7BJ/uHfYKtIRjI6oX1qi2GiXuPhZ+jHnmdCHi8TXI3HQYgwEsulVnAXM9NduosxqXbPgcua
BNKvAnebba0u2aP0eUp6ycIFnXzLuQlxZM82ylUkrzcO29+I0oHB7oLyUAioqeSodwVY0nb7U5xN
iwb4UORQV+UYCs8gsKhgbr+WGzzvcziVmIvkLnpAn4u/yLM+Zoyq6XxAaq82ziM3ghU2vTCwAKLn
LJVXKxggjkYvcQ0fhzhA7kUm1jRdE/O4XSkl2LwptLo7F5nQ4wFiUoRu2O8QOOW2V3aTfyskRaqv
VxwqTuJK3lJczhQoRMPZpk4RmhUXHT5usyDF/cOii6U+0vv6REwnwww5buS9TpSRQxaaXmnjfe/8
3g4kLIZRhLK5qFGC1k8Cjy9lx6FDOEaOaUofW4/Jwoo90atmLeH+W/0mLZElKopwIggXnzB6UFCy
hOAduPNBlJyX/hile+qPMo5KGDmBLrFhY0XJOCM7VMQuaazBLDFjQygQODiXL/YDLMgUdHjL2Ooa
JPn40YTx1WjqxL30QYwWRjRpTkdibqJJ1EfHHVUqUBgTKhwEIII4wd3ThOlVheEu+TMW9aqkz1rJ
28gVrXKjAmHEvUk2BfoogBeRrEtcj2AlsnCmtx/ZELHgnaCxR6Uv4KnHw29VyV+OVkPj4Fi4HhSj
GUcawRtXONMshuMKE4jB393n0soLnqGXfWYBrGgoOBRuzuMMOkfGEygXjECgwsqAdQu47fDS1r3/
QYEzP7D3TeFgQ8s7YNDvgrvzBZxQMbyKz5XNO5L26NXMJcBleOGEfVWcUjistwsCoPv+4Vl0Actz
LuDa+4UT5YSCrMmIC+cQgc+uAR0O6bKhJtOCFGtPhkasSdpD6RG2MwsI62gUBrmIhi7pBlJJX1VJ
UNPwvt6RAOZac12qmUcKP94qR7Cs/eXs5alA32qrB+CV2aHvvkXtH/iBH4jSJizayPDM1F8/yxkb
RhIGYGVl+r5HlCr9/+T2xPCvpkmBaPUeMEQ/TUm20CJi+e3tc+MTNxaBK09GBd4Vk9G/iFEVgt5D
CfWlb6mZ5t388UUiaRlKoUSNZflYwpAFZcEFNadJh5Oh6EqYHGLGbrFow9ykSEbu2gp5HX2y3nk3
tKgCVIodtHJTxuiqH/lsNN6luva8q0oUFjnPRi5nDRMwbKHzlcv4pzmOTZyc6NNCwcNpQxW5y+RF
xVuVeI+eTRV9sGajKJCpcwBCTm9O99X1xB30Kc3mzdsPddZgKLrGmZ9W9f4Pvg/Eq6LDn/qmkr88
ehHInGXV6E+rHnoHKq7R7ePv5ipCdIrcfx+9VVC4rbNvmDN6nJ6MillnOfiQEvb9uLb7SNUAGIDi
+6efvXTDPzcpJdtLVFlFEaz7jJQseJdqpEDJeO5Qg2KEP70FXaZL4qD6jgWVzWkqbrRZu2JkECxC
Q6pX2MU4bfuiCw8d6oipNhNUP1wTcg+eYW93o8O6ByxZEBr7/t7+WpNGicisavUOJvJxZ1/XZpG0
Ag5/goRLAvYGyRXYZJGvYDUDIySlgeElOehsm/wv70wuDFGz7WQ+x/LGYiVQnXKXuyVshp+GxsKM
Fh6VBC9tp5LIJdsJr2UYQHbr26V6LkHsF9o+bQ3n/JWfU6NNvo8/GZY8G0RAcyX1woAMASLU/2R8
aEK1Kqnkc2qQp4NLmaTXnakHJnD01dD4GBR1o76sg9V8Tm65rD+mfVrp2j9vf7J97wyUuC2BtVnL
MAWUBZAu1esTwRGLS4Nfx1FvkDeYuQrkoFOMtGZya9hhRztBz1SFmo3BXxiFqpHvm4QL91HRY+Dd
kvrj/68YuHkohTq77Gp716OzozhQhpV8DHn+6F/t3Zm6dn6/a5xsGrmkiQgtGJqypLpQcZuBURTV
ukWZOWigkGMmrPLrtLTuFyxD4ptXMO8727P9d3eEpL09Ewwh+QEB8w9QbXoNDEcYMiBrtdyztd4Q
7JAg1VrK7azDV3yBqrTUXdHZe1+qBikiTKUU9iOMFxnjoQ3vV4gjC6Ml2yJvnWPkIoKsyOLeo9hr
A3R1dmwKqdeBSbGaQB8kZaSEy4ihaUwdD0nU97nGFrHglHqeuSU5A1JrNwL5HLAKXsdV9cxXOWkO
1hNyVm70XmGGW/GaIqdL9OcNxLNZMQwcc+vn6r4pAC0uQ+2CWvvG22zt1b3FH5gNsvo34uvB8Vpu
lxJXsHYg4VawxgvyJ9HEYE6qwfrKv4H0tJUcp9xn+SVO1jOKhhcypWKk4/cyP1hBCr+j3kMV08wa
WtavAAyGzwPl4KUkWdp+9gAcARidPKhDfopwOhYi7yIJurDYj5NRvZyNpUStel12MD5fUNVugvF1
JYvyJBJ+T1KEhMBR9V+XbTQhdusEEs9aKIzf0dWXO/THUtj99MNRXqnGln6rX7JTVzveqyF+xLgD
Iq0RG9Ir0B0uEEN/I9sy0WUlAQdvEIjIAACgPSlxQujdIeoMgPJ5J7NBzSsHU1SMbxPK7ZrHHe5X
/buc312Ges4kyrnF1n8rvicL8Budg4dJUk5q9xsuIxq0ymaKNJ2mtU3ZHdS0N7yqQAGt5mx3bpRW
qQnB4UMP+TnMmgBy25oFSBhHEStcnJ0Z1DWulJiArK1PTFCpnLtR/PUzlGDVmxcZC7RqZXuZEFlD
dX0bqFV0gEYdOG3/ZKNrvVWG0enKIU+A16rKfoiJVUPQ2TJ8p6rEbKD8MFvTbkoQQgdK2llOX92O
lb49M6k0sRTPv2vssNouBUdsVoLyKOyn0IXe4GXYsUGWsx4Ni2+6RF3uu7jVmHVXBp5HI2NdwTvt
zTarE7oRzI1+AwkT1hu2Aqp8cxU3rJIbyLxk6cY487nNGow9CNX6IOmDHPgnZ9g0gTmjSpBM3x0C
tiKQj+Bnr//yJngn34rb3t1pizKHSaDRtzEArrtgkEyOf7kFIcTRmtcV63xmbm31Yo4EeOwTdKGV
tNEdTntcWzLyWPjSaOmhzlOGKQ0GsIjKoX2hECgs+o/ZcMR2j0Tdwo+wkpFEnNkWu3kYdWZDEqjz
oMARNIrZXhuKomL2vX71SrLN9778QX93KsZQML1wPuhxlXe/W7QlJGSP9IPPWNAXXRLkcx3Erbnz
NHa8S1YqNMjFCOwNHI7L8B6pFBwTnWd47Buazj/iHRKWI15SGxDrAdzDiXoWWJjFEHT+A2gJ4TTp
KtBtdks5b5UrE5WRHyHPhr7NkdcdZ6wwH1JH4w1s8fgTD8+VEKnAeHYbYjl6Z7xxoR+ep7TAgi/r
8n3qRlKutyyE/Zk19KPYceaQFxmcGkwLK6KiOS3M4dpjSOpQnlF3g2zBHdQQfJEbFNZjOJTLKUsc
AO5FvQ+2GudXoMq5BDhMRqpJdPXowvUQrD3QLdpjpsmcoIcq+FbPZBGEXLA038P1BHnnwKLd7OD8
iiTUwiZ4C9z5fotFPS1R8kxhPheFFWbMombk+f9/oV5yzVOrf3JlSfpOzAhjBuVqwSfOaxOiPAWT
u9wIirJHIqQYrudm8Eqwj3gBEy7+wxqe+GTNWLAD4q1CLXkM5sBvkPDbQ96+gwx1e9N9/d9wK4TY
RLpP6gI8gFmMd1Yj4Bg37L9B6T0JNcQXUuq3POedSrQMGcx7mJr7nwOPNoqXSNEnVn6e7GdIct1X
rqO5BMfuLe6W6OFWKK2MqRdvgBVbwtELlAsMas0wfueIYEoz+giQ9+o6647GJ2M6fdwWKfdS3EcQ
7Z6aIe0EGVk9iRQHWR9qGsxOB1X9xeNolXf/yUcBvwjYBOy0eYWNqtzrj39pcAg22QOSG+X/LZ0b
eXSUSxcfz6iZbQjverArTHtdb8Y6jhlpAWPMWLZI6h/4TwQ++24+ZvAgCIQfEfOaITg7dneYL0ie
Moixir7XUzQsXcmGF3qvjKmF2kiYQI4q5nT74u2fYDebzcgafcZjcDleaMpEYfs3GpsigQzuL36y
bvDCQLl/m/KfFn82oxhlabXmfbcfN9u4PBSwR+eD9rgFJQcuRyvsP3J7LOYBtpf+n/SMgCsvTebK
MYLXxwnlwDoSaxQiGjJWJFC/Cxiorq8124E7MhYgltQbzbmGM41sDO2YinPQu0dXDEPXadCWCsad
pl4hg5oMwxkIFLfj85McvzTTmm/kpt6X8/Evf+sgYWcWMByZohFZbRBGdQ4fR85Woy+GcHB6kZTd
ogNgrLq6oCcYN133/8g6RB8zHIve8vb9SOBBBwXX6DNtgJ8M2Z8CfiC0RaJ2Kj2ypICc43ViJpvN
h+6f0utud9bIowH/kE1wG8W8BEM5TMV4tJlgJflDT+sPQBv9qm+KKL7CwB2mIK9QtocLPLjeyL7e
TvHqg8Ddo+M3o9UOp3wAWWJ1wsb+P3QvhcXH9JllTZL9xRGYa7WK9heabKtuh/qHWvInnCj06Hu5
5bXPwC/MNNq+yzABXgmzJ14TJ4s3e55O80mVpJOoK+iopePOQC8Yqh5sk9T0eBWWBVD1wzEZMM1I
hbnshDe77eoolX7CNT4zSC4cLCcfWtkQXcVJ/uXmTG+mTGUnbDQHuQqmW/sx0wUq9FrQL1f8k/Lg
L8MqJDYfkMmJpVe2/hueHHcoAFVq0MtXmDRH6DHINLg8nySz5zynhia23+3Giv5TAcRECMrfojcV
yMVTCd7JQIb6TBCCDmwPF0j373FyTnLHVI0YZ1cJZUfyDnyqz6rbb7CKaIVTrRGWg/qcYANJK+pU
my75xPyYSzipeh0fLLKYCiLaYPpWfpWWu8GLWOWVWNHW/euNBg1hm52hFpREnKAR4RqMiDObnUpo
u6IsNP8OeJH1Ao9td4hDdsA1bv0gQ2Ess2yrnRTtqBDBRRhXMfoX9H08cmmotwMaJdS6gckbwfzR
3Vsbe1S8CAFoFJYeJ9oJHbvsQAKNL+68peoTmMWZw3GBMNZ2BLSBNI3q1+gT7qFNwX+femn13bqb
HgYQJEGHQmLmFDufbJBjJPbUOiaE5DORUCtzkdj6lXlUOh+ZuKwY6XJs5MNxgjqPr+jkfQXBfJwE
8ZGnM22BTQMwIPfwBOrHLGTjure46ZJdLijOg/glPg9rxZqF4P/krm/HfJAb+L22NnyFO5qYMh4I
jFdpeNM1T6Jq1MDLJhXZZD2YfpCa6OyE+5Q/1ucQGzMw0xfQB5GFmU32ZMLucTNtMtzPpoLuYZdw
QVNRa8DFVLJAqOB6VZ5umj75UpNF/Q+bYBOVJjRoG+UD6wCVR137Cinawc6b1mojcqPsQn/efGTv
WF5R1n8kMn9vsOJNvPZnY4GjKPt+y6U64l6vv1QwTrWDj9r5dz9O2/7EYK/4FurU8/cRfPyCqMMg
aWsOEH1uxcCbzOIf4EHDnqFXFlOK2/ODxKVgbeUuso0XzF4p4LB0G3T5dIozgxIsE0kJ50CORJzq
ToQ3zyrtPtp9y3fu/IedEU62SfO3AbrrtDIfollpQ1Y/QS6Liv1g5p9H++ukgkA1l746VH0lO0db
zcMLPzjscuU/oz7bKW4VRKx0Mubhf0Ir5pKHyg6REOsyv+bqxPV9bUIC8sZdpTSEB2E+7QJBJV8z
2mlBf4hQEcR95yxNdalV1LIM70h8Pg4Wiji5EWrqamjld77XXTGgtHCHdBX7IafRiE6t3f4hzsUU
PqsKUUO+sltlIy6hAI6NIqK0yPqQ6qoa36eA7Uwb7ooUudy3M/XWd5J16HkNVc1bfAzxWSmguzSP
kYTvlZCd9EUPo8qN1ArActKVqdD2K9IVuStKOq+i+4X19EU7U3Uo2rJnxr0Wm49kY/wzXyd6IwMT
Kb7SMWk3LiSSv31S9BZkK45nIKXF4beOHPnwM0RpJl4WcHLdCc2A1hgTGE4F8uFz7B5VbcjD5aPg
grFCFNQJY4JkdoZ5q9CGY1tafnxn0tUms1TZxRrOcNGPh2Pr3Lmc/NtQi+EPEp9i7DlsvzEHpr1S
zBddcM8KrWpuXi9NoLfLG6TSiNLbh+jm20quaVUwrKAEWBxD3ueZeP8ybPT/UVhR3mMk5KMvtIy3
9cR7WZmeBjiic8u4F/6VPhbGVN+tVbu/j77Xs6URMF6Rr8nTqe3TGsmGxm2+ncUn+df438/OnfU/
MBih6Yzg9Q5Wfp+ENOfuNG9niCScRRQwtP28C99BeuhILeX4AV2UyxY4mqxJe0dMnNxvHQlatwRL
eSArVCNaMenwxDS75Ayg449/IEJdroLkk7z5ne9wTBzrG13dHcWrNYzs+Ksdeixs1le+AX6/Llaf
aCsk9wLR7yX10pyZyhK/OpbRDH/X46E4JZ/callCUtimTHn/sH+p/MY98P+TU6zO/OzKeVAiT0ph
zKrnk73NvkAzDbjO/t9j0I1JB2wWxgtkQCTgClxRVQEFdIgeL/TQPGRSgNl3VeznDs7qpm309XvM
4YrmuiFkWRIG9JZ2lLfvHlNdPNpXii3WDJPsaEWaihMRoTbLix1b4Toicp4QRawwziw3I7Du0M70
y3zA74Fyt/K+eiUnGeIQaf7Wx09LqQFRmZJxTw0ivo2JSrC8hQgCYzUsRe3nyUzmhOhRyZpclFQ+
a39/SvwwHY982i3kkf2TH/bUksjkoYdyDdstYjyprqcTAZElnHs0r7leAv/v3YnA7IBPrF1uZdIB
6PQ5Ot/jBp0dYsmwnlXIP1pU28ibPwwVlEaHUJxe7vwFX5TwmjuLMW2Xdt3bLN1n9beF+MJ4yVCT
FF395CjOZBK+7vp0OAXrkpwJzIuJxjzX/8lyH90staT8F/4VaTyDrZb2/sJE9o20FyNCUp6tgLhH
HzOYruDAw7VXsrbpCpufakOGnucosZ7kk9C3Rd8zpuymh/GsW5d/d1P3ZSUASsARUySgrYn5Bjwv
oz1j6BbbmQVbEdEYNpSMvJ5El2oUtu75ED46/oqCqnk0KLSTQpYHZHiy4R3EvdL9npTOpWECw7Kl
+Vb6CshaQiVVeAPtY81RQs04cySA4kP4UaFCyC3qWXmz7JOJXQ2bNxB6N81S8ApT0lwGMjq+puRL
FF9wl4S4iB7wzAve60+1TKUln/hQuHFD3vBCllJT+mSqdoxuck+9p/gafcBJuie9KWAbBh4CiFOn
0z1OK7UBUeI+OGXz6wXUIr74T9r/D69a9kQqW7uLn4zChI133foE4zG6zaCBp9emtYD9r/xFtMqT
PWk7YfUDWhOx42NsBWz0z5fkroYFvc3aqMFKq3VGUoA/h3wBaKG60EwEnnB2JuDki313LRfqaxw6
r3ZAjmUU0LquVS98t0nvhh7+/u5DvG/wSLwOwiS6inam2YLVg2wqTA1doMvVVI0MolecxfBO9xGC
mjPiD5w8gUvkeOHWwl9LzavfrSzWQnu5bq6ufUH+YvyuzsusSE7MZPCUfrS3a9XttLl3r56k/ZqR
rc576ANAW4rhBhavNui3xQ9tE3tcsEdfJD4hTSDXmD0ig2AVQiCF6bkqAMrruPOL08VPBsAo05FF
YkcXmsw81/jzLJJCB9ApH19Ji8cS/ntq0NT7FAmQefhPNqTHOwT2HTVf4ll3zWrecWrLvKlS3/ce
yUDzUFb9W+gHDruM1A7wvzPrbAJqjIMBbfM8CmCco2cfDwqhK7DMAEyGnEEujtE5J5nue0H670dV
rKDulE5v/AoUV7hIh/vKstTdP9jHRvGXIEU6bNntxGlJzyRCho1c7cmv0n1o9XVwvkqTGsJwIBLM
bygVeAzFNHaygCvmjT+YN37NEGY+DKu3jSYNx1jYrsR2CuaRdtIE/RE7kms2Zlau/ToN5Asjsj37
dRIpGgIsHCbGvRXjjRMQOYh0imvN4ZVzKUaHPmISKX99FX8mK7XoMqsn0edVy4JVWomDg4Cq6+6Z
L/TxaGhFiPTSLIYbxDQ/RAcldwICy7KaQrmtCCa5JigiKk6HvJzl+ANLgEPw+f7I2jAn/Wh/QMHs
2372wlaaZHJnZanYQr/iBzZbir12zxjLBKJE1w6boGBqYf8YQwuqlJZYMH+KduR3Ox9vSgXN8ST9
9JWVlC6l3hAE7x8qsYCLjQzDtmDF4YP0DdDitL4EkqGLDiLOB/aJ58gMcdkHgakQCMcdbrgyRmbp
GN2OeLgDiZIfe+IPR9hwlJjmsLqYX4JOX0fRsunkemGF2T5Ws2lzDPWUU6D97tqwLA5iwCIguMAA
IbRsh87/UpxUYfYa9PSLN5vhydPXxWmafs5z5xvscqbquJU1M+L5Nfw8rIyoUUz49bh0GdnwkxW5
X/m905B1M2d7wrSkQiJH8jdYIbu8ViOum8KL5R4lmS506RsQdk8hHYPbkm/ZV219eYokEqaLiL2w
jIYHY7xVL5DfV4GLaLg1PGBgRz4rqfqZ/a4eeisqai9hK+Ch1xuku+hRKrCgDQpUyBlp8qleIeTH
jBn3QPl/HFtzWn9C8HEj52F8xhZN8AWmUbVbTePdTKKcf1fqbTnLcVYxcEoXLh6VqYIqF8i7l3fH
Vq5bavnDfWSasxkpT08XlhlB2b872a+TmZQO4d123BBY6d4XLcwvO4lV0FBp2bUHBdqP9x/oEuO0
s0so/9VlQBPO8mWI70sM6gh5KtRWwPiwF4CA96F4YL9umKuS8cx9MkmRNryTL+KwBHtl/gajWtTF
X92WFuDn1NaC8JR3T8iT7I4rkg6P6ud2DeQBuZ5MntEoedqcXh9SYGLH9oIl4ko8GPJjLGb2BMKi
qQOjSp+Z3uiuyuKsPfoOoyWdFCVvpsN3HqExtK/sAD/R5RQZaSY6JPYo+v6rzEpmtimkpBW6ip+G
WJP4CDM9y8vvtwCLmXb8sNKBsM93HNHSv7Gem2IdLZAMC6m9VzTfAXMtfLRIzcbfKAw9XJGytP5N
tiQT/6Jtq2Fn/ooOKE9oEjd0e0BSRsT8JceGx3gnqU6VrEgfUwy7kGjrg0PWVnuyPsNYQt8Zu7aD
Ca//qUrV8J2dgS9PMaK4QegToZ/Hf43ZHV5fyCQ/1Sd46FSpKGhPTnDjWnIf+3BK2ty+0i/d4I2L
XT0LyfLzjqXvSi61KY4IvNIY2CnkdL0KigtRjwfgebmag0D9tZDK7clSALI6edLk5sFYt7tZGw26
bktg/RhuOXcc4EJ4Wr9v6iHXRbMN7EEHTHn/0nJcCI1spfKIR/e9kSfyS2ECr9E8vPrIcqveGxy3
cT5hmGyxRRIVkr70Aap3vFrSja8QZS9Njp3h356FPnSZaSVfQ0bEaleu0vKIIW0IKLCX+ptWTEY2
ODdtDuuI6UTbj5GkFQ+yK79ZexYvTdjVRVnFfXtOZAlokipFqltp0ZAp28nU3hiR6MVNqqkGgiw4
hnXuMH1ZHwSx123noOgElUycLHdQvuCHZbuWcOvo8LRHjjJkRA3xznAOJoaMO0on59nI/m9HmHxd
GfR5Z+pymOYqumQW//k1u09dHZZeCk7q8VjELNo3DS+vT1WKolDJKTILXnAIl7jM0/Xpr4ypn8Ng
9uz3GdXT5HOtyhZmavxa/eQuugbWm2o9sohzBihu4lw9FfHtgNVs0FiOLU/HPHb9VLsq8VZQH1P6
iRBszyKOv45SDqXpq3rMsB7sToRzESprIk/MNt02R7NZ3LaDfiAN9gEs/QQVNwQsiSvOTOPP4rov
pQifbfW5+JL4xVeU6inOo1dHBpiPm83V9+7qAugsJvQjq9D6LzjSwB9zR9YTYXOGDx6yZFMP5e/E
XoVZHZygE9vOsNcy19z/XsMysUdF5wS79nWhXgQHCWy3kapUaxsz0WlB1bYk2NVOWOCpFj3VP8/2
ofid3IV9Ah7wU6h0aL3wb5sLNNgBA6HCP2gP8Men4OxRnQsO2cT9LmLdlMTFWki8BZWVNeRVRYBd
xOGkhfAuX1THUc+LEgRbAZbMBlgJ7Iqa0vIF4laLgJf6WcgRILIFrcc7Me4CJjnmSQ9c6mdP+XWx
rYzbDm8cvCnaknW6y6PLsm8WyhmTO5QFFUlx7qtWn5ogQjPt9MhsxwzIVzodTmoUes6WGEmWUUH5
iPPQeQsYUMEmWcGPHK69XLVN2HpmexsLSbA9LLwySpcp/d3SuSfZZ9kuzfYZ7gW1bY++OlxqyHbN
qXdkgqtdNnp7zVlHnKDKYaP4wCGu2ASLDbUIA/7piwqRzbFY5Q81bHxd9mvxZpTzdiCvDa9x2C/e
EvmKPMhDbNaPIJw9EpKseKE8vOa0R6em2cmEcRhzjn6kSTk5GmpRTNENzDIYQ8Dg/u39Cfjx5guI
bhUUcAXTmSAtqnDtNUb9gcIJWQAfHuSLIehpAusilz1qzcCmsULaHJiwEbMRQrGdDNac0M3wI72a
RQGZ2kEnljTro3hv3rCnZRiqyfr/pDtNj/o+t+eyz6S8fxOYak5gW49MNO4dcHrzvRNVMrxaPQhn
w5ApJvc8t8PPsZQi8XDfoR+UAfFKqDCJ2vHpXRNkY5iypNSD0K6QvOmfvUkrta4VPD2xTYzFk8IM
sQg1XqjbuJ499V+INkssI2IRLSFbCxmU3NDBjhlKn5rSxTe6YMX485tNJA8kfjV+qLFsQyyM+xGI
s8PvAMEpc4CaSPJ/rv4AD1v0BgveT+f5Pch4m6WMctiTu615FKzULtdAAexa3wQnqT+JQEVJEdKD
m8Bk5hH9cc0kXTYfDmHKN1T0ww5szMmZMe/H9c6zMP6Q/Qw6Sqmm3r1c6fuRoaMc13WSmJYB6aBQ
aJvgBGkRP1lvxPlIv4Up0z1wyPPf4Bi5667uxZ5wunPokJFpTRNs6s4vdTPe5X1ouS0LtOb6NDQV
rxnFIk16EcAvm6OdepIWAsO6Ik8fSs8jaGiEWo9oeUwaBWaCrZ5AoZMXsGKqpneulhhesPajXGhh
ji/jmHFpjVtBi9yzpOyZI5pfMOBuG6vq0FkUnS6O4ZzzOZt4ht3hXPnoIuh2m0D+9k9XKEWPMNfg
2heYXgOvMrbu4rPy93hGXw5X70ouYjwDDGo9jF5T7MhaejGIHqc+a9pU12UFYEVSt5H9sm/jBekF
i8MWZMjbr2KflTrIm//TcrK+kFviIagPoSmF+JIphiqp3JzoBt8d/mQYZbtv1fBgq64UG7QVaij/
rj6k1aoau32bfl4kbYwyN/GIvDE3t7ikWHogl+SQl5K//v4rKtFzOV0L7Tuis3CIYN35mN3N+vVR
/VrLS92Ga3tUzoiq6Yz2y0YOYKs8gF0s43Nd0rSXruGwqi/yjAZCIGQZ/rHMG7C9XxPK3Es2EdPk
V3RHLkTLVnYZ5K3J66SolOVNMkHqNHXzgseVbsdtPw70pirvJhjNS37GBxY3zvwKO3PXbkf0l1w+
5kLy6BvH0DcAu//37ISkUCtBIZZxjPdkTNCYErWfvV7TKXhhVkLTk7wBBQIzKso/u0a92XzdClSb
8RkGourRx0R4s0GNWBafGfv2uBnoCCfG7emqDU5wXOhUA3mw6xetVcf2fm9BXiSwxFUVo3Ru3AD5
i+Vn3p7q9n3BM+O70RYAZ9dNQqnAN4LNF6GtllpbJJhRclf4KnrxJICcwzJ8z48UnCmNKetPfJPi
VjcdCy8VWFXor/NExTue+BCC4ymp2e8+iNh2GDVbWnS+EQN5RiHRw+DKeSWbfA5t+M/FUDCVGxLH
bI+wMLTmobr/Zv66KLdEMygc755xDU43VNMT04fyXkR67Ua4B8C+xaOULnYueJxAWVWFJFP3OJ5N
3Db2c9I8/pH7NTym8B5klzwqWzUh2l6e/3Nth+f+uMxlThOl8RAwvaUCPffej4XsM7FwUXZjhjmY
L1NHpS83m4xEIe68UW7L7crskPmMA4by3ngzeHV5tEUWTAGcURPJb6Z2+TAfE1dRAiv9SUHYuMj4
Ba5bfAuvMOJYxVQBNYinqlZFb+hObwPFDqXBmn3RpKPkX92NHNQAbPRxdszY6Q/k388/Ee1Aac9F
rArBoRFpve7pSA344iJ+QfB8jHJHQ9Q53cfqDEZg/MRq5vekuql8y76GrEZ706mu0uXm2x5B6YML
VflNJr6RWmSURHv43LHZHH0vgtVmcI0Q2sPQFPXYZupjUkZ0Vm/ajD5Rh64E1X8fhJ5h0j8cGq8d
j59qwKC3waOajJ0LyC6kxyQzLRgrD4DUe91MwSrWREQYQaHL1rf3ew5wa9RIIndInyCjsgP9YP5u
Vy9vG/aQ4d5uDXma5ldSDh8jP5+vweEkVrQdUDQQq6AWwFWm+YUvP7/BKMesBAfS/vSk0y7tUtUy
i4Kvv6Tk5DauTJrO2dOjG2RxTzh+QVMJzfl/tQdPbcLG6efN9toLkdAICDEmzQaaFg4sAkO+UeWr
va6p1SpBbjLfCrzZdhv0g/ggSnWY0KHxnlDfjKNcXJyaxL0Hcqorro3zhLTb+A/NV9jBvtykWOsa
Q9ZKIlkg4V9F400RFxR08sJbSD+9zCvZdirjgeNW/ZQDXQOxw1ghvkt6SstokuI2I+8X1I7hlArY
MMJfjtWSpbgILtbgnpS3555Xy6ldI1gqHN/IAZDhA2vr5wIosktDmoioz2brWAQZ3cM7sOTPW6YH
IAms+KmrnrNif+KqZwe3q2DEhGRR4bPcALzp7dcyFK/Zm0BOY9bpCP3R2mkSxBO7anNsAuH7+TQd
EvyMML8lTyE19uV6/EIlk9rhkd7i66cbB0GFh5Ahpag6+t00WG8uebzXDWIfn+6/VYDpiNNILDtI
ptkYf31qChltlypQVCXk29IauT3pqmAaAQYti8YaFgosDbNsf/hWseXO4+jCsQiGwWySvL1aiO7C
vU/Mue6q27zPiPWNsJzXoSn200zYzHg+fKBufugQvUbu0VW2Uk8AhYazHDch83mENPHt240I6Huz
18SH95KBiqk2AAKhU2V7RK4oZgobZ6Kft8gd5wj8ZJMxSR9Bvctgbfd4ehjPNU5fHMxQZKf6M20Y
dr2oNthJwOG7eCd1uUcIsipcsSw4rkc52mTOV2wAWnY1K/TyInpBV8jHDMFT08NfD0edd3LZbQc9
HrMDg4YsS9XRsBmpte+QIOjx2I1TFDSdtg8jQPZL17hSw/I4qA19aswV53amdTLTydVCWK3v+T+A
CDcz8MwaQYizghjr+4rgWablPL43Wuf0BxqF1ZbVvo5U6Gt3YERvR6pj1Op8+kt5JiSplkBUuSqK
+W+SSAOJJGtnuFJWrCZdXrEZoCFnCpcxdOMY6Zqv4OLNiZuPjPgo/YgDzFtji/GPxgteKyR3LX2R
ELyOv+GTRCbevbypmThYVYDrnh1cZkfvJ4LXU7SZ1CcOqBXODKEklaM6fd5uxUlwujy0Apb3KHfH
Y0nvbTVzn/y9WKrTlAZoz42ilqB2S9qQGhd/F/26b/Z+fIpHY85pkcRm4uf8OjkAuUEysolWwHSM
tcas/Xdj0OASdYnhXabXyrz1incrrmpuSy0h4EePqV4EeNMEESZvn5qg7QjqH+DQJbNAdP952yWt
zcPSfAA6EFUcXVGx/56dLgxw/TpjmK07nIfQyl5tXzYJYG1YUUvnawXs5B1MRh3gD/aZx+uU/7tY
0kffx3mV/FaJ58A7HrOuJ42TJSHtOS2pNj81HHvvKHCsz19NvVveVX4zkkN7K/xcrm6iZ4sV8pyv
cHq4yDyjNwN0/EpUj/a4n3WAFpxe6jr0QCOo1eN2zCpApP++WRkL+RCeTdVr+JpmqV0U9q9ZUh2n
Cyi4u/UcIaNEg2XxRtkxlJRla2XbXAiAilazUcx+DtI7mgZSEsxrHc2F+P9syms5gyNCtjWhswK4
7ZV9adsDvHUdk1kScs+0Zyb+gHPofyNkfCIDpBF3uG5/hm6uG0yghWgSIgQ91lyCnQByPIM0bjbf
D92v+Uhmh9ZNC8lOPTnryRj/vpjNgae14hYFvgvTwtvGSUoKmbATYBNXlK0yF8VNR2m/sYQqF7wX
EYg4X7fvsDPGAU3Jl/6HlMUZxEz7khAG8tt8kh9R0J0gtTN6MNoJ7JxlhTZE9luNAAMyJPudrAbh
AUPPUrg3fP9jJ9XCrtt+JYXX62CBtGs9LG/4sd5os1JzjYBnyfRuU5WL2v4hM6JTVaIznoEEzi3P
Qz61yJYYl8cYFAXqgHVSKjCNcqbafcH33h9ZNKwh5PbabbSrg8S5pMNiymm9+2scwXgMaHd69kOk
h9bNbKQgu0Y43pZ45UTJiNup8n83qR2gHu2wBWpPRWpfRUBMMLTZd3F9r+ZFZkD+k4pRm1VshvOU
jbFeItqCxT8iakEdOUIOvJi6VW9CJeKH/JAH2K0fm5uw9ekan0wD2wtmFDd9C3Sy8ugyDrqkMw1G
0lgJbvmw0ZXNPm3qwg/drB9uRmsRy4hGX+EIRPyylRdWlHtxqjpFOmBypmgeFgTaGGfyL95jjllg
A4YOEuQKSWawq3XnYV7yJE1snQ4w1pXWi29717ET0WM07C9RaEDd7+C2shE/eUBF/S1T2cc0CV5m
YDsJYsCxU+FV5pmU1ENRnQ6v9WXHcbA0V2S4Z6CPWYFd/lb0Pzl1ya6sb8Nkw9uep7UidgejxRWQ
S832WVF4nVlGh38Vh+r++7c0GexL++dmfW5up6oiJ7/nleAJ3sZCZJQLvpUmQdYbtSZX/3r9tpiP
LhBFhRXvQzkCo9r7yU5zHGd5hpb/SbA7oNaGpj+od+0Sh9JfOPm00N7dwUhinaQiqnJh3kss2fUB
Tqkxb+M6iLITRrFeKj2JCN/oBOgYgWoJsEWLaaPG4lJxjErWYjhFdJ0WVi+9hMya/EQ3XazAdAnn
A8xVxw4f/vqJnT/tTNUWe0M6/O7ISFr+bCNxOKEwByUI42B3T2x1lKqAalyHaarrs/9hq0QHKTXw
vH2EkDnUfnRDHFGB+/dwJ0FRrnv4hx0bIHc5QYIbppTnFlWt9ZZgm5KjiLsJuYMbIxazwgntSCCu
ccVFF1yH9f91i//SShfPo2hGdWleeZQaj6Bwgznqxh+yYxpWDz5tawsP8IbA9YHT1kNt6iAw8Da7
lxVwzm/9DaMRnW3SGmpKNYylJQW4N/D+mKfrQ109aL0xvnfOgEs1dtXIqiQuU7IQ267EoQ8rkjy3
7FY/ko+UL5jPzD32fOvdaG0iu566HyjZ9+aZudMBpKGBEMNkovy8hH5YpP2dT5tJ8o7QIPYLfx86
w/PYgeyZZDodWQ91qvo71/c0ITJxGjyx/w5zvHbo7RbFdwJ50guzRPiGHH+VNOWi9aUhlStqEF+L
Y+HNDgEuGo7KepPGRn9MSdwDGrEcPprfnDGilmEDQ9fPzkD1cG9d7AvVG/hjZdz9lXyiYlpurk19
TrDWAGg4lpZyYdrb/0Q/gX0OHvBLj+BCnFNw3RB8/OgImkNiRE3PK/V8mcmS1SjylS4UKCulKI5F
HAcPURAXlPQVNc6AY1LFkYmtLQL4hAPOuWpBsCzUFkCSwzbIROLELnUXE6O5DuAZ72OEPh7TVUNh
1MMAGxACPti9txVTF7ZJdJ+ERVNvpARZiA0I6zCC9BL3UiU3488TPrvweTsKfxpD9l/K+K7Q0JOg
55Nqih391X+JpSn4JkGPHr3myujQ1eRXSlluj8AEMU712VqTq7o+xfsEsy3RxaenMBsSS3GmH1zz
gZ7Odr8ig4uYS5mz9L0cUR383JNxrJhYnhaQsQwhOud8eaB+ysRoilyVT42rPFWqQFDzMZYTZ8f0
tDm0QXS1cv0Q/rpkoWMe6PIAUCReYBiKAT6NRvlrSN5TyvpT1/l+najgxciRXpoo7W/2v0lmuwT2
sOylateKMSlIWML9hoSoasKZZS6GrdPZUliFUOMh1m6RWoZpxdcHmcyhsm7S4dQImZb3FDGOwaK+
cJC7LKlfVBjhKKYLyr0lbLrlgvQdALYJIe6KPCFfMaSpBHP2QETxDL63v4dV4cv6dJba+LgrUkSV
7EkCGtu83RhcTYWtHGIcCKVSyQpf3o6iSIWEjyu6YZ17WPlnC6DzcqqD9VZg/y68mI/FR6RiaXzf
nNeKP+HUIaWMwUAO0QOj0Gg2RxP8j5O6d23hOZFT6vkwz2EHdRXJ/WO52sUYq78Ia+Y+7uSBhOwK
epus+yi7Z2ejU+KI1I3c3FokYUtvjpTwplA8WoqIcv5CCcFuJa5L9hi1qUnJPuq8JEmbsvt4lQaZ
CelFvSUt5WokQ19Zdp4OhV/S8ofhPfHa4DMd4YN7jMSMPRU6S+ymKXDonPApFv1ep1u8+vyV8t8Y
8QNcIstNDPxUKz+6HT49NrR78OzYXt0jx0PwcwVyDUFMXFUbtjCxCxGqMNBQ6Qn8kJcNRjSruZ26
TOofkmkF4ZBLT9wc+auhcmzAOnbNtjatLeV05RAr5461pRUb+vLYx7qpmSaT2VaPun+WGNIhNzfg
ygMDT80IdCFAT+8gqrIOiN/kT2e8vOn1DAE3s41lNFTmAH7cC7xtVSI+CV5NrL0jJI0bmRXcY7dj
YRVb56W39YTOdxN5W6kYeG7zIkkyB6tpWxR1aw4H5gmcp6gteQ1b8PRasI4OTUxUbAALNMC9OjOt
kMJ2IgBj5DqCtN6m9P0ur6mLP3NpPdMWqLVePPXufY3NBBTceGGtsgw5ri8LrZS+Gfkk5MrXjv4z
7xvOLnO+lmBAl+tz3sZuGdu4qq4QBSZAH7aR/615q1jwMmjSLP+5eC5Q+qC30soVqU6CPHvE/+IL
PTQpO8BBjW4W5W+lDPHgZpSf/Uu/GJEGJ9rgm74YQoM932OZ1dCIrgZYv+9uIQsLhtrhg6375nyp
OdKOUa6fR1/FiBTpUfaYUj2VgEZZV8MxVmnLMlDs2E1P3xjcpPWqNTX4rxFWrfhzz0Vs9xnTLdSz
Tr7UZmw8sVP9lrE8ImQvVvWqzvyQjiS5oSw8sIGVIAZKt/zyw06xWlD+5/uiGxIn7YdWeKzdwiq0
a71TL4NptZzpTje71A5qegH8QZcoMn51OkT3qK/mrkBHNiDYFHAMrve14r9nc6Za+qlfXeFVgspU
XZ18LCZAHq/8xH6LW/iuaFuvtHxg/A1BWK4AIYwcoXHzTUKIH0AMRVlc6W6mI8EN5zrz06nmhgLe
fyBMP+A56GFs5oofex3ZqHydmyhZ88rc+GhizxZhP6T+J8hULXfpZi7eO0k2sX097VQCIs8wpUFT
EFIJxDqcV/Yu+iPNZaZYDhxJFXaou4Zyy9uqziBcK5unSL7/4D/96furlqo1DfCdm76lOcW8aL6S
3BOd/sotQ27DF2OWe/R2rj31nYhbapSJA2O5MBKQB/WXD0n8MpypuV/4fickPUowNG6kz1DzmG30
NGty1zURH/F1JIUV1aQIgpNigTWg9UHiF8jOcmC4+qVJe2nBQmlWupCr9VVDxsFkxCdTZjBryxIR
d00ttYGoTNkkKLgIRb1t2Uyui1WdIm5JgJzAOAjZD1j3E57YNNIJ/7Xp9V4FiBVGx1DVWmnY2n/V
PEs238aDoWzXydO76zuNg2OnRaZoo0ltT5kTkubDNcQGj5UPggnlzbEmDUjKPSJsDUDXWaEcpebr
UMN/TH7FAeQW0if9U5boXLZVOjgiIxh6H4+0r9biTm1z6HNpEHsxj1ABW6iCxU2TFP13grzgfacN
BRK6bwiqbq/OAZSx6jjRi8XfE3DQnTEIuTOFarYBBMKWa+Ef0yrInj/BSapQKVMzX0SwGO3bkigy
XPTrppnSqPlD6s94JnDp670oYFqBlpWcRUOOXuMJhVcdih6JDySew/dS1B3xgBbxyVjcDXCfWPBj
IwLexMuhdSHSbQM1RyNr8GcPgZEQmVttX2iqfRBAVM7iZxOUySxHAIL0Kig0Lyhxh53nOVLp/K6L
eIWny3p2HuEWhr9DX2hf9nmiIh1ZbKNs0F9d19Hkuozz9caE1l4pUPx3huvzcKw83Ku7hpcTJoAL
bqOkvQemoqfBtX3AP10zcHtE4LtlAVg+HWBBwry0TZn1frJYL20B76x197x4M++NqTzOBqdP+dEd
Czk02DqdVCodp5Z4NIJO5Hw5vVjCB4oKRxo/3E350xcgeBdl4mPYXV0ZZdZ7Q9OQHhX1rgw1SKJf
VTk9DCVcvVpfrvzw/gSsP3om7arztHh7RgXbN0VfrISC/BMBvbLFyYj/38lO9zgh2opsPA0CXwm1
DFVPdRFcObD8WMLjfwOEVCuM7E7anUwh5jo+UwjFdPdx7YuUQ3xbbzfeH2OwTZGM6hd/6UFuYsrJ
eH00/m2UyBXFRGnF0fJ4ApuRW4sW1REkD3MPq6uUH9J7tqqXbTeoj/i/eU3dN/qpdFnaNvkEZZmj
dg3lXghnTXVTF/zGZNySlPC8JIwkysy47XbpkIGWC7QzfQ7xm7W8EuaeN4tJ1+8z7fg6z2ozqv/J
+VJBRCbZr2uprYAjZdg4pXzzLApy10BLfq5aNDYMil2EFh1NToHGiVQsOwGiVuNQEw04bEW4sUyC
HzO2hKpMmxC0gTqouwkSdNH5z2ACVU5gZ1SAGwwMjUa0ZqtpUDhCgizrP4o1b+xGsYlU+Z19+oQL
gTKdddO3s5YwcmDN+KjNq7iMlpXD0ix5KGfZR8mMFvPrwgcbDfXSj6T5deZBI+Es7F6t97MlVU+H
jFXWildjppMs9uLrYdLbAS2BpctaE9NY6bvWBV7u7iY0qeeHhkIES2eEZWS18zmiQsZzl0wpBTFV
R58mMFSAooOWbyIYeu/j9vDHIglqqCuCY37q03zuQXzLfBHCQrTot4PbcEX0mcLPEVciDDakh9Eh
MY5EdBLUwopQ23bBDAfui8T84yH8NTeZsy5DiL5aVTVvc0smPw3vXbo0Fqq3uu7tvAmjv/9qjN7O
J02gyXQV490vcA1pDL2rMUgGyXIGPFWoUwh+A/stEBfrhBJwRxhiF/VqTxEqk/59hga8RFVzJeRV
gy+nGVsVtMKPAWYwSYfeFjS/EMVlx7T8Z2tWkKbp1QcaH8T41zYSuvNd5cWOTpsgqd6iOXxFtpL9
r4NK7bF9XTrwUTYBXeznX19nwJWXVBjix92GCn7UIvLMs1C6Pgg09MmUB/XkQcyMFYL2GDsAmDna
lr4hnBp+Vslm3Ld9eJp5fujXkXO5xftN5xppZNJO/Hfu5ks6dKKpV6k72hQnIqCx59XHE1gQ0qpn
nkq5KR9X2mcFG4/1ZRMKNCqA3LmviCNi8mCOb/vKFOBFJ0W14k+86B1UO1EfpFBsrWOuXhDrQRUP
8dyBSoWzJE55lPuxQSZuY0+0oheEyGBeDvtwdn2jgFFSjiX1RvFck9Rs+1/B5afCj93gtkw5HyJm
Rl3evWLQ527AV8s3sztuJec4jISTw04mz/OPcM8n0BY480oNDMy5UmdbrdARDEk49R6ZiI/zg1Pu
PuTScEYB2ro7YTJL5qNgYMO5tiKRuaDEy6nUV3KEBc3+kORfQ4A54Z75kE3kKjeEfgjWaPWvFbMe
LEBdU4Y+rgtnvdvR4gElz9cPFoFxE3jOrYxhhHrMfeEPu4u8ANSYgFG6EWMX82X6gTbFgA+2qfjQ
eXm81VWiNlgp2ZcfEEohrK1IzGVCCK9IXokUDj9ec4IN85OMTDoBat/eN231pxaVn4kwCAjEMJdM
aN3jFqefYNfcEnFgzGUCJuMxsR91qUoba5tnH+ouycGuORSOBKEGiCJYWxECmE+hMZg/9bP7IpOz
/+y7FN574o5P3qtGWiU5vovSJkPSAt61Bva3q5G3+WCISJfTlY2Qabb7PdKAelA+KX5Jdq35koPX
5T9mb1jbOY00KdBgfvlsWPyeIpo/1aUXnfMGrfFVe4UB60WHLoXB5VpPuaNf0AasjdTvyx4+Lsp1
Uzb+8RD9h/y0fjcy8aRc+zNsMyC5cKe+fbH2XaEAs2MFFDsRQIf/y3zVm709lk1tE8ePxpZaLYu7
MSWtERU7XHWWsofWGSZAySodojGRC1JS0v3o45bVBkaoQSjlnII2y0Uax718MIr6W2NRgfZ255T1
33i3GjiVJXPd/ngB86/wyhwS+1HFM3HP7J3fs/yMuqgKqeSYXBVlF6WtSJxoTK65YIJfAUiWSgza
b053EhdigKa5WsL7cNXLSe6nOttge9Fw1uylUb6G4M5ZcuyCEghmt80IKTilFMeAlk4fIFs4fPie
YcrE7Ua88AoMIgjA/oGtxSqQwnXUiOuJyacZxkI51KmNvIGkKVVKMFSRXtNUO6LOilXJOmAHhCnd
JIIns/U+gQe1BqZmyM8gJfpSaj7rkPxX1gwy0R8305hbvLPyiHJPCSaHs1OhaTfAGR7vRaZUjIE4
trBGpbhPtCSBDT3CJ1jnFOX+n4+vpFvO5Cr3lONYkvj9k1IcAZNJJIdeSIzkg2wkC/cjlFNPtXOH
szsSP/XICHxy4mYWkB3dWdZMbX2nOp9Ua6bZtbLF6AXn5WmPLE7JuXr6ncycvztsXE/xTdgOVa2J
muWIhtUtO4HwRyk6/gqXKb2YOZQMlSQ4tKbhHEi+zdYxSCYFRT12R5+yHLrNLF5n4RULkJ4nU+Xq
xcgqSFMsA5OVvJaYPyZRS2NbUhIZdu+pKFCX21rwbb+D6ryvHZlDdxipSCPZG65SJ/4s2D6sx41Y
/3Be1J2NezVj4EJRrjsH5sR4MioioICpFbkqi/+Ug8O66JdbADQcbBORA88AyUJl+SRmKHVL+QEP
jxvk4BZDbmDkEz74WX06cy5zIozxT/6PyAHD2M++8V48/VbmDreJj44Ndzz9/69ANQFXDM7JuUx3
RM9FLKbIrlBcra60mA3cTe6SHI2ArmzKyTgYFgvKn3N+6UAdS5eZ1savG9oO9m0qWTpxkjB5/mVn
I+lMUASj83jIO+LCHLpDCEnPLgeMaTLh4eNt9MO4MRSf+OkpgkRA33QBu1BRUiKRFU1ZilFpip9d
AbD5IO+3NE3C8jXof6i5UlNW1ewygMrN6Ei1CHv29INAez0FwhA/FJXQvPBv8geSviu+Pktu5Pu/
nsnWIhUaHc9xwthetH9yyqejrG+PYJT134Vd6R3QanFXmTGvZhlUjQILAMIEboEsn3WAf5nvdFvc
P18hxcwelmpMqNOaOAvmcO2boUR5hjxVRYefNkjB0vDdWOFyAKjq4bWx8VBZHtMqrfbGH133NaSq
jhUyciPMInjNkcfyQkM2Z2IgqS9JOMJiwzD6b7FdajMMWJ3MSFRoFv+Uyz8PNJcAXGvB/KEExRvL
PlDQAzfU38vCo5fjrjJaa5Yh5nd59CCfXiON1fnlw1F4mSfAq8+tBFZjN9dl4JFdAJ/Sr/IFGHTH
nH3/45+EtO7hHl9pJs14sC6TIhApiiQ5xTAPJCy0iaBDzbLOE+RRTLpBTf2lixH/iPTSY6BHc8Kd
gO9eJkB/oRwDXXy9QGdE/OOt1TGziMCrC/Cgt5EhTByqT1pVCISW53oOG6OLVoRCB7A2QU61OnWA
T2J4pTf27CGL2KDQx7LsV3FXKgMQKLyYmLWtnUNFSDaIqB2AavfJAeKADJW+66tXT5S6ro/g3L3D
q99fL2J7FhV576+BueQRmkDrzgA0AaeVBcLGXwkc3uicjubmPwg+5s1bkpxpgbpGJ909JHgKGbFt
vVQ1V68ThiLuxjrdtlSd5qJoS3wkVmXhCnWWjFoPfqtCbwx7oWgdEnfQdxBwhaNRnIhwUgZwCJaq
YffTf5I8ptKm6uPJHweGb1WnPEcxFJfssoArStodyCa93iwlTClgri1UiCOGM8E2jH8yd+DlPUYv
1S65PRQyc/W7UvV2uu7FOTNFWwWhuoSGKxmfF0V03fuMyVZvQwDxhaGFCwgoOCiKUgkL/sSLAWeD
HEW5bJrBF3z5VRbi9ee7J5p1u3DlwswdakpDlRZI9Tnzb/RIQvmQWQRU6iVtg9NDWgEEL+f/tlGG
7R+n+Flw2qFmbxBn4R7uZwYQpbiG8Nt7+KFl0nLlRTmSOWWS8SgHTt7DhI6cNScV3u7g4Wi3YnlA
yH1Nkj+L92Syg/Ku6zOu12MaYN+CCNPaUtbl2t9IzbX1NaptC1g68ZoXgPpSg3CfEKZ/diAD3O7X
T1LRuVawxkRTDCa3gt0moD/qpRkqJmycDvO4G2i8w8NRS0W7BWDjMPC0oH8F94yzpjvJmEDNHbHQ
VXjckv1TTrMKdN5OaQlNJrz6kN/fkjeHkAImhsXR+29o9WLcEbiF949yeP9hBXsb4BN1Y4jcP/XJ
/p9p2LA4yRGtsaUeCT0U1HaH15WYSJTFERV+WlwljSA4ErAscB6SB3Ql1YRoyOCDC2hSxJM32PSi
KJRcaToEi7/Z2WkBUjucR+EiJI04ELY0DxnezxQD75s5uF42J3C0PSBkEjnDXyTnBGOiKESHGBtd
uOQNaZtTf2lZYL+JNsVnGYJJSTYdyN9lXEuNFqB0Tlx0AQ7ycmNlBa1CDiIDvUAFnLg5r7UTlrYK
kgseafY4vniyZ84uzRLvcqRjqMTVswULbmFy/xaauvACgK40AN68uOpqBXyBzPrV6KUO3N9fRt1A
VUZGLu90VN+qCokuQQK5/6bk5GjotXH551GQiUj5oTMngxygx8DZuMTry/1IxKOUmqCmsKudbyrG
86iBH8X76jpHoM9I6XwJybfHvzM0KtEJDLxGmqw94Ykuv2LMXdTB+/163Abj85TGRGh4dR9O+SbO
NZIIRUWhNYyQg3HdFvOCpmbOIMDnzMuYJH+31C5GT1Eddq03U4hKYxPeilGmjouZ8Y8cqtaqkYYz
8xwxHUGPQALAoBdranocMSTnLh7BG/8DY/sqNz05LQ+K1TO+P4HM9M8FbBdXleByf9dkimIFMQuA
OK3dgB+98D1fSclCj08NBrwfyib4DFD0x0iLTFAsumJnKVatObdHanyFkvEWIATp2Rjv/dAEp2gn
i/43ErywzzlVSizE/znjhdKRmtDvYadF6m+Jqxh3TGM7CrF/8zcPRlQdOrTuOyVDtebp9xOdIHE1
FFD8yt+c51CtvG/7hh4cb1G3xTJzG532Df71+qV0sgRIPSW/o5v47M2kcmOubMXzF+6uUYQ/Vv4D
CW5j+SvBI2AMRYyuEpqffXHTcnc+lghdcfaDFxy/yB/c0GRwQFbVFM7pOxpx3hedWVhjrEx1tiPZ
N3ZSAxvn1AkpZI1TuS7EFhxAF6s3GIV5njvpRGoAcZhoVZ2Pc9J7dQ37eQmL5h1wgC07Kjik4caV
KAi0daH2gjjXHOs0y5l06DpFei4PueQ/OYg1uoYzTfKuwwKCGMGp4w69tcpM7/9yq9maYiysDWe7
wzFD6eGsijDf3wxie18LpC1mK6F1uqDQBJmlbmAFJcz+HeURdfk+/lPOUaUrLEK2P8u1OuuEC5+d
PSbNWg33PNe0hos3pHTYCKLI3l1spp3GwfHEs55cy7UEDV0QqwgX7wksgkzc/aJ7Kjzcwd0BtKzU
lXVfncxHXeUEUVcJHRH9SByUxVcswNaU5UBeo5Axew/ejrxFeNF/GjIt70X4uqEduHJmDKs+fBzt
cz93E/xsKr1yAnBD731YwvicyTdxTG82T6N5+GoLYZh8b02ZGi9Wi+FhswFi90vP5EmyALMGTkQ7
hxJgnBi7IrQbPqwpyf+qTKsB2clJwfHSUN1eUDIo0im5GZiB44LR8usI0fXD6hUfQRu7BJiHUZSn
/D4Jdv5BL73o4ek7fZ1JvxDHcy/FpgtYbA5EdaaDq+/s+PMrgxRnW4EaEMry3yx5o6KVCRrEyAZf
GNHFP1uIIMb8A9ZFnTFTgZD79OPX/lf0DXTPpwYmGas9p2gB4k10SqsJ5+aQTsH5wNjv29wY1+T1
MMFtT/k+Bo/rYwC8O2dkH6UnlSe28fJMk5oMR/OIEe9N72DxqkEDVU53tI/sDxXMYLW416dD0ezh
uspDHXW9KorwKhqld5FyYGmTIgApMEZB1KJ2QYvYGY7WI/5E41i/csiFvuCKIkj3H3N4ly0G4eRu
+2ifes+GSEQNjBC9wcUnKiZ9oSZB7PqSrsI2bHRrQywjMQ0uoOPn0eIuxy9hXw5FJ27ct1ez5i99
HucgGa3FhUBdrqfEGCS4kOkgOGK/eLLrklEG2kQomuwG5y1u+d+YpZBzMotvwVB1dP2DqeJ9TH0x
25uNK5PIjjCP0bVKKGf3LxF0jCv16m2cVD34kU2/oPKILztPpt/V+wLlB3oiT+NZqdk+MfVKGBOL
1jL34TnvXiXgzcdifdZSexIdprdNqxaDIna50UjfOA2AQUD/UZKO7rIDQdhXhV66dviVcjTc2F4o
DCx1kVv7GKPRf7MsbtN6/eX+0rvGHzEYvkr0pM4uzvOmq0emHU/l2nfg31qvxBWVigf3Mc98nAPr
qxTvebbtvv25IImQqfsbngmZM/oGldY2Cz85+di4WVx/vgPWjD72AxP65+YyBQOU5+ypS+KGFfGn
ccDniXdc9/n/6i0kXMV72Kd8xvSBS1ikZC+c0xVDOQMUUZ8CvV7mR15PIIyHflWLmtJH/B6g+F3z
Id+mQRxc5dU+v35mPBA1tdULPKWbYuXpIfnvZjWbTCp8ILnwBs9yrH6W0TngEFc7Ra5S1jfW9JRZ
smUD1891hTBx0pNHL+Kl9H0POiiyKsjA0CGhlPdsKt5bmKQr3xwAHr8AXrUvZ8cuu2jZYhSDLM7V
qBmtEvRkS/YxnQHcJmWOgm4ikRoRJRat27YNs4kKSt9nYT/0iwJX7qmgdtzID+Aa1pp8lyq0TQKT
zpdDgA2Fd0n7yim7DVm4NKRJYRG6Js0MiCMnqSFZl5Z1JgwQidj7yM9R78bcVtzPnKQ87JXdcElb
p5b7A6dUJ2ixzQuS2mGERJMHFRNiLp9zM2TP53C28MOog5ATm843xJfVLfoxYxy7qzTs4t2KlqKc
jYZKWvXgmu2lBALna9K2maJlJ4+L6WjliWoaiTgANm0tiff9ycm3u1JzzcpX7SuThi+R9iFUWRNP
RAY6VYU5u3jRNBaf0K0VOr0rstj/bWIbZUchibKMTLQG3eWPQs8ubNnIPp/Rw4+kCuaaGTrihisg
qcogUxAh5k5P6UuIKssiBAhwqW85qQtblQeFPXyPp4wrbUU8aqwG724NqAFp6GzHVHBlDV6w94uw
LIZ9QESK1vH59rx2YYOxiO0jajHnaT8CPuC/VG5eG8kXNg55RpnhRzUk7CbazqrnEgbMyt84POuL
dYP+YOOTGtWTGHLdEnK2AZLftVJB+NpRGwK9z+wfvCGWgdTma21OxBpQINnveWHCOzOdrg8KYj5B
L5uzr6nBa34F9Jvy2dnH1H8G14e1snFjGPZBUEIIvBSD2XWZiKnsQLxzKHn0Slz3U8PNvL18anPQ
xlbIT3CuaVLs0pJ9wW9evJD/ROjt5DzO5YbHaovGH0VHm7BJh25iMWCibpYySL4sQyDfJJK5E3IV
a7kPyRctoE1UCebaSRonaVr5obNS7gkEtJ8hTzGo8Y1C/nNJ7aTFCXRy8b1/zgp+sbxSEhvsS8rc
sdMAq4nONFzEr5jXoIi+E7DS0/BAvc3+Wm9hUJN+2lvwCMUgg+9g6/6S9frXn/F4XpvktVoKaTkH
uhO9Rn0nQZ4puJe8bssnbWUoKEGqwIIChpePYuuufF3hG7Je2n7aPrjjaq74Q3xHdNi1+8d9fuRK
JtaAbOrxpwgrTz0k4finHSzMqcGPzYs/fxY1t9ds0yazXwwlUgPDsdOE77gARJZYE9RqRwZUBmQp
TUHW4F06Dh6KQN5+6PjYq5U5BvJde3gmvgg6jOnwx3ePlXaT8rcb0mCPa/7yv4FH52LY8vrd5qHT
ZSa4GAgdfze8LsypaeQF3xt9fNlgWLtxzk9oMbPr7qnRehqdoMwmNbOrBE1J8Vj3K28+XlvZWFfP
HZ+9bO9PsK5F1WEyrlCFm39o8m8BdQCDBfnRIETZLXOD0J1+PFmKx5X8Z20/6yDBhMHCMBqVpLRv
jA4GcgE4uzQlF78q/9bhPfsjqI8NQihdTVi13FPguqNVJdpwbbT9dj8s/yCbKsFDMg/ZuFw6ekIs
8nX7CxukEycXNnBLAYowcRaYHhCcI7yhIiLq2VxlMwZiC/iq89uZLMEvFDD+oENxqjWDSuWEtL/7
7/rUkSlj4rT4MyfMTuPiLGJN2c6zz7Ic2cB46JXalpBySsX0DRDJ8r4jrLzU+jYW17+IsAXq0i13
uQslctLNiYaVp/AtoQ0pNTbu5ZDozQ7sbYLC1fvTKmaoC1L3zR1n5O5jilXrmTj29J1kngr1/vj+
wbVCLJOQJcgSNpsWNUnkIR4sNMqhjsHmzwM8Awcge+BElrFhwa47bVkwug4w3eyhPfSmxFuk8R9s
yPLuNp8fquw2sEes/wunI8lHoBen1tQPBWsAFX4wpt/kEr2/zCFtAJhRlD7XiOfMU3RP75KxNKLz
YaZvMz5FanM+XFGp+bfHHo4dI6yPbxE02ZI6XjuhoQeS3EIeg4cteYEmodztjbKXsgvuJo6D1rDs
Uxa7OHuax8fp9i47x5UQG2GBKeW1hEwRDlJa4eYmeVoqq7sz6PlNJPribDJBmQrY6GEa5RUdX0FB
/HigzueKwOCfgBn4c8abwljMpirLVKkXkCziTRzk16G1piXL6lBlToX8qRohFO551wL0mzXyhy+Z
qp/RjPxssWkNcD9P6MIGVH0TtD48eYANbA5WEA/+AZqH6tl+kFOKGfuyjZss2Gas1y88HKfTl2z5
p1JJF+FC1o4pVR/rV8/dl9gTm0tWMrHGkkGdSy7BDL2Kcvu8B4HZRVUvLM+jS1KVDZZTWXtZUoZV
S2WG+CLmcEvcqtWjR+BoMSdI5ht49vymdP6QYkNbO8f4maePa2GtH983Rp+F9koeB65ktgvHE6CX
iDYNVgBB38k1ieYrYFTiS+cC3aYLVEzYvMOfeRVAcKMlZdZ7eVnlpMr/mT6qVt97mNH3RZ1lQHqz
iieVfrBtrUbnICoiMUUoIhvANEGDAhWhv1iIKG55oY09JXsMJqMxNaKJlXGp/GfC5uFM+pkbyAbP
8o4X23riSco6wWPdhED31+Ry1hB2e03lO6jeIt130CoVoZPawqytTbIQidVcUH9G/70Csju1iMSM
pW5PkyOdkDpa720KtzIOZrdKsZ2n1xMYB38Hq1/VmVSWZSmbaohSNzZndTVukWOxFAKWMzMG+bDK
eNvtjYET17D9uQmLoniO6cPAOeC1Ha6tTWdDWI/MZ74AOQnGaPeEinkVhRgX/m7WmJQK4/ub4S1D
JQP+2ibLUI5PJqzzc+/FLuToXt1SscsUgT7V/j2IaQ/LbA1CU3lyRf03K9cyIwwBd5W7CJ1vlSyi
UlhjX+7sjloFZJzsSQ0suUnhSlwKiz+DjvrkuYrtJkE7DgQMBcka6VRu0B7IPoNSzEkMsgG0dpYr
wmKWfsegV7nGKVtQneYT9KNNBi6VZw0zJ70ErXt4R4yoA6pRxRZuehKAE6sC1Hl07UBSwLVXZKrl
lz6BJlMigRncY4KYll54B2SP8EheIB6Sae9zNF5bQyzZwAF9Drr2AJ3POjxdaCM4kyp3deLBr834
R1iUZmM2PKlezE6ti9UaDCwca5fEq3W85Mbjhwx3UG8TNKwSV2LngA7X3Wm7OmJ6iYiONbIozZFr
0RE+0S1AM7Ls86p9gy10l2FCCx4DAyCe0ubHxJgKyvQOgOE8jJg7DBFznF4tJj95sxJ2BWv0tzHi
S8H4RDV+XAf4lZACoZLZKmQe0UzBOgRTjxP4iOqD0ufYLg7ey/LxKZaWH1FLbYe4uS4doCfu39jt
VZ00gHQz9+QoXCoabb9xGTUKjAfrsBsvayPu9zL+biPvaIp36XwU4KHqgcHBiGf9VcFWqDY8zNzr
Z8lfUjKfzeg1zNSDFj+w3QkPSkPfx6QxPf0ZBCJ0xZ7vEIvgyyC8/hkizw4yA45xinaqgaXiZgmG
gqOxNio9xzI1wuYsh3jXh06MOfAjNY0HEoX00zacaanwcXVwaJFKAJQkly/av+ft6ZUrmHE3e6pd
G5lJqawlXyT1Pa66SOomDPD8JoaM1oVlujEbIY23+p6AjKTpU8GMLOcSD/rtD98nxYkxOeNNJv2i
wTYIfmHa2u4pAR+RfWNDhA1FYsZBArQ+TQKUAQPNQNc29D36ciKRr4EWS1WZpCAs+t5I29w1CUlj
4N5ZRWLmlaHCcBwHgXk/HFIABk8Dy4RN/LeBBATo1wQCF5t1jA/F1sEp1vDnSX6KqX58D63gYQ3c
qMZwkLzZQF7fYjWTYlCHrP4k0cvcjDnKeqTAHVoryVeMkhqPWBIMdIEg31aT0HwwSLquQ+LWVubw
q5aUBVcJMl6LbHTQ1f09GbT3rdI077EB2RnnMJB5Mz5bsXpos4ITwnwycaNkyXQV9CBXwJ2jB74U
O9UywAfK7QjpJzbbkQ1HCvJFLmbb/+YIZLh3yYo+vEF/mz72a7lNb5F5WsAS573fnYNYZdfCet+q
sOFE20QydHWUH2vhvBdLrlLoSRO4/ZDFETrwFL/RRchUJQNZNzglAYxDaX89hQJ8FzdS9Qo9ng3y
69ypqoHyAPq62EN/Yh45699Ynwh8btIZl40Rx6FRTWYIi4zrVnKz80Xkz9oVAdtSP1pnuT2TsHCw
sGQ+2IBVK4+w9YCNBbmpdhD7PLMiMrhropp0JHSxGJVT9//w9eBUbTNjy0raWTUbc+9FwE1/KmZm
onE4bsJReR3cdJ2fQiVC/H5+hmVlLIhTcBnQYuPu1Lj/cVvaWCfu3IRF/oYz8GH6SXUEEOG34p3t
Eht0SsRguShelk9fznyH12mddHSyLF9LPW6ZUu5bZ67FucQCk+yT2JkRDqnvbtLDEhVjH+obrbb7
bPLXXuJn/FbiOEeFQBq5f9HQSSLTBBC2rdwRPUZR4CG2s12QTZrEgjoY7IdrSHDXk6vgm9Cu91FT
hGfhZBSab819d1JnbXwyOEcoIvWEr7bcWLF8j9v1hlx+VK4oFGZqiK54F3htIaG6EX+4vG/3CcUg
BI7rhJy0ozppBcUeJboi/v7C43WdIavcyYH5sreInkDjqQWAWVSrcB1MiwW0UYK+MTRv5KeMV34L
hFnBu7/2Sbf41t0LTVDPFnurjlDVJIAY8sBqBv8YDZQl105Nh3h7+oyZxg8q95slLk2Z8TrmGyIW
MGG1Yxs5MhM0j9esz/wNYGKCoQDD8I749n4S/wTNyPTNLqSPY6nV3irRzjPHV5bZf0Z2zQLuoxUu
bqivYFPfIhuIO5lceS88uqF/8wadrlNzizuXb8dLgxHb30zLOaFyX2AXYQDAPLy0dtDKI86ZByT3
gE/Y16gQjHD1PYCIwIqwahp6+rg4C9/UvR58GhE2eFE0lNHrwTPBivnOum2sLsCTS2kjx91HuzOW
tmBPm8LYVnSfc4cONl3YAp9KKNA6BLBAcPKiOtyUF8fdKY+tb9vpAQ/TyT7ITaOQGepwD1u99anr
ftk0Fe7uR8QCQ2Qbs/p/7/uX3n3pKbObGB5iTQQfJGElgwOxhOIFoSVOHf4S8922ZhnvKMmlA4zC
S5SNIBqDQxABX+6xeNoItbZzYyC/ovwj4FueG0qGSkEniqwPiwtj/O+nLJixYPn96ljiGFsPwX2E
exyNbH7Kgqoozsn88azCJJCpsTxbiNWrnFe4fKwKrQgB23K2h7w/33m+e9dETQA897hVnQEeCnst
sMEyWYplxwZAMn1QOQ327rlAVV7HnXB31jXtcdg4Pud7IyUQsymTILOdpSOJLF3h2xugIr8CUkju
x4I//wJeTKUmvJd9FtYerxP//JgSCi7MMeCzhW5d2YE9POLx1ingx6y8qljJU23xmYz3njb8xHgj
WurEANdVYigHzMvE7n1nTYgfFfl72J+Uzt+u2S/y9oYoW4vFPASU6lOCmmEehE3410lzE+MBXuS3
BJ95tPLqWXtf5D4aPXM3fr/d3zN0zCv+HPUMtqrNCJ73DfOFp8DsE6XWpPJRrT9CUSykWm4/7uyq
YMPad31rzBZhajRPnNEhqtUZErmo088BAYuYKea4f7GjnsxDIsLPjy7xkYrEqFSmeEbZeahEmqZx
O62XKCiN7qB3p99SV82F5I3viu1t4jujNTglwkslRBel9xOjfF+PRgoy1BM52QVL6S7R0LC7QSk2
oJlhL8Q2D8bpqv7yUuZWVAbKAI8GX7vnMez/LHNJ7tZixxpp+VG+wkaZdNIUxyvf4J6wF1A8KO5v
MYgbBbeADFJbZg8JIxBB8Sq3BGReep9FpQdjriaVgf5lysm5ohijPXfbunbq7Q97yk/sDjC6VAYK
9xXSDda9j+TaqX4n5boWK+Rh547G2zNwniRQbe6qZ7IjILbauPSrrGSQvilT0sJrNbkVBqV/rt+l
QLWq1wtduSb9xld1X1O5ESG4eJBNIQ2jbv4GsdgMiiHMNrErfoYeRIkGvLQvfG5W1T9uI8n1/J9L
TkEnA5SqDDScflF7YK5/QEc1pMAiG0qn9MYRuU5tGYjw7U/EAMD6K4JT2Y/MrCwSMFjDI2OrRu8G
q/2gc1Fc8SsXdAPPDWWo26MGTzIkiQZqdtmd9f5r+0eVYKrmQtJXxZDHGpxSMXwND5N17epY/EAW
PSHsMTDtJ2kk3aSzLjK/UTmZ6aY7Y0KdJas12S6WYpk0FtLXcRXCNVPE988OWGm70Vt6HYP0WIiA
2mK0IV573g/31+mH4XBljGx8IWysQV/KPkLCvbs927W/ePUcfphkwJ1h7zlP/H6OVQfq8WmnxeTZ
22oR+73sqYLbvGWno2rZKK0CoZs9nUWO2qL80d5XFPACvSNhoJYXlUjIBDd+mLRcpY9BhmFNM/Wi
9xV3Hyxrk0nN8CmBL5owBeiXylzb3rXYN07Ny0M3lIFy8e2DsGyQ8dStfWDZ4VKK/LOmCVC21sE7
Ich83fPaqUM3+i9KbrImIKvcqHdeguwZBqTo4dRIirgzsXBsWYTLLOaiTl6PK61IiJK9Meu00Prb
rJuQBfJ7rRLBg4Ke2OMdXyXerhFZFKhr3o7LTWz/AC+0Yi8+Bg+TP9Nt2gcZXe5T0BVwpddmP6ZW
8hzyqS2clbjiAUUkvKBZ/FbG8cRP2ZYpyczjvDAf8/Zg9HsX6+0isJNeP1NE7AfjIV+0W+AXLV7x
MSwJmix8hihyMnc2TWU8M3CfDEmOX+xrD/OWwdC9/MLbOzIv1GwxH+vK/V1uh7RtEsp9kdjkGTFv
3zzPod1aVCkZvwcUnfxc4ty37V+v32VFfrKRWGrrVMhuiwHTJTUCbTmyd+7qnEy0jjXWbrS1/awy
qi632HGkFYbLgpPx0fQSsVv7DqLEOZGQNW/47bpyKfWGOxd72ZWgZjGfz6WAfO5V4MQ40gI2C7vS
gQD8zO+PKGljK+Qina53CKbbtWLW92loSI8vNdxclo4dG+EhMDk3AKTp+DSUAqxmLCogwDjCaTcR
0Cb9sATUvnVrXPjkiV99D5gt0t/4ktkiQQD5FtJlSqHdiwTe+HzZYCQngqW4rks6fBlxk4Z8f2VD
gZOj0J3K7xvdxuYNOcebiVYncd6d1GUXZTtN093i0zwOWBZQ6zziWi9c8ZMpgY9gzxwTsId5r9Wj
iW3A3I/Mbrd0zIEd5EqSdSuyETXVUthkcOK2xSYM3nVMF0AHTKaYqGvF6srIVbxU2+ALxzOpq5Ba
TiH3F5OAwUyxsNXaPacHFIAnYhdMaJ1Wvix6eyoZE1RdISBSQRzWlNPn/uAuLyalg0JryY1/Leo3
r/8X2cEeAnsfTDmEXhm8DqfgBgrtvff3IP/CoRmyBrXgnoq1lmVr06FCvZWGT/XJHLhBY/cM5lUk
TJiIxCOPk2kQCZvkioV5CEyhu5lIoRiPy4IRahHfJI1slEKaBoOIpw88SXTEIdOGYjq4dko3Ksnl
4vMXoV7DQJ7IsABkMs7r/i1+jkQuASi43eIG8hdQAmKF6NNux+H25kZOnx6RHLTOolwDSm10Hnzs
BnFCZvijYIKwEHCSexqwiMbYSjb2wMtpG9r4KMey2gML9OVEhcPDkaJUKM+6N4oWrfB10DNPnrOp
BH3PH9IqXXeUx5FKH31Bv5biHw1nO2wrwcQY8Cfol4RU+f1wzHsGOSghKZ/ER7nP0pPe8ZNU5wzm
I7tAPNLsVeTd9WJgQ+OXAF+QhRj5y7u7RjGcofr6nd86pRiHgwTCiynds8oSpviyKfcyvV2ZGWoc
M7y1CwZ5sukyWukGdEjKZktMGMx2hXVDzumZNVKTRRkDqkt7YRi8iWgMzYC3SQ9V29cC5q8oRNFO
EtJsdkTlM3Bir9cSPBFq5JRh/ZRkc9ZafMIpCGP+o22ualk4y831Y3LXssNLUtEQtqeEquA9P2xZ
N+QnKS8Rx56uG8+nEByt0MmGYo88qHDUtgsZfUfcUOJ4LlU0Z+lYAV4ktigzs5Od3X0OnTgzemOp
JtxUy8si7dOBg1SNxTKNqD8ikR7iVKjh7I/kfmVhTb1iWq93nSmEQmawPQ00zP3vO/FbuhReaU42
52ccV532/E3V3mi++mBaiZ4pJNdi4D0PgxzeNUFdb/BlfqmXxCTvxXEspNnomJMv+7JlBEl15Zkr
UtsGEwo+sLlrjSFDX2plRc1PQPHiLovRM5rUyZPUM3G9KWPmXytB7pfowcd8LZd97XF0CuVCr4Sv
gkU69YV3M4U95FbggbpqupD7j6jy4xFWjDb2dPxFMXpKrzOWyJ30Oje8Se4Rn7/PXdFWta4UEhNp
kiG/hBUUTzWtenPG48SKAymGAVRkeXnQmUULXAlvPzSUdrrfwMsvXclYt0wcK0dTR1fbiXVW8Yuv
rMHL2deHwgrrvf/3sH/kgF2fufQE4wQ2E3qUN/t1WW/svt38bZhr4B+HX3u2KHhoRLlcoOMW/vO2
Er9C4ZaUiQZaBv3fcnmGkHIYWVl2BNlmqf1rlCKXQKe9d2PMjHrz9ZEKcwEIgx+Iarwg1Z16Hizt
AaC1gp/VJp/DRT/4MIEvwbDIrSHIndbLxP4I+F2v048hNc6vULKMRNf7O3rH0TZj6pAEk7ILm308
OXjSSi7yIsyBOXyOy08qaOWPOuWb6Yhm3TmWWD/Ljo7tjgdUO+PrIvLOri6fDTB4rQXM+wIDkoZM
37YTnlfsiN8CQoCzvM7ugfVP+5QEUtGeHYbZ5J5y6Mx3nTmwmwOZ3ZbCffs47S5FUUMT1KcDDr5O
Wdu0ODuOcIuqzueCJPXKtFQdDyQh9UmO+1sMwqTxcoIVFxCh8aBN9wW5ff7b35vT2Snbrij4ZuTL
wsseDZL74k64m81XVyFGWQ7T1uOpLKfD1orC/wgU/TNzSk37GyCn/hVu6lpUPO36xGwbjy4lYlUA
YouOaOgM+TjuPDX/zJ5jbPeAJs73OQYQ9aXOZHx77Uz3kJdejyJuewAnjo5uwvBBBGO+hCgPhh8C
55gUhvY3rnRwTi5+hhseOqKWfbkibMZl+xINQxGzF74l05yCXdwdfcdPfBIaieIYuvhkYO+nx/sC
WAjQRFBYrpIkKYwSFhwY7vYXionzJCu6GTw45IvTSW2UreUhkVY/mV2FitVrTUD8HnoM/FH4Fxtj
PB6VpMexxX1IqTGf2gIR73Q3jamIcxp/YmQJKL+XDR2hZntMb00IV0VALFApW4YRDDN6PTg7bpVj
i0MMJBhdnYdcgiyF5PyiS+M6AsmtcbrvDyedMzsuR8GE9MP9ooj1iQtHhf59DQcdWXaiM/drsUXQ
RoCN1RrN3ZaJiR4d3fMBvyOcg8dpK6rkRGdAJKCm9vwKS9JvOMfAAAca44l86C7tEGkHT5GbTp7l
1fobdp12WgAT6sFlr6BlknBvytPeWcQ2Cvcj8998lH4N1K3kF5t+eKEye/P6qTh6xaaZLJIeVPU7
K6HjszxSPEt9E/lic+7qm6E33rHrLwXNRNkq6/aFkLSk0ApajiXc+bDmJYaxP3G+kHmoT9U8UxJR
8W/5fDF4Kwd4wccFWunHz96s72vN7+RgMJ1rILGo+Sg1fjKlr5f3ymqoaUGLZplZrh8DHwb7MsC/
hnUS7tweDXl/iS04rBwEEC4Ju6rCP4uZPI7XeMTZtRh/p4lsDMYcDqga8Z5HEnZ5Iu/vh9DsnIQk
9pZ0MS0I4mSHDC+kN2q4YfbYRrJJSh8cqnLCZbr190W2iMNdszxLKYvV9VsEcHwK6gsLbrICqYSx
y0zJApdIY5Jzs1Nuf4U/B4eJF3gW7McWrAzTiaNx9QSJ105QQmG2sKjU5GAG7REaucE+1A0v3ViI
FY4Zua+Vt4cwl3kk7g4UW0QO48XkZOyoAT0Ha7hWczHznhHysxJyC1eUgCVrrvAJpCjNVoYDXrps
pCCOj6/fepo83VqZY1RNR5WGTy3GC8M1RB4r8WERIEODzWyP5/XBcEWeHHlN9YjYtN4uaR7M5KCC
w1MC9T8QZRejbBuefwdvF1K2zqa9SWsFIVF16sLidGgKmTV5jT4Zhi7ySzkPDYbYABuLuspkdGWZ
3hx5oHoG/2ZhigO2LEHdoCsAyd4gfrY9Euh9dJxdcGT2naBk5fr+VJGoNmBUo5z9Qa52zbwEjUf/
xH2SiWYFoefKXg3e/zHw29YINGNSoWt28cDcdzuRtQ03aKLW/F1lDDEqcnkLEccWoO0G+b28BROR
XCBeuw8dwwVCENKkQqDjGZ89+ltpKtSuCw4BX45n2kljTkoDnsGeU4RtlhhZXuooQJbHzB+fUqQC
WZNq03WN1OuSOaVDvB81nHSpaOoJ5C5GZmb55eLAfOTf4hy0miqr7Ai7mI2DMJAPmMdUPWH0bm/1
OQJr6qK/PM1Eup/WvhWTM7TfEhzKghLnn/eomhA7xR6uSBOanOJxH0whGYbGZhRurKCahb9HRRAw
VyEuHxAqFsZ5alBYf/3yY87Z6J+Kdoo1k5JqdVMjhkUgzvbGOoCYF+4OgerjO3eoCi3QMRa3flEi
GAElLBm6a0yQrEZjBYy4u/oGBUkZdE1DXxNFqCMwwoo7rs1F+rnve/LU3VyefSkPoXTiq/m5Qxxm
N8Pk0uYjsxvUdOP/oNMLPZUENAPTAosHLMuypNYJJnGnYpU5tR2s7F9Z4USLeFfCDH5SjvgfO4WB
PhHsQPrDoQDOvX6Zgrkg8hRwYwDFJf1MZd/gWORvCqAuppKvt3YT9kiPEQ6m3dXIqQZCJDqFAXk7
wbf4Mlf9/4zuDzfWoBAdX3RbBHWHAi/ZaeZLM750xULkk0cky+wwjFwF2PWKs7aU7QVChdA3o5DG
Id5b6IAdr4R6LunJkeuMUNUr5tZIpI7aVBzYXAjNWTWxtgPgCivnqfCSU/++n8FSYAwko8AlMpuo
DJx1R5AGhJ62dsOEicCJQWUrlslVOAZoNftt/MvXnXmXIQx5KknngTN9rj4sQ+iCsGXRYQ8UPFLz
g98RlQ1J7gV+fO5JpwE4iZplZ0wEVSOuJn5oRj8p2M1aUezKJoiU31/lbGJYsWfIl1eB3iREBWhB
c1J9yhxRYuWckjq3Qxvg26wQLxhnF846p7s0MbtPknso7jB/5btYftBvvLd2n6YHhOXjOctiD1kp
ZSDF1sYwf+/zC9P+jp/E35fjmWs76Nfcowpw6sCOFWrF2/Ob2Fotr/G+0uvvbsvN/r4ck3EzMY0b
1Q/iX7mQbySrJjtI0lfBPgjvVRn1Dv7pckbbL79hXYloWkPF7uE64T4W5RY0AqbbB7dD5XF4MK2p
QOmhP9jdpeKVgzV3/yiigfSJvFvfl9ofg49qxUHhPEWeAUcqkcztUY2GTm3BrUqzMpM415kYp0cV
14jP5BGq9maXD7l5Hv9reRkRmcass/zO02YV/QqVrOq2x2CH0JnQSfzE8O4cCkyGDTs5PXLgN5Yl
jSr42Vpb/OeiS4BUTcG7DUKJ+/qf0LygrcjOZ8tn/k6Ca5Vw0uHXBz7jyurW7P/3djPj+ftFRQhu
APo/p/t/lf+qLA6ycuJsFIasIkGUce3AADyOjWtu5tS7QdgdZiLTDXRnuZPn4tbSs47KwxCwRbGF
oI38N8YjaFexx5SDOwNztFFkmhRN3f621fG6DSXJWW4aN5U52Fe43wvS7GzgfryIFM0Ek5TtOg0F
xf1FR7wZ93jAedzIYijccwXxqjXslXrZvRKS/dRJMElYMW79TBUHjNVqGCef0qUcSA4/q8zY5tUr
JzR4Y/u0IqR6BH+wblEy2pG0TvNrsdc0WDfhV/p7HQFwYyzt4GtDp9xcGf5wnjwtfsRFCaDDsweO
a0o8349qTck8VzkyMYxcUG9vf80UP2g38IJHrpAfzKlis80Rn51WFw5BL5TdoiNONurpGk1Ud/8g
+ZZdCriR8QVCWdf8IUCAYfHhw97Fo1JLtZJ0qZOSgXHNdG9nv3tcHuEc5ACstlw57+0+81fFjClB
5Fel5fLfa2qxcJMkF+3cS7Tyt2r8jVAV+zeL3ZFPnUTtdDrZPJUcJq8nL3SmxVDFhEah5G30c48r
42Fd0N2Kq2PCP0qovIKgkinmBm029WPU5kHs52Rcad7bPsAzL0lAaWR4EAzPWerJdcQpaX61G/48
5o1wl+pTx3ErATV3Xl7nBmnsa+ayhQ/+IEH9WDTRLm3n1ND9U6JVWcGygLPpNTB2tooGf8gYU8bQ
JJHK9mU6bcvSlQ/qCX+MQHZA8x+1XiSN/wdzaS25cTqFTja1N5lphpa8pzj/7a1C5PvAaaf7r4KF
w4dHx3MVR4E1ynbzexlcpfJ9gSMGmgZk8lRGpAP23Z3ANN7zzkN2Jw34+AQ/gMrajJ1Tz+NfqYAb
cC7A6nu+mU/F8qlXOwuCZIW28Y0yiDPPDOHOJ6Qigkg8ucEaPjVJZLB++A8TRr+vviN/zXUr0BI1
JBaCgYm53HKZzauNbBaaOIAYiPQKRbZGZYLaj6kvxRHzMNdyU9OIfTtopUZcCbM7Fb4UD5Febuhv
ot8Ky3cnlnADgXqwwarlOCZdX6SUUELr93Y0OplPueLEw9S/hRt7BJBX/3Z1oJgVPuhXly9VDW1Y
mTPR2CeHlzxvC8JoW1Xc6qYASP34IRzWjLQEu54DJg2r/hINubiS1bdGZYXGAVrLfg5ey9fSlAo0
i1JgDj+/oihDpmcQaHSfUBVME5AByT3eRI9OTm1xqssz0JOqJaC0drGYjIkQV2Tjel7ta//3fGKs
WHGulqMjyYguB/BXKfYQYZQ+QgFfRoXYyOWHHJDTyel/yNRIGZcwcnpmVgWuCNfLnu1/XkJmCUYc
sGK9jmnnUiGP85L3DjNVOfs5aRZGvayxQcENNGrJIQFPPpWA0s8hdw6/GMJOebAhYoIJkoUaTbb6
F6UrTHQVOS4Ac8lT17TrOnRCGZAd/e69cIyccNQOAwvZz/vDVsiyh9f3eOpiAHPLyV3jcDLKz+NG
1qxNdlpOkCMw5xtWgjZ0lu56nN37pke7IJJrCfL0M0W6avkYtszb1FhFu38XbeKXAm2/BrwTW4Ce
V9OwBbzVUIyuu5dX19XkfrI/78qZ8E7ZRGbWMNLPEgI3GMZi2kDG9wnRZx3RTvOItO8X5NMmWBpO
JPffF2w9Rcx0oP7FM1asDvRgyRMrIdinnvsZFvOm7aGhGalrBsdzvJhHSCsZnt0Ks5O8wrni3qUH
LmndLIf5Z+XrVkbHS4F2nbQ7+2UW2yIaP0wkRgG1kA+aCt3T92FuYhObp/DV4JfzAiioc2ArWLLm
nUlDAtzt4nAuuSleuEXzP3xnq88yT5Ra0MV4y9zN5yiXxVRHltUlxMQeyR8UxKE42iMZ2JMmCe/l
2KC5FLR9EguVPDe9KN6LD1IYAfs20c7qdrKABM08IB6naTWFz1cLKpgPf9RgOs0KFdBSaZLUynH3
hXX13oxoogd1eRWASSvpm6CBaTo55jHNW+T8WOAmaVvlUPjZh/tdRGjAKNxSSktlej2UhnsPh0kw
Rn9Jx19iPHrlSTXzczOQhAo9XD1a/I+SKhpYTD2HDTz4EWrVYRL1n//BYpPxPLReUFYlYa/0PP1Z
iZiZai9pM6CKP0zzGH+rr9baiC8ahZSOeePL1Pv1Zdys8WD1FMv6XU8/fh0DTY0Cx8pFkmR+fTQS
5fhka7qgXhPKhtAjBkY5O/u8wy69H7evSKcsecpD8EC4tw8qWiJQgdlN98yc3GLQkRWs3JKXouSB
jMuBzVCgP1H+UKoySj09ffm6auoqkgSuUll4Vz4USTXjbVUzkxxY+ovUuONf22tHtNhIANYZQqTk
2a9a2m7gIJNHd2mCY5QfNYJQ4FJYblavCdQf/6O8SLTZGIVIyqjCQGDhrbuJlqQ9IaW3oq7dRLK8
SIjsdh7kA2M14MSd1BSqZ84l4t3NomiEIu5AckWHGqep/zOthzklqXYhcstRKVGyz64OpigV/vDc
G4AYHDmHmm53+p711QXquYolAtG2H/g/sfbHz7DxBPWsRGaP6vr4IxiunCFMKYA+u0NS+CTk4hp1
cpeX72t5HM4boTHXeyImonM7g1QH9rLRFVGZu9G917cTnXyGMrnIt/DrsnGjPqWLeAaqwArtQg5C
u9TM1REKiSUm4+APqx+a6/qBA51ypT94ZNiRyrymGjhYrTk7+5/i+zvglyomt/M2weaItF1x+T+E
idEHipZj2aK0vPBiSnk2sPdIDKE0h4vgwk51HA9ypn4dU6b36V14DK0ulm4nXH35iYPXrlM+71Rz
PwyjiHTPYEDC+ypiMrqRSdrxM6X19GGbQuDU32NcW4vJbf3ThND/ZsK8FXh9rg8GRUNPQQXHpSWY
91hQpSXFlAm3+cU6rzJ1kXbRiZD9Y7hMqyri5TYHCFfAKHWtXD62bHE8FFmoFtcfdLdDZlTxW5dn
/LxP9BztpH1l3tzzLYrF89uCikyjUi5cJg18K9pXY29idmimciFr3wNFSyseC8lYdfUZAXKpHxjC
j1vG5C1UUGjgR3EfvZdzsCYmzBCbJ8YEM7RLFstiz6a+RfRRaPoYXv1Dr/Y/4136+Ke7lR3WiUk6
nq9M4ZKCVpV20ihi7YwIC2ivnsTkIDs7+w4H+R6gprapJRMy+QGBgmLJCyL5oba8rX5o625wy68Q
XKHYlyI6ALfbAOsELwmWHfA178saeilGobx/K39/WSe6iyYbFIKAFVVJYvrk8TR5KlTNQeRh1qdo
3uKWYJsam+m4F8vuA5e75BneQkFrDBRE64nIHxa3k9HcI1kdSO9OFIk/55DOzR5ckK7j/gYA2Sc4
NOC+gk/UPWW4YPbD8BqQtEe1CGu9eIdVuBM3SteXU83rM4c9/lx4OUsrWebpig4N4peQUauB4Tsz
lSGyAsDViXFPzVBkgN0Tp8EDe7XFDrJaTbhPE+LLAqnn5CdJTqN2NJhSokmxLO390fcM28xfLYh3
9aOhpgkZuBQn1jnnEqbHAwPUg1dbj5IBBnORsNNwEhhZAeOR6gVkjFSizvQAz7OusSkAciLGg1G0
mW35VpBlUUALQS/TUprcM1CradwCxJS6X8hE2ItNPA/LSdBUKnJ85uW5821jVF6ZXtBF6F4czxcl
BNs8ZKJcUiCuGsC3ntI2AzKw19OVo/RyvPUJKBMINEqSj2F/F7imzEvNqCvUq9P+bHNMCNqlR4pK
CP637Kt4gqTXSxrYxy+jRA6viU3Ej4mz0mjQeHZCYSB5EZavPKLCOM2TlFopoSdYA3kfBJzYg9yn
3kcWPY7eWoaIBEANJ3rsS4Tn120xeEYORWEa2M+Eeu8bVaAbJAnHQepArjyZmfho7xqEO57JyIaL
jUJCELiSn6pPuRdAILJO2wAC9h0szXW9ID2oWqVkN60jskyBwYZjSoYdiB2xY32qIvoeDNy0Y57u
UuEux32v2UxxtJH2Cws+uks5xkDHkRuymUDCNNoX5iKTillzM3pAILjlrCbybs41Bx/Y8FJo1pKq
hTM2F3f3ngMCZqfljkG7o0agxvdXaCeaDTVFhlROElSG2XfO7kCHb2kbLlRhHiYXDLL77PpRLh/D
ugoTOD+RQDk3XeY6kWIupu9lJqKi1B2bjE0Fw/To3StHuWvrSMflbcyPUMJ9jsqI6lGjkow/x/ag
94iD03QF52KDj494CLRO93MP0ewStqdsj3+18ZuJ7kR+v+ER3+6J9R7/WiEFrU3yC3ojZP6oOhP6
PERdwSiEsH54IfGT/P1OCV85NJNE8BiOZHojhhbSifCgSwBHXOu08uXC8j3GpgzjbZSRO7KgXj8w
0Dh755jsAK1xgml7zT0iKx9sLJZeGdtgIL9Jf3F0h7yW/UmygpWWJilbN1xBhMWtnJDbpNno9W+g
fD75nZ0g009FnDt4lnd1v+DCCg8gmRifs3M4HmpfdABD4i4Ghn7Hf/LFuJ5fn5VYSejMAT7f5OwV
BtFWgyt+TtBzBIQKgUrjBg0oJ8IxhLRm9D+WpNh/X/9HcDfmYoZa/LUjpOsJwithZL2TfpoPSGYk
YCzfkokmlHSNKRRF4rsDVJoKl9NRK1CpGGAni+BZDccc/h5ZHI0KGsaK1lfWEyG3WX9YYH4trgLM
xUEb6zJJMAElWcVpmzOkSv2HXYZO+8upsHZj1G6K2lPdcd+cQKGPonYqKYVL5Gf9a4pGgor6y1by
eTwDJlqjoMFvTy/v2BbujDD6K8ZVJh6bI4YtWFQbTEbtq12Lg7pvXo2OKQXfmTHwrPuXJJiwP5Cy
Y4wjLPxuNf8btSJER4UkGai5CBZ0HbHoN5Q1+ssDQCpQUSyTyzOyy8pgVNbqtHSb3Kx2WrYGwvW8
dMtoygFBmKDUAcpaLEuxx7h6cGXeWISf55v3vP5Aeda/zgZZNzYapz3lqBM+rGGVx2v0bvujo2xw
1ol29+ifeGYdJJ+tVvdzF9heSrMAClkUDkrB3RMzOXG8FmYPqMkH29oBTZpeRgKBtkEvjHovCH9q
gYHFZqFNRGLRB7PyNXskUK+bJwIhbtzT41Q5RlqDI8Jwq3x5I0dlBBJZZIcmhDArGYyQKuCNUuGm
0cYVJeQ7bvYF1uLZRWZD+UT9ae6cMZh4nFjpVsInxUi8ykj+TmfQSz9pGdFTT0WS63FcX9CBonn3
PMMv6UBC3Ff2PZ0gM6cmxfIvBZaKhLp7g9uOBlDqpFxDZAUaWpZtOkNDqvaEEBR4gBTdI9a1qUcj
SkxKbHBG+BKzm4x96tY5+TYyDtZBWMG2ron4hg2y0LAWJ1BWIgzy4K3OgUFOGTKy/3q5azRZ0gJZ
+VyoDVz5D/XGyuXwE2BxiLlQPi4EYy6cXu5TuhjXR5hfxKErwgAr/3mT7QHdyWEO2miU9F4zOuuf
5Q2jad3f1WGrwoEH/d6PMnI6s2voAM3P+rZDNphCNjdyz/doQldMtBKORgIYSJTaeSq21oLnGUgb
PHadjCTy9muVXNKgf6u1KAS0Ea6y62G2UUJQP+26q//bV5i9hnMFzL8oJjmuZKu3gZuXUUwUCpQx
nzI6bWdAPjSNXBmIxN8gsSRT0hofJOa2lf+svNTSD09iWDl2v91tJcxtTACVsrr560RCwGV4kuy0
Lqr/oNoZW8rZzvOkc0P4wRn8ZAPiq+pV8lbr9GuHOvASJkbqg2U6ICjuCKFzyu7kvFzn4DL9acXW
lP4TXf2/RPPtvsVVcVYNZTPcVVYwumZnYQIGM9F5YVpk7NHxNfiHmj+twA9UuzY88yRBsdALYWcp
Ab/sF6SvIkkDEV2NGNdAx4Bl7gbYIxi2taMmB5YdgyxpyvF8zgtJt7A5gZ4cSyRm/J7qMyyMDjdr
h+PwkQy78W6FC68f8ysPMghiBZDp8I5dhn+YFWV33siAUQGrq0Hf726Xs+Tr96WlGMTmX7D++Gvd
vqisPasAh+csuiYAuOkCkuyYEmFnfJSp8/rxssDJa9ZT9dMmQlAsCGyCqUdw3CrrsgmWHFmX3BUv
R7Mdw+Ztj/peiwkL1HuUqv0bGVtB0AzaefQAL8kJiD3gVw5aVNs4pI5j9F46dd7xyYLApgpDEiSU
sxxDd0UDxBVgdT9NE6ssgNbyEx08NySmIszRbmyZB1VQYra6dxWWk9ROuy2hrAETWaE4+jLeDZsO
EVacODpNNWZ0KNtCKRHWpr2X+bTFdhRy29XbaOHHOpQoVmM1KU5MErO2/nlcegVz6aon1cp8mUn8
6si/V930ujfbVjDLQqwTRwOcO2w+Ms1D928xPeJodiKF9K/PEqWgqaboipiTOtKevnuLMk86QNmW
Vcvfcu4XKwqtyVfu0U5KWnGdy+4ai8FPlE6TSj8vkn+ME6Y9u9FxHyryCcvIRlaLfduoJ4efYLCj
EDTrqXQG2XdOVHpcO9FXzoINziPEGLyxa4SobMYXAh94R3zJmMXy5W/t7zgk4j26R7bUdrd0zT9F
yN+oHBHh5QC593SJYdheV5F6hQHQhlzScxBppdNPu/vsCm7wlf0L9f2SkuFjkihXbdqjlpuR5iJn
nt7w0oCvyfKofVr/GmWqmB8ewd0/FUtu5r1AqGwO4f+n2cjQ9z85JetL2RJtC0ODGGAVrOeS3IUh
OC+mXOIlpBDc2+Y3DEU6hfjKexVumOWjwVUeKVw7ASm+4aQEMgkELfD8KNOGJSkoYnxTmJe9106o
Z4cy7E6TO0rEVckzVM3X6BsBzv2NemeiyDTKiosWRvo2RVFzCyg8gTHYxtZOB/mr1LpGgAPxJkNk
H5Pp0nVMQKU/QaTB3jTwmpqjCv8MiAbsjqTVNunDYqlv6xTNbMeFU6GhRtupenO5V92OXi62TJlx
W2AMW8dcT+BMphJJCgjFajT1zU5zgbl+WxJcYrK86B4+QMQZti6pMrLien6NfrwCf04A5DD06jA0
kvIO5nKByjkqTc2SygO3BemuSIbfJtvKDEbO/w5jaP/rP1zJQYzWdXmBanTZDW9xDHCImyrV45Go
MJQmu99iHjN+5RckHnn1D5HYvH7DBd1Rho0Kdi6uXsN2VPyx5vYEAgAyQqZEehLKoJ/AvoBWswdC
PKOs6CUvD58DCEnIGkzjk6apDcKHnj8xZRq8jKG11eC7TQFU/N3KOZE5OwmHXrFnkY0WZebcoAX/
wk2zIbzKOWnA+8qrOQ0HzGpOtBKg8+cc095UjWoZpi4KgSWQ1NsazXoLD7/ggqWKWo98JiFShdej
en7PtbXFkVX8cvCz0LA5NaaMJ2c+QVznMKhYkrQ24hxa/or51qS5YfBIhPfmGfDtSDi83oHuT9Uf
SB/aEcoNKKZ5TAHc/ki8icGYeg5oux35rHNVXXs5la7sBWTIKk/jGN67HYHRwrBNz3ZvY1lXJSdF
Fp0RYzSxKXUPzwD9J6tgMdmpYCZIgk6PBPB6KQxYW3N24L1hALZrAzc+SROAYOadIB2vE9oDl2Xf
OOf6tDWWmBox+JqK1B7dTDYPR0DvQBaL6idpdT1tNfKbPEaLh2I35vF/tVvT7e28sEve8Vl+bZc2
vI5jxOy5knvqRj1gpp2FKE2LVvYn4or2nENhwrHDHJg60XRYbDyfA887HZXacK7EXIAkRBg+h8HJ
C2CLdvPhyNKRzLT2Rs1lnu713kU3skEXmrFaVsq8vWjgi5mrHcsNgSmZwXjuDu0LcH8A2NQ3g+2v
rIDxjXfQF7Pec0QrOFob3MvWomHlfzq4fmGYPFmNvQFLNNTHCY87192X+vBwsnNMMdi3alcEv+Hn
FgdCo/XFFQzcCw2JTrt2DtVPaQzFt9UC1DXrWgG86K+Ab3t1uKnP/mBHYVwTdkTmMQTdYFjVGALh
mvyRw0sRdRMxwPFqgZS6G30nbcBu2awbpfJmKXnbInZZXer63y8VkJUFt9mVy9E2KnQuN+It4vDf
a19iY9th8aHz6QJ/VjDOAOO3I8TnUAxsECEEVtUqxgQQlMLCcBaTWNxOQPZ2iKC7B8G4qZsr/3/q
KDgK5ZfOnitVpUs5Yn0DnTdbLsDBbV4eRtGRP/hsXc6XCG5xq+93fht5oRzfZlqraBaKdYB3u6Re
D8fs54nup7fCW3RHD0Kzsn7/jaoBazD5S6phjgqEeYIQKwDydRqt/xKr0BDWJDg+JRgcwFLGXXsm
7HD0kHkG38+8YWCcZQBcjFcg3jBjqW7TS1Kr4ZibQleWqQ0N/wq0oRDT4RuPSfRXXEv1gQgO/Jc3
w93QALfSPdo75TsJLqZ0sN79POUX+Fk92HLiYlOP+9xbuZ3bqMJ2Uf2z/SkPaNwMESzSA4YYwfya
r6i98Aeri6IRm+NQ1bNWirgA4HoTa2uIhYEKF/mbyhKFpeZwhO4B0ZUtA4gLY4R7VqTLwYdE5K9T
XdP3zs433i92jEU9E2b2gTuIpuccRabmw0g4iao/A3ieOE1KmDZvskJKa0TTjO258A2l3YWEFlim
/0HRGZkvHjVCSzG/UTApci38TPJycjj+4nEcvzSpSeqX0TeBM5oCZh0JyBC94otBFDMdZkrqBrfc
9VJIFvkPPmnWzDKJZKdJOoqxosDO2UeZwuMFaeCW9tMDPpoHlensq2/tKOefLyyfqCK10XOvcuhV
Gz8KnKd3ZvRUkOrYL7DwXKcb1l0VIGiC/4kj802/G/LXTJ4mVOU698hPF5H8ltoRV4slYSZ1lpSD
tYJWmDTMKAUMKAnd19bflEScBKneGcHYzGRJJaozCnKNVLSFUb4l1PVofyYGlPdTlM9BCLAiQFYx
5dP6d18BCY0GS5UPwz03C2i+7C8ZYHkreX0CoO6pdQciWCVhafMlz7eziup7PBhlekmISZnkRzGq
svOMLXFD/IKVq+DS/ZsfgsXQ/KwIG1PsM7IOYDE+WAjMcDfXrWCVuAiE535NKpDsM9djISIgPMEG
2BnEEm8OLxVsxgjHec8SgRzbwmho9KZ4/5jZd/u2GxE4IwYfG6yt4ExpFwZFXDfaaDghoVL3/G8Y
wloYEAHyYVQSOB00F64dV+hIJAjPTKROhQB5fX7fivbN6YFW5xzzuGpxAtVu8ANABWUUrBwU8XnN
3r8Sa1Wqa4BpFROlPa6Pc0NnVrIzTmRP2LGzNCojcv9q6fBIgufQiflJQtHpmLLtdV59FCIWdV4R
NVbo+d5EZjKmTT9oINoQXR6bvnRgfY2SlUcAMDvATtR4j6FVfoN3GcBZs8d/PzXgShvSiXJmwam5
kVKgO1tOli5b+3KH224FGXtgHdPYhVKKzSNKFATlY35ZxxthNEeWrUEUlHraLXjnqhF4Z09ahbNC
9qCsLXkLgBgFU5DzqFVTh/Mo8OcQL4Fvhw0SCMeFsyFteedmlz6uRU17isEgopcrko/aB87RViiz
wnQFZgqy6bb6iYEICJrF4mTHqCHBO7uQqCC2EUX7QCGakL+nY0j1eGfVtjo+m4BKYrOhcvLF2AgG
oxaqC3GmqrB35IpZoTQIxE/P6YJ0UGJJd5Eg+uF2fbW1d4Ckdm/6+Wo8PHunhVEfV7BZpY4K1kpP
tyiqvGb/wvtSzbDUVrC01OZGj9Gva0F1dx2OfbSVAvulFZGhhRQBdKdjaBJjT/1cfh71WWIDRKBP
tK2RYnvC6iyqVUA5QFv2MdAkg+CprmjB179Bq0aDw2dqSmzGhgvMq8vgHp+stRmc44WtACJIvijU
zMoq47aNXPCTefB6Zl47zfRgixG9fD0+fWe82UTUfDKNvfo6iKj4kP7OlbP+kCPBXn8kPv0t4QaA
jOGQzMt9B4Ov/LY1fGHreOEFwjFaNbez7Yq+ZoSpVWlQaEyt/0IhCUvFMTt9QEaEjGPBft3r1UM4
GjyXu15XiUuqsOb5IGIKJUegcDb3gpkHzZdoGQn5rhZNTzKYFRC/xKTlRh+hiekz8B0Ug6jl/sog
AztSR1LtUJSq/8Atc5/Gkx+3RhHWeFOOOSN2xmEPsQJqt0WikeHTDf31Us+eGS3Xca4+gFtMOvNb
UAuMAdTKPtXV5LS/VyCQYrNr8A8zV48mUm5ye/AKwb3J8pNJvqxCpnW2ZlISdgGEfh5Nd902kdMV
W7W3iXo+kBsWrvXrQR3cD5q0SUqzJ1Pb12r/oUHnkubYYIvY0VRLKybBQuMoZNTAagXM4EBgf/Sy
WNTavPFqy+/Q3efYWK+1CtKC917shQhMRFqV3Vgm55ebK37pykiPOYKCgUFk6+Vp/ve79xO17Oqn
fNMOCA7ChStauUZ1qVa3cM05G6O8BUlGGQu1vzN+P6xegGOty7uAtMl7xxExVI2ZOGgMOVHXFYop
61UIqlQh8nscihVYRuWW/uGH9M0HNsHV1ZQzLtwV99Q88gRjTrz5QiTKOk62Mg1izcRiwv2Z/uw7
Ey1zM8i8Nzd6x93VelkCz8/7XZdy+t4Pwip1fgxtjCYLcKjnTDOEE5uulaiN4i2uEs8dw0bz33Q7
pfr92FKUbFzP1YBWyTsKinP69+MevdJzex2a6AQ+3U5AFbXRLM7nvQI2dIANyyopY/XtX9O0N1fz
Z+NcZgp7Feaef0/CaxK1xOCctbULcsxpwoofuBjrGbWDkaK9xCYsT8cjgD1A1ZCuCi8h1N3dw+oh
7P0rBp78HUDSguSKZRmep/OQcy4Ic6OSHAZFZWlTbZaC/U0XDcsaC1IeU1yT89Kj0EGTuB7sVv0J
O0rEsr7UEwauv4qcoAvptGrrJBKTqtmewxltXGvA16bEPHDFdNZFwKYFVztJuxotBqwPeUq9qLFJ
x+7L1yxwFNWfI60hDTktSNc3ScmocTaNWwX6HK9I7zOtNDUwOwq4VBs/VB3degcc62EbF447PGVt
ASnvjQa746MKh+qrNl+DS6fXPu6FlilK6FcNLTLj8Dtk/CqvekmE58/6A+zVMkJEhQuFgjZmLGEb
FCO6p8tDvAdkhMW1++pD+1tH3Wvc25a6oRdAMzjZ9bBtERo0NV26dI9YSuaHrgJSqAUKOy3WUvDq
2AxfUAJ76ugfvZfleZFfhcpgV5pdXCXPNaiiDzlwX4OKMHjVnVhZBpSNrOEMSgTsOgfJzmvyBWil
xYGwx4g/Z4GFrNvNHzJxUg1HzeoSuRtHsAc2HaYOuYH+NZ6NFPvpSFv0NU4fxEuWi/N8/DcmexzI
9KHdm01QmBdXqq3/ebFcAf+Ox2WveBRUhdbmfi1r0P3e7uWAqfebKiopN1mHLsFnu1V6WIAS4hCn
NkgR7eZOJTFM1I5Z/Fy8rsWzZV0a8QEHNrceLWrd18naFZN159sDG46iUZgm0gyF+EB+6ObztdXJ
Zf4ibHnM4CfXYYGyKTfCl6lfN2ggEPlYoIchey6wBBCq6kZpv1sx53E917ivsAbO+W0ZeZWZzxC4
de/SBiKoQcNQMNvJLHqucLFn/Lfa4iDCqjyPtevy3e0nI3T8IHqobPBNUWWdA28fMMwizgQu7Xvi
FLLd7nFL5ywkMoQ4p12ECEFWn/3RapkTTrZ/vaYCQtHwQ/IJXymfatHyE1BvAgGqYl+lmHhCwua2
vkI3MPystsZYBRA4xJJoOiACEfFeqZzUdwbX1Xtv1IpAe5LLqKKK2824WAB/t1IsXjNUdK7olndf
XQ65rJNc6IvS79CsuIhdFiF+YB4nQwxi/CLwSY2M4iBle8GNHLmXmSxt9zQ8SwMhoIQaMQZuUc9g
1eBrrpt2aUXiWZ1v/PN4ZZ2wHI8SfNFmV+JiJaEs5EdJGcpzTiLH3nbg0G+rNteNz5RLTSq7VMLR
p+kbkcXmAa0F34KJ3uG/ICWFxBMlvgU/4QNebN//O78M1D3+ljWg2CsxpGuOanuzJGWwOGbFTC7b
+xwhDvntCxft5BTJvB90LyB2r64i3QjnHzG6JxCpH0MPjBd+qw9O+WFQevXTB9xz0DE0ylYYMiSa
Ny7v2xbGtNg/JyNCjPeweCd9iXTbNwSkMQA7QU/VbGUUI3UNl3FmzGXKrDMJgcUuoDP0IMfp8gZ8
sY89Nu1plWJutv2AMcs4ebv0L16M+XqpzBxlRKyc58lxAoAPAxKgU4+XDcLATAIsXVZVla4q1+NL
YD1gxQl36QiFBXqha8GdeDKLO1PVUfS6VUG6bJS9zXFRntuUT0HSy2Ss8Y2wGxs6Ob742UlX/DcB
/yO6h+62+E9A9C8kDvdrGaI3NMvGzS8QYM5i6xxXp7b2N1Jafp6J3zwo9VayWW9Za43hDsoZHpfq
qGsX8tkyNxt+abz34tz78dVguUkBSkAhufETfJepaA8vK0eRDhDRjsqcbJMzlQCb1rXQezsgzUEE
P1q1WYaXLLCWqUqlJ8R1wzyQ+jx7AtW3n11WYag51erqd0xZGP9xedbZhKqL6FsMQODdXFOS8Cxm
PMvBdm5MFXWnITCbyAMsAbylJkNkFy7XJdP0IhCdysWT/Lf6Ls9y2T4Rq+DH7zRJv/QdHEZztknI
Gd9POhZr1yHb1Ym66mihyjP6jQPT7Uu1TIa+VkfNm/nsxMuQ5gzGFUPUOgFrne1EDfTkZxZ3VRS8
mR062wuyFqMip4I5g0N0FEvKKatKpAO6zbd9EbpXRNB4NWebQote+DaCZicYohQ2ASOuWQBR+LBM
ri9aGzKT1tMOSALjLEe3HBLOjZG0eBdMvFuRM2hP1t8vV8PN2Y2po7/5sUqf9bW+pFAvKKlNcJPD
J1MGCxJAUuGP2ITWlb7ym7CTy3/ctv8lYmslvxT5Bd6WSHL4pH2A0KoQKLs4uVyOky+nN+b9Jd7d
6DsT04oDwPJzoDLE34YJIjszFK9quGlqU5oAtiOTfM/23Esy6Y8UWugB/b4BKcdV9u+A30W80d52
VieVIPOgQgXIkuZTeupJcbc+mu1iItlPX432DJzCHYNYfie5XY64FPE5omR2vJTh9knAx3sIiUrx
G8ePtLEynRZYHkp7dxNHmXTeJ//ykzKA/6BviYS8mds4yyld903yuqHPywcbmnfUThIobc0WL1/g
U0HMWbjRtQYW/DMy7/4v2i0YT5rtrYLGmzUUlkqy3owXpfQiQhpqAMdqenr6mxI8wROe048mr5wu
zU0xVa6wV7tZV6ioBxCrh+gTwj8NVgKPwt5KbC1R7IgKCLxDOWJx8n3Bol4tvb06sgjdIA/0UeCa
f4Q+X40VPk8nhtgVOtAvi/62E2UOR6AD0XIPZ5w/cE98YCE/E/XCKqtyEUAYs//0ggUJEf+dulpD
SJzDG4LSuthKY46PwfxL+4dpCiO4ZT/7ToH2qJmyy2yt682JJypcSdwSeBRJOUOcMm+SCtytBtqc
toOTkP8Q83ymb5oxKkkcAy3OBaZw85NS7LV9Yy51+eSqhHYEVdYjhH3LML+xWwSePQ6Dw8muHlnw
O2vx8/QosEqhM7zR+43gB0rMuZa0OSQ3WmyrILy8zIfyKrH9g8yc3SOdsP0SN/a/HFDNi+LVHhMf
/gEYQqBPiNLl8t16oH5olUvRzPzD/BgWCslOidDErPhhLr3jtme56Xi4YzKsk4+AtvzPIePHuxTE
/djsN4kwb1lLjqtsqrQSftY4UoA2eSsmCoGQN+nus2fxfqlxkA96IdNhIE0lk6cPtwf15VDT/9yn
8QpShBbfG7PHaA0cXatWnBypkfs0BTP/L59BLKHtqvipbnttC11Vnx6lhs/bRlNPZeHxy906hqnE
5PQx8C8BdPa7o1N/2E4G2TsYS1doWv6GRy39l9hE+fL4lrDctOISRxifo+2pJ4n5XFJ/zvt5BAIa
BJB9Ulk5HHGt9Bq5iYfQVkzLerJvKQpBW4gKIjDlDfS+vV9h9sCVcE21IdF45gYpGtunhIWXWW9o
Vk2Uk1zMSZNXMrXSEBXnrXRGkTEN6UnLy9EDn53KRyEzPLKgYqYSzjhAbyXt0PmSsZKdagaDdBHx
Tk6w+7mz5Is/VktN1CcKyrriFZPbow5fUigH7/1t2U1OnkR+o+VPnA4qzBJzv1gXukD/qjyFJOCJ
0N6I/p1zDGXWOmZYUb27faQFH1HqQm8D4SSuRORwQaWNJE8vMVun1KgzRpfUuj0XPdvFYU7pFpCf
1/27n+nNx9h6VEL9AxXMHUcFaf6sGmFQpTI3UnuUTKBEavSHGdID9aVO+t3qnjcCFRRFFj1XLJF/
MwgrTTGF01g/pi94iADea01mpRGuSK03WNriwQLrj39SxPyoanvnRgf3G9D7Lpqq6dZMyJ0Pe4+A
ftfDcp0wtAGfrrUJ9tP05pJr9wPRH8xgjaMclU2/UV/2X8LPjGj6kC9DzmsHKzCL6TNYa7NgFHtK
FvlmInQsYlL6/emhOznfEbi2v8aGes8nDYqGWSi0IeHMRl7hHPrpxyEJ70zjcUt06KfCleazOJ9U
XghXitm6i6YLWANZsBcvCb6s0r/pv88H3bjTw5fbG/LdMd9tsFgiQxz6dDUWCEt2BqHKv56Nict3
o4EglsvQncMxsKamAx6mxfq56zi1oLbiuOKVsgsbgANcYAW/oEgwJrs3Cfn/QomA2eRzN+SZ8JBR
tpi4fHdj3VDOd8CkqjGIevYd/uGXgYYqfADQjvGTdhXZWxW9duT8YNA3GebVPjYkicjKigTXjw89
U87Gq/tQ9oHbRXOXl7s4S48gjfk4kvokixQyIC6luhanQgHunsLRd1Jxu3qZszr2D8AlCJVbaqOs
RPXbq4rTgSvudpRa2lsRMnA1mrf1i5Bn+gDGym088OHq3OIg9t7cSQfUsNGNmP957QOjSZxgE9x4
2viorG4z7V5VbShatNBZp8mhZ/QIFgzg5vcf9mMLIia0/wiomXnsCM6UNEjadECPRTTMzxA8jh+F
rrB9QSQZwSCtprPVpAZ+Bpmbp1CO8ZhEPFbnzi0dzGFb4UvWjSXoADw3NAbP6DlEElgbB/V4Np+A
vL5aOikD9gWyF/wFzqRVRv/uVFomRKm7pGVC6rWPFkMO7KIOaIJgN/ut3WrefU6Wb3pw4DzmwOOa
HzSp1fXbqIN6oFay+fBNzhqDxIz6oWGL5lqNcG3EKbxA0ASRDNu2+cGrw1nEiiOeSfbRjXLU6n+C
IlcHcdizdlocQGqdeeKJc7xZFoT73PtAukRT8HNFMz4b170v+QtpgnPF1Fxrrbwk9imNUAOM7hf1
Fk0HtXEeE7HEmL3yfv9KQGn27TrYiv8hTkWDqPx3soAFKjJ2kQ05AhsxZ7LeswKCnZxzau1XyyAZ
zR4oXUIG1atuIYn5Vb/lsW0gq95nkkxGx8rUmGA1TsCU9tlruBHEGff481GscjXdk4mEbl9pFk/h
S0C1Wa3mG4LmUMhW5fGgNPW6WxerLIH9LcYtfwsewcqTnk+/OiTyjq2cTvzOpLigRmGjPmcNq6d1
1gGXAFRzQ3qWyB+XBq7nvAEP+LKWZcgNqHUxiO2Bd6k8QMsOka/Bn6fYJze+JHt4do289KPBMNKq
Flie376xJd0ro5G8NGMFenNLAz+Mc9MdLeJGGr8uLyyGBYx4yTC7yZSUhpwmSs3MmRkXnsGOk4M7
oiqDgw2Ehcp4zHkluv2ytqZxwGRecE29yruh849hN5DSO0Ol9DRuRdsMgmN5gr9KDrJMYiQ2cJMj
UkLSv8XE+chk2uZmH9bd02BLmWXmjLL3TBuus1LxTLSocEOufSE5Kd8PnqbuB5dkvz4zWguXoFks
hP25TcLhk8CINMUlcvycsu4PFao5Uo1EZKLpfs8AeDN1AuuHQaGo1em1ZPMKFC3eJlQm5nRoGklX
sGfgDshOstb+Ic98UoioaMg7PG3rk+vHS1ALWyAsEYu5MPWxQsfiRf9svdnM8KXIBd9h4PHzISlQ
jjELxzfgwG0Z+hGF5BJaslTGpVbwT4XZ0lZ5rLd832b+et0CIPGU9vBP4bM3Rj8AFw/SgLUHneGd
8DQ8oykRCymMFFohqmKZmxxvSO0INPSwD2XNCOy4AIL5Bz/tget99zXJJ2O48orv4roJoY1Y5IJl
phxCkWuYDb/rPgF+NNWJtBKyEUO1tYR5jFW1eegkB/KKgOYJrijTvFnrqeLVmtF6W7U5IhLIZjZq
5UmKZY4w+jpOe6QP/yyHvkE32G7KRDPBf1uSU7+4NQV+layDaFufYMwe+xpTkpBxtT/okAxHoKJr
hkF/pQ3vFg/cf81YTuFUYf7RHKYE3dqgTVmLdVpaH2dgvynq3YI8N4vTzbxt7geQsyJEOsOfNgge
e/XcNswNmJznl3HeNrHi4VUp6vptQyHvuAmbZfVU87zMjsRuywj9nceoNK8Lp6os8U6wXo3NAmSe
bmIOS8de5MlMUlA875bnMrdenbllWFoio/EzYay0Q81uOE7XY1BVh6ZPq74k1CC5oIgm6evAm3LV
FjS4TCynz1gNNB6BqpaWViUbZUymIZ3v1/u1l3seLfuSKQnFwhd7yux//VpHtAbOyTLZ6Vx8QtaC
UFNxFEMWK58YWx3/Bg1yhGX05Uvea0rn4IKf0ZP/K/tuVsOisJJqcWDaJUWDCcsWkLhz26gz50FU
gR91KTGILs5DmZD9cztoe12T8tEH11pVUrf+VI6Ux8HSz1B15jvMZITNErS8EoI21nJsf3fOcbhw
y6N1h52Bwk9L+EIeBWmskL/8Iyv7/QNnMtQ7ZQOH0m2laHE08FCIkSHclvVzy/7xnxBSmYUYhdv5
sA1fY1oGt/0gOXnhYiRhIgPTHfjcTLzIATCHgppCzAa5WHoKBG9FNJPC0DxcDi3Hd2CRDEzyDoPz
4ldE39h1r7pbuJWe1S0xg9tEauheH4AL60J5yONpETobqwNBXBcKSsVAHcca9VpmmbLBeJGZ08ds
XBj7vGDuI3IJwOP4RV+U2hZRC5GsmsTcJSUej06DREEA0MQu9wTIbymkFXem0AI3i1qv0qH6BZzB
LM9DTvkeCgjrgwoq0N+WnkBBbToVBTlObbTjEkIlVBo2hlfFCjtvPyhHnL11QvOtC2P+zeNlhBdY
Xoe3ol/C74lfUSvBBTDgMhhwRSq95d4S/fbcs9qEysi7g6BUxpblC2RGYpjgPAe8VtoOEcfiIn/3
QElfcv0s+6EjKsLiXjieT0wFfGYJ16DbIIyWCyOrEJlkiVVP4C+T4KZZrTv8ey+Vw7pMi6rNoEy6
XlteY67AB1cTqaBd4m9FyPm069fvUMw3V5eQ9Glb5+2l5kDKSmj0C0zqCSxgVvck0QZiHq7Iq4Id
7pXdpb3RtL07ba2/KUAp4jWqIJaxDwQWoak22YjVzJwePaxq4tGsVjapH9JJS8u2LGHqc4W5Blrj
zTYJ5xK4zJOj1U5EA+a+6+pg6rEjL4Y89RqWSetjllPZh796Zd+Dy/7uPZITZPygW5rHykFR2xeb
49/WeCNBxXdpZdUIH6+FY0QSR7ZkZOLOzSjeGzLI0erskT33B8J+R+EA5UY4GMkihH5zw5CQlDD0
0IaclrgO+l3C1KktqQ65xfny3enrjQz6FPjCwVYwC4GXBI+u2O7yfaNMDzowIVXLbN823i8E2h1I
XsFD1sRXc6ztLDxdcgs5Cw2n3u91JqkxLKW4hDO9T27N77zqk4AaSyA8LbWJyJExTGhB6Tt6mWVv
iiQ76AzZihkfAao+4Plz3+v9QHcY91e6AMOXCP/iftLcinBkJs5OrXOSOpKKIRvh2LFXMGYVX8W8
auMQPsbkr1DBayCefhl1Koo4tYD1N11+U0jUUOeDgQRA/1/abb7dtQmVqtwUxzzI20RgIqesTI5x
TB76FSYSLU3qvXVjdI+iDFgPZXbtZidG0FajHugiKOuRCgjDNoFG5OuJcDY2/o3+z+NRccNwZhJY
ZZVlcDkTR1/eWddapmouWzZ1ics0e12IMFYPkLkyq2xIVxh0l8poIYg47icDyZ9CYH3B83qgXfhY
ajFJMJqPOyZcqp5hJC7UeknPhSSSItqJShAghYud32UNMkrqA9WAFDiliTVCLTl5ZDRMXp6LDJFK
GCMB9nW2edgmNpDDAoHcZceMMediG+7uQG0ZU3k0mzX4uyXmhXoGHlQfJUNCekqUHHjElmltqn7w
C4xeMnGQupdC71PEs84JIH8haHOKlXeDUv5W1/F591pUb4sAK+ENrBY2J9WN3x0gdzBYgcAnuP0c
IDM10Di6+ipDGfgcCExSoRECauvNzEqN06jBZYnDR5xq87dN+hfcAJNgze8/1sjQc9L6N8Hf06aB
KAFAn2fz8ao13FhCXk7Z5T9FZzZID0vRbDJGSS2F2Duhu6eHRIWWbuLiRVukifAmcnouFrptCYth
UsSqGCV1kNDefBYah2InkRCSExSDsrpNhcCtmBWK7GM/ICE9zPEnJ8nCBKBx+9eIJ6wGhzwGtp+8
TUWpW2NJc7Zry/0OMiT8tBb1F4JOa2HyKNcEwqThtMwWut1wa5Ady+8MR5YRKZX/ykzcjF/F05Hr
JblV5HhkWeVDbLxk3T6eokuJPlxkPTqblLHiaooeQLzJ3o3JOB3AZ2UB35xIU+yD4bVez12c7bdR
cZorDm+CPCBG+vIBCdcan+TsIVGivhKBguDKZowkCMS0pNzO80CL9U1j061jTmJfaDw8qtgZHXrR
yHp0wKDnulWvKmSNPm1dhiQRqEa5l3i0eqbt6zIxO7L/g31UG6S7o/WfRiPiVQp3u0Fg41Q5Xl4q
NI1wG6Ul7xinG2yykg2QAaMi6Qig9fG8XP3acAjrx5xbFm3O7dJzOumzcb8SSxkk6qmqPFywXjzm
qjyX3AgoRaMRw149K8EjYJXM4GV9PEz1wmMd7mLhQhYtZ2Av9r91yOvLZy3B8pVYl66ix2mFAyUX
VAjUGecyApGSgvmBr0XjLV1e8t2nEenmtC10W3h04jo9EvmNvXaiV5dnO2goyC4XELXrGUxXMigr
+0mh/MWiyHQMCHii4DBahqCFODSGqRET4tZKjz1t1oe6sjmPX8yYtKbAINxYAQovAyYj1TfRDC2u
wAZT6d9UABRG1EqX7UXKF57Qg5YNhSBfo6lYERkXGwt0bvny0k+1l/kxjL6yqYa4R8ovjuLkLi69
+sw/fQ5ACsy596fhSih45KSbL3WgYtHL82wR2HUpC42BxhetGqLZ3TVtkP3Qg3kJOs+ihN4ZAEIQ
XQnJmPULH8uQAFzDvqu3rc9IuL2K7Wvk9mAVanSwIRxZeHSrltbi6ESdkglHG0zccjoeNp/21E97
3a3ArVbDRkN1Xtfq1G0J6pG2O3b6huLamdA8AohgRTlb0olLPGWwIZ0oxffS2G11DuzajKVznX8q
sFTYK6nRDdRZdK/0KDWKi8nRDsN97wzLGEyVVcExWdP3gQXROTINf3Y99/0s9QqNHpeRxnh9Ggm6
PzDqnVqCqjizSoGzWoNCibGllAaBxa77tJQ5HxupYPQR9ot36nFiSbZR3EbivE6XJ64/LgC3jiIx
UCqdtE4vn9rgqqPOqBq/GwIkeyZHgR8fhWOxfrhxX3tti2G15dpTfvlKSUWGze3h6Rv9Mb+CRoTG
boM38KX8gXi8m2fnADBzHxXi9xXTCMg0lhR63JPJITxmu6pPCUqtWNeKu1RFhobQxigiMxZUneYp
h1XXF2xtl+3YLFv5ekgA6xOnc7s1Pnm6dM55as1nhrwoXmpTlC4samWC5hq5Qgd9pYrX7JWc9aF0
lo44RIIRVco1fh9rhWaIHhOhy8Lx8EwQTUN/+lDNU3+OjklF2OGxhGwnVFZNOVA5DCffHJQZA8ap
XQ6m7igOnk+uZZA2Itg13nbXmK5NkTEvew90+R2+0dAdJtzio1drqVB6mwpzD4dopq850iRe2LAI
vi2JGH3+IHzA4UOxo5XJxJqY6yejxD3x+f6Fm/gntfU7N7l9mj1DC2Bc1X0oBpBYpI857dvoqR3Q
QkhdZKTo63pYrOTWbkz8PLFyVrDEoLlSSSboEI3+U2aGQxdBildUToow2VwHu/QzdJtKqDn1pTZ7
qF3zL4tbww51t3S+Mmdu2PxZl4sTgCAwbl5lQgkYSxdpes/g2GISUVlRHikBjbPW4gUNtPI0DQ+H
U3BWHRnEiSpZPnGx52yGW5QwdU2mhugYN0HDyCrrraf0TkXgTZWMX4JIkTrVJrCHl1sIiB74/D03
JGHtiT7HUxp/hfVkAe6/gY+ZXMCntIWKpgV6b411Jf5JdrJKHTrbWdIp2sKhYlapzBmCCfb+n4RM
bQImpPr/GtOKp7x6g8ZEpy3Zg5p1RMiLUQaaMKVi5Mp9GKXv8C7rw8QXQe52SmNnwFIwH/Vg0mVF
Dk8n3bYYkY/8g5qTa9qWYKvv3EkPdQ1YNh9ccj5rB1NUA2A3IXoFDv50j2UcEUnS+3JfhDq5Rxn5
PG4BlOuYuN0Ip9RuDjOXuSJ8NmUpidyAO94uNS8eBLJixlKuzHw+7h4o638xOY7BrI/P9Sho48ob
3+hYXT5rGHMuDHN6xnxnwwTOyXaQUFKRPbHj4/m110lr8n7vrl9x5g1c+o9hYjW5rjF4py49C6IP
D26GrWxa0AKO+T94OJgRmlBKS3mmNv7O0SlZ5Ou4CjNAuiSZUv4OJ8ZhRKdO5xyJTBP+tD8S1Izh
IBjyuDBfbxPqUH4B84j3zG5tjzzQsRuyvkE7KRPjr4+d16YC4XmjPf6rFDfRhZn7XvHZv1OuxpCu
YikhmoqZFgUK53mDoMf+FGwiUS9N3nYgrurIPEybrttfn+0sjgNHsvPvFGHrZvbWpHbTm0KS6Htd
AaNSyu/+qM6a6ZgEjdS0KsXgN6BIwFnnoGxuhJfQsuqftDZRZS6WsohybcjkZRNFsIm9vA/mjc/W
x+BxTp1Qy9qumgCHYXnHr9z2jpEeuZkRw3S6EgAiqddbmmgnYXL0E/Cw3/QI4H+T1MP56ty+ePI5
CLUbqGpWii3euGp/OZWSxeBy68YOc00wpn0JoQTSmbqycIdTK4pendjY2rx2UgxF9nVUN8lJfUMH
2+nR58FwGSQDsdzV1EVILK1C2ygfhtaNFA5fBppkD1VhjNLwqfxGXN3v0WnN5fitnVI5kwHhRiMp
MoJiaWv9GRvMCFdsAblwXlhbxrhiIFl1gjdQBHSJRdmiZcgVlYM+BpMdooMFAMEzQWApmNO+UxcJ
Z+O2IDHViMVcg9O+ZA2LTd9WHpPkQ0ptCRRyefKlSR1FWaUovjZlRBJ3nZ3lZRbzEXJamzUb/rC1
/xSeSQCBtXTlSqOM+EuRxbRUJ8NvTLs2d6Ec+Z/xSIyWkQkq3TbJXo3W46HzxTvYMVXkx0Bqfm7t
kEyZZM/aP98rgRUvrBi6jEtt6eIGMQORTdvi2LKnabdRUTSCv8xa/zl5cUsv4t1v3VJksuUAj4J0
QdKWu1FLTh2fqiPPP8xPyvggWqiiu28dcgPACURO3d+UCSgO84QtQO/dgmpUwI51RCgWSXcHFN7o
iX+5N59pTkoB0s13/cROwxFW15yCpas0dvI3cdwyKS+10QVRECOVnPNjktZtrzWrHQuCAxXhOcLm
GUuc2xK5Q3f1OzVyJBbFBOdDWJevRuwQsO7VHsvRlZSAzZjT0XA4V8jNh0o+z6MORdUKgT4McCjt
54+WJVK+ACM6MpZoQnNUylNjyb1j0WxyZcmkHSlQcXwzAHW8W9HY0b0Es0iZWhNp2vN5ROp6nz9n
8xpvuSMWCD+GxImwJ78+oSK74ZU+w8eJBYbzsepa0ov7fFws4DJmes0rdRyQwVAjCcbwemPkG8XX
LnS7d53DpZ6Eg/hHgrpdfPdX+rrEePTp027+IrvS2XzCZ+rUSCRcF63v88k6wdOs3Y2Y+MLH1USR
WI1g/0O3eWv/MREi8dz19+Vpu/syixlz9+CpiGfsJwXcJKqM6Aaalp88bq5WNrAr303cMExeOWIb
FPmq6YrAEHbFMtY1ZJNFITTwSJ96ASkYuQnS/LDKbTy5ebQm2etA0KCuMBFQK4Jvn2HKxRmvGqRx
acygzjJ8vhxgFjX2bjD/8JuNFOZ1Ix77vHbF9Z/qFrwaK0uXbtqb0JaOSvvoTak7DU+jb6Iq1T3u
rwkX4oCwFByv9FEg7wIMvmGVWWhf7fz0EUsDGGFYTVCkJiAOxI3rZ2BlEsJW9OkXt0bUn1dAC2Y4
NTXJQP7O+AzLztu6M1x1rqwBP0A3q6V+P2j2XxezTI40Iw1bG/v/d1noxr8IIjPhmUQmo2hYGZX4
QtEknjzhMT4INAmSU41WYL1EWVUwJ1xW2p/uamO22ll2XSDOW20YMfsEjuEaC7nl0J55vpjlqP9r
sOPK/+cBFpa4Tvf3LxEBK7UDEVhE3xfJnpbS5UwlyZrZenbmz7yGu28igETf9vut3UcRCcfvOELz
21LSJiS4bN/XB4STsQm6eBPDz0MkdXUsqtBMvYEc16frEHTpFqgn03AcnaxWHuqL8vOocxgO82Xe
gtweg8Dbu6seBzSp231tJydxu5g4tj68DophmRMlfbTfAGEjpeuAXpc95KRXK1AXxOuz+K63Axok
Zcv6XF05mXpzGrV192Z+e4SkbPI0AAsQGFs1IGtKnUXePOPIs9klVjC4VWCVge8x7VYaTiSb5STt
GS1oKRVSIJsWdBRVG1SDq6oPe7tX/dO7g5K+xhPNRWYGHvlh4RCDjlOA0ZOVRW4znlDDQ9/xp+vR
CR034IGZSgWH2D2Uyp4Q/mQBWbQiV+VmtiSks2A9V8DRiYJcIuE1UJ+nTdf4hdUsj8Kll2BoWpU3
4VPFgQPNk7TXYH5z0to+o1izNiKdj70oPzpPw/a5Zxx2NAjK6qT3uAxAbGixCl3Wg7M1xDyYa4hM
CysSEkbzPdu/nn0T8z+5B7OCqC9QVvGXTKhLU8Q2vEXz7hzMLuH+pQk+aZZYsSCkB0/FBuLFrDvS
o3z4HGgvEukf6ubWLfn5Whoa53/QdTntNcsCja5rY66a7ZLbrwjb8yZKAxpy+ZNstNI0S3zzuuqg
1w72blqS2gnP20kuAUBR3+i6tx9kESVR6XkQRf7qG1Ue6fEIzMVhXUVJREd+bJyqCN2GeLPMSIAN
SurKjYWLIC2KUUzu7F3O9LfM6XIbtvZrwsoXhmtL+Vyr4Hlnqd+Klrv6yadva6cYr6QrUKvJDWOs
UhD9I9woJAIQbXTS85eiAo5TZcb8F0+2Q28nHILnVTGYHlO+KZfGb+Aap7ljp9w0uhztG0xAldmY
pIWjKtZ7omiKXJzdvDALRsO+cRs96kBRY1DMv3jt02mkT1QquyZFssaPV47TJW1VFWc6RqFXcQns
HroMelYW2KityccmJ4i3y3WlTCXB9OfVgU3XkYG29Myge5IeM2a9la9Bbuaeyy50K0GcwTKblxcJ
p8KPFdPPVUX05ScZu8vNkmOK7ktPcc2qGnSx36Tm4cD0VaTyfsCKDSKiT8k8jHwpZedlgOivcEaO
NCVTvSV9oLsWqYZTMDy8BkgC30rtvR7TtmUtDGVz69ViShT4MWJsmT1yySdUxvFrD0QIItmGTqD6
Yad7JzQAmS1I08vxKALWemeshIZFyrpxewMC6h55+X58IgitCX22njQLRMeMx9AR3j6SmLxMCsG4
G8k1Pi8D6FRJZXOvAx/3Lyy1FG+3dX++UiOLIl7SmDlRc46ocaWPl0KfAEXsi94GSyhaZmYXxASQ
QYljrXjx1BWdLawDPAvTFScnXaOoUxu7Duy7TlGWAkdILlYHAZztvemXnX83Gb7iP52wtatluOge
xje8r1xAGXAoGEOQgC4N2TXxWcffd5yIHPDfb7GKz2JbdxLPnPi+GwWa+t0CYQ/QPWf7ujPI8df/
8ThX1kuQ4jR5+W6AjEYEpuRlDvbUP9xICy3LO0hZ1P4E9t7BaYezTEUW1r+d+SeRLkzWGh+uIhbJ
QYT6/Lp7VsbTL6NBHtQAug3vwIeBUgofwV/I1epXYeDiUlw5UeE2pVc8jTAgFygmH20apahCNacg
jG+5Z+MgMk0Cr79WDX9qGapoIVnuUJg2fhjyIp2SRqSEruzgJtHl7Wqq/8L6P7nliZ1brgAnVgWo
ZDMI+vRWHqLg2skjGv/g9ZUTxPPMs/zZK5Fev36ttV7kbdGIuNlH6wR3b0feLygD5xnLIgAaIqpU
adaQ7yKzBCRNM+HJm4WAPeKGMUfbmd2xGP4XR2bLBT+9DhXihBsOoLQgdLm4VwR9S/ijaDHYFPH0
51m9OMSdsRW1quuqaDYQXnq0rikKHiVaMQXr6ijSa2iwCCJPPhnCYPq4VFElLOLfg3ir5UQS5l9G
k5mXHtKn4KQ6rv6iCC3+AYOpa9XDaZUGHsRI4+f+8VUVcqcMCfoJxmQ3hjccRncmrS4Qny5JGW0E
95sh2QKP2xoVE/0Bx1zGpMXVbeee+gokh8njQsz4Aq1CpcbuRLw4IPYXBylHsABC4cMal7l3ZGPV
oWKbQlgdZ7ZqUaWfkJZmQjqp7kc1CoD8JD76jrvmaTgz8PctL4yferFjTPzoJHF+Y/IzIiMV9DrJ
WoXFmEqOv+J4vDS65OmJKmYqUSLo6G+y4twyp+rUvPjHg93KbqUGqKizD7SaRYXEAMLCiJ+z2QY/
oEbO6KC33XfKW1xIH68pZmdFCLur4e31ZlplqKtHycxjp+gdzxWUwWgtfV0LhxRWI57iLXYnCegu
6e2Tk9i3Hui6mpBUcO2snsfGxCzmIArF+j7Qt4mWIJi18OKd+s83KxtJCwew0poFjmZU9eBuM8l1
qTvND1jscYgN8Yw2+Imjj1D9Ege9U4RgwOv6Z5Ll5mnsNnmnnW+14BV4wx9TDx+ESMyHt/iSm945
qU9mYFFmXmwg4IvhuQq8/LXt6uc9KrmsV2txPPtBfN+b1SEM5ZgNtPKkU35UyCxA3uLPoBM+hmgQ
jpc3cLo5JMyz8LL9Q4F0U/hv8Fvpk0AjVkWMX6+qo2LJecX9N8vkA20lkqRoUqTUy9g6kvLqM9d8
ylUzswEqIhRbiFmPm4xonsUQth072WIBDb3MDr8ELN1VZpewt9t0lLgC1hZyTg/iCTV1GCLJ0J71
sspuu17IJR7BWi3U1DbK95ksVfCnC/V6n+Vi2xdZd2R7kIMYobm2xyEnWNRZMwshEax8t6EI7v6e
T6HzrLbAZEQNbfzNUqIl43hHo4jN4oYRc49Z2zHreB3+yoM08y1YfFUMUOeJX0lwD3jg3cDQ1mIt
imO5qu/o31rc4Xi7IeNLQD+pQt2UunPLMmOUDQ58jcNQ+oBQDgddfmp1dlLQbN3Pa/y+6ky/vk/S
hn8FZmYl9h6Yv4R9sYGA/zEnJKzmr6RHyQKSvf9TPRuq+X7ZvMc+Qi6s4BJLZcCDtRKNEEJ/QRfk
jBnTO7cqZHHJ97Z8BF859RubQNdY4ciGiUPq51iGXHLRpHMSKpj7bT00ah28IChHN0lAGn0dkOkP
E8sLGZPuNVr6IBspXkzLavx9zJKgJyDs/1jQJEnJn1dMzvucQYsj77lutsU8ENUOZSbMfxUZ53mv
kzUafxVg9rtVxETD5ThpXMCCDLg5qyeTYAFdF6AqUGFiolOg3bByGOPEyRP7273kAWqiRz/x2kKw
opFTRhz9k0VQ/+U2Uo9yGyu2daraYKZY2EDsaBoAfa3NVjQVRtrUG60j91m0BAVCqUib1/Ud1C+j
sqmtsiou9avsVOEZzrefq/XuHwOPPT3ZGhrEkZu2her4r1Zr4YQ5U6+kJ40OLdtbXsPIwVyU2e6O
Irc/vZPO8UINBDPjn1YkIjjwdZNpTYImW7taQZc/elqsjAK3F3/6CuUJnYLtkINj/umb+Z88xRD/
yYPMHNfYYaP4WoZe7bfiRYYnqgB3LkMii+NZI8SdFcW5MyvLoiLRUKgNJwN7B0rJrDQaQvy+Gzy2
0I+ja0Jr1SROa/Djs3lV9lCnJKcSLvdeHrPfCZglVD5U8pRmvCDxIgMjq0yVhp9MGuVRzzhLiEYQ
xF6dUeO/NH76sfDjEUGenQNpXzNrTjj+I75/ZWmgu8FwjL/3G+Hw/Y7sVZkWK1APX0duUcFRSAbu
dXtmwR0qDj6go38s8CnnCXHZxzD2daPhxpRw57sbUzM/D9JcRRSi9S2zPZJnKoljK3X2SiDXaf/S
BTbNr9H322wVb9MndBLAMZcXxfDXTG82P6hZvlFKTdz5oW7sk9/yhjvMoUVxkSg/dWYderddLou0
dJzqBQa2wHd2IatQYULO3rQdFyLDy/nGQlbn+QpDD/Yp83UQy8lU54PBPUIzf9QMSDImtrxDF38W
6bUyWw1fhzoSeCTKqVbTtaJHcb2UuAa7x8SsTgwwRL0+l1VQd+0D/+t508RdJYZpyqqR4hvSwyOF
acS5gN2US1ln/WuXN2Gf+QrXBIf84IK7krlAEKoWeDfZi5frUD0lgj4/qtWXF7qG9thPw7tP/O5d
PWLNPaNXQQY9UTSvxUDp306Gv7YIXaquA/Qyk5E5LktH39qiJ2J/jvjoXeuj7lTNql2vNTcjIdQq
og+hkAGx2WjAQ/Y/mD3ndyDVG40Ig+xZuklWnHHew+zYd6JbqDUqHnfrqVmXBO/rBEu7uyEhyRJs
SNRFin1XRbITVl0VINJqnyjwM+ECXSs701Bo9MYDAAlR0py0OIUDK4BSpy8m9WxS421RdnsKvE5P
RAKpG5t2G/xr5PbEaAuBAn5gqtK6c1FQRNXPgYgVV+SGnJPPYKJ7KSpQcgLjEhgePkf9J7QevDY/
hfuMD0BMh1oKtrIc/lyNqQAFe2Si17v15UFFRHsXF0NHRWUH5ITX3jMETwOpBKdhFuF0XkwX/09x
aoP1yHfR+nDRgdxdhc7AMnvbcG8YAFUetVc2ctXwlrfgr6MerEnNsMEx7QaU6qokq7w9lmAKHyYW
2E1llVGi3iTQaKRWv7zOoze4s3EmAyc7ZKyynD0tG7Wvm6Y+V9Ip3tBzLKZIa8BoJGULte30LPcC
97m6tGvIcPvcjP2kDoFMRqEfgzoUonOw6KrZ4tYUqzq7BfLRJJ2yc9xizJnomvEhKITglksoGgC9
Yd3O9Ausdd+u0KPLhWsjtzSyrE7JrLsMYRMLArLzbhEzfH54mdeqPxG3PNcz7+0Kj8QwIgHVowEL
do2zb5KBBas1bEBUxpV2Hjk4X66DT6mVTqCQCHiCvaMTp3Wp3VhD1F5xYzri2kwCs00DwCD8sxwP
EMxUQNw5IKDXqq4pR01RVDb7Q6vdMoCBzNmxXtTuljVavxH7lpAfwYHSvcLsDgMBiv9WcVqlhSYa
GlAxqaomz9dDXVPmhKEXSy+O1nPOonNu+bvAQLi5lt8nCCDHMNwTakCjwgEevgF+G+9AH9LT4mt8
waNEzd5Eh/1oddhE3lhaqf0iRx0I8CXT3wflF0mHJqApwc5zWcntAcDzmHJwxa9VqdweZavLfQXi
cpgR1D/73shwbIIeF/4H1ljkQbFU2dIHNSFJySpiS7kOl3eI0+C6sQbPq5f+QVTM/FHZGjG4+lpO
H2gzeyT8oJpAZfGQuyJO7BciG8R6+cmHb0TAM/jheOCIfRFqNXi94NcWgLursDDY4zWfKqQbWdOi
1lw11mdzFAnGz0SK/yFAiGBF5uQYp167fJ4RNgghrGdFlaEgh/N0VqbuHQNBy8YGRxGkHsy+RLrE
UllNY402psi2ZyD7oeGOn38ewDpRepsLCjIkLlx2/zHko078xQPbf5xpj6pw+FbZy0inkToWM5jE
+wwW8oiOhgsKKsONEU8hlq2zffEryIFjxg1ewmApQGBmD35vpRyQYu5HFoZS2kDLTA0/FjgprKHr
HNj6aC3T5CrBtL9ZaTkfu/13rKiOgxq+1kvxkuk+V+J0/yQP3Ok2u1YQ8JukB/wxfUCFNBHOG+zm
3kYLzkJk27Nc/ricriqIAjGrnQgPKiKiBjkVPcogOtCnW0jJFe0KlAG9Wee0HeChzhSE9JbZCHHo
Fk7MhtveiRTBePwNVTLkJyw3u2/e4iF5af3zi2Ar1TNcZwKewgIzo+UkTnbzOw6GyyapURwUqdK8
hsworoqMIiesJ460yjvSuvAnBNZ1rEEsNZWtTi2OI0mbqKE8I18sMtsKkeAbk9NvK7LiGEWCqyHu
bygXaYLQ0W8ADXNRfzw+8Y/R4zOkNi9zEMFGL4eXazAogm6mdDcxChIH2cZq62HnSsaFtzbTs8bX
iaq8lKWm7vrN9nL/XU85U7fJauRSOL2RY4m8qGzrF4hjVPIV3ZGR93yRaMlTiQnFznmOxA6cGDAu
FkamwnOBkFF6Zp8PmycSEq0EHyrhiBNkidF0RktHC1Y6Un/oeU5OVrhuJgHjrlF1m3iHtq+Pz3c1
Sk0hcAtg8tqwS166c8NRqr801aXeaF9L1n4M8y0r8cp2OhAbl4EMbVnkcrUTxvp7t5U8pr8ZP/qM
L8auIrP21ijqRnuApXHIEdisYQhSB7Z/Sq72N18qDQ5UnAzbY09APt9IXWaNvVZ2ytusO6r9AUBP
klK9D+trdd98glKB2REhjV0AQwwqXpiOJoAzJKE1z88adYxyhPLsjsRJ2VntGujoPNI5v6iqyTgR
hjjRmBZ4uXiaK99mVzGZGjSVRDhY0MfgsUFDfz0V2Zq3bsLo6HbC/SzMK0QxVGwV93COCASVAxZz
uxw0l8eoTksUa9JqrJaqPiGZVPZp6vYBACIx1ZEuvTch1EOPYr26ir7P+YAQPAPTUbsH+bne8X4L
Jj5C4MJc7gBkYGRvlXlCdgxZXnXB51oEZUyXj8qAXKu6/M/ZVSes1eI1IgFC53UdPH94biE1fd9r
5XybDmej7BG9/7tmra6rKZhvZD3TtNY1te8YNZJq30WnePhrU1NqgdDq8YVRhkM6smOoqF3AgAsF
/UYcR7FLFz8rBdGFsvjqOky6wvF4oFppm1O2GP4XJxtSgHhJSSkvUYZ50aybrkGRjl7RL9qQ6Yka
pVbjSNY5W803DOz3qKFzIhT4vy5kT7MKNvw1YzXJbqUSFJHJL43i3oMet/G8Xj5V5Jw3J2Vc1XhF
J4OovwQI3UKz0CgJDmvJk/1zgCxIGbxNbtQ4oy/vUZIFhAQ3/XtmsQhdkR45MvANMh9aO9KgiPR5
sySP62SxQVBT3hmTyhLPuiV7FkkIt9nz/hXNYlCVVgGK3onSqk66QQVmSuuIBp8GNgW6w10722t1
JZb+FffKktHcttOzVg/5XLLkLfbsPsOXL12WAeeSS2gh3yeZ327CyfIvfSaCUCgj0glRcYkDdxZS
4iMxC+h0kx8FxjuluLejZzt5pahG+o53h9o7j1YFaIvhX0+O6oVSFsgFxzTVZcxX+cxXr2SVmxM4
u126h06NpHNKASFgxIbwHBPSrA9Jk9KZMXiAB4iHZMZgRDQs6c82C1kJpKZ93eSgrurGq7Mf+Gre
V/P/RjCfQnYdTNa15GJG4te+7LTHF+WcpjiI1kUHu6khyfM6RywfF8GsOkVFPfRT+0gBScxgVt6g
5KKchqp/6fqQ4zpaVWlGeDOGhpa6Qp28VBUj8DGzBFwQ5swwbqkcj7ry+242f6EuKKyEzFPN8z81
W6a2LmMJfpWWeZMnJd652gMA/lXQXRUXV7eEEvS+wz2IOG0a3K5Xn+ZLi2J9Pcq3SeBDM4RT0FC9
39QguA8/FOIpdYiRJkiBV0FO8C3PpVg5SNhloPrEyxkemav8teGOSTN0A9NAZ5QmLXpc5qTynN5x
4mdcyy/QrOvMxSyPirMwpWc37cmWNUNphUmM4igy7wswHM3Oq30hQqyhYgFOlVUPakucjXm+i7of
txms9nWSLBYi2cGEtG+nhfuOSPEZU1bvFHH64jPX1MEnG/8xZgwIv/7G47nd2cEfE5AraDT8wm4N
JUylnIghSZlfw+kG64XU0ahQFLtIlgp7sZJQKrf2Hlu3U9gu7kPGtUEQYBbjoYal8cpWr+IhlHKy
FCJpRQToehzIz27g4fmyRGeQZBOUsI1gukxllU1LNtA9eQI6gf7ZobaLJVDKGwsrHgKg06viWuxA
UsN+1X/M9O/SFhJhjxGbUkMBbempkY76JbUsWw2N5otIIcxvHprbhfzvxtVi3LZLalphlDLmwrR4
x/AtlKEvzEujPmF2gqT7ZhUVx/TDoO9s6Fi/HxQxtPZVxwcS2i/71aJuSzqI4oDfN4s2ORS6ZHlk
wPi02FUEOgKsyT//Uf+kqElOtEx9PhB6sZTGgwA/SeEKjJiVfKhTbA4EbLSt8znPEwV8QJ6f4Q2V
Uhp1OQB2xKaRK8jQrO/YixfEIyPjAPTYLFaNUDEUygrtDvgx5UM7Bw4JuL7WxV7SKEgDaNitE5J8
KCerSjfJVykPKqRhbC4CaFcvZQmSuZ8i3Axs+vDqC9uOdOgbQkZv9vPte9VC/GN/mJOYNs00g8Iq
gEEIcsjtEOqRBtohYaRDJYIvn6bl/WB5hwI/SCms1W8eiaXj9pdp72VVc0RhzcFJ39JyWNzu0j3M
uL+PFvZFQ1/ixWEQHIF/OxHS3RxFidMRmb7i7LLhtHDFXT8WtffC72H9lHHrRT+Q7jPqjYZthxN8
AkXrF6q4OHemxtEf63ZZrCCZLtiNrtZ5t8/3yOzDhami1Kzt5PjrEKppx2vdx0nZWAC8WqhIi6qz
Wj4nTNemYaY0upKRmTRI1mkjuFzTqOgLpVwX9b/ExNcm+UE1GaI3VbN35P+HaRT9ybFE/4bRGaNf
L+tGH3hh63ARlgGLfYPnh4Ik8F+Lrr6BZj1LHQ/frp/yHYOJABLfjCWH5duDxeml+ryJYfR3K04y
R+ZZqVx7YS2oC1EhuV8FmM0FgsIPXUsck/P9LQ2P97WRNfggoSQPg6dJ4slurzVfjsa9a29N9wHN
IK7XExm9dT0+RfmcJ+TLPOHblEY79azJJrNfHk2RoYWHTsMIdsAMOtAWBpW9X3ZmX+fbPsCwnJMy
rdLLI6B6duqjNjJqhUk9DgP33Jxaw9mSsH1xnlW0yS/sa95UvVlRhlU+tRzh3Ft8dB1vBQccNtdj
NkdRGoP53mXkzdJAT8wbwoC69guHOc3xRK8lxAFrjQ2jzl+W971gTmJIvAnq8WdYNy1KSghNVnYe
fKWl+PGP+9g0MiXv7UepQYsKYa8Hqe8rFVPCt6wXLrmQ/jvGiRqHO4k6240Ywi1vQKlwOU7ewV5T
I/T4nyiAD7PS8aiTumVKNRd+fZvtloCq0HtXBAarF3QN+UafbIIkReYXnow/WhF39+bt9SkJfmHP
6UzisAhI61fSzQGu1Wlzy48ObXvv/rw7cnEUp0niXKi+xGGER5B8aTvBm0/0SjYaYAneA+vxSPcv
wi6RP37HN3XaGSTZ/25VBhsUmJM/fYsWvNME0chEIzY3D9bqb6gBlyvKBkgK39UBlBzFrf9eZKE5
NqQj1X38KNYWuMpw8Dw+sJoF+5fyBE0d2rCCb9kBmNt2qsqgj6W8qDwzGZ+mnyoElmg3Z2MqgErD
CIydPmrMxUZ/W/h59ZYrb3y1ZeTI2DOrNS1n40MVM3TQWXQIvzvybP6EhgBe2mOR9ltKaRmp4l1O
cqr7w5+I+8R9/EUXSCwhkaXHTyCW5I6ycyps4b5EYOcjmVWOhIfuUQ1wBiTh4MhI3cfALC85ZMCw
Kwo5MseOuXNihg8oSNNABqFB5uZlJqvOEFhFdehRhOUSBZJ73rxpH5dR/kCK8YRHXWw6QooQzfsT
RjnDqxx7nkAZGlnuk38+GysjEeTWX9STgwOfYE2nNQl47zX7k+UVxUOiKifzodzZx/W6mEy2Xgsx
gIPA2iGKf5DskddZD2wqXZ0ielLOgrb1/D7QhesVfuTqMDwWdzXeOpwM8PM5w+EiWtYCCoKNOqCf
INdqX2RIQZBduPimjzI0vms15krWmdj1cr3YHKn70tdvPtHIDt1vt8+wWG4gZXbkgcwynQ3E4GUv
SQypNXKikBP3zjwjXgjI6K19fJPCwuV3p1xUlN9nOU+0jxql2KzfgEUbnKyeQlIi+YuRh0BeGCCn
IqIVbFSmX1eo5s7u26s7t+udW+cgBc8lZFkfrfpLtwNpP+SrlSbh4xXrvW4mZDhV53ryDz7FjIeB
b56fwJgBONhlYYpUkhJpk4dhil+S8XCrJbDRnUZlOBZprFWF824l9BUl/tA1sVMKPu5lxmZ3+kLm
1jTRnnnQkNmlug2VOQhrE/2IvSGR3CjNuwH7PUXLMsxOc1+EF6DKZJpuwkQ92ZRTjhhh13rGQA1V
p8EUGTqS1VSJDLkGXocIZPolxa1vpJ8okgH3ix3rNCyBbhH05g3/t+Bd0e/rCZXGvL9woMUuFdS+
aAhl3BCk7sdmPqh5UckX2wiO0BQEOknBcjOLnulBAY30YIm+SWe9kWlgKNnFMQIs5Gh+BL6yCKaY
sVKYh/hoZaWRQhgiw5R2Z1ygklZsikj/DbrpwLB0lOwA023oDkoyupowxCpCgnvhsbaGFTGXwmPH
WkUziIQ2axe7RAU7cQDmGnElgt7NIBF1anuIoJfa2WHIKDI0sCbFvcoaPrnzPZbeADfh8Snb1EdU
z2PfSsPWgj4l1dzO3ulxTeJKWtvO/ME0LfJy55wagrjsdZLK8TgIevWczvItn36Uk6w7j7yPVtG8
CdtzKvm9jcdzQZ5v0SdFHKBx3MYiKJvlyBFq8nrvG44R2ryM+lywpG1A43U8qEEo48kWQv0M9HJE
nEOe4IxL1ydgMKf+R7/0zbwVu6pCx4JO8PFLI+x6XXnvFB1Rk+IiS0X7TyVhFIHa4tUbDnHrrShZ
RPsJhLxnFi8yoxEPoHmZa6k6tQq6qr2cBTqcvWfLLsOxS9ckLNPmhZqbL0kTVq3rwLeU+ernRCNc
Ne0U2IpWn6anwlpdEjINfZ0k4Rs9gc9BFc3m3mQ+93Zj2x8rftgnb/M0dFAr+YcmMcmr6JFgfxqr
er8iHAv3IrTHo4gpJgJdmmcnFDysfxDIOWa678XRNdcbiDuBMBexcNLtoOcQ1MkN1HFEFPOoGiXZ
tPatd2/kf+YlWf+jpuMkAiz62C8cZCPtZu9yZ+KFVISZX/o7XrIJY17E1yyMVZWSLi0BWFyntBVf
lFB/rUT95YOvTey+BrBBzESdFLhcLFt5PVJM3lxUfoqxmrLERSt52014/JnoNdJhwSgvSS3QwgwM
k4/DY8h9ClYjrxc2J2PJZvU0MZsh7q8Llt/m1Onfgg+cBc18oIi7lOK0VvIdOq4gNE2bOn8GT80x
XX7C+r5dCrOTcDZ9LHB3cwpT6TFtDqnV6ic48CYHODTdCar6138kayDSNJo6POQ8fmdUfQ53DjDt
FTWbwwhMxQRApeSpbxsNXmcHZHDoyD6MmzC2ZorrRJ3hTe7y1WvqrVwDSqSOonuvsMNkMzSokt5Y
7t1G7CO8kGqXVuD3sKEfjsp7WuhyTnmGhn56Dp9P4L/i0Ck60t64o+VmOCF4XyxJfvz27DXXoa0p
GyE09VL4kQY9eJT27GJX7phMffaQyxXU0X9Fz/BTirwgD19SMPL8xbtcTM/z0DzxI08Gjt2FIVyl
/fkJen8o+Pn3SswQXO2wtst1cKj5CnGtjXlPny1IqF3QFfKV5QdRG0w/R5cT301ACz6R98Ea4qM0
fHIoO/3WxiAqOHHGmLVjMCq6FpfX6UkdosfMRfJkhS8Xpo8SNsuyqCLOpnP1uOpVy6nHdAN753mT
SvUnykuGP3fZX0BBRTQ31g+Xh/M8o7UfjmPXrMEVGpWThhllGy3tXLlgAKmhkInTUfGSCo22tDR4
J13+hVjNJYuj5lBk+Q8rYLGVurs+aW5yxgWBrrcM8DQexyxT+5pN8esNF0TM3uDdNSCNOWrGErEl
WWXsynPoomFryZKMr4BJwWrj3V5SKpSqq8qABHAPy1zgCCH3iuSEhllJQn+ughF5vGrlsSTUQDqm
0+Tek4iWyii2FUAvqrGEqXGCB6oAjpUk9qEmr04NyZuUTSIJ+Flk2QJSu8e3Ol3h04VeDZomF/jQ
4HTvtPZRDa3TnKgVpqkaVLQMcSek8MbwbKE+VWVQTacxWNxCycbm9hWwmSyj18tJ58PxORl1a007
YGqXLW6k2zwscElCIwbuE7XML6YEtaEzLFS3vz6BoYcRLTPHRHGQvk8ym7AomkTyHgb/ATqkjygA
EzrdaZyfEbG9ABIGVKm/8pdmnRsFe9bFDE0yj+ndoAsXw+f3HUTL21ldLG/omb4wDF8OGE+Y3bNV
YzLi7oPQp4w2opzqcSOVrW12gRNH3/wMWAhdBLGOqIjWYSwVuURE6MnCWCJH9qG+E314x2bKjg5Q
YtueDPgt+TUrGDZXd5lBJIG3zjs2/JqYnqYPYMy3/yhsfWttsQ6DDT07EbpMH1fOlWxdwAhsQWZt
FV7UN3+STsp7JUV/JnL2MDeSMqO85gFLSzNcEiFpIJ+6lyvIMPhKyuzUs9D+Dn6JzIx6fVVozVuy
3alUGg9q6ZeP4fOc+sXLa25d5nqB35z4EZJoJug0tGX3fF0/JbDu/ZxtQ/z2rAM4dU6jkNeFohLM
9+DoeOsrSU7kUc9UDHeGAqkNnWy+M/72vyB0ycSk7p448yixlYzQTq0SFhJuMhdYmO+sE1W8ltmo
Zu5EzuOEUEcf4/H6RygphwjmmXKsniVhyxOI/X/KItOntxlMLSu0SsNnNHPo7I/wlX+rUXcQvuAB
2hMAzqMNXNjuYfPXHhU15CEf8BaRxU/B5ihEYDFY76DkKKFg5pkfCf9bc3sdQ0IxBZh/3BJJAPtN
k8qCYAL0SyaVforPilczl5JXfFh8veZlX6pqfSTp3/BE9moViOeJtmi4nHKxyY3KeF5yS4aJneXQ
jbnXVXjD7NllooKBpBCN+fqCl1+1P7OhoFhVj/1MTqwnYHX74gP4SCQ83TuC3D+gMtxW6+1RSRd2
HVmtn0NT0hZR+Kq3It+gilAgzo4F0Y8gwVDqxrOrXV1G2y8EWjXuYkoBE3SHxyZtCne4P8n/7jBK
zfPxk7QR/BfmE9wjSY9qeqg1bbhqiDQtZra+JsLlv03WSlGayOpgddqM/Jj/jLlPCfhn+GIxL59C
Qq3GXskwK+0iOVC4JeLUJM5exyIiFXnIwt3XyvyDTy+ZBhJiG7x4R8eUj8MZ0Ne8HBc6mf+YCMWQ
Ys+XmFZWRb8H/Weyys2Y4xXQMeWaYkzvTo6fWoBe8NRhO2ZmaWvSUKV9dj1bQRrnnNrcUs7IAPNk
7BI5wu523X6c/ZAPPEh7q6wp+raKKKGzUUpxkuFZMVjiOS3TyRuS457nFGGD6enIEwkKFZ6CmyJB
TPAEiOz7D9TsSNNfieXEqXk+W5OpswWsJf5eSwXTVW+irD/iRnTDOckATX8sEYy+gvd9ziF3+I2i
nAc4t4d3MDMxLKf4C4Rj0VEa+0MdupoeCM47fP+dDHgadg4C4LBuVik873rUeXuVYsAwM1DllThQ
WoalQHRLrzN4xRMd+6iNtgBhL8H3HDJXwddDmSLE5mGxfsh48/PFDglwjjq/dOP4/abOqLveuIpA
zvF033j//C5i/Rr/W2PrxATpxVnhaUI3Ek/JR4YN4/uddz9qENevmaLWw99tMmhWv3pJx1nm7hvD
0myoBWMThHskynowQVySqIz1c8Fnl1Sn6VQaND0s9UNVAPbcmVi3+m7Av1mEFw47SKBWtzcE8dkO
ukFso7p+ZKNzfbwhtm4OChIYgytugtgWyDIXuJnT1CnETivXY8ZFQs4CI+wv5HLp/2h6HTo+i3dV
+o5CLhvPNDRZpwooWNBfoBzJpnkdYc6l6mPQiZleiCnqO5pcUFD/BQDTZn/gyiXzWgLBDHWgHucd
x38dxoF/tOJUzqtj68fIU6HJP3tqPpPY4dgUmTq/8XDyKPL8dua9R95rQac1EQa8qWpoNlhVXe8V
rcCCApFBApe68Ax09rVjOxr9izXgMBSXgrzN0l6IAfuTedwTFuuBHTjcc47S+Nldfg8WelyZ2tWM
bSoIjrMDwYBaHdzePl1IMYJTf8LixFrHtWFW9Ll6gVDXZauA13kzFquNMso9Kk+jsQnqacaFJ5ZG
K6sIM4y77S+FQe+1/ARVe/0Cm2jwqk1AN3qjl0WCAgm1qG7o7rkoU7KSBinPTVdyLJtygS+3n9yo
veRonpoUUc7MbH3617f9pYuoO9TtbHbqb1MB8piNOjl0YXIKcyFUN7yt0ZxoRzM8GiJrDgmKH7cz
Y9yBXdvasqqaZtGnMYb8RorWRHCgN8FhqXlNjiY2DciVinjXFpsZ9lDB4lFF7CwlSqutxlAOW+F4
bRUYSKw6SpEM4oMuVjQKZkFoVsn/sht88PlTLck9m9QMZj2TJpKnyXygUfpv1M7lekCHtfFfnYVY
ZWH1I++vaImQJmRoNFzE0gK+0cfPxnr6n3NIpVQpFPVsz9/cd8kKtuHaE6UryJVZj+C8xyqSajoW
pqoGnEP6YnvTBeTpk0ygWy7WBjYXoWItz0s9kg65T205QKoCC2fbSXnWjQk04Uba8rtZn04ufDnz
wCj2b15N6mSpAb2uaKCJaWtzAjyDE6aCn2GgBhKGD6lsvFB9zxJBMP5aYZBJd6At9sE8Oubx2mOj
Ij3UoSuB01Wo0G5wPZ/278U/JDkpK2wyucuRdc6oDCa8ETawsWHGAFKvvQm+cQw9J5g9uAQ6DcqJ
mRH8XQ3UIAM8apZWINSt3N4Yuff6B2HTij9WyXrqWP4m/cI+AieP/dNcie2hwfy2jruDzbOPS8GD
eNFZ+ROn2Bjr8SDC0/E7CTF2MXCdnjKG8kB9Z/UTS2StS8OqSKAjd7xg7LmJhLqYWZW2FlMCuJZ/
Ux/pWKmygdeJfzREnWGL+syLLtKBhsOPDer8r3T6ajfkqgevBQHyX0STW9bSDfobO3YBzG/m76dx
QqD9j9nfHH+lQB3nlM5gw5kEW8Noj2owCh1GjYTs4ajkAYwkQ2iyw9bE2UDiiUrON0mUBOkAgzRb
mMwqwyC+TxAgOrlTjOfJb5lyIP2Gj9MwJO8UfygvpJr423Z6MFs0jtM+3mRkdNA8EGSZRaYwU++y
k6yyoN/akLi7UnT7rCge2f2a5cEY/frq/lJnr5ribQbcte3T0ClBIuxC/mynJ7iTK9rw/TP9E3ok
LuLkyhT8jMXidlfuBGEWdtfmS3kjnF9TVD3cWJFRswkEBCbr0vwb2dD286fZDV+AOiFPe57Ppkrn
ooAwemwHt4TTmKr31XEmqLANwXHiJHfD7dnG/Ab2hNm0jJw2B7MzfjgpsdCRgJcLqSh4y4oGOeT7
kkr/6eDLqmV0q5TsNPpFA2b6wd6+dOUYp3ag/eYa0xQzcAvncyi5PzIChZz8tGcz+8VSf1Pot2eJ
YV0UzCzfRzWrwsAkwaD5jrOWUJaedoEB4KP4va3qb4AOOtlF7Tg/bm28iwLuFZ5HMmq8tMJERG1b
OehoYSZjdkWb5k1CLtqd1hukvdGP5WHWDbfT4J1gIPfCQQ5sBnci7ATg9crlaiFAM4DtnpcYQowt
9MaIF3FN3uQwuQIJfKnoT68Vxftr0hMKf9T2H5dv7Cvs43C3XxoDdlvec429dSBP+cLRcAonmZ6k
OEtGVWZiK9okkzFMse/l0DmuztHpixosTyjaXGfc8Ge1UoPIV3w582ksajrKTQQALn7UDYhyG7rZ
mdU6RvfkDkFrE/+IJowH1WO7h9+5IBPjhv+aBuAg1MOJC7eaJoSIkZqQccauIMH4rxl0NU2LWL3N
B5H30oNwaQIGaBSYnNWi/fLLupY7RZp+KnlDmc/Mnk+526zBcoPHErAe8oW8/clK/8sRR84lPyRz
0xF046mJeBMUcTtUYgU+OJUV7asji1xcKhyxN/5cm7Tn28QhjrprS147ffgbK1iY4hFd8lsOzTiA
RVoeXmmg5i08haVdB2W6Cxev11k+As2umTlq1i8PZzfonrHvFah4U+lzRUNTkWLeNaZsn4vbT7jG
ChzTviMMujRFW1bq8tyeKQDbpsIIytm11GaJL1Ft+ZhCg5eYwXT4p3YzWxJe5VyxkGKiKE/zTZqt
MhjvbCxNa1st/BGhU8D7gnLoyjoBZAcos8Fy4skKxVNgiJ9n44GtquBLmz/XUaTUhtevS58v6cXP
ovIbtSl0aZm4QMgMWiVMWgcrINOHH6Dm2SoB+9BisPNhxLJXeGRDs5TCDzhL/Qr/eZjSWlftIcO1
+9BGI4Hp0GIKAKwvJhYqUqzwTMWvlH/iqbHuRntagap6jLXlK49ROJ8bMobZ6IaYoveK+AkZxZPM
fZM6zid7waOU26WVx8/YGoWlGTezqiiiHEAWnR7B/fzdle+XRDBHLzQwHeLSH1NZ2mqiq9wFlI0f
qv3Z+09vK88At+oUYOFRMTaXqhVKUZeknyFQvRaXV1S1p3sAQegw1cBjOsBnum0y45IWfCTCkK6Q
iHJz+CJ6HfxIaDSext0baCgRIz5aijks/1H5PphAh3W0KKzVg5dTO3/9sxomQKwYhRkEmz3+70z3
44ovPQZ0oCedxuDd/adv29uBaDoTYttjlFhxWRl/UjpUHmtlwISUPtZgEqOM3gp8c/Mtn89iGVCI
T5zH3jAZaPWt6LFxXyjivTwh/DGBMbM84WvxHL3l2KbA1IJHbBbdGeDEibFaAC9s2bAZXRDev/Od
2QTts2gotf+PnhGTDTkVJ++Jwwuvrsq6rLkrIaQBIPrZN+TiMOUgbXyHFz/1nDvpYJLxA6ZmG14K
DaAJS99479BkKkKIaoDo1S7zpAYtQQRSBYhZP/LnFoq9MPKnlC36ROSMLJoJZ0I8ts1ZkQFfkW0Q
Xu2z1vVBS0uyk3B231MDXgNsHVmy/yJaA1z1IpmLXZltOzcsJDGpuX9pblCGldfH4PLOuJbzh8FZ
uFikCibAMYZegJ2FWgTnbUVDqh0pnEIBwnSYm77Cqq+Rq13X/ZUVtlqWdzB5hBuzQavSP5Xp82G5
txj7jcGutEzQG5cPP6QIBXziBiSAtr/X13ojIhQKW0fNomhMETXaP19mzTM37/PF8A3urqPpX5E/
7TLVg24NgHwFAweUoE1NsvpbvgxthMQtQUCnLKNcxPlcGjnr0N9FKURFSxDjRItMAX6PaR/gUVqY
mpf+6F+O6bt3PnVLCijiY2VvsdRjl7U48PCbOOS/w8s2PI0qKXzUmLYmoraSpg4rJAV6PUr40YIB
gqbpGcUjH6uYeWpoSnNKXZF2G3nKiVi9wzK68z8w/Z7ogv5XBFqGUGsjLZdBM0Gx8DmGFzeeh/q/
Bw8XOAV9fz2jmLqZ0+jetUFWOXNoeIGG3KG0BfNPzc3BwYvAxqvdHW7zBUS4NZNp/CEBoFmpJLg/
hdgzqvTTI+4WOEhPRYreymacVwiSrsMc3SmYhoC0r+TU5EpwtaXJAHFUQsAQGYSH598yaMSXqhkm
eVgBYXLOBqtTuAe5d980FKebH7pWpH+3yzWPtTcow0g4sJsVNJ0HOI/xdEfVl1clRvwXTQeSMjc1
FE50FGl4eeKcoJWvBwL8fK3lSPFw/0+V0I9Hm7oWNI/dl/8uiY/Rjg4JokBTEzFcFyN2LcIszZaA
0WnXSz7Nzi3oh7dVANZ2k3Nm4TrtF8kcciBHwCqnsYiSZSPHrAW5mavz5f+8B9HX7YhZbCaPDyvK
srGUFm+57KEjLd37mS6gFGGFbbY00pK+6xEBf/jXkcPbCdv9S4cWYZpVyM1B/GRoh6N0aSbLJLU/
bfg5VdIt+r3JxezIBirAZeNU94zkp5duWQm5fkmDpm5eKq9y39fzFKCZoPwiyYmZ54VKVo05b02V
ouax9s+PqejNJniJza/gLc3RSRiC3VYOYMHgM7OhRvuqX3+20f8AnmSA0iuSlzmwu4vCsE9Ye5kv
lAK3vP24rbtcD7609K5Q/o1dNi6ZqSpzmtnc+KnbT19aSkCvwhjhNtaTL+xVnnfDTdaE7QEJyYLi
8orkqm0fMO9EJt1QTQUnKMJD0bH7QWZZdt3u+H1m0PDD8HMRH/G0WjACTKta1Pqri1Zl3iW7rDyV
5U3LHkTkpEJGb2EZA6n5z2y6tPEbaNoRuOOOmUcXMbFMsDO3j09bBkcAT6uU7RA/PI/geGZRSHSs
LmrymBvq7Pej1GGRnpHINUa3YKJdd1JdfdsUzrzTZbUWd3tlBPXvgufCQzxaOL3dYF+L0x9rhgAs
9KwiQmyVfxV40QR1eCNPmm5V4w9tGBa0Rviu7cU30Q8Yn1vBfQHhkxOiiadbRfiJ4YJrdZnpiyFi
1/bZsGaR+xAxRXNLsZ5otrqeQJTzqnRHR2gI2khBZ/yogHG2geTVPFJBcTYrZ9JGHej4GrDcOFRG
U2h/ReMT+LnMgF0q8/zubkwYM312R1bEwsXBzzamUBjvcKmNHL2W/Y+t26mX1Qb56gKNngrh7Vvu
eubPYiQDKaFvaSJst8kG4Ps9sjiw5CSH8YcR9Gcb8Zmzx9m5ZsXS6ooLS5F3bl3nOgdCd4lfpdNJ
OfBa9hvNcB6OVQzrbBpAoVSbqbninIaMXumCt5mxfqU+GHcQiDRadwnjlE3Hsl6TFJ0aPeEsju3A
orW0gUhRy/eBLTEcLDViZkzN5fV6jBWPdFZRQCNSu5LX/UPPfoJwPV179yLsB0WoLiH9I8IabjAN
oBQQl9i+1MR+N9mLs7UyqQW5Uw+JGuBDP8ambByHUO5qJFbdaScD2Por3/1Qppf5KJ/nfzOxJTev
ec0GQ/urTewYNIqou6KiaInfWEVDDKKHZh3q6aUZphAx1qizskppX/cNn+dRR5pXfRkKPeJ8wWYY
rEdsjp8XT8CBb04jLbifYlJDN1UXxHFJtxye6ppNYvQLxJN6Y9EAetnygGQNPH14gHf2busCcUKF
ChColRg4JC+3SvraA8K7pmQnqtZnHu3OhRS6IctiHDK02I1PJRCRW2bseYXbgwwekoMinjVNAevF
CgumOdG5RB3mfwcvMZTT/NNQTh2bW1zGvAynSiWdWr0ILhF8KwynGpt5cITUXmbeCTNMrxEy7gr5
bA+7ke8bYvnCMcCZmNjOZCCqL4X1zAP8/o3+JbHbAskUrelzwqxMYdB4DJXnxfL8zDYllgWjg9cp
7Ay8j4FE3s9Qvz+Y5BOqgTv/WwbflFkUtFyGO63UmmT9+ROsobcU6Deyd4qSwOFcOTmoD6orHFxd
PfCT6VShuNshAsJTfWJPkz3ApJEUR2u2IUlfz5l73rGg4bgWtXblsiuSAOIOaShIFb99S8CrUp/E
+vjdTxyVFouclk7BdlSnEl0uau3RH6EuiDBBk0aW2jSd8+WnhEsJ3EKbFfXRHm0qb+po7xhUWMpX
atheW6rKoUVIg8UJM2HJ9y3Dq0mg9A/6iUvM9d+Mc1hEzTWNR5ZE8tFnT/YzIK8Gt15oV6F76aq3
udk+GRlzyYvCSUU1xElr5FXYYQf2Otl890B97XunjO0N1bdlhZJc4PG54pprRPCYJ31bm1gSJlqR
dPHVFJpQr635GzdMqbBKjn5CqysWsbwHOtjkh4+1LFm34SW+DHEqYb4RR27R/XVxvwv+UYiaG0DC
Yvzn3ww8MvJj1rS8f5o4mlM8RPGcwHk23olvhleUwjw3r6611kj/E6ghbV2hoco4LxW4BRo1teur
lNOu8TILn8zWAZTtmhxCz57n1WKTw25qmJg51gIek9nyn/SYodiVLNouOBcgAo8o7rNdlwAWFaXA
ZxKEQSe7t5kKG6pW5EH9569iSla8Z1g0A2mmUShtt/3sZE39tg9OQd134n+RsYgwPK1FwPjVBrFo
mJgpoSe0AD/NM5esOiN4lC1JyXfPEVQ9qFfR0MQmtysg4z5H2sO9lpmNSIuFnrWLJ2o8HaWcIbye
vt6nnN7O/HgZvFLz2wD8q8Fn39UfqdnKkY0D1H2Pq80BvUHlvC8oRuEtv3JP2R6oqIP9kObSwlfP
ZeoXOOeEd81JRrMbrcBW8xbLZS6ZK2tsbOCpkeoG8c7JiZBoY512vo5W+f2y9TfMwe6jkZjrcCf9
dMLyYAp8nx0n9EPPnqF+1OREgzyEyEOlHcWFuSECVQs+lSt7dxGuOLo/6BtzXvt9nNXVYFRBoqVl
5LrZS3INElvTpNkgovJJEq67RFU0NKQGF0IU+eZFP05URjuMmhNTAdTaDLjiJwhnlDKPHlzTYxSM
v36NBXFkvjGROCmbC3P3+v+JKWUc2EgcjSYbajPbw6TNMqItRmJd8bFoaS1EsRw1748AK58tRuen
02EOVG0FeieEKrFTNkaVfkTexk6TSpWVv/wk3bGC6cO7s1JS/LBMjOBIeb9DEWRsyveNcZ6i2eKE
gRuGg192WwbSBanS7/RmT8NTmHL9pyCSl40seFVucDqerx+xu0d55so787PCTZ8eHeisvBHuorXR
joFTHAqZ5GDA0nvKSP+Sbc2Zsl6WjH7DATYlneHuYGDnoi3ll1w88acTiDfaupz89iuwhDIAjaEV
QIVpY5bbInATJb1TC1IMulO3UPV6CNciS3O4DW/KQ7nwa/N/1pAT3TofLtoy+Zyps6CO6EJP3U+U
zjAVopI4Uq045IJOZtxs0RxDEE46kzOli1OE7mTEqOMU/PHHUPwzjNxoMU9OjmZP2aPI5L19o/WL
8dswLkU+NK7GFhzttHHrBJhpp8PHBtMNHUWB8F6F0ooh3Abf1huYVQGjutxr4daVbougNQ2DMoYs
sECugJscFuwrBPZpi7Z2sId9h52k/BVNVht7Ec4mavgZ1fH3Of40gH6hjYazAi/K6601oFKN0jgI
re3kUbWlc4IXf5YShpRJZRXYgHkZvoWSVl9BtCmpymlWo/0JKm8Q4T5eVY7Kf4cIGuH6tvGSOuUO
lbRVTSgOiweCujjBO4Ncz+tDCxrItPtMpnKXVh6ggCQ1hpOKcqP96VoBvuEjuD8b+BhuDrTLuT82
aWgN7A/f8I/4vwJCA6dJj/97rCoSVwIbhnBwONVm0gGAyflVKxnIEH9rglrUfv2+8JWekVQ82X+t
oWkebz7J6tE36a7g193vWw6ztDWBd3aSvWuKhnNlPjwTo4+jEJ6kQmYuL0cCv2QrLwb6hI6PHmed
7g7mlEwj206jBDWlSVrTpm6OW1Cg7hOljQRLLDRquf5lYKclKUrFLvITiHKNvaYWWQ4TB+e6TkjX
c+TvdTqdS8fEYNZ38o7yg1ydiEhDGxaZudGeOPtZNSVpAC1IFAy4kzRw1/wheYAIGorwoK/YpYfY
J2+sQUL/QdG4umMtIswNHEUgZNwtIg4yHYlvw2Zvh4avXZPujtJWkZE8RqyKF21cHmK1X5xmlKXV
Gyk6TJDZa5RDGBG+1WvA7b2VJOpYQX/cfr6YrMEby90kwjToEdv0yJJLhaVkck7inxq5P58kEodM
1krueHkrM8ze4fxTx9Pelbwg90b+rKOGNwjCgW5TF2D436kkDnzeGtfNL1IVJPZvQuOhd0KfWgim
Ne9S0WbQxMHCwnTFqumPjZBGcMA91CKPzUpizyGQX5cW0BzJe2RYVtUMRYjJHjGc+PI9S1S2ryQ9
h0QIo/i7V/FA6nxrJ8Cl8lAZEiTgQ+djvaZr0WBAoUxwr+VobO87rCqz4Eb4fPcu8U/U7ZKfVtix
O00qiAIPp3HZEu8AvSmYGjoooarzZo56gVgfdXl+sfVG/TYyt0U/zaGu7mKQ8FvKTtAUhgVy8FU1
4B6Y2wDpcNYaz/jKraI1O5cOmwEgBnc9YWnAaZDXl4YVHplR6witQEvxAskjhV2UMysQZRpHTj0G
o83XbN+0WTNjbqcrB79EgCD33XPiFi4uBHZJv/wde+59jVyobTToTSR8PIjmBMOXemeEIlHo3JzA
Oszy4aXG7nsuOeL81ImpGcbJViJqiSWEAJadHlQIUtdNbapiWskRuBh9eYlztll6U9Tvs45JY6ny
aLrUVthVFeuwh8/nP5IfGSGgipvbSobDXCAFTdjsS4a0xGPZl7/jOoKZHVz1WQk1C2ZTxVoSZWvq
l56DcoyERzVpM+Rn7gt1s92zTp59xWAgZ8Bpq8t1c2xl8KEGrFkZEjpGbALjOiyizdWyOX5K6f+W
tAt6wxOecqj1pkwNLamdClowjPvu7VHS0L9Y1nU6sG4ItaWkc/YbgqSi9xKhEuoq85wYfaMwsDdT
4AGapVEx10GMwCRklUVAO6cxL63HN7a90tCuCiY1rq2rzJ8S6lPaoi9Wk843jpgpRjZR+0m35v5U
oZBObBAsqg/56kohI6hfVDKxTlGXHutWXj5vWd1lq8irY9YKqgtyf34mi91JXs7k6kuGOzhdrnOy
0wdkD51FdkIpkmMEKR+19TeSZNmwEKaiyNtX0WT3DIOlcN+HES6vdkI9/nqhSAZjs5NgtN4Yigt1
+sGRuubdgwpqrow7eFh/QlqzN5NNs8o9YQSpOR6JYBYCzC9ojNKQYS7dSSMd786scB5iZTtmt5Da
VcN0/WDrADJOdUSCE1P4rS9umOEZYvsK0DPCaj1cPEW014+rzmZIkxxpAamwcIv1xW+Ad6TbTuJn
i++4oNwZTQxjqyfzS2yGYtk/a4Tvvn3ba8QEjm2PlN48mCyNMM25AqrzHAJvi6ZKTPwbUoTICpUI
5wTCVZddHdONUNYEJqRNo8WJw6ip6m/QtmxX308pHZ6BQKWwKB/G0JD8dfJTfNChF6vuaKes8ppE
dmZQBl2dtnqZD2HvNChZJtx9hdNS1nLiSnY7zR3EBKkHnZbYCrCE3xD+TcTwTOekHpegj8SiO928
SBl2QyZS+WC712tap5yz7P92AXuPKezfq0M3cPd7OeRwgxuFYbKNQpltI4I8bwMvwrdZ7U3fXWT+
WiPvrLw8pKWmeqho7wljNLGZzf4kUCk+K1uDt5KYkDvZ236WKf4b59PJ0xw/CjoL3qInBgmku4fu
OrOTz+YvxOkMPVAWSznmioP9kC9NfbO26UWRgaAGbPxSb1Am1xYHOOQWvME3hQHnc/GqDmnXoUzn
th1YuOcJSWqO9R3oWXCr0euc1+rQ2GFiizKP4ZWLjjsLRR6oRm8R1n04WZbimQwMN50l5fcOHFDf
QG55Lox2lGOVD0gUdXdPnWn74l+UNlJGjqJcTX+BhNkuZlWTEZ/pcfNz5h296np4feJIw4DBoGE1
E0dJ4gOSuX/QN5afS/xMgIE0P8QmAK44FByk4tpdFM1FFWqKCFNn3w83OcsuVgqcvdNaS3+Vgppw
S7G4hBpO0VfJ7Y68O5cS10BcEPj35NyB9agUtxEai6azP/Ty0znbZeOMqAEi7CFPIJRpUS2/hMrX
9vdUHRjE3NCcba9+3tebwlsDxNPvHXkTE19e4UTTapFo05YffHAy957gtKpbe71ejOMHIO2dBKOT
UJR19CCx8GoAv/A5nlnfO0a5gcj4gTzedBornZKTXQIeO1+ZTewKieUJAffdjclX7NVqpHw44Xs6
nxmPIHO1EF13OImN+xYp9iobzPrJbGZyLCoz+mmn5dxcprhY1WhYGcnjAL7vL6jOyWLqTdp8Xy3A
fHL2S1Fzj2xy+24ASr18UKlaquBPAablU75b7QRMDxYe3OToKk4YHdOUXVv8QMdq2REhrrMV0Dds
fChyBYnQ/bvtgp7XFkGNFoqdOpcrN/zq+Dn53YpkYwOi20EUhe2vARq8mcctUkB7BojLMLh5sTyW
hcExhxZ313Xjd8/fihi05hHYr0aYlqzn+KS3qQLC9t09r7COETu3FwUb4jGkBP6mY23GgGeZrjVI
x5GVTv7izLIdTDG7kQmh2OVnmdln6FwmlTRsyRgId0Rz/KHNRk/3BLYu/Bk3F0UhduDaEBeaANHV
yh9LHVCNGa0k9n8xlrI9jg9nO+jL/zO3ZRraGNXOgZIwPtVpxBfouc4TgJwNbxg01lhmQ8T6eA2q
CwI5xN+lU9dMZ5+AqFYv3d45xf6qrKFCR8OFfec4DXeQNYN3ta1ef2gAdi6/OtcQEldVPBeYsD5r
5M8qzYjb9ZNCPEF7CfQJQ1vMA1mPWdhbhwviBAY7U0fJraOWSXfhD64ge8ZGCvpj0W1XrHcSxTi9
1+MpKcXnXSszK/S6fvbCBQ6zrIWxv5YM9pjKemnMk44Qnq6KSBCP5TRC4WXFDirgRZ4btCEj45sd
Kdm1cjYAVuIV6dZf+vKKwQAFZcWKNZyuGd0/3rz+bYvyVwS9AiiufqSOS94Jmlqs0inSyQo1WVki
QRB6Bgm2prdvItB6TVK0/r12zRw+lSo9/AjVzLsZCB8+KjfhCSNZyVS0wLWTH+ZsDpJYVp2nrY2Z
ev0wmslWqX4NxiVMQqC2zvznF9YmdCcdDK4Du5m7bOqPstpKKM146v3Wd8VzmxY4NlBtKimbxAEq
9/ghRh/2sVHMeRufi4htPX1Y3GYIwetZX+/KXb5hy/pAiAWjfAYUPBtgL6RQrpM0TYRfeBCUsOVD
7Dxvsl01t1U6T9ch7JgOLuHuRQruWfeF5g5PZheP6jJSmYMpVc0/jAuj62SchqZppBg1+IRgd5Y6
s+RS573w6vf6EYBGqonatowY4h3fbURFNTF9joAcnLs1t7JTJBwQcoVEjQTxS/MJhqM+NscW8kTf
SA+7JRsOufwVdtP3YCGkLw8qnHpi4zO38Bc/yP8SukNmdTqcJ0ikwZSafKgX7vVCIkZMM/kigZqo
ffATX0jS+Wr7Ri7PpdLecxpTTBxLn7nloNg8bwVQtpglRDymV68J+0pmwoJDHApqEmPnACpNXqjB
ooBdsARI33Mv63jNHZ3z9mEjwr3i0n5NJ6BWpk1pQ2AuyaI27kbFxs/7vj0J9FeXtRQH5iqL/eoO
chPU0y3WbaYqL0o1tgCrD2am54FJYL1ZO0hPme4c/jw25mvzjq3tcFx+bt/VCTg1zxS2+P4jRbUN
8oRKQ0ogyqvsfTHQqpNPR56TFR/EppdiyjdB/x/tKZPlYMDpzGDHB0erJ2ecDLOcWTN+q2jEnnZn
SAxQkBn7V8GTBF/4YMZV6UI1UU1GWfTQCgAmFx6ztK+ICTCprZfq6gIbWxKwkNZv6aHIf4BRBDGH
NLXJy/fS4+mSYJ6jeZBqhctk/SQR2JGaJb27Ash3fZafltfXiuO24PrjOn4f/zJgklZFWNlEsnAo
Pk3rKoh2gTi2QORCF1Qy6E7KTLPyTheCBJ+P2CgTeeOpEcdJHNgrbOrF8sFuDMyqHPR59CYVbuSn
oRfxosZmIw2vuDX58tjUM0AK9yUg+7LCwS8RiLFhsw/kKx5ztl4dHsnGeA7buxk/OIEtABeRuN12
roDECxWIxefLMOoasiREb9OxXAu+7CBJQaA5cdEkFnlZxdY/uJ2Wr3Dis+LgwWn3nEmR17rDJGQR
mBhLCSLIhLZ8BqcK8kbin5eSvYBE7SPNp6sEcU8fLorE2KWGTVZs2cGhh3zIootPSRqancwkUYLt
/5VBPxBVHccygcmHYv2PxdXvIXu8PA/ti8uPFwVmcOR3qNN7+y3XKOiFcSqKhRdgea4Sfu+TTliX
tZ8Xfpbni6Tt+n9pqrZgT0rrqVehbpqCF+oHoaS+fkAP14rPeQKXyyedKsc3ZRwOPwythH3cdNVn
cuVaQRVEiBfFxUJ6pnXmyZ/tePT8tos2PoAQiMrp8qjItSNnWkf6eLhri3zYi0sGlXX4LU2wn/Oe
kTIh+wJ6lrY0/RHhG1EhQn4TQTVAan1+mnhxeEF3qWw3UK549Dozc4y6cyyNx2t0p96g5KurJexS
1Oy6h3rRfUBloiY09aZaJMtKWPqnfZC5P4cM5+c3tBfSs7uPv58o3uINXl5kVwobx9NVuASlQkpt
IXH0Pzn7YsaQHQ/qzRV4gPjXJCCR9Whjuc0X2Rdwozkb9LkQFXAqMfRv8wybJ2jOXcPO3QvVmN7s
BHrC2rWZw3C29XG4FtnsL8Frxn3+ZphUgYYrl7lSRIj+NacRN66SjFJI5GAL/WHm+EDhPy3+zD68
xiTWw3lRWoPdGIbPPoNMqIa1RVPDTdmEXlt6POioMEgov7ba9XdHbEV+vVVLGgKUh9Aaxe9NSI4M
bM+sVGC9VIF736lRlp9UaVSk+4xvTF5levM/+ybLSQ66h9uTuDjAIVER2U7SHJu39IV3yGg3zTDC
YcwuxyZEpqk7mO/26CX0jCrDlFXBSEHQAe5yXdiqclat59H2ZxGVklzP79Fi2B4AhXueNBJ9Ulmx
Nk5sNWcxOA9Q1NlCSBuXKEx0xeK5Cte/SGnDh01s0eiYyuNs49VRrqUocZrKQ7e3AxAh40LWEvVM
CVZnz/LmopKm38syV8GD56ujoWhIyFgvYJ3XgPlQzyxz+e/o8qeQ1OgANdhl2ngEK3RYiFgKb8O2
L0lv9wqXiMGGpP5JtpeaTsgOdV5KOp5g6DMODy+raQUBnssIoa213kie2jvlZYpv7U6MwGWE1I9R
V8I76gkXlh5cS6H2yuYaI61zC8HeV4xJc/okKFFWXgKiY3Xn0/MvDYAp91cwXZSmgGGHzzXl7k6S
vwyrVv4nTaN5jmc0VM9gk9jvqRsvmt1N3X3L6fGIFzCWwfE3gtybrHCZnkey8/TzlqyMTnjpjcqx
ZNXk5NvxoLwm0jzqxK87VINiR2PN/93RQdtd0oG6Rv4pipTtgQB78+iAoUE05f7bGuHoEtPQy3ey
wK8aBRURK+JyCSA+26j9TwGXQ1HteHyaTDv1v/oRdXuVriUo7GQQaIKkhW/EJRdayCzBJ+9CkZku
KdEQzY5HxvJbQbarTm1N2ItuAPnhthRIVrD3YWAwntxNHobRYCTSnifciRnny2iVWUPwRYOMUHOw
WiTrn+wcByrpVYTfbMjKjMnAt88gFgghMx6Ih2KuASg4jQJZl3KAG1Xt8qLqevyksW5BMRZiyJYQ
ZT27SFncTDZjbG0VYS7UfIyDCDEs0T7Ttas4RTXew+EMyMjxaGnUB1QTTVSwJv5UQfsTM9dgbUxr
+wOgLeIWnXTwtizap1jMEeGc1b1tDyQhLhtNdv8Kjt/OUYKrfYstQKNy1CvQsnyeXqIjSR+Fn/rd
himpDl3EhEUpR4JMWv42VQDAGH6CjJwDL1DCT72TZHfkBOjLG8fpwN74ypjCmokxi6d2x8KOp2ya
iCz8PiWNJ8t/UmCTa306yGgT8FHkkMgsMY6vMkNtKyqigOxEnZrOdbAlDVM10k6+XfvngTX9+wLM
763cbLTi1tjDpEUwCj/2U+l+G136rjkuubwXJyJ3OsdFkUbC70YEQyw4vBfuBI13qiuDUgWxUiJY
P8iRuRWxnFGqPQ0WgmkfUdxFzkflGkLDUlE9mtuUguUtRSb4/EPi9NTXdyiOQr0C7COy/Z59gCqj
XO2v+F+9FCag3VNiqz6AOkn5Zm0V21CSrfwe1MDi+B1X+ozVnZ4TA7XrS5D1FPkJdlPrvtlZKZpm
/UYnPbEnHtThQ9EM4kQdVQl87jKJEE4RgKDaQi+S29qAGsrjQRh9o37mML89O5Sk42OhcmVKzLNJ
H6aRnPoZfQ2Tq9NtnaTeht2To23JFkIg3lIugynw1hXi883QD3mC9lv4hzSzOMu9FPhJnVY5axiM
O4F74+AP4j3flRykqZrr8E30Zps8kF6RTxfysiTU2Tu9FFXSVam4QEINUAaPsurQves8NWTYxAd2
3vOGslTJpPeVUP5omnkepRVBNHcEQTXSMO5zhEoFnSmSK0q66ZZotBKcWDwC4SSTNAtAlDQkKIT3
nv0C83vIyxzw3XOFWlse9XNJITfba9o1gmo/3/uayLciMvLBC9IIydKCi0nisgZxYEUg0xnno6uc
EhUIac7Ozz+GrDwL0iRjL/CA9pX09ZJ5+cq6iXqZyxSqXsX5TdzT2nX8D9QKGPBBVr8UJCoEyNPg
Y5lr+aP23jQRm+imTnqGiXDbbVtk2kwJb1Ph82SOgeR6nKpyQfTppzT067SSL6Ykaa5viW7wxidU
8HTXLo/vAdBETLlLNzZK2YR3SlbDTiP+bhUoFWHwiYsET2gwcYNWTa/rTyVVnLhuNk8MBzVFafM9
A32zUzbj1Kp5640WaPLNS9i/8n8pI2hhTBzijcKh+HMLkd3wYt4QvvMPUmeTEDeO3fE9TJ3PnQ6G
ouUFMPyijuqQx4NBWaeEEWOGnQjUP2Ct3P+meHtXK7BdccVN7GwTlojLUwrzFQrzUB9nU/1PlGlW
YAgnftmp9X2DHckQp5TlAeX2cNqv5OVSngb5rJyk6daGVfZlKKXSN6A3GcwcdYCFfTwhV5GPI9mT
fjX3Sthg5komEkrrB7DRUXZ5Spcx+pJSwpDMECspGI7dmmAls70whPJZIvJyAI6DsKLprDGpEnGb
HtZENP0fdDnN45NHOJHPI7xMeAxSLNDYF8MpvfIioQAuLklK7fhNUm1bQs1MGS1c1JOh+IDNyyq+
bsN5tHJ1yN+CuCkDHC8oFvs/A8QMC58TZIec10UYzFWQU/Fz/06idFl1fWSe5CeVNYVLBZ0WU5XC
LY8P0AhWiKKE/+Pia3wNPaxbonT4g4ptNTLfMwfqYeHEcX0AuHuVZvOShMOXmLwuIUZrxm1K+rQG
ggUTvLGShogB8bLfEXB1tj6BuFAOOgoYC0MVk52h1ynICjIFPH/CjyONBud/nkGo1IafqGk9gZ2y
yGZTIPBoK9wnrvSQ5QS4RJchUbGsX1Y/cHMWzQwzTAwThxdxD5s9PBJr8Z6WXpkdTmbv9y0b2VTs
Z80Y2gQ5VXVSFFdlggDsadtpfghXHRn4EDd8yPvg0Qbur28okgAlOBi4LmZ4sE4GPm2uiVGXTr8N
hJOxOx1LGc8eTxaclMdsE7NqECc9JcOW1aFgZDoaFp3pvr6DeNDMlylkIPe4R2eFRZADhGMXPG7Q
mPYeJscoXK+kC+ZQbLEJXTZbyp4m4yMkD/DlnfTkQF2nfjCnMPOqBhbRJorGzuvyamtoZm6Ln4Yk
2CLsk3TjZELozfU8IAIp4PZ+ZZlse5T0G1yEo9aTuokSWoCCLwtWR9Icsrz252wPJ4EqsUBjetVw
+/A/l1fx7/99ybfqD6nOd7ton6PdBtVwwI/IBJaH7Dipq8cyFLHSKhl+JsNGJuskRYbOl6hrv+25
9sEbUb3DE6c4CkAKfyEGShHAzbTCOumiNbQteH/CSsDoC97T1dpRpGnCoAjlX3QBctWB8UdtMUsj
Mg+vyBpeijAUYGZKZJKJ7v6C/+5fEwEctpq67fzhNlOQF9JToltLekGatZrzR6wfAst0tH6TnbgS
TFlptM6EJV4kYHl/34j6NV5+28cvIDUtKgKoYI/O9wGdv+HPkuUa/5OzehwfvKT34urUVz+E7dYS
TmiCqJjka+chcjJ0CtGUXebmQa+X7eOU7vSdK4Y0YYUw45PZUTah63Dm2A/it4qgAA2dIPpGfuN4
5/c6oLEW5iq69G4IOwGcAfRQQ1r1B00wCbXfDxylwIKFPxeIlnYSsogfSmrvyYsAAquEOdNO5fFD
+svkBSSJBnYhvZ4/RBYMVqicNBllPzZAfWFRIwK1BnhI4NQz+yFdUnDmebsN9srggDJGRNoVZo/h
IeTQFt7uvxarJxsNEvjwxTMVbq7exnCsVvPYXD7VizZq0s4FV30DGtMNdua6J/fn6HV8+TTeQYfa
ZGWYF+3r9GpdijHyHuE7vGphBAqS7knr0IPsn4mx4oVjfY2iQl0Wp39QrgvisojhBIjKMC9soOt+
Ejq7b/MpqcBQtOqnmLXNzglXdVtoRiHWMVNF5sABlz9kSaQH6tQdpDTAqvb+eIWJcfvZi26bSvxH
FbDq9jbFlgMS3WclW3D3XQFdpQBHrYj7KVNimgqKekpeBeureXej09jSrKh4ZMq20R+ECl8A+tOF
4VI3wOHbyxF2vXjTq/WteIHRaW50xlxNV+so8IUFjTootqIUV2HT2TufNjsCvDaMXW+iXNso5oGL
znpOHHaPDTimWqzR6k+dLV+iQxDTJHQKpUhAs39F7SLpY2XiE3+8mMIHzNfHl0k1fKsmiIlN2lhQ
bOhMCzyt3c9RMsCapfsgXIFvqPSOkc9QrhdpbCUUP8cE87Kg766h+7o0gwsO3lKuKNITA4suOrW2
WQPomTrHUv++0HwW9M7HqSGYAFoG66x+vFGpzGsFye5BTqZhn+FKqO8G4oqLGu8Tv6wNHen5DC/c
ODVgjOAZr/wJya55nVSrjAGagLUHVNi1GJCQjTKqTTMTjxG+2k4dcqgfH1VBC+johOOUy0eWn0Bz
O7Usbs6TAcmZGM48Jfh7JHfnjvmJIn+xPdLv0OMX3nH1d+8qSLQ9rZwnbcbbwQuVFHh0vLx64S0z
Vz6iynF3s0evN+qx2dhexZiDA3aTRVZXTFC+lQJkL3PbjeaHpZVgQyYT0Pb6krnyq2mprtYz4WF7
/fdRD5774v9SS/YtRHetcxvqT/xTrfncII97mSG4+/Q5hDPUKb9sKXm6ymythPsjNsPAF8uiJQpP
UoWgQdeTKy+Oio2Cd47HNr8av3RS/9JY62Vbj+XGR/VrDiHaYCPH9AU3+UfHJgjePH2HXxR4Z+LC
J+KSRaPteio98m9Kz02i0vG4ECyUgERHtO4D5aBTZn6efJQPyObJXYrYJ16fkyQgS3yK71JnURjt
Mh6XDvQ6XqrvXY0UYWsr6CupLpubbU6aa1bp70cBYkMWjG/1sdG9GEZdl3N3HO427RfvgksfR5zG
4Zp0ZeEtkujeM8egVxS4mcQvTDPqTRtibTWJOtqSHdCrQ5Tqb6IvHdl416T8Q+sQ53rr2U2Ia6MZ
YrGrKjpvodf/lnFoGDqPwFbu+3rOCqZZ7R9JaxxyAP8kiMN9oW3vC+Kn3+AJ1/rwb7zzqyFxbW5I
u9P0GhOAPVxPBdgynJTdgObuKKkklZfuNRyUv0TgPUqoVXjX/NWAPJFwic4yUKcCJ9qWX/rjiq4P
bVYgtf7s/rhx/8Zfg9L2GlST/Qh9RZZSNfzHlkYDa9K1yNkzNXzmA5fYBOIgY1+zof44Fsm1a/QC
p8UatgpH7LWWmu9V3b4DjFWR6j6hRjoKVSKh2FsrRyQ7AHwk4zT2P1m/WKtiskSCX29EkNQMsObT
kPVZjjK8od1qSPVT84tgkTwof3ZerRslRe/OdNye10mWJxgK3V/2ctFG3TbdqZ0waiwdGXDajSzm
seeoNr4WJTL2J1Jf708LchIXIo9y0dG98rFcRZ+kaKoWXEWmB3gtqxmRV3Bu7mfOLA3y8WTjb8mb
4kyiAcHunaEObg+R7Syy6UjOWwlSAwByBVU81E64fwGok3vigI0loJICVil6SPw257iyxqQqxN6f
jfecBYsZvwVeiFAJo0e6b7+s7tGgSMH7V/Z75mti/f5d8U97JT3x8NqiC6zuPw+IX4b3Ar5nr1xo
3UMJxotAJPpgt3b+ERzNxuVp/L2wk346JrmJ+pCa1iXpIv8BqSk4KMPe331QCWH1kcCBfwj6f3Ui
YZdCu4Y3rY29P+BcodiHtasA7Z1ZGAbJsE2ZqInrMSZsST2QZQziJNQv68JXXpxuiZts+O726mDS
nL/84H4S2aC/m2VfzARBNSZpLyFu2jDRZZ5TtaZMPeI1vFzG+dFowMREnr6+wdHbACphCrCFbT39
F2LyKzR6UqJPLWjqngscCMB3mvGDTRaaQhN3RcOyyAtehCWNBjnKvoe1SbItyhtlN9URXkcFSUHa
TxO9zjnanhf86Cq3LkL4PZSXPBdKddYQjrm+vG0FTBwqDoHtVMCtkjIvOjh0wj7XUKGlWb/oTmvW
ZlGqeuMaqtfh/bTKy7n0frCj9q4prISF4j9Xnhk7vaP8mbBOUvHdjeXTf9RKdn3u/3cA5nHAXfyg
d2gRZTgKnw5HzLiVp7mz8Mw0XdZhLeu7KSKacMaT5ephAtwvaxHnF+OHRyZdUX3dtgsVwe6ubXNB
tDsGcWqSyrTQ8kqOF8MF+5CgYXYzUlpe4OQ0ZI8injFmgzee0GPBDkYllLpQUd8UdrSO1Uqg8PQm
2+4E443KCEFaocT+gf14hEUYcHZTXRBYUw8DqmL592eSe/Yp1yBDC+09HL+XYrjDHrYqDK6HH+vt
C0oz6iBB3wChXQiiStbZp/hlrdARprkUkjRmkyvJHfrxCWcEvdoKaH/vVf2nHho3xDH3qmm/aCLs
7CmDuq+TG1xhKbtNUQoEdXVwIrsOKFZ1peBletO9QENxFGD+X4ufppfA4aOMAxbqPqmyzoGsGZBD
y1JsWVPJimCFjp4SdMwdeGo0WBA06LoKnIKCy9rp9ib0Uie6yNDaNi42ZJD3vRK7pDOEWhtFdS6E
BgUeUfu3u3D0c9XN8fG4Am0vFQzu9FOAEEPDuwp2DA0h+170h7bJexMXpo/OmtUtk8tZ2bFeO+y2
Q5SRnkvuMwbIxucMRMzvDi/wh8nMjaCdUqDviW2JsMwbXqcRiPkfUpWkvqyIycfzNUjnJM9Jgd/5
/V4iXslQcjcF7G4xZfR4uhtUtlWFOiikaaACADgUWTP1e+UPBlnhVS54DkCe+PoSWkesJ82z2kv5
BrkSFytkNsOmK/sPyJxMbw39048jZbZcm/CUq1j/zAWB4QOlzwzlhiVEnazzNfY0QsdU6xzp40mI
3sH7J8wbFsu0nrpoKx0/Z6iy2HXTt5w0b72rQ4/xSwCl3x2VM4p3rnclJbT8mfGGx0l+flHXlrTr
zy7t1IIG7WVidPVZA60dgeJwrVN6R4MfvwYlAaScfZ3QiRty0fdjJvpY256MLVaxGQ5trTl5eorb
paWT6tAVK/4q6lGY2984nm9Sp+A2xwhDK8tZVPMk5Mu9BDe595dLzO5fr+S2acvsj+ISW6ih4qDg
TEKWFbB9HQDtTVZ0xz/FuZJweRrU0Q6fHV66cX2X8L5dIrDE4vMQnqUPVbbgBc6ILyPRNt4FO4Xq
SMFeByWw5YuJA34V+aFj6VggoFcQOSE65LExfnnEk1/oVg7zxadnQuEoRYorlxv65AI4f3M5/qPM
5obDgHQHFcpSlq7/YqweIPyg0ddO+uIMN0t8di15EOcOnIUWFgA02EEmF4L4WaVhBE+xJd7k/vvx
6N14IRRundKiHx5V5MWBgbPWoyItZHs0Nks0NIpoLQ1wKX317BiQhT8DtuHgi2MEhaFamLhmE7G+
H2XuV1UCn4GR2K9l4UNBj/akq+2gFqHYuY6HsgKZCcdf2PYFoaxdXTiD3HeVmq+vFeNFwafvZ3m1
9IS7qsiM8Gi8RlvEKO/CbyMLIQPS7YPC8Ah8I7131n3SePrZzqQIYHoHiZyl4jqZzNHKDJJDwYg4
1xThwI/vMuJE7IRFqbsCY7ZW8o4qD+DHoRuY2dx+b68eJnV6JsGHC/a65cD2mIkJ9lHOw4px9btf
0YrVRvesDVg0BLeBPNu41zncpQzFfLxMgzf2iHelLsHFNyI34VH03w/K82qY5sK+ZNttr1r7Bz28
DphC/cQ2KV1gDN1Xi6MemqRunt13JQwHyW5dU4E6cYP0cRHrH0mfPSxV2GddaM/8o1PoStXA+8qu
2+HXBKA2V8U/Ocd879XGLK6ihMVzM2Sm8Dfv6mHSqh906liudZeoVmeZXWb+Ht6R9YReDqKX4ilx
KONt40XfKurFsb/h/eYsHNAtNv37WHmHo+WfzuF8yRn6jnd0lIc7ropZ3tTeHP2u4o4F8Db6e8Ov
s77ljjWwi57TSQJbvV7wgm7Y8aJgGehH4UA1Q7K/O/HywWI9dbJghpIjQTLXLlpgs+7oT1tpnd5f
WLMCRTH4NkAiM/HmsYGGOqsLP7d765/cmSQFHd/IHWfmNqejSq2VFpwFCJYxCRPpVa2KxH+8uFsu
/dc7vEdw4hUL1pB8v5FS1dwAbLUgwSQqAe+6uCZewO/q+k9By7iKGi/5FV6XS+GJYoeyV3zRR0a1
sQgw8PG3SGQj9DIdjkB5fKO4gPtldNqP67rZ3kNDAy2W2TzPGGJr3A7BX8C/QvHfpsXeFGOBKlOC
dDrETAT+Ss8lMqJ6ZGs6FAhJgZHlVC7GmQ4x/OvbfIiWT6OSuJnQ/JakPLqxl0dwY5bnJyw0ottr
TKocODDTkI+a9GG3V4o8ui/nxSrZ/PVI3NvH+LokwNPt2haSMqbsGAs3PaOUMkPKkkwwgrrYXT/t
J0E+vhtp7SDuIW+bN1Ip1VmFQJ8UxAv431SAoV5P66Bvf+Y/Am5fDahBlqjJp8txqWpUfmrSNHsT
7e/n6P3NVYZ8YlNt0iWA40N5n/+3/rduuBUssZvds2fHt7FfnpdHGOTF3yRV0KMknHrXscyp9qTj
dBBzUomc0f02RTuhCil09BZvBRSsT3DvxpcxODXGRtu1CKVLORLLNL2CukaR06J2Jiv35J6N4TBr
VJ9xmKNjMxR2pQlri47cr6BwPJ5CVxahPdDeAJphnE6FpCaGmwGj7bVkNoYhrRtj4HC4UPsRfSe1
VfpwY8y6ByIE44JURO24QwZN7lvLRs8HAizoaHQGpk9fj0YtA7VYGl2hUOBTPW0lzmY/ghGuwJHR
3l0Pjq/L4rAn3Qte/ihv7x9JY4rN9xabvL5bQnsj90rXDd8MaFZfRG0IUWxyiRuL8KsdlrwtaiKL
KDpyEyaUuR10m6H4tTqkqrKrhZ5Wz10kmbZ7cYZuKN0NeCqTs2YkmtEbO5O6032itATc0wBFzRHy
yJKWKSQ8CD0RYwQmkUtDLiQN5HtFlXxLOBEZLYAc2N6hnDKoJQiGfCafdUC8U0VXhhwTGbHfr+KL
wXMpCBo1wN1Ii4cbMavdvBr1Q7z8lTz+uPYHFyUzriYPIt0tdqLno72b0/3qebqLjM0qIPYZqoDb
Oi6NyTedXNTcF4mPSaWyq1oQ/uaYVGbFHiake7D/mq7pGpvp13eYW0JP9jmgq8Rs6x45r69YTdhk
5zPa+Q40aMdvMafgZIns2qHzZHxShxcxfS0QPv3ItlZy1ELUzZEGnhB0vbLCaGKbGXPF+BC9ZfUE
BXawQrhPfszTLVcCYmvSGSJDIUH8JotIF7T2duerQEIWvTEqIskvLnLdcAzlZzEBZsMQ82xC5Wdk
UcWmPs9p8aRugzSVeJ+t/QqH1LWG5k2lZsdNfyIVNkcYKIYKkMsAVBscbD2q3DKMze/ZeY/RhvPZ
xwijCH1SktguMsiaI5lUO0aIVSo6H06Aen35Us2Cl0Syk44lV3meBNC+Ki75N+8q8KTXtkT/9Aa1
e8gZXdjeg21WiU/xKzjVIlFZyrvNmxKZ6FBoM9psnaA2neQYuwHMcfidBFzG74zfswuv9hKKxiYC
VzX81fwcl3MxFJcGjSAsNc8XcYX0jJxnYVYZwlvn561xIAdzx1vVE4nidEYkOR4gQj2SSfKc2g0+
wBVnz+jMO83pYhTg0cFJAfcXElaKd40dsqqzegN7Fz07lvWXl19/KiQqzLGa4Fb6OKNFkRuDMhdA
hfQPWV47CA+ubTueUGkswevkLmDo5nVxvAgIPv7ex3sBgZwf9gLTblhV++Npy525E4JT8HobQhf5
oizpykMq2Bh76ucRf91TLZKokAkdy+R3/2pEu17Uo/vsHMpGCAlPZXYS8iL2U4ixc7GjvjG4kKXz
vFU2eKrivTekcmAFOI62PcbggZOhyP4N/UMqw7cpzrjlnmMPx4Xa0TuZ65OQ4cfUXU/gn2qQfGPp
rjkpYagAGa1WVYpF1HV+6IbtpCP+9ST7X138a7dZTWvqthvKNd8wuOYJ9onRTyNKJGHlv0n9HhEo
Z/BeaTeCAyi0mWDZiC3ARyYoyccvyo/q/CK+FsbEJOacgYrRrNRKdHhw6H+ej8DuPDFpg5FY+j4b
PMXo+QRjogbbjco+B4v3igV/UZH978YwieyOYizJZkP4vHTJY4oLWPj0DtGw9FcMuOamvW7NBQr6
/iCGYc0gPHt9p7x2GaMg7q4Px5H/4a+dPlMDXCjwAtt6Jy12EBrLUCf+CSeQT6f7/wxwg7ywrHM2
sm+nCEF5/JBwwWXS/0JhTkKLTKiDnvNqGzQMpKdVpoEMZc9zH7RAYmZ+qucEpG4ecKY/b2IJxJRi
EshPa5a3LVlFxX5g0vE9hzi85XK6fdQJDCTUACt7xnDzlyjDBlAQCM0mXs4OChf0sNr/eVKUAHge
Zp2yl1GtvtMEyt8CsBBOzzeXP8vBcoW2jsXnuG5PSstabX1hYVlH+w0E/YSa1ZnkYQNcQ2Uoc8tM
SAiIEmhuWgA6xGLmy+kxg29C6usV1is/H5zFHMH9uRIYgrMc6LS4IQwA0cKTuYVEL/3SCcoHXeQW
kBzRyHrplF4xGuJM8c4VSo/6BlQbzlClN+12GU0YE0FTeAinfSE/n0cRuBP5Jz+KAvOPeKSELQty
cHJOLm0aimmKAUOBsfiTP60Spku8SzlCgsUhqohlMwIxgRC6V41vtABpbJ1QHMMwPbaYRVuti8f9
lSLmnvIGcaXfwl73sb8S8ReFvb5HLtRU1Ia6RqOWcoLtjHSpXs/av6+xQYWY2Jcvh8POov8cGhNQ
xEdZz+QlIOKz3IGhAm2yl0BCDWEkUuIwnzui647/9dk6JHYVDvsgT0sAkEbew7FN8AYfvOYhXNbd
9AEhzfp1vDacbsDdLzDLozTWth2HwDwK/ZJVEVeGwO4d3QrPLhRTbnJeQmmsLDQcXBUHQyCJ5Zrb
FJ2xcx16fpFtqgMUGg26uHoroYRcrbXy9oBDtEm4xWazITuYl7CUKaSqbMSPdcKR/cOYu3m6IGDB
ul4MsS4NSoXJw3H9lis5xZXzoubio6VGGr6BGPLPZD03cdpfdRnK2e5j9AiAWHlfJdeyMMWPooWc
DVDGzEfezhaEYKBa3YiUPfY1RbyJHms8IiW/eNcfRzw1L2KkDhVYnBj52dXaro0IitiQ9cAcNuBp
xNciQDqXEt7VKu4WRHBCo/BWjLFPHZwSeV8f19gYevga7nNq/3otFT0xZQvPb0wyCI04F9vOhwPD
WD5rokYC3yhADV7PkDA3/wlrN2mhMR9/qS0RRxTmv0JlVo7Xyl/chomAT3/IF2znFZMgfLNTaYE8
Y/9ty58bPfAaJ0Kuihki6qviFgP9u6CrmVXqdxk5fBnZsR/MZf6lPfNnxRGA/h58Yx/pgsEcOswZ
37N1Hjfcml8+jo+yRAPsBSR5xXnj2OqPAW+SBqchUDO5J1AROUBihZCVRXSDI/W/ZckEOfVjfeEc
dzKRYT3gjiyA79ClY6dVOmcetjpY6inzqbFWTleSHRa0mfx4YWpn0Hui9pLAqAFs6VMK4KRsvaMo
FR9FEmxb+OkvuNAlsg8vLNbvQDqe0kaLxh/nPraGU917Gf6nbpmn0ZvTX/0TtsUgmvoySKwjDHK4
74It2HiNXKxigrhd2c13Cx4lxyA3kBeco1sfTkKd3ozWwUaf2DDgVXDSa3W9HKyHNqwsl0yPMWCc
gQ1+vsL+cRWOvwllkYS3AbsnFku7KlCVeE/sI+Cd+/WmoQOJZcJHYRnh6MHr9AShJLF4oGQv24s1
vNrnJPjOIWi8ENr2UeCYqfwxBy9CpButTdvJYsUCeDVPBu9hx7kj78+JZyYdpt797BGh/e/04kHA
U5slD1It0z2bPQruFNsrSbWmMzCgKMz9nwIVy/IxIkMkNVIon396XcbLsr9KIhKX6zL35vBQ0wh0
qTKb9d+fI1ZGRJyV45YpqYsCAOObRUk+LQJJ9SXsSjiZN3NtWhEyYpHkSt2ELWye7JwurnCcKQhn
kcqwuQuFIoB7RHUp2jQibkId3HUjViu8igzjF7ZcHfjHwhuTDvioxHzQFzMZiivTZP00l/nx+8y+
Y/o+HkNeUyBdpifzppuY/+AefeYv4kD/4KwpHDZWDteJKNZT/yDMzQKGDhd/HWGp1tOYaI+SVF1j
GDVGUjzruvvSSJMBCf37qN3csW2a69l3es1DFEQ7Hb+c9IcNP6wDefVGN5FN/fAXguhNDIq9TUV1
tDoYjwXEyad+NeTIvZCThFVVZZxMAAo8gMIk7EGOlytw3/uj/w89UOUnF3hd04VvoocliHo3Cm9E
93m0WU4K0yWpdwaCtLT7IrU+LhQT1Iz7Qxt9cVqItx7lW/nKGnkvI/tvOwPo+Acxf04OX8iLSnJv
XIIWv19YS1yV6D28gy6A0dw3Z6uLbBrv3N0eYDK+eIsCp0Gjv1SUN5XHlVsZjgndGN/5U3YMSH8r
/b9MYuGgM9FpM5WLqnOdV8hDW4FQGB8TUrSEpQbpj6H9HOYX+Mkgky6rrWkLW9Ify58supdn/Izp
1f7X3BIiscfNUeOmTgqPorSccHlO/MTJdOCcEHKyrIR6GZYvtLCZ3uO8Lyxro4kUfbtoFm3ixTEM
dxRjZA2FZmjnsFyXI5C76qVWo0RHF72Hjt+p5+2fNAESr4n4S9RQ+ZV+DbR28k7TPrrVcCrVS7hT
Two0dfm+ltSndVh2XspQZK+8PvJanrwaZ581IWYdxMEpbXaiJteabLzFkvyyo/1ONAriFeJ/WJi5
NGHdUvDkA1blt8wCS6lpDiN595lm1a+pZrjFnnBa12xE9xrgsCObkZATXcYNOWy6tXgjiMaR/HEz
tv14QCL9Uj6nLiFIiJXDXAxHQeETm53MFnUvHmo+m0omuxWqFcWRmng8bkR4Z8PB3za0N4y4rx57
nmTLCsOBVY0Wg71BMvhuBvReLEi5iMYZVd7gjI4wXMFfRrMAv6wxqjqsDOiCC2UjcBt3zkxAIB3l
hBOEVqb+NDAzCTmGANNYfBMgZAYVWWI+IeVoJ3tvliYEtGUqk1Nr9o4KC9oASjCAB0MRI5JrRjvs
AtO8R/qq7+4AUbn0+8hYpkXUJS/OlaUgytraYlPykQg/P/zVkWvC0fyj0r/NoSAw//AmZJk8djQk
e69qrf3kig4u7Kfnwe2GvAnJKEn9bwJjixFsJbbkocpDzD2wVBMjw+KIgT/BbilfxwbNDgT8pGGJ
CIZiJLxn6/qqXceGkgqEbYFdicy2mdYXcCUaSQaYlzkOgRsFaLwfbs3BMaWsFkbAbCWSx6JcxgQU
Q0IbLCQfD3LpO3SKRM4uVe4QkhOzPHI0XUOVlF6HHcIGoDmr8myHzcQWLWtSjqKds4y2Ml1Gp10i
/SeWM/1+aRqXEbIUh/sTF7dtzudX3dWzQM4VKaGD66OZZCJfDzblMgCurmfcsaMtzTXbs2n8hSr0
piB3Hqvc3HG/3wLbSDY+YWANJ4CgqIhwW03z0QA4G3eOVJGLNv5zkqaUNpHLUA+WOLkW8WUGe09p
GAhU5Evda8tzhOW3a+LijEcCbBYZboFtg/Zl127m/+tcdChl4yLkS4bSCpEZoAS4wicA7vTUreI/
dNCRdPipu/peygGXZYYzbWp84WSb3u2wFgQi8VDp8vUrkPMQxKt6gAadQJrr9MUPXNQwG2Nv3VZ9
UzvwLBXbjQQ2KcpmXCp39Z2nc2UWAsfv9uekq3S2Sv/uJlBMzKoh0ND1lRzm+3/MFv+Wmv4GmN47
1y3G9aj6oGuiG+Q3QQ1mASRfFfYwZIt1/lekh4yLyjYSfsNTB1EVufZ3H1rkOgroLvfyDtC5Npr0
i+0AWpURlk7ao5OndJk19MkNCDQTo5mdzUYLfjwF3RiKc9gyj6vINIR9xWzFweIftNlNT91pdKXm
w6LLo06ucgvHsVNNsp84xM8SbNnVGzxugjQWIdM17d3o9UIrn3mGoUdgLVee+6Y5RhGHOt12ITLM
79lmwdyRWFJZtti54Q8uyLQpfve/ZazTWVC7Qvac/tQP4IFlN/sLnzkh8J/7YF4Pv75XWjY5Je2n
QmyTZxkR4kTE4AS3BWoai5cbRUwN7Hxm8tPDnZR2Y1fPzvNRwoW2ntjdHJGv1Ti6JewCFhwgH8jD
hWssyqHCkGXFhtEXDTIuo9YgWfIgQHff03Rv3m9UyGAa43UBX+iXJ1xfjLWjCD0/zaEgQHScyxY+
mhIs5TDb47H5peUHecUQwRR8QNxPhJeddIBtzH4HD4OY7cGEUxAopwdFx68lyvjna9gaN0X8wU7x
Km7PRKUy7deUQjKpcff8KQs5UU9X9hbzI+x+yH4+P6VRknFNzeYBkhjdU/b/PjgyIpxDRRM0L5Qu
kZV4r1U1o2HXhWFcyjjgxXTifKz05Z+E74WOdnYFFBGnRWIVOY9RXd9K3DEsl0xz7frwGa37ZclW
5UXjxb9U9bRSUSdSCutX20bBqLbIoCDpCfdnqFO80RPyDR5iillDFjtbArCK8IjihDt+QRHW2Ilz
iez0QR0i5ExYLYZhVM/BDQ0hgmqQAdor2A9upLSzbeoQXOwN0HNz9omTfsIDVl9T7qfkG0wxp2dZ
Nwh3TOSMdegJdw9OzW7mtLbXhEEzqmBuuFAjOSCkwpqCsEN2RYmKYrmAmJFqO2bxZTIqg7+pGxSU
/K4IbX13VMsSskzG4rsNC6I7+wREsXkYO2TnHfGxlZcXA/5g8DDu+UOiAi2gAaIW4MzVpzUJ6o72
/M8cgrOgsFlfQSIi19/qhq1l3KFAJ0uNKbsIPUD5GWVA9/dJmvXFTAn1PA3KN5CJU9hDilQ9yAT2
52A1aGWfeU33opRve/ADo9xBc8y3sBGSsS3LL4cUQ2qM/q1/lYHF6jA/G3JNxYy77LH3+x8E4Uiv
kNKeNI4s+RiJY79hc5iJmfHly6UK1oc2FPlt+lyHpzA2V6zCKmezsk2N/BeekXBO1tDDNucEI0s5
H3Z+cmcuMDZVmNaex1SRRCfG2189vK1kkxQrRCIu6PQEFeHsUYpBm/JIISKymu6oLZxFbEo/KEff
cM/yRjub6o91jxHw13oNrGoYKbsUzSk/7aao2hOTvwZAFj3ChLEjKXKGHV9nV12//oWlu4MyHKb9
g0+MQc3bYoLjXv2KNao+LdsuV8nv5pP7YBGIY/cwEe+NMz6/aUzM5M1TkmkLI3Y4l9QI6HMoVRLw
mTUj64P7WXxTvcYl+fSm0BZJSo5vVSER+V6mS5aaA7xfUcKePvKupduPmSUueK62hH73V2tAkyu3
rnyMKPguWdzVXE6B42GCwYfu4Q2g9YOJ7kpPrpqfKm9WNFGuOAcXysBlMea5pdalLE2SsA9HQo/Y
mDBFiXJLd5KR0jP+NDKu/N6u/ZYH7H0/sM1lWn2wWUoSVvYHwR4Fj+aZbEeJS/m7Lx1A2H0yHEj1
6N230CbRraJMJmKxg8u3GBmgmxruS6pdtp1pno2/t0PACPR/XE2Am8QSWYQ6oO2ceCnXadVwxu6z
IOPYfXitiB3684CzzWek/daSnLbtvG+lpDOyoioIph3I9PY35pD1sJyg97cINaoqzxli2P91nE0K
F7eTjsLCCTLPgMa5AXhoMkJ5OSHsInM1RCh2qI1P0IZWCkeOWKrO0YHFDK9oBd2un+h1lWpqfHA9
L1omUYb4pWxsY6mTnVxH4ktAq01c2mQKtCLwhAU9DcWaoeCx+IHX81pg0GY1+82f9/STdkIDr2P1
9I0W+7YXme8St14c7I8s6pXt4Hsqg9Axl1Rf28o5q3rqxJuoSYFOU4LvRhc9+F/PmkdkKll0AAsf
Ls0D4yAlburtr33dWNtrX1ft6UzgiMPkt6KZJ0E2BDx1WRd8lLMbrhTyjRseYwScT3KC+xLGlF6z
WJWnP/A1Z9gPAzag1FhSv2jvbsGIE1m4aQkLU/XAYaRuFPL6IiIhYmMFbRlbiTp3ON25jYLyqz6o
piolI7LFfAjwMHFuPNqluIfTRnnFwQ6VyONi92XBJ2pi+X4JGdnYzlrBL1UlDbHXNQtOMh97TiRT
X/agL7vqfGXBo2C8l2mBWsYdhbOFco27l/FULUlVCmRKr38X2smPtWkYtExMpqZdfSHU80ChZYNF
rqc7TNHsP6g7kPc4lobidsXX0VnZ6zu3opuQjaSx7LNDOnPd2FTs200WBxQkiCurWNB1GrIUzqZX
FHQyItMQys4td1Sm+5T9B/qyhnWpPNdNMmBzX70IKVkOTRDDPDt5ouxX+FnXCDLhsx5HadtOSmQf
WLSP9QkTNVHJjDwLjiUqFvUD6vhGpNBTnE69khYaINPoYFFsSRv+tmzpzz5iVGg/auk9ZiwPuxWZ
f/QejfbQxYSbXbfSRRu6fg2Od7BsjThj0yfSVs+tT1u6gmvRQJAqZnuHEGj82AL6l1qH/wEVmqeg
cZ4KNldlufDEZjW8hr6PSHKgaHle9TWyE1lp04JhWluYqHXFR99p7s6WhnfXREKBC08KJmRouAQR
H4wjMPSmJSOL/+OvZOPD3intFFzOJswCfeqY/eecPuKL96rILOHyo4iB9e5gTlvyAafmDmVCCyJP
pLBV1TtU++rI/QexAhTu4HXSlyBjHCEThzlR4PgADao+mHI1Ueyq5DqQAkyYKvWV4MxdWLq06Or1
guWXqmFkFBoYRJE8JMz2qjHp5LQ4504MIqIT3ZBp8weeN6MsXDR0sDY+6GN4xOI6urn7Y7KERqCN
Hz5SYIqRt3wSG8z40xvQ5rknhCi57gIgSGLSuu/RMk/EkVeTpznNqJvSzWdU4b/dMUGeCBt96mma
qtOy/ixQKi7icChWFhxyy7LAtDkD9CsFWlh81W9ovYePQsphCSiDuD++xE5eyL9lk9zgK42NErMR
JGxPpwg51G85AECRV4kHk/5RfMPqgI+hpcG1GOgE4TfO1O7WNvfDiFUwUPtEgC4DQfmLXud+yHpT
op4qVhgj4ZOsHrurwzOMn7ZIVpm44dVN3xvkK3ewZrvFL+Takv7kkYnmvhlGE3IZw8oBAnR8JGQl
BYbbeGvrtExTWr+0r8vAMbUnoGV6/UbyDFQx5HlIgv6GdXUgy4Sh+exnCoVFC3ll6VEHsiJMYa2N
t6PWXpTN8FUV47BexeB5/tejgEfLwsp2W7MYPokdrOpsQaQNo+SYMQYpTSBI7Pw+g/OCXASkoYti
kvYUZS2LlUjfP/YpWPVjx6JHUqvCd+DJR7wdrrg/sLdrS9sfixVGltaKlv8VVD+ogLPWDHYmJMKZ
Jw3OUSG0ShQlnBsqtmVD/fMbuTPhBAzygBfs+uuNBfBiNccIzkYkaqbZQEPZHRq8O6Z6MzDjpIl9
a0Oz80iR9QVCVddUlazS6/gRqo4cWOA7iRhRDgUv5CA3Z2qBYXkFPD2fiTOKUmBRvKrzux51QdTC
cQ5tMS2IRLLi9xuTO1o/HJMYUGOElHVCIHaZUvtmTBxURFKh1fcL1ljeu5f4SdgNsL0+bfVKiTGp
4Y1DIfBZexqGZlBY4crlq8G5U5BaOh02FiJhSEq1PtLHcZHi+9WAj/WsM0UN85V5mm8dx8DRuUS9
1n4Ep2K7Mvue59s3r5lkH7CpioV2MMJ/qP5qIQUH0mUZvuRiPEcYMfkp3dt2NoCILATeTJtufY7j
9o0SczMLg1Fp4lquH8e/XvlAX2ZcRa+IbtSe2mb5JfMSXyqBsdExk+MBFEx8W3BCPmjvfjPOH7G4
rwb48qbH0+KR0OyiZl7i4ZbZo1I+0nBAXBvnU3KbvTyd4CyiXHaflFEWYGL53A9hW53kvxQLhrN4
XSUChqvqfbx/Y2EwiuUWvx4j2MQZEcaccchh/F8hoN9SHhimaUVyaAdL0n9pc1Bs5vyF06b2BjKy
UOo6qHGdN1YkUPZr4eHR2XPSw3yuRAPUE5bW3mVb2SqZs9F2L3dpBgtuvZ2+wvV62MM4/wDoRC8Q
3hZv2fLb9FkS0wga7YxmTwvwDlNu+OWiH8bG5AwjQDzhLpH06XwecVCS8MQrCAc0maBPC8janUMz
swMDTuSFz94IvkpcgtwOXeVS+EjG8gTk24dN8T8l5DA0bOfgqUjo7LIC9JGr2ErdpZ2X1W4jqJ8a
MellNDe5G+twUPnnYcHX6MJI1kJyR+OBxbu10hzEm04rZ7GJ2PASkflYsquE1b11+5KDMnDcaRxj
qC1zq1CYcT/S/wNyk7bIej44pT3tcVBMwSTW0MMmjtPZQ0QCzr0glLYz6tUqARjhesSd1VKmH0nf
Zn6eHSvR8yfiO37+M4vqJDRhnBn5Fu55jAQwCKlR/s7SvehkecSV+SmQvLxXWsTYBa1iETuGIM24
rn0AwnbSIcd5bHYo3WKaPJxAIr3O+t2eMDy3PJZ8+lMTvoqyK5oitz+OmESDV6mgu0GM6lzO6zob
B2wOU+xDz6GzrlXJ7DLaCIxIdlbDmhrEsx1OAWYBjx3r2D8yAtUxFkv7YA7sU0ySxq0P0fJzb+db
HPV0RNAIFRPv0lQo9skhQV6WmRaadh85/mIHLvCQ3CT6cFyx5nB2MZybWeP/+dCZxaj3UEq0ra1S
mDDWzbcxMErMh4ddwUtsUdqsZRSYRlmBaebAdAHBqrd3kr3lWfiM5fEVSFI08M6Ntw3Zfo8Ej3Wv
6VJ/T2Nx9U1t1g99+Fg5CRUGUaRR/CdJulcHrGzaypL1ewn/UDiKkiiMJWR43BhuFw8YOn3vJuQx
PiObp5LL6JboF2guNp0qiS9Qn216iUZ11MDpmYSykl3fUoypQJtkNKFP3uNYQyXAOAV26qirI3Z6
ayZ9OUFB2fNYjS4kE+9EwxF5Py80LjEqAPVLiY55eV1Tij8UbAa+BSx8sGdB2HRCqwmwAi0dMJLb
7U3uaYqy2XYx41lIB4dpsyRh1WCHqx0s0w/cagExxHUO0qyggzEf5uLcLwwIB486izoS/FJse/rj
DyIfhQvLQeTFb1Dj7gRksrHlD4wFfOE6q1hMSQAUaaHCFO4lWdLCJX2apCBB72+Nxqcz7Bail2iU
Qgn2xEiVya59v21myr9LL0jEyO/H8r6S9+yk1WbDpSXfuyLCjTp7qemWoXAF4syscOzyvxhaED6g
2Lo0j0yKbpLHikGcRdkq9efR+xKiJ9YB+Fuof02iBuqQCaUUTCMKi/4rp9waisNnWHa4UIbKdqTT
G/PV66/BmDe4bbKVJjayfAXE3b/wpJip6why0j/nJMtLZuGx26O6NtO9PlSccEQFY/53B3DeceEA
zq96cnFGph4KTiwCt2W6ODHer3qLI7KhKa+d6bCbyaP3Z8WdHs4oodqxG7zJn0fd0AAgRG/8x4tb
dghzRS0XgQH9G00fEz2qlnpIy4y+y6ZrrSIr9y6XB8MdRtaTm52jHIofANhZswQQPlZaTZjFnqtk
wLHt3mzxKVRpD00T0GuD+XkInrAvEk2J85NcKw93e8uhnD1gzb94wqK28ChmtgeyM8zaMGrAzvCS
5XVsM9g9V6hRaxI1SBslZO3XvPsuZgRaOBiyecWbT0unswSVjSbG1v0YeWlTX15ldEMud0vs5acl
aUGEfywj8Y3syepUvZylMW6Qtn0j7HDyZNA0Kww60M5v4U08Y31zSJNoebQGvYvIaOUOhC+6UgAI
1xLNzSDY+Ea6iKV7GY/V7w7kyB8A8ecZskbcI3qwMJAe2ck3QblL52Gv/yI3AiUBUTD5/bT6ocak
5cwGWFTVSYEi8pWTBpdHeuaCfkRzPUyuOoHyb9L9DCOTrX+MkWN7J/d1KuSoKsxc0PLPqcvKcIoP
h/4d5Vk6Jnz9l8lYhSNdXT5L612v+NmwuDowqZqBrzMkP2TWs6lUVtFjS2nV0QRsUdqS0aGNQYO5
usBdg3LJkx45ga35e6iwxSaHvUF0Y48NZASt2X0Uv3uS9CXR0DVDTyp3782NBC/Y7G6OXd7yQX7o
Dszc4MUnoCXCdwbVZ+f0PBvol/Nk0DNL8Sx4BOBVLheta2v1UvYSqUVKR8wIC1cjorSiAqKvDNbe
c8oAzXyhYorBlC7CW7eUFoxqfk8EyL69jJmRhokX+jseQK448+7//2ovOkEboxcEmHTzah45EkpX
yCAt3rkxXLI/bDUKVCMyzM3ibJ8bRCcCg7dyytKAylNYPw2ETK8AH9E8sSn41HpZsJgmsET7KZfU
2NBNDUr8Ld6cEAWeWHoNNGaSzZK4H87VuuEhTf48Pk55vSGcplgIsO6lxmHaOwLEYv8mf2WvQrWC
p1FpOhUv8CBJOXnfonnburBgHNURAbHGKMdytIv33Lj0MgPj1ERiSDlVAt7RRUpH43WPuTUG/07F
VcCzwXhbOZCF98LGlFD47Vt5jP/Xm2h1brWZJTZXITmKfcjQWJLSSe7bwlqcI3XEzLmTIdO7Znga
ddoF0m93QEu5l6d9g7rBdptAwHtKAvIlqqnqSupBfX2IThHeUUHvuwYFsi/7cejnmrWsLuJr62yq
dmowO+qK974UC3obNpFK2tvC3Tcga12tTZb2wz+KW8IkHkQWiYXe+HjBmMPLHViO1qTUaVnH1nGT
BYFPOqKBpYqv2Qu32jhzxO/zdHIqRznr1Fr4LBqJnC0R+UmgiBjeQ+ZGOH7iDir3qISDCTBrVP66
HEnTPFdMDo0QS2G0I+lQf8mANXruQ1QDA6tkVPy2kgkSH5NRTYMY3ejACmwqIb1x2XUUW2Z6nRSv
feeU5z1wZ3iGhFgaau+hV1/tuLunQ/eMfMtZaJAo308ad1sa0a98l1kiek57JC1h08Ow/4eIAPuR
pdAjRkp7b3sJEtdolFdj21SBBlJqQQHVALouOULcAGSUTiVI1F8jr8PBDlTplNfIfpdIYI9MCuGm
78f5lXelFoqTFrJF/Sn+/xSZmWA7CrQjfu2GFhHHPzo5VarWaFj93v0Ax8LWVFqm1Fl7mH08b8OA
RvITedwvpj3uqQ/cQ62tsmFqH5xEt+3Z+wN5HKeeS45BbHlZhvtUNmqzOf9cCW+4gCG+ZetSaDpV
Kc37QzzQzfGc7+1NeWAsf4perznEbIzyAe4YiXicq7j2c8nwQmAZMdK5E6WQJZJ1Ps7jJQivs/G3
8AgEH7KGCsGsboyGiTlQa4twiLDSg8wxQ6SrjNO1RMJuAQIXEI3p8p/Pu25+panZAoV/n4L7vtWH
bF249L/U/uSv9fc7tcRUOGc/lNd72EMbDRD9l/7orAg8vPudEii16yh6mY3Ig19mTQ02ZL8D5hZr
c6qZYIYeVwM6GV6YSG7oe0K2Nw917bx6+9faYEGrSOaENkosSJLl6q74KzoXvF1m/0ZLt9rJBYDY
uPmcH2K9f0YpgVutJQrG6xOQUaTBjaZzjglksaL6KmubuxdR66iaX8sBmwnpsqQEIqhWEWY7b96E
+HJbvRFLVRT3eihrYbyc4I9mbEoX9Tf/d/tUdqOkZOEDJq6VU/IjOi6RMDxtzp6+lJPMGEKcRrAR
pbSnRq57Ee1rmBx4kHWWFwqCu83ugj8vzgE5dMrKtdavIDL5Bk2CaS1jr964NipkBhl0KayMnF4Z
YylVVdofqmd82PoHsmWt/SLCx+sjnEdWdRW2Z735g/19g2OtzZcD+mhae5AzCVI8Yv33qspA51z/
loG1oOotZ/ucQ+eOImWWKBVF4Ze29CF0/pAQe1bgqOrcUFP/9hFLWMSpFxBkQsgt6HT1xazQ+klB
0WtWjJk5atFosTlWnKoD2W8tF4kO08cM2NrLnVV7iARqLi3T0iMEObs+Xd8SIt6PcQjUDoAfGDkw
69aGvyQrjule7BdIGO4NcPu+ebGrLTV+JbSArpZG4xkpi8v+IKAnvAiHlQHhlddBM3BrXnqb4KJW
O0BH2dZ/n1x5ucrpTkhjxMlyfiuIhZ/6F16ZOEaUZHAe34E5SUDIvkGqhKfwfPvPNqKcKidViG+G
qz32PDy0efBSoDmTCn7X0R9ByijuFi65ZCbsaZnsW3iEI/mxM4A/04Y0+et+eg6g5jf3+PEA4y1p
dP6xD2sN40HREsCZ1Yzqkbta8fRGn6Kwv+VjAXEda9lzk86iiI0xGmnwmp5ZtzFMqeW25J0SnIMy
RZdkcBMcMMP1vb5xj00m+6arqjxQRwdbDiferLd5FcSI1wu553Iopr7Q4IaoTKnj741Dr8J0jcGd
VbOhh5RPFSTrdy66Gj9Jv/NiEUr4tOKUBVaR4C+Pgrv5/iLiU0vGNisl1MralIphJc4404vPFVsj
X2wi7A42LyGpBEkbgIlWvK1GZ1a7tmzJlCb9Dn7imPGiiZZ1x6PYLEW3HF1CgRJWYYKJhVy/LR8R
EOb0ZDYKw9WJujluEQlUE+c2cChJObiGeh7Iey8cTAW+9mDiOnF/jOPq46KUoGzOXolJ+84J20FC
osFQDDR4Ua5ngQw2+SOLRY6bVWfGQLQulegczoj6GPK55tunPyjvoMRiU5BzIoHezN8Y9iL2UfUj
axaZY0tUSX5O0tGiqKsOxDUwUssnFWo4mOUbpYoxUp0jevyPOqtspxjlfBkQiQeEpQirHTVvRbZ1
XcEik1RKi7dmWPMi6UJl9v7bAjLSqR6UaAwPvcqS8K0kSNp7CPX8YmJ6giEstY7z5y6QMtqDrOMs
IUOxteRjVGI5WesGL46vLz6oRF3WY3cu4o1+dx3J7/SdxZaXwhzPxQaEKcTpu7n/ae1glLRnSPX0
KBkvwodfM6RgWcpo9aPZOSuOqX6ByH8Ls3wGxa+YeSYy6Mu2KXzTEM7XB8dpbOqrsh5OFNYasixh
Gy6loH+r9LwKjjshDAksGgbmIGHYFL/0qDcaypktRIE5IYLRlmAVHSW+y7fdUw0hOrNeu7Iu70vL
FVptvcMMP0a1B3zcLRdJdgMqQZPCa1Xg5EScISh+4MX+7FEuIjJ3rWT3AVdQ7WV4gMtidmzgwK2k
J7+THAiIUbquutEbPFDyeCM68pvk1WMjVpG7t8vR+USbARx+kyuDOprFAURuuP+p+tYgmyNTr3Cd
6O+Adh4tN9MBtixqwcRxBMpl6hiP8ZiEqZ/hAmeQh3yn2pPGoMwUXBYqkRlMHV4U/5l19SMh221i
DeeeRorjIc96LK9jPA7cAuc2NuzXLRmwZrPQcB1zWVzcSFBy1Sp6aqQUBocjA80V6pn8BEgRknnh
TnL+DLoXmrfB/hW/L0u6vR/Z4M7mroNJa+fh2vNpEgpsH/1OJEufYu/aXtgbWYrAiY6X43IgU957
cxl14JgXoLjPdyTah7e6nzOjXoQjyK2A9aHFDJI+nHjvcB/RrWOfQNy46YKZjwl4KQ4380DgIbtB
cdF9c5X+rMvqMXnzpldK0YZKjFaKOVJzhgGNGrjl3cTBRPqn8rVF2/rhfx0RVt1qtmTa4b6GwBvU
h1NNfIyAS+KdLk4cz0o+ZDQWEePbBAu7OOg2ubqvHQUdzTlC0tspAJS0o4MIeARBXK3elMUZ4yhf
YuAT6iSPqxD31ItBr3A6NamdOyPg4+/06nm6QgqPROxg8un43OpeRjVM2bFR/uvztROa4nkFbLwX
NwKK0w6NJB+FJqlu49eDSRi3dtHH+1HcdAK2juSkUE1TBrHNOCAIPM4ge88JTbbbZBb+SPmiDdNw
A55XREH3sCw4hIO/v5RblL/OP/7BjROOfkdiJ07uqyTsUHVEEWrZhAFTdXI5vUbG9713zKiWGtg4
TsrYtR0B0WiixhCf+GypGr+gCz5wYIA+ofeSVGMCEbQyKutRhzRk69Jk7YY5m0vuwASGgruoXnSl
d/nmEdWy9n7NE7eyfsHpdkIVE2Et/Tx9iPqR4Dhey82fs1DsNxR4leRgyAs0gYXw36HPsZ7lBIJ4
WUseOgjQVzZMBXgzQ0PGa1BAsi3cPTpNNE8cnT/Y2kpjmpvxr2Ajwx0w9v5SiYLruhFf9CUT9lF8
nQrgwOfQTT5Mg+4jAp339DsFiDeupthCAUdx4LJffdR9Xuh8ojesmmxQq+exTc1Gc2qiH1wOpDwO
Zcf//NnFQExLc230lDeGkNLiJlZvGJbHlo+GN6jdQFGH9LaPkcGKT6i2Ekdl9OCtRA7iHaTu0S+2
3sACu5m78bgp/rvLT82prMrAa29+cGWBkPetvQ6eRKlyhPzB+tf7S6knJKtv1lX+3kGSmuxjR2gK
YIEyHqHDElkNAfGjJ/rUhqWPjKVyYmtsQXiQHpBuZdn4RbRC8vEp0H3Imv4xinX5fZnMWH5LAVuj
j0nILzgoX1g+HUuMwm2XV0+fpnZYlMTeBESpgpnJP8HSIMV1vX/ZcXbNvFx1AI82i+M2YQ/55psd
FJz1K6XmNFfmuPYSpgZfMQTW+dFdLa4v/uX+Zy1waS0jLLsTexthn73CXe4/eV6seTnFlSdb5S08
fUh/2A9/q2jX4nWUEu4kzWbywwwCh4x3DtIUvF/huK+kc1EMhUXpmKN6RN62p4a+xfjj8QETtIuj
1YXcjg8OrF/dlnEFmtsut49DfieEhlzufy6+DQVhRj/su6wAgAjsTVAWxaxjcHLyqE0V7cnqatdt
CvMuPaJJqdoA2l/L9QTDqBkI9IL513nOkjdwMUqw5dCqPTta5QI931az0gckIwtIcEQzVLvBsfin
c6xFU+IdZNoZo0aC4uOODODaDl4cRG044FRh7IPEb/AIHkED4exHxsnR6U6lD9as4qVRL9/Uy78k
YXTW7DyHtjGtMYASZ9V1F1GfY3XsIb7Sa4DJZt24Ap5FnQ5Gy+V92DKV7eW5WCySPzL2QY2xlMx2
DzYdQ5GjMt5ZBP3vyrCp0+x597z9hynwvApc0A+O68JaUdes5CLLjyZMjgdGOo2ad8ibYWUDNBJI
Q0l5J8SKpYAAv4fLyo9IaGG0hO8kCEq8fMhOdbDXrX+YN3AiZfmn7+JBsG7cNM2pg+fs20mIMXsR
3YtUrfa+8HLXQU3vZqtu71sHjkUh1elA9wbdsTrloG8lw/34Z9/6yuJAI8OdPV8dZ4pO4NFJrHwJ
6eVSSLtxcLQKjd+QZomb2OBy34Q6ssbA7pinq0oA6Kl/sYxk5k/5FkSdqc2hL49wa9IkZe97welU
pjpSw2aUe+wugnJ8WDFAf804LM4Iu8U1AOD4nqOstcvUK6TlVa0q6o6rQH4BAWww+PBlgGAyUxM4
eWqOSOKLaDsyCNwCkjbFPV1Z8mRN0a5CA3LNeVuXDebBzl34UAvnA1FLTCYmyMQSFV1baQ9RYN7f
DdjK9Sexc3nmlYY55aK94qVQoc6RUzV6I3B3kwP89UBmCle7RFIRW92WaeCQoclD4VCzfBvdt6BD
3kJ8ef0KepNsytzwmWSIHGtIypIk22xwC7E9ozTQlR+1NiZLN0pA2tJikHBfmNCbbH/SdQPMehv1
pHC0R9dnVBiMSQLeoyvTg7Hu31AJFiFv0XfcTkRtZ2i4e/kvLwJkVrULyxTe/0VrPrewjkmqk0Nh
bvpHmE8DenKWNIitdzS7vVyjpkTVY9Ku+lBHsiQA+Zcum4RYT+808w6JfaZpSGf2oemI7wzdtzgQ
FxXmU40FTl8I9wSPPSGsJngzz9QQNa2JbeEwQk325/DeIPvEfNHWR0CchuM64xfNtCC12qNisMyg
1DicYV825yjs8F28bweaixLwcfiM8f5EYR6MsNLWAGelCNTfSXI64tGRL9P1NptURyG24wsk+BeG
4Mmp5AEawXHlIdNn0RbpwseiBKsgjWStJqClVtq7Fu4QApNDSXjA9cA3CQ8z6C1TpKTsmm1aXdOt
zUFAN9wxAxjy3uN9J49aqDO4bCtbi4yNS3rPE9Kn7RzPRlRCRUcsLZ0DfcB50gnetRAQ9Pc1CuiQ
Q8cbYkLDZml6FQDJko9VlZar0SpdaOo0w879LEAiV9UBAgBs2zLJVScZIko24mwWExYG25Z+G8tk
L0XjvwW0zHELjPi5rOe6JXDgz40HDfteLxEYUn7OpOBDAYeqIzD5vGglv8PnhCiw2/78Ma/dDcHl
qHv+g31IjEgPFlDbjITisNwY3cdo2Ifz83NUCOdpNjfDU1CYrnwoioa5sPwtjgMlgaYDCuMqvpWj
h1lvrykvjMDswFaAJzP+vOo1W6OvxcLO/fvgZBcxyJtkl1TSQGn8VOmZXpVI3c8paxm6QOv4A1fh
Hl6HLj8hYpC/m0OJOEOO1Nqd1vtsKMzClg5i90Nvbz7NdgQBSFMC1nUJW/HBmi2IH+NgNjbiw8lB
rpDm7getyG0eQlJ4kQcPN9UtHXB27o2Ojndwq/HyRFgA0Ad72wy1MSGzee0sd3xygjGk/J8u2KVk
uGvACHXcikyxXPL+LnSzxpOFVW2YWauEWN/0skxQ3Wh9/OKPhSUImd/5jFgLCVKALPc63sUTrCGJ
kT1rdT3B9YWPVzsYF1tDRIYGSL3e2sktwMYp7dDa68oos4IPGH31Xc3aoLH5dTXlAG5/h50deDcY
0iIzbArdza4c5Pa2nLUHLy/0ehlFK2ljpg2ylHPKz2YNHkO+BXcRVbNFFx5NThNVh5nqHRIJkb6o
4wegZra+xf6bKMUF9o3GOnf9JDTcqdSzkDYtvI+yFU+c8wUCjIQlKcMwOw1Du9O7MCVI4/uZGMU/
EapD90PWe8cHSgGgEAoHorABvSzBmNCCKEnE2SWxAyqMYQ6Jm3fFkHMQSGjqkLAiTNdukck2UOOk
fHNRzMAZOUK65x3jhcQcjpXITED9t18j/JZW27u0PY+XwwHRVtrJngrTZ/PjCkl0xktg+M5x35i/
RZnMyn+hQ/447TAQhSKfd11kq0fgRJV38BxGvKfLelE0OUOvVswVCnv4SSwdnRpLCBGInOaljhs9
vjAOeWVcnOxHVktn1Ve83bp0Q4vs+tnVFxxw0pLTMTAOXjj2TSe38XCCU2+2DStxhnp6qldTWwlv
Ethge+D5i+7LNZmclqTQGVj99//CVuSHMwr4vp5lFtm64Ze4nr6FNBHnr+HxYJQL6ykSQneOCTKu
5tQu4bJ1bRprgnCpWazPxesA6lEGeLcGrXrbj7bpV+Zbr0lP76iFQIGtYqhgAGaBQPSzKS4aMreE
VO0lhTT95ti5nhkxECgtHLSV4w52WQnveIAK01dkK3zdTOpHo5GeIIhwlDimTpa6Rr1zBETw2dj+
nO33z6TytKEeWSa4ZxrojrSQlan9X1kNyUUyRRleaIYsRw6zk01XbuJqEIqc31JV65FdqJpA3IL5
7dk5NEfowZntwX8A3jaXjnwxw6KBg2Y2c+pg4yWDN3PNeWoaITt2VDH56DInhRwx4mfTb3gtlIgm
1NeGHohrzdS9tZOv/uUtB2jAWp4F73AoF9enI7BL372qtUTf3mtksmAtRldBtwMnIxWgSJ8PwzQM
yfqwPubc/KpoGa6hzXY6GuyLbY+b+POYV+wPlnv6MGO8O/mctXYuWfeLCrXVphT8y07ugOH0v4mv
SY1x1P+GO76J3xEd0rcRtgcRz7X3N6h/455PKG9Vhxnu3ZpOy2xZYXaS8E5/J1sx7DI0pid80ODO
yvlCAIkusLuqT5/qV+oZlKl8jqLBFS2DWxQOeALWe4k3vJQPHNVLH8jcHhAvuws0Jcp4e5k8lv16
WgtU0jPfkdN/ERMXpWvnM/YmwV6VdDvrb56AD0hS2Bma0jma5V7qoFRpq178YETHZI+KbwQjzap3
9gWIWHnOvxnsJ8FltSIKgLWruzyVt9spqfwk5HhhJygq44NRUMZfRPoT+Fdrbb72dlcFGsDF5RAd
JFHwbDiVU9D3cooYebNsGxzfRuV6QKddSO1/mMEwrKR8OnfjrO8zXsyANON3Vv9iLTj8L5SvjJ/c
VdGp1InPXbaFyH/s4pqtD0TqQ5IVJClig1UQCgFYzpK3CKKz9rDzC26LnVUi65wQTiI7H7T5cPli
Smg1ai6ML+T3phGQdgiwbVt9aYY2x0JYTqAC01lLMmhyTUxOGRKoh9/bKbk4xHpytB6xTbCP3Qt/
ILWu3k2o/AE/g5P6O4BY3XlErKUUEBjcvp/tJE8+MnWfbNr6T7ytKPYOzl0k/QceV2izEijFt026
FBEYRUwCYBiiNbfvrG0h3ObnOv2VhK77zqJGS+0I1SXf7IRb1zHFncGo+McT+KqlXMS7gW924jxh
nEzfyRTzmbP+k1V94kmH681blgM0Hnp2TQSIZt97PNMIc0NGoWHcC/aTOv8sha3wolh7/sFFyPgH
IhLXQdRr9Wu/aOfy4Om7+WwB8/izZlNegEyLgEwmGe8QCW3xk1xDkuPTaMPTMnF1qdA+uG6/4iQv
c/mQLBpmGpsXZppeHjAdtu0mWoLfJsoL3yIBhb/AON33A0tqjOw6IIZsuap+TG7QqD3qUeFnpXZr
ApY1xfbfDH7M/XP9Iac5HMSZoHdzvyCgxVhSK5JjCdu1NHPr2XPqKCJUIJiG+wjwEBHszkWaGI6X
1dRwikYmpfszmM2atxw6Wqd4gJS7BXIdaDsDUl0uiUbzKQeXWaO6nY2xJwfn0sfGlFG7wv2CT/0d
4kvY5vRC8KI3szzYPam1TYhZu1SAcVkCl9kUfjhVBkk9R+j2tMjOQtSjYsr8AaVsZcBVBUOGiNZe
A+5SA/z+gaw6ngpcVANpahy7fCUjmd2iLqGKQM7o4rnzEqpHLRFSxXMIz/Dw5kOf4L+ZJrNseejv
mLWpNXJcfetFSS8a0e65EokmHJLgIejr2snr/Jtl1aLeaM6KRi2obTaS3wQG9e3ZkV2rtoIKtwVw
GaH00OKYnS4aIPQARAhmmjc3cKw++6gQBREtbsIGr2365tsfgE7ZHKfRzOKqjRp8pcQ7TnZwzubH
X/Zyl6I5I3mjZPSqD/BlFL7MoAI/kC3datTbAhhSAHifGQ4VKWmz9IHYbthjK+7534kWQj0BxHUK
TkarwxDIstU1WbSAntAJLpu/KaAcpdtbZs2VUG7eBViyuDT7M8xQGuwTeioiJOhWy+uSSIdRRRw+
Uq4iuAoXsVpoWdmVpB6KADuRGg/Ae2Tp9hzmWphNmEc8DNkgbohUtLWOjMDI/wAHhST3zUglhkND
mAQTY8tmTXFNtcKYYN8j8UJ0M/nX9avkat377O40vCurU/FhVDNV7RSiVqpKxFRxtg6tCoiSZwK9
VAtsjMGSJ8ydVxceLBCBHzbua1xcw4558NORUWDOXfFgMVmr7O4S02z6mCN+PoYjykAQOcd0p/+o
M6bPzfYhziJwBySM8zNmRl2Wu+hzbuA1EsSx28OWxaZVa3JMefsbHVPiKHtWVMVeGcfVcbr+Sfpf
OFE6tSZWqE3dCLmExV4O4kEXhiWIKQeWcr91FzpaLjuDilrUcfAKMFURF+tkJ+guy0jL7rLKSns8
UHmbzIu9KrjSLOhA/rAgMJ+cZJG7pb2eUAaA/AWFb/nsRwF2SOLVoxtusQEY6JU+0wD8CfsBqCMZ
cS6lGIjRXZHTA4c64fHQjdZLuRFwT1NhjasqOB3pKSIqkgfrOU6hr9sd1TgKVg/eU8NYqcSiCFiS
1TcRo1WnUYUnNzoTN7HmuuIMNoWhNfl++xOLVjFN3XpzI3fCVMhzIuCHWI5CtwUhS7KpEkz/5Qz4
BU0imYoKCQu6dvZvgi4zl0Nf8gT3MFwUsHVuC6ColnA+t3WLxQFAU5i23PgOLA9/S8mSk5ApiUk3
QB2cTgmTbwfcX/4nKkXVZ18R/aVQntt2QFzZqFehL7RHuQKkaaHrablv2TI8Y9VbcwcX6d9oC25Z
moO0WY/GZU9ZaU2OCUKyOjdS/X/vlJdOt+Y1dW6z7EcsYWt6YJg7b+UHkjxuKTzH2JvRwHkygEvH
I+JvK4vWQKKtniG7++NnQR+gTgHl8j1djHKRnERq4NPJsbEzs5yjkrRun7j5u9BL8iX98Vu2gIF8
o5tjhAEZ74W/A+nYVZtLW3CQcZCnwynEl7rdVutitkWQx9F0ky4/IuD05VdgZue6GPUvLb/8qmsX
YHKV8beyN7NCRS0dUPI+EsHBoe33gNAwGWDV8kbZM9rH3FfTSe8PpeeE9uDDxRZHTf21IktT0o2T
YaF26Iszq4EumEAhWQpEV84gErb9ewNNocQ0U89nIcvTRFhb9U0EYBPfkiH76gKJyDFnSf5GxvXI
l40fq8AZ1insvjC69/5nJijYhoXkcQ3rOokwiIMIw+HbODLQJ5YoY4+z/mIfdFbrGqADooeKg+8Y
t6ANj7LZML+4VTG2HLPFgFM1fBw2rUJzzPYHk7Mjoud3f1AgEGK9IsA4qK1XezFwwTeuPSyBzOM5
Q6nvhA01ll3T1KyMRJxQ3RHOarJcYbfYsDELbbFQ3sZe8DcDWkjlWdi9+/h1+D0VLGphzyxCXERs
aFVOjq7VtTW2WmwTBMuqS7ttaFQ4OzK/ZpOLw0OkGATsJ3YEtzK2EpShDsGja8VjiNVEfx5dYSbN
WC3RT0REWbSAlBbK6Cl9zBB9YywHtYoUl4fY6TBh2a/p+XEhBnkMVofdnD9SuPqCUr2M4Qpa8NEl
yaYO1e+NFekF6RWR1Vu1Ndiuv52kfnZcajV/tz5361MEE3Nq/TyvKwVbwUgbtiV1Mp/leaZ5k+Fl
dx+zYRd/SDmhjQj5xyUa+fzkX2BZuRS4jOxNqlC/H37vmaIwWBJ2w0RtHx7EkTvDBAqRqLe6tnpH
xkl7zD28/ZYvr3lJzone2Ibt5O3/8b0l9GuBigp/Vg6CsWoW0rqV/SvHseLG2s4EuOgmKeyTVjgX
oWvy9e7jzauq92DugINsD8xJqWjT/LScooT4tpXpkOb2NC/YB+ECryohQc8xNSvgz3Tt97KRSVax
FnXjz5q3w7JdwbXoogB3IpCI+GfwufguNhrb+SoduR6PR1rVDZ+0vKsbz4kzDoyEKmp8JK0ku9r9
acKvTSCUqiOyRtWEcjrZtx4OCU/gxHRh7Ne2K5pf7HYiLc3nCqy2qiZ6QR3+QbyomxZocIEhyxRS
TIhRfWTB47+PSwGIpeQCW2+c1Iwplkq2QJfRbnxogHBYb2YA2kzecRp0LNSP79dkrZn4AbPUlAwT
g/EHf0tU+F2gET45y1dxeq0teYVBxDvVO7MtuBAkKqaiJ0glfAfRJ+o87gV3Qg0JVt4nq4OUzW8z
qlR4wZDLnQbRM6a7sm/Xa0L1cX1cHegv3WDI6yZZ0qJD1PsHjcw3Uc/yHqCwVz7ArEF+NGhfvnwH
K4Xs91NxAu/2uQbLb6kQPjFh+U+Dq6teBcQmtN0rfwEIUVV/bFI9r+rDaey88clJlRUJn/JokkPg
AtB9a3y/StLJVR7egN0boYiukKgaFuce8FczQuwZb+lPIyBOVAXUKZRiR17B+lsXhqzBN4pOoDX0
E2Z+MheT4ToEJvEmPLUE5pOPFavzeBgpjct6qjjILmYWYuJHCDadoeBuEgsw21eoCFQ9toWLlun8
RILRuGhhrVRBb7HdCicaUSUJ2HHMqUw1AGZL8UhjPUzdV/YffIK3VNtdqAtiLUc8oLq2pJeoSl85
UgYJ1VXTsnaQm/BvAErMs1Qs+V7ce0OgO7Arc1p+dRtKD9PRJFYACaYldA+x+sUkooTxZape193a
9KlZ2bBk0hz0yncfZHq4eehED65YtzfyjmF+Q4hJJIdNnlTq7CLrix/pJ29S4O60qlMEU10rUbSm
R1/sObeZYneaNtObgkSHdf8FHOt7jjMEDSJaAb7+P3ysT77tB0Hh8fVmVt9MHcBQUKuxhp1TV5Qq
F7lxRI0H+6JlgihLCXPmM9i/HI+arjjY5Yp2aGn3OSXS7HcVJzfEcG/X0DsbpcHq8lfpUoHzvH/E
0d60Uf5XOK0bbD3v1UiHX9cXAqBZ45ke/rRgXhxVovdgfNBKtvfMtJFVxTpqGXtUd2+dUZEIKjxH
PpOmt9L09t7u1mRdvvNm6jE19Webxb/4D13l6y2i6rpaoD+qJeNLvESGHfNWjYUFhxKLYZaUqghH
CNBSLYUUetyBbySTkluqkhjNFnxWdAM16Gfz6aHi7pinYfDNrWLcgrhavH3clS589RC8R1zcsMlw
sjfbBl3UsBatKb+HDSdQKfoLv+LoUJBrE86ktfaEvN6IXicr2+KNfPlc1g4PUxgxPUNXPchj5amg
FUAzdvqgOAyeBWkp7JnR3Uq6dE+hHLCmItq4EM8pExJvWpgZZrLquJMH0vQpgKpxszWF0HlQWNG1
Ptv1cNot8qV3HYZDaj8k1faHkI1PLOTZJZpxgdpUb2z3iuPMcCTpwSjqdd/YK8pouOriqTroJCUu
IbswA7EYpjR/tZD8KB9M6YDA1bJ75sKwu64psTh2avQnzEyusBN3vICsAKfjZ/WSKEK2WzARUgT+
KvN+yN+sAzfma9Hklt7br7nyAyIaae7NYrBUzmEUzhk6xN9EfXWIPDMlCLl+4GNSbFV1ikX49joF
kvtRupn+elCXB5HEcE2C6EuJ0EGvvpOs8n4ptClof6pLFZbS0Jd3L0QhwVXgThiODfoZO2zSZM84
0GtJlggdXt7NAZscsczgza1LiJV+6hhQsXpqxIKKQijSNhafFOMZ7zKGl+h4e2W0kzkvwEqiPWGR
Q6u10gNRT0SO8Jp/YlzYJBr/+bb21UaP/vYl32337ayWP1j5clD8bB88D0jzaxjRJgBvDwG2PpsV
OIU5279dCyJEzP7YCviFDcZQDtTxzQpacL0n4rptc+BMSaEKzrBwife+9tI6I2lMjL9uonJcnbDq
FuI3dGmpT7MYsED84UBjW4L68a1xZlLQ1hpYDW3pMyt3SdlrlJ50JPs/NiM5vaNj28o4eMLIl9pS
j2qlHLpHai+M9ianfz8DC8J776YNxC144slxPNLdZCnIVdEyUbdQ8yaOCIPDNdguqgv0XcHIcixR
XbZKP6CdD/9HFNRBbOe/R1C4AOCJErqaFeb98Bf+Rtvcaie87bxDoLMgCk9oJqB9HzT6DbDbNSGo
p28YzzOIOkYxURgHuOIbFTIWu2o2eKvSwSX17FHqJQtJCCqYWQ4OeootOS22giy/HtIjeH9D46li
OwDSUWrDEYBcp8Yp4jMU4PANX0PvIxn/RDvb0uLSQ1NBU+0xlVmypPtUDrKpUbbZ6gl2VN2tJ0i1
MrW6kzsHQC1PHXxBtYzHhiUfP56AFbIdAPyytLooMrS3kOGLqv4sGX0CuzvTH4Zn7naN2XQJl0uK
zlaFSHcIWKRqzNYDmwBH/6j7SBH5aBjpYzs7ApbJV6WieiNFsTR6QrpiDr4/wwg6VdrkY/WWyMQU
kPiQwJZsyj+U1GKeQYCdcsA/OG2kxZWwKXFqZug1OQDIf6ckjH4925HUi+B1htbnn6H9ob6UjE3L
q+41gI+Zt6ff5IwCemDmwTLUr2KyY+U6VzfqIdC5P7Td3H8Ta7tlwncB230d4p2o43WUfcWd2IFs
5knzz8/QPWBwfrgUTNymFJRYrqvv8/HYEI6FRhElyXahohjB8LJ8JubpR0RTmPGBQcoaN2f0sFxR
cJDIvTSNqNhQW+ieP+l0xPY9hg0yAlHyNJ5Q/X/qMTS0QF9S1mSwZXqDUiMM9DIOP77Pb0HgvRy5
GAV6VBgwP1dPK0J/QkOlTh8xGoZEWEDMcfT2kaghx3EBxUYfXShdsRDLI7HrrKd4qY9aRi6b9NBs
7k/+UMImO3EIlSVhI3HVXhiGm3ZfYnMrY8SjDHtVb67SFnq6KsSuymWu9iLg9RAwd7VcI82igNjF
SuCjmoLwcLK2f/vRSoOHzmlGQOYmRCGnAIy8s3EfW2ErtHYoU1Oca89ZP59TJhshZ+rPDsSCFzEX
r0PklEYjugvmdJEeKHX/n/B8MzkGfBMcJHySlQnod0XRVQp7h2RPxaM4zhdtQ65g8CHy7Tl9GLe0
kR3s5qgbrnkeJVmX54ybVFucYF4lP9yesqovPx5iXVMQRZGc3jkCTf//c/beKqP5BCmAM2OGzws/
c1AhMBt54DXJuwX7m598z0P4Zx7mkl8UIxiEBT5+/q75iSPns8gZ6CYTjaO/jROQhDn+nY5pF6wF
daoEq70qjzB3KpHVz+PrKY70faqz+10dcjNx9x4Uu6xkA7xcWwsUvmVn93/QNfgHP32/8O+aefZW
ppBj3XQyHusxIRXZrURtAEyCHfTQ9vY6/2gb7b4PlimDqHmdR/xloHUd0TymtcOMuyfUfSYGvigN
iutx3st1QERNbNvRrKUmOiX/BkG9usWOzLJplB7yIJPbs47xZvgISIKglmgkescSck5dIcLDIp9i
hwJ7Au8H6dFRfkpBNnivENEUBNbatj019P/KJRhzP0TezEUG8A7PEY2y4tIj8kjZOEAGiQR1bAZR
hZrFiHUfVboma4U8OF/wXJHpfm9wGrt8UMeKwfWMCK1eZAwZpD9SaON/uWUXb/QO3zugdYq0Yny+
rlZVjMyBDPEKsu1xN8lXzMQVB+hBamqX+yi6x5Vv7VQHcWrFUOu5cn5v92n6NryvMN1f/RpWjUCr
M93MwApisl7hIo5vtYU6lL2/JtyAjOKBfTRvL1YKbMl16I8ypzXM2JlxULC185ypJqJLG49lKAD8
ozs5YJnHlix7i7mLSwZtPzLclE3y5+J058RL49eQYrFHKgJJ7JxEmfui9Kh6fs3MLf/6i3WJAj3I
iE8b5DRT6DztCQBOOYw6/AMZEO1kAC0ABSDtzY8H2qNJSMXyKA/EoeLWoa6k/TdyJlcakKMPRX1o
EwWs8ZO/SvTA7OIZklPw7qmKrE+EHWcX1d6OakEdJdeCjdOGLKGP84eNWIF+YIyXiEqEUdGn8g7I
HPR13jnS2YU08bGerZ7ppYMlRcwquSl9DEVVQehszWKivap38omn22K2dIlkXuFI1Cl0Rmmwq82F
OfHeUXtj+MctoQL+Jj0k2MMEF4BbxoF0MZgfT0MPKB4C/UjpK/cYwv0I8GDv6qx1rJCuveHEQnVs
M5w3Wi3qRpawU2CRowk+ufZf2pG+QUXWfcuIWLtUpMvEHOGjCrqhPE3mqEWdvy8ezlpfFM+wMHEV
9AEYPrjH0+UpRbey/WFVlF/w5MZGTawJRCLbck3KFCuS9McpLePLe2Mzg9mCsNtudRkc2csuzNC5
cnmlQJ3dxD657ZdrmpRZFSjmt/yX7YYzVBNC7eqte+1ZmLKQQ3Zj8LnImsXO6DyvNHYbGU7Qfrmr
bgQiksH2x87LEnbtt5U3dPeUJqjjZa9DIOe1BcEmI6saRN9IzVXrpAEdpyCidVA4BvfFqfoCU7sO
c/t4bO5Y3/r4Ow+DIwfUq+TBDBqZ85Grhpcmlzm4OWyX+A10WOwqQhZKvq+FnWLmeNOwivqoCY7C
myym/geE59Kl7hD3tYXmtnMbMJowAy2pGpjJbLfSXu/twloEn3B6YMIgmpdf3lvQ+uEtclD5i+M5
vwSDi/L9OjKleARog7GYn4HyjMBBnlJLHICkD35NXBkv6xrF/A/IqFuNmsvsxwFp7TBj/1A4IqKj
fWpRvPaqmgQn4pQPEnnYaXi0AtrvgNkbcPhXWlIy7QyZpGL+wMLrDa9NFF0r0VzAqrx78ywCSt76
BBi0gRarQmZDImXW9KK7hs+Vz4O+tPrCH2IENr4HnGPRIVjA+qm6Yq0felsK0IXi5pVsg/ONnaqu
D9zxXZCPDmHYe5MnvAfODfKwbg1qLNU1CczM8C8MQPmYprAy9R1ZpD5IawMV+oaLMknQ/Hyfdo+D
TIlDZUcBgBrZrRXB2++UmT0flPSeqq8tKNvYdUMGyL/VuqVP9JlskK+cXN5YlIlmmHtaqGfrnQQI
fBP/4RH1gX8joReOd04nBi/K/ImhSDHiQRN8iAqtnBZIZrxKaZ4Bmjd+bBTek7ROovDCkUBsWLa9
VDEDlr0AOBnvEP6MKz2YbUuPJVvT9AG3Oul1xSF8kyH2IVISfhfr/MXTurWCGtNy05yLprvTXKFE
Qv66tpvZmKLXtZMPfHflH15MP38C38uDr+onan5nCIEgbAuNIfDYsowPEli3BydE/EUm8u+pH0Se
pDu0ltF+T7KErqHWbg7kPJ9ntyCpD+UtMlXhp5VY/uTxEdmYbEP63OMwBbx91Otqi3tO02vS0TQA
+z5nuu6xJdqx4H6cFkvOijrjlGtvXHbP31TYIaaxuR4/WLTuVGVkCsxdySVu+vnFElusTNi5KEFA
ZQmN669zqaxfiu/J7z2KBQKjUr1hU8PPxY3xBOOEtDToRNNPQzojL8kepriFWHVW4TqdeloX/3UL
czUlcHd2O4pPhU0/0JlbUiMVFGO0phDVoPYdttjn4XEYJ3EkWbxNktOcZ9i3eCjHGrc3wPk34ek8
3QGXFxKy37/mPGG8KuSEXywvlWTHSqOoRJ048Bb+lVp5erNHYX/kRTtv4SSJmVqA9PcLYn0tFxcU
ioFbS1+u4ZLmeYrf15k+fJQrtVkgVu/l3uoKVNAlNH13NQRKnbN9X0pBdwaJKbS4PcFjUFuBytVb
fDblOH455pdzAv7YIdJaSIqiYYJJn0eeiI7jPpmfPstUQTu6ENR2upv0royHgJTdDRL79HJr7JPK
gGz24TRJZRuwg0FOXe2KbuK7wTPTymrurv1VQMS1VGWlJG6aEQdOVFnz9Mlpe9MNXjy0m6r1DjGN
AeYHXBqSeQXNv2ilwkkj5zxpdsvTpRESQcrO9V6fJufaeJGFfbN27bl7gu/GSPkMazPAqlcveBsD
stZI7WX9Y+NZlDJsqTT0mRYHukMuH9IVYn3RgQv9ZffM8mi4UB7jPAFX9tPsw9QYwb7dfoFtRBZ5
nRdmK0M3whpUEG9L4XrrIo2CTY+CrESJArD/SC0kxDLN/zi0KEqzTIFAvr/ncHVyqHJXIRxl3oN0
MVDYAAV1uH7zU5RnLHPP3daIsr5sqJcGRmvkBeUQWCBuCUjEID26H4XN+nxemn2LlGAt04kaYS4N
KIVVMQ9litx80kCFOOYRjXSo/TisBToRv9k1Zc2L0ubcM4e5KaB30KThkza0WMp0lAOOJrYYfXk+
UnUcP3+Br3gzg5xCb3SR92quQ3Y7qF7O1hUj16K9FDfE2ZO6hHLevmoLtyhh169NVBwJ6gC3hm6O
zca7Uo6t8Iv6mh49xbAfrScOvlIV6vfXVIQ4bhz3ijXi0chZa5e/oyjNpZSBPQmZ5vK0gpRY7mll
A2FY+gVwYGfU/4lnJC4vGpdq15s3G+tC1yYGhs/QY/L+XGQmu1FBqEXkEG+kYOmGCLE4cyzOjUaj
+xsxs2iifsEJ44ZeQZ2Tfuis1GiGb7bdUeM/a1LcEKoRnUbffXQfUTaB5Z6Pd/6w3lNPkcYrW/dS
3Gaw/mVLb3WwRogdsmyR27NiYMqomcIO9MVIxnbtFnu2td5J3sPwbZWH8I9Z1QkUZ8syyzNoFlhC
ONvsk7yv8WnKT1HJhWgp+qkQE7EBf/sncIdrdLBtW7Bvy2qwRVBoA8zZJpl10FXU8fn6cMMatZBy
n4kf9vssX8AVa+i7aH3ugvYQYlwwZYSDKRkKzy96gFBhyFgvnAqFjTL+hBp3TtxSG5ZTiFJd7e0/
TeDJt/Z/+KoTtSa2ZU+UoIVuITZJjrjwwoqA1VNq+Rq6bAQEqQ11bSN8kPwF50bwre6OTCMJQz3/
S7y8rySayIYrKJuchfI/F8fQyFPuPS574o30K/K8VeuWoOsfZKn94ZFgexQSlsJfteYfghh+6e1q
SapsmzET5bJR46nFzkCECoE5OCtwgFpD9M9hsuyzoCcGbxyAlfp9Ow9ADYKL81lg2gI0CqzrGMc8
rSoB1LvFRUlaHuP7LgbSKVMwdgs1ivdjaCQLNdfzzVscpJzlIRoKgywmEBC6SzIPbBGkhz8FiXWh
7OUpZE41PRmyxdSB8iv77ZKXEdJyN1hWdKnN1GA9jalb2WfOeOxaq4oA55nxdTPL1KqWzQ2cqAla
ay1V3jHPg4ir01C/x1nfUDCY4D7G5tD2gmxLAbclcpt8VEzdBiDxXcbZugdEazhdGc6+opJJDSbb
PySkdqu5V65vzjPdvh/luRcWIRIkgrCpghZsnTP3VzkRggEYpmXFQw0wRanwdjxT2tYsWEIyUZly
G/mMYcG1iugJpRw+PwXtVOpQBYUxY3LF9pFddRo7SA2GFXfUUqaDfrRIb+64yz5Hy8PfTDV4XVda
S5/G3EbvGEXAzxdH5mC2TALx9CdIxlyhFDPHNiu4H4ep9FbgwCoMzFIcLCOcCFuIbvkJBh6m4JoG
vmzL691yO6SouG4Ysifw7LHAKJzxt+FJ4WeYMBq+4kK4fId2ZdP15E6vBQZ3AlBSoscA6QEIR50U
eegv8ZDXcLwHVufzClVq1zlZZb+b5aY70au7gHTNNSvhFL2t5YD8LSDcgAjyNpzksLDQMLp/QxtJ
tvqpPFRcVM8QQjy0IONd/3yWPx71FFz2/UhqouB1tYI13+N85AAJ97cFW8v1D7+/e9O2vWi4MUMd
/DhtZCFM8cZNPmG1FKvQs3pjgoyvxlEbuOK6mV+h6HvCIuW7K+pULtmFl4bK/UMC3FZLxbeSdWyc
5k5idmTp8WlO3b7E3CebQREhlRFmMXTv9uWX9e7TgknyD9SngQqIIXN9e4V1MVWkOgaXrZgLvxxP
4KzsfnmcyAhdV9rp/saUqqRu+JrzY9UVWr3OwOtSUP8ghzvontJMkzc5EzldNsk2Y3CEt2jfpVLN
N26yXzzKW8WEm3yemaw471lICRGd2fhExRHvcQAY4dz5A8I48rYfZLNkuvx+o+ZNs5BVR/NtO/Ur
ZbGfK5TdgnajCAVHobIpBKi3sCTD4o+0hWj6OYEQGPRbkasRDFuQG7vptl0RaoMxqyeNIk2WCKuX
PymNoRbO1OeCRwbqT18iRHUTWPbz2U5zq6INk1zdp23Su9HHQGdab+qrqR7B3d3pOvwIdcN+vAdm
1CLooTTcauSmqd+IrF5cTR+jTc99eg02YHUoCU8JYj8/dz2m8S255zOK981kgVlRWt2Jsf9uxE5Z
NwFcNL5Wznf6Bc0amXXIlwpk0O642gSvr45gjEYAczxEJSpGGYuyKW114UucwP5xK7onkZtp9VDh
VJtWXvDSanU+d1RgDLpLetyD9V1AB1Mtp7PKbh72QtyHTjRHCRDVuaXs7LISaLDXfIfBd1bp2w8e
ukfQlB5XmKvWQvFopEZfgOGAg+ZWMzYrnePVIZ6XdJoKI8pweq8u2sGPDpyO/w+xL8Y4pXuHuLso
Yk5n901aABeDqxkepH3xtIa5/PyQQHuAmnDuge0NGf9l20CwFzPpgNUmGnO3iTs026je3ueiUZVU
5b7b/4HlXS1DxhML9xsD46L18HaWN4ARKeMJSdRuQR1ss/UFh69fupl0gaB62j9B7iK1zWPzFr3J
9G+BK3Qgnft9b5cP7J2RGgto0SwXTlKiXQnikJy4dDaAW6Y1kx94sshHhK/iKWfqAPlgT7DX9Q/Y
mt0Gk4hV0AaCxJphltHPt3Zb9EL2RKCGAD2UISPeW1iR3MuPSi1Dceoxh+zB2OL7IxvrD3cWd2I1
T4IIFVjcxf2k9MuoOTyc4XKlE4IqUMmKNXfk65masNRbmNVE5SAF567yOQaM7tyu5WDBle4EfK6J
41bQFy2UZ9UAZGjiLQbkF4RMTgAby3fiYDgYwXJdK3jjq4SOqn08X00NrIFzq+75/jahZsZafKme
Uyoxci6rUnt9hgXJ8xJ+Bo7mM/vAx6+6J90mtg9Wt6IiGwrwtvvjvxxWh2/EzddAW4MLUEqjKx1I
MFj9IPsQ6QK9aoAudQrC/y+WHbrPLUN6t6Q2OpTG4Zb/od2IPKhhSKRiAS5mfSDWpY9uGgpGBVx5
N0H/bbQEx7rMmdteuHxLOgt0Xo4vdcY8zprM13+/0kN1hhOlwFoNUnslrCitUJre8RP/UfvxVIuZ
QPhDXpWJOiTOptT0fANMV6UYO3kqfQicfo4C9jVIaJbx0JVRWzrGShg5+L7RVnhL3dx6bQX9gVkY
gKKxod6zbif8h7til0husP8/5rB2IaJJCP2tZjykeug3zCSRJEhPl3y8prG1NEgOtGyVxaCOk5ak
7PA5WBi2Vo3/EvHUViuD2MZ4yMtCLW68N3e0dsJTBnt1yFxLLgEAISSr3mHHh4oSUeOMVNLISPUy
YjbPsciqadP0jMrNCcFCezSQrJReh9JSartXPXYIbMzpw0b9dbX2HiuBDc/A81ZslEWOo+ySKaib
Xf2hizxLTrDf97+CZZBdzBviXTQd0OW+I3LOLDM4mY0UBh5SqOlvNcztJLH+0gXZUL28UKdfIxHJ
iJOqlX33yph4ORq4PNYha4txmKKc6bxqpXThlz1N5brsL73BmNUQlqYyv5VcL4VMpaZ0KGkjBOSA
lUkWBn4xbvngTlwlKjln4HR4l+OCXgPo57mfbWuOaVFzmnCWFFvi+4yGr9A0Fg7fgsO95mHhAHkD
Vn5ZvYA1DoguY/sYwoeCVhw2QxM+aGGK4Wl6jxRGxl4AJUVtR20Y/rT0KQYCYL3sA8xwx7crvjdG
23LBK2ieeNhXJsOZ4CYr28GxY4IEBcrtqbWENjKAKPkCJHDou9mD8PFI4oFwPpzhFr1qWl12udbt
9KDL9fiWttioErPJ+430cWwj/iNUkULoN4Vch7Cg94kpA8Q47DGw0kVeQxaxN72eXsUGze2CNyMq
afMwoZBBTKPBJSI5qawmD6qsYuFCOVEqpddRgZFEFx9RpBwlCQEjPE9R4oFD2l34/pD1eQJQfYNJ
t4S3+U7fX0gvjba0l2+cfukKx5/9/iCTSEO3U06K4yAYMenqnqh4HKD2SwdbwRXjvNYpexHnjeb+
QMRHaHeki0OAZDIGIFl4XsMLEwBEVm6+8tko4tJApGjIAKrHNRIfKxL+e1ha2Woq7rfseUSslT7c
r5+2YOkcFnQUOZCzE5vjOhMxzf7o7KOr35OpaH1wt5/szxA8FSRCWqRDotijvOizM6cV/5Dec7uC
hNIw763vlbJhowIZI8dxLkoqCIeUNHrLwXn60osd6LUdgGbOtNO2BdyWoZdWgi60+G8M3Ecz+XMK
3dF69XZTCEjX5DmRiuBZFWfzfL/IDW/AIucPC8JR8N98oa6MdHI3kVqJGVAClQZ8we/kNwrZLW62
ilcdl35sPb724dyfkeg5IFwfnDjw9+SeuKZEkRq4zipKQ15540Xjf9hSuGi390qnFkOlnUaud0wn
5DSKj2xr2qjAGgSinWS0Rh3y4t5H/p1383ETWkWKkOwUWOWqE/k9LSPKb/3y9HkFRQitA1jc3Acc
PIgX6OSe+kvDrPvLUOFx962EUn80F69HAISP2apMDuiV4tjQSo8cxNFRb4cwS+Z8FLKM0rmd+7Zn
KNkqUynVmLoF1IXGQoQNGiUk5BaTnYMse6e7RTKMX7zgVuw3tr/eh8R9dRAZVYYqrT8u3gStMWRs
7tgE+F9gJRov0i4oRHav1Lx4yY3uqVKdRLHfk7Y5oVY3OU0JUzAYbF2CwEOArnm0Fu7dmyUYpb1a
52UPhZ+KdTdRRk/nSW5jsjCwjJU+8vF/naJSyMNdJoph1oqZV352S0R2Jvc7esWFWZT7r4I6KT+w
fJQB9dJQ956OalSePstu/4LhZoFZ2o/oBN8EhwoU8xJM3Bax/OMBF6zBHh2jHVN22P6tTigs5Dpq
clzu/XAVJTbSaDEuxnImFjIifD7PpWHFU5EXXQ1vmQg7FrFhbNAN2tB7I29RccV0POx+D9fLcWw0
YYs+Qp6P5SrRPG1lTx9DdbWRLL81KrFGGJkJOgV0utdYj8Ck16bjO1Eg4onyUx3n0kzdm1F/GOMc
g5kp+57Xt0rTNZDxHF32yzez8Y4GsgygDXaHnAnLmr+Wg2IU0MaJTu3+QhLtbk7sBTJdttWha+j2
LvhJ8DOlVUUTg/q4AuTr5k5vseHSpLqfSmNXqrC9tmG3L2/eBM3UA3dhzzGcKBWzDC798GAsMEZ5
6rMycjPFUmkYXJGmnzVXku0eA74a0i4WKnT2IUhmML/EltjP5MBI8/l0Z9s020U4uh3QhAfpiSBX
N2RkkoYEgEM4GCUk0QQLpC0q5EKa/m+SXe+bRiF7S2O/nNkboBsTMzUJU+Oe0qLQic+ckjEAn4sY
sOb2X08HFjpO8BmzVUi8FsN2ohgHqDC3JxQT1c9XgS3Qn5FjxCEur50+e7LkLcAnJEqJ29q6foPH
GZbp9QdBzy3eQG4PZIQPRkBLnfNZk9mR3wlQhZJsM2N6W9SAk6GJc9Od8q/pkCt+Oc/UJjjbECYw
pPBWMQJdvIKpYI3zP9yCEK64LgpUAS05OpxN0QBHliNGER4ug7oc9egDXPs7YXw5XB7uVwCjDPgY
x2B6CfmO4a6fjHvFQfNIJKXsIjmP5PkyyW6urdcIuIje2Bm34jxn4hVPiXAaTsPs0T+SZDe87BSG
VL1eMZ83/gShbdouhXjqd4dKlPBHUBvpSVa0LzcosCgS7oIhh1jxKF62SWXicjZd3q2iJmyc+2zk
G2Y9xHOjwltATCaSMGwnn4FvHaIZ/psJvT+r7ok7hoGvaSnn3tCtDZQxaHgqOslrbpThzlTQF9f7
LH+dnb3aqtThDHn+OPpC9CqV9GXaxewVQQzrNrSZV8BO+lyqouJmrlbczEZkt23tGtAVHsTdQWr2
3u16SR6gSgvInEnQDfJTI4Unkuy4Wz19z07sR2PXr2IUo78rQ0XRQgjBdiMzLiwa327mq5KGuHKJ
h2P9M8dHYhRqs4bMeVv0MUlNbHvVrPRRE1/02u4ePu7ZM9vBLRA7Uv63/ez8CrCejS9QkEH3E1Td
gqR4G+wtwJOqPB0JsLP/mUAlyaDpRjPD2alwFEynU+chz88k52jAJQ1DuSYtGgysjuvTp8LIHOjC
dNJTVXFl3voVuEHmo3yvM4AJlFl95Aaeh49UPPbBHRYopCtSHdi5UUsRzxROeY7rksNxlE6iE/K9
3H0+F4oxBrMqxyldc4ST53qYGBnSX3pN5rtz3Nqrtsr++rHjvNVMXcH4BlGIo5yUZa3ezqhWXnN0
zFFqCwxH/rKiJUPXhyiCLzAdxvddRvGSmcJtk9OLDxZOYXHYvQNmkICcjQZsj3+zsV25OUYO2PTP
iiJkuMMf8hfAqjDYA9E2JF64dpkBfI+Cl7nnLvBRxF+fFCuhBZDxQlWpfopPLGgqJTE+n7bhGicU
ApPuTZxK2mSaDkgGCS+GbQjwI3r/UDkVf/sAHliLeVPsMOf7fTAlPTMIOmXL58TbCSAePCPN3d/X
sqs6or4BQrdsQVcBO2bQGMiR50vHV6Y+V4Vd19mvfsFfYv0FapKkewQV8dMFmclc8ZSEp92PjAa1
4Z3svjMFapHqG6J8BFqyB2JOGv3Zk/+w9z1rME4aPVFZ/AQOrFuZQouCuUQBoBTrkExWSKdiEZ+C
J/1zoX09NvylCwhvHVoutbIdMlH7oe4qkis/H3bdzy3B1Qtxj1qGtWcxJuABGv6a0JNKlfN8JCAk
iqFBfLzPsgobPjBUODtCqNjtZ8Tpv04lkNI53iT1Ph3jy3pXvXB9kU2CLWHhU5KbD5gqrrS5wD4Y
jr5Pn1Va+/wiRZxvK35O0STNBh6lSJMGazb5g+ThRNQj5runL8CZdmRnrgbso73sHHGsJbRjCwnV
85brhctPquywsUq0DgMpXfHJG3qEaSeohJq2Qk/smwbM8xs/SxRTQj0flcOzXkRWHSaI03GiYah+
ts57FfOZMEeYinNVBb9UHTbkFmA5GAs6VyO+Q/o1t1DIVwj/BclqXF45Bv581KuzNYFrc8ymbNXQ
H9qrlYDAHoBHxt8uTKJtxvyFJYtM8N+xYhCrqlxGieo6NbUcJguWhPdcf8+FiWpMjSY+f6CWFO+O
JIu55+x7eFWJCH1DSUaRJkvWW9KKbR95Tdiot6axOXcS2eR72ELBebVT9r72m70fm7KDcHum1qBo
scTXYlWQ6npnLjTuSp2ZOp89uCMkTJcAxPJMNMEEJfV0Oxfnn+L0JZFSmqdsIeiKQBLh67uHohcG
wy9EnfyLXMG/sXY2BnGoM0QiUFBWRNqdP/Ae3cD5+070W+ieq2yIZTemwfGjcX3cSyC1if4SeUrs
6U4a4XuYinhheYRTL3TtpZyaZkN+7gnX2gZJAaYqnuLcfaQwLO3CqQvqAIRz21GJR8CqdqgwQ09r
UgB4rXD5hYPp5bbuDzNMnTu6kCJH7rarpTAXinzoNqZlYSzOtx+drodVH05pzZYB9JubMWh0lh7e
CLQQnKaQyW30nxhgu3900XfSoBU8v4MpgrNbc1Wq7EXO4WkccnpRMOc+hXx0YALIcC0Sc3LgMLWv
VcwCwaOQTJM1QoFF3QIUu1E3EF5UOsiYwwkwgNxBfQyZZXGoO6FZf+FZkQZCcuAZ5v+pPbxSldkk
WrymxjFp67by985LtgGPyvvdbUJPzvlHm3WYcgX/notX1siRZWCzzgwJUW9/Lnjk1ISUg79sOc20
TRCCu2+5WK387zBdWTP7ZCHuIBAxnxHoVLS6NAURU7Gj4yg4V+Bm23odqIQ9OVi8ZNN+yzTvTcqe
vNW9CXoDYF6G6F741dIG/cVybiAeNrgC/ECzNg+RZRcbRLBGYrs1+mmOBkaWVimJ/PLfSeBqmeLE
MJcY/phVXxrlNpA/T6hvpyerH7xSN/0PH3LOd5dDLlnRHNs9XnkSu2phakB/l+KKAfgj9pgd5ekG
s0Dqo0cdm5YZGqEevuuF1m6HT57MGLiwjUz/S36TTef0oyXSPmPYjqtKPb9uFpLPNS5CWrp+Dt5j
IDgBq1FDvoURA0QEw99hh9f+gHX017lAWKX9VyPZpFydKNoddCY8t1qBpMPkvEMwkQQbTccUm7oc
1MyCatPVHzVJr6MuOI3mbEHXdR9M3yWbp+qZgIwzXYNjWmLpFkODXfsCYANEULXjMfLmdBU3n/0s
gnjAybNQs2AuD8W9eNUmNjTN1MZm9aGPpVMJHAfVkYbD+HFDoK2KQXqA5lbPNCeKAyGD4YZViO7u
5wtkEFo/xGUrNXYbYqgP48c14DpRSbe8+wgXHEtgpzdocwnbM/zGKTDgIq6YVKCYQb+qY9yDw3a4
2G71ePwdUZ4GHDia5kkvsH6EPQdaVEORcAwmndoLVjYI/L0VwvsF8PXTgPd5aKyNBwuPm1tTN9Sp
4ETj821d7ETGFais6vD5LHP+1vFYNa7egzEkWjPLxUQp8sGtpW6LpWZwbwW8/EPvM5yTkli1/S5i
qBl1vBnQfQMvtC71+i5Hso2aPQiy+40RyM1UFOd8GTynjTmypxPBbMkuXA+vWzXnWEbZW3idmNo5
Lb/lwy1g/lu3TRr7YURuiBkMolP7/8aQ0RkRj5Qrt0tEL7jSUhE0G70rXrZGAbHNJSd0scPTJ5AT
CTtJtnCVr80Ob4ti3MS0bjVFfZIViyAnySjtfzchcJuMucthHgh2bb1ExOBDaZtmBq0iPwpy4wLI
Lx6CeZL8UyU3p6r8/pSzb48iKcDauDUJsaBE6V96J39bme2xFMNeB9NYR1muHXYMwhveiggej6Eo
kko6W/bah1dXgA4NBGcrWipgmsi7KzZnKhiGw+SFFifFQlNblie8nm2A1o6MqsuYvJm9RlpkVWdx
2QfXU5Ggg21IcXu3jeOg6OLPe4jlHR4cT+zfUtes/lXSLo4GvawZOedMqnqEd7ca0L1diXokl5df
U0VALKtgdQgu9XxARyfZ/dePlmzs/grJAXeyU3oTst6mwyVPeYeK6WyITMT9t6yj4fuVQglG9EIu
CQ8pvKSdcN8JzRrR2xXdMbYxrT6D9otYCWupjjL6RjktSSi0zPP1i6dTDbQ+aAqtpkvpA+VCOX8r
PFisdcEmPsCrBhlv4PIAK9/cguuE+smnhDtAchw/sP0gnqKnAes/ldaNulWv72srqFaLh4bEVRBQ
zpsnjBCrRViw+rGwHyQJP9p3cUaKo62NdxLcNqNEg5EMnuuPqkA5QOM9Mg59SS1cQNriwJjCVsLA
ZoLTqPvCoUzSxIEFPjsu/F+g5qvGh9haAYJpYhBVbZTIJX9/7bDMUNe78VL0NGaVgYOHjXdKHGy+
Vi5m815CGRBReV4dBi1/NwdB2sruJTa9OUDE74j3WpZI4O0pMkANbAm5H5GvoGocGYPKU4+YQgwd
iiNkzx1cGz+NhNHz86Vg0RjL/HRxrrpoGQi7yEXAUd3IQCVM9XafO4QVqk81sS/A4/Euqjw+A6VS
TVXybmZZbJWGwqWQ5W1SgJAtMdLwLKswUSVfEmJ+Kuei07sI62ReNxjDuu+oPaksGxGlHGwIboww
Uy9/UaiCbSNloQeJ3HFwxSREL6/THuhWgXxz+10pkWIta6kbqr4lkavs5Ec3sqswtKUBCe1G7EwX
wBI7Cyyi/kFatNgGAFdk30ZHC+bDwc4AsY7bujhc07h91/wewgzqX/poACA3Ho7zlXQPegRWudE0
ZfUXlWi1NvY5fEGfcQXsYw/3KDMQ2ox9XF+jMt0sfxqbYpHDdPHOiu/v6ywnZlUDRbOGFuBb/kay
8EWgt+KKlb5Mqk2xF4h6DtVW+ug0RhxILsXCVLRBGct+ScGibSXymf6J3poq4M01/niz2J1EW+QP
fsRkPFJbwPgUg2RY6/J6TLFcnzZ9AKWWhIRYmVlnfKOE2wAgxd+02LA22DggSdKZSGNjOvcotUii
H1cvDPLPCFZz24I9gpXwnlCYzy1IFx8eqqzY0+JDHaVppwqBX/PAxCufAcQ2MKxJl+hQv+gqy++e
qy5/usVvZJsznQ4At3i8cCfZGf/fnpf46NuszCn4rj+nKcQ1FZUqYevgPEl7idT+SqGs+Tmu7VC2
xGR6FamH+IFNqjaB9eiYe8P7k8ZFSnocTwvq+2N/DqtZ9h6qrb/UYuyNybaT1oLrjVd5pom39nxc
kKvsMruzv/hwKyeebe9eWbYYzca3pb+Z0o31w6sJygYJ+1wKpNN0dKkB5pqZWgCKshpETqUG+ymJ
XQu3SyUIq6Sgv4dBnfUjLmYq97jxEJ1rHVWQ5iOUnj9ECcYlC++JzR+SxEZRglbrUYMRqP0Nx7o5
qQWedhKqsPu4Kg0gEI0snCNo3pZrDWhgKuKco0UCox5mIKVCDGy7lX62nd6h4fRvdr7vqYwVM3qC
W/PvwpLTmP0C4u1FRDhPfoHLSMHnPKBZpvJJXdh+BBsjgDKtz+Ks8+C/qwE/NQr8K90tW7wKeQOa
znHhGmimjNxySVT7hfNbufAy7UXQKfAJq2AdppQZkzWwi3jnTTiGs2KufmBsJtK8+eC1NRAgxSUQ
K2I4bIUGeXOAqzN5V2nf8V6dYEB4FCNsuchqqHfHrN9EsXLE5YckTdpzs56f7oeacf+64RiXtnnP
RA/2R23wcWd1nab7JEjC5DC61XzD7q/r3gBTI4tVwnDcis8I/56MqCg12ppbdC22gGjlCzl2pDZB
i9KI8GOOmq5NDC4xC1jqZxKYLiaCm6nfPmihyCpefYdoKghGsWvQ31ZZQ+L3CLDqFSPgwXXUMjID
0yowKCFEmJxrabhBwLjXyRv6iowJJp64n+LSJy0XeOExPIWUPzX+IkC7l6mANRtScXFbEBUP03FZ
dJyCJYt6bXL0eibVNiMxyYr8zTWLrSBV2dpo1D/e0ziFvR6seS3HqEc5EUZ671U7/ylUmdP4wL9I
VteUJJjb3aBWof06n7Tq4tGIAYMBpYQFRGqPXiQPQGlzyARuSaMc1cNZsH/DYxTyVRQY4NOxIo0G
Vkg8pRDED+7YJmDrbPYmx4+IkIUV4OKgjVa5PoWzIsOIChRwy4qN4P636O3yXlNDh7PM+wy7r/pT
wQYGRBVRrcijF3bswKWXdrOWhLcwWykTVYcGu3yWmruZkg47Hl8H7Jrozlmj93U9aXsO1jDz3ms9
+Xbq98mDgZLFXOD3ARhpRYY7cCx+9wyt6OtIT25KLmcOSIEXvmUlRrgPtjmKkaE4EcdlHq6tek0L
DpcUI5a2uwlq8Gy9wfEAkHjgg0iGBybiscvX81W06pTKm+SOVkKgJokKNIR7joFvXKrLmvB/UC1U
P842hkC+2v3dMKQa+AyBVbFBDHSCG9+rt5+gCiRmoltbyvldvkCXmsAS40ezsE4uqcpMVa2QtECy
c8bSjVK9YzpB3yKgZgvhd8RuUN6RFnNYsAdZNs9HnSSqa73/WKvRhK7+cnB3grKpT9KgPURJciNl
80woZlDdmHqPZKad9TlvoVvSG6HEAxIDCw7vVRV+laLJhZ7iAuWwvczbPIIZ03qesedZPF8N/ro0
e2PnvgUFZx9nDX9+txv4XwD5kyU/I4QNurItYbfr9Ts/YW8YJmkjLfUT6ThwBC4YEjWWF3gTdTul
ATYuGZfyHREHrDzc451nb1gV30rzm/DbSQkbUfNYEeJEKnTxeaa1Fs+AYPWWfn61vEXCkO6CDUvu
67qaKsvjq0GfNXVukv8QrA34Jo/lba4mzOiveSmoj2KbsQlQPSAdw4hw/R46eWbJ4rp5gMEL0gML
dgdAF1iP2RC7YHbDOHn3KNrHQ7e6kcKEcm3+VFkwusfGu6VaPsvcg7ZxDLnQf7ZWZLunCpXQtRg2
BtQp8d1tt5mxFn5oZMOs2K6uwBs074+gIazYMWIl+RQy7KupjxpLC18rFCW9nESiztwBG+K/Yb7v
Q0Is8XOlSG8ErcHPpTBB/WBd4PChb+kDpE3keiNtjecvRdg6w/8dYw08x45SIpDoLiAPzQ3Fqfd6
k5D9OnwWnwI5cVpcFf3TwxqdAl8B4OTzXWT/DOaIiAXjLP/4fPwK8hCCwFIAHbsVpbQyQgq5Ehgn
tv3+uFmYPJO3zqoqbVjK+M0OmeH6iQF4zVHzh1p+gWQ5PKJu6oabsqYD1Lkhw5ekNA+jIbAV//0A
RlbvTFbZ75uuwZuP+0g02pyxz3VYbkfyRs4SQoaaekbbKxaoD4BqM4rU+3m8dF0UdyMEPse1yXCw
2jLeg0uRp7dPN/WILjbXCHBrHjZMRMf+QwX0LnWWNDlID4e4B51S0oifyy6apzvtxwXw5g7xTF8i
gqHsnAfDrAqd2NLF3pwrhXSKhdGkPg2zhes2p8PpI+0pdHGIB423Yj9iCXAcjyNPpzC+692xZh+T
Qn4/X6m8B3SaEXYa6ajBMD8V07LtpK8JcfXmf9k4p6iBmz3YP+fEftiZl8eqs9SBQYHWzDyYd1wW
2aV3TLFKJCZd1JLdZ1c53i0ABTNFOhKKLKAdijQxjKfHFyCgnIYJykHzC1qqfadHQDLeS4MKX/Cg
IyLIJbl/TKRB1/xurzyKIDg3z8ErLhTy3RQ2PWPo7C0E+bXq1o5RyLOHcbtPQGEgdBtHuLIisSlV
PuFBEhBxFokZT1qiS/ioxkjRru/QhbANzfmhpuqc//2YoRkcytiQJcyY3otIYDundsqHzDwi6rXf
x92lCtnWdhpqbmy4/mAvaVxp0VIiIhJFAHfQPQPrHTKrvTFliQBJ4vcZvRszIJ2r++V4Jo5oLoSX
7PklWEDXGhBg1Cx5UC+vrvDWH2kVEo8Nu0LmxVPzlpGBZxqBY1Y6+D36MzHIpAYoQa2qcBi7hl2x
ynLrPIKuZzJhimKL0m6z6xAHSo6VPvK7m7Zrq11sMEdLbQj12xYhz3Ih96vnb9wTdnLES1sdCosH
0ljPygPSETaTbjW+pFREOcCnrr5xzYv6qYV4RRyxVyOkXXUSvy52GC7RJKvrCxn9SpZiF4szDmxB
T+YY5jzd/QvotuF0BJfyl+bwTGdsIUaTsNXFcJCTKTRwbPyYVYcX7RM1obJuE1NxsHfhYuEazhQ1
3ZWBT/EQXnRn8dMHhyMC5mdmE5ygKqvWRSHo5UIm9q9V08FQ08pq5hgFPkwQnkwduo2LGBcOV7DL
Bm5l7+i652Xz2Siy4jivABRpUxlSsrzS0vg4LCySwXE+gHuJKJywPwLJbbmrANSNDiVK9E6908hw
qKUPCwu2QE/pW3oubkY5Qv22bmvx88G2OOW3pgiVFcQTRN3Yu/PYdTU4BmLSsMTdu/duq1OckHj3
2WeI+btkepbkxN8wEIJFf0tZT/tneOQ/WaB/1cvLKvX9AAgKYGmo8RQpzQwY+u6is2d8UYUOYkSv
sp1uDG7nQpQIVOc9jwojGwnRbBxWgwKygNUjfLmsTA+BOnOm6b+KZekB5LiNCQ+ck9OZwo+0dTAv
4Hy+UfKq5cF4YzQL9GOpR5D2a5cI9fwm4J0EbGPsjinVf8qrr+TtXltkaiApSYFdDxn6FGtp2vHI
x2AlqT/oNUHdT5K9ghMTP+y3MgUEIu0h6R+3JOTx4FsgKNVAgrhnmeNAUU7J7A8ujDOs16DZozfS
Hf/DXzK6QC+oZihGAmgOLE+cGBaZ+pplhl73uWocFTxpYby+H9RvFYhhGMmnNCdJWsRUyi4JBQKk
P30msYzDqBRJIgIB1wkM0WcI05L4dfM9n97vp45VNX0Qobz+PSIJ6r6vyZ+CZ79NQZDA51fjh+X8
T8L5rfLE5HX3XQoiOkiteYtCSh4C1dNGSTMDI7RCn1XzNrz9yWsCi8AxgRLYeLj8IRlT8zLUE7Rb
EXU5xe+sWqd0e8TxHGaJn6htgN9yDISTe5ijRqF9eRuDt/w+iWQ9DOYowqtEZIubn7r0AjRI9Qae
5W39X9Q7NdpjHdxUsJp4GRws+7fL+hCQz0uVsy+QY23XKAdkw86S95Q3oMwkarBvi59TlgRxyN5t
ocumXP7hmCvfus4IqNqHexOnSwR8dNQthh9kw96zI83xqfI1R/zlRB3QtcLfuVOXJOaWj4R6HlX3
iXN79Nu+JPuxU+kLZRirMrIL06HMaQFb30SiXI4kzFBKnLBcgFQT8NDgrHvPZqjVr7NB3Qpj+9f4
bCzrW940os/S/X4wM94+tlxbV53MphIgRkwA8QjG1xlmqfAg5CFFyYcOw0TukGSsoyzJzhkJvcI5
o8pNGrEEs8FWN/fzl8+WK5Ckt0HE2UhAulA+b79v7ckKYditgJtHf7zI9iAObCrYitzQPhMTdYxc
q3MEQQrHU73UM9N1IxRGLiZ751ECH1RCmP7EhlLr9VeYWigD7nNYOUnozjVAfRQlDDMjqgRV1YbR
Z2x2Qvs+YRmaFGO31JeDXeTZXJOqwJy314rKSMFayxlA4X3ZPerMhA5u59OSFC8ZN1vXbQp3VAw0
ZwBlae28rTOohXQsSPEwS0jvhLCcRfDKLiG+iN4KiZCw5th29DDag37Vo7VVzHO8i+ZY0kgGVRD5
cZSQOpLZstxZZ5CibJc20vPGljYMd2A3AScH5Sf2wc4OxPetJ276q/e6/RdzZym3Ua8VyQq+PC23
MGZ7DbLurcEmOYuPO5AHF8hCLWM0TFKYJWgWprHIEHZOV9pBJSLkvg5b/bwkdpHzt5J4+yzaTGnD
N6oH1B3GCZCYM4xfnzAkO//Z8VS4Ks6EGWOSJaP39NdIrvuyWkvYXPugtAZA5V2r82g9Kha/NeLT
1iUzn+f+Raavgo6fVFoUTBSdc1zSX1+8w2b1v3hzcyWbIZvDhrqz8xbrFsBuVaWryGWVyXcXgHEg
161s2zlOwgLDVNJsLCRYEmj9ohMdpoZuQR2vpFayM9izWCJR4d+94LFfiEOR+3B9Iw/Lj+B32GZZ
6qdVDzRBiPB+QCnuOLa/29JYnoY+3ch0+q5SKrED2mU0e9n4XwH2cKHHYeTdCu9oHj41I5yRk63g
Be/nMEfrUeQWbgL2rLbmp7Gw6l/cvSth4g3Cwex7A4LFkYD/I3xhwGoDSplibOjTAtk/9SHfGcxr
CMCXjnBnr1sJWnR9PB/PmbG/WAqx1OIi03UEauXWs6hc97k5MqAMLMTjf96YJl3J9or7nLciqU/l
10YUl3iIKA9K9MyHUhFSZ/WmzcbbCAmQi5vk1DTdKoTXNsR6KxqPYQK45vSIdusk0vuC58bb0qSV
zIcGDX3TF2gAdSyJjy0FN+zx8X7rdXWJSycPhNkB60Q1tZc5k3EedztAol7xDHNmhXhkea4znkzB
GQklKdbUMblx4rWOO7CN167obHB4UogkXoOobu+8mT+USguJTU09vR5nwG35qbJnQRUzz+2HX3aZ
GlK7YFwtLGOX4nmqw4WnrF84ot+20j8JHz4ggcmiJCXKOEPjbosbREMlD1Epwv2zNFy+figyzrBU
wa4Woq958aHJzKHIuzeS3whRmNrp3O3v5jaoU7jaPs7TcFtKvZa7mh0mtjBUe6JqEOy/wWs6WiXr
fV3HWpxYjQCW2n8zZBS8mS/pH98YpCk49XpzdvVSQp7pC7Si/Qj9EjuXnsyBUAUpUL/lLz6QixFF
h9dkj9fcV82cGe/fEkPPB24KbxgP4rNwjN/sy08qmyNNeaWYsTgmRcu7XfYd43zHAli2NeIMJR90
FAKfGffQ9lHPpizn26Td5nO+0sm6M7gi+AA5vpHurQRjzl4psSr5Jt2SvwIQY9Cte89uNsDncJcc
lml3+00zc9EAbcWfr2+e8ZheByFHQ4USkzOYjLjEyPNeAhmZBy15Z6+7MACPHTtwJh0zgACmHeRX
uFMdxD4m6rBxFdgno3FJ/SDnFK0f+iqygL9eB9yUhkYeg6nmRwmMgRO4ij2eGd/RAatfAk5bQIGT
6K6CyLtUhOr126Sfv7GyVg2h6pzgg0L/iEWJlgqrSM0KcPiNhmvXn56RYBGpGfOX8eDybyU81vA5
zjH1YgjwOvH47MnI9oK4r0NOwL5trsdk0Bxgn3DxwWWIxvp6dt2vejh5fqhj78GFRwHkQpaN0Ct5
0vx9sUfuPizPVm1XnEwLjn1oH/hxZGqyPz3zV3p6D9nJ++hrIGz3cjGgfMcJ7FPBzKYDEqY5yNoA
b6WWXFUl+TXJ+KhGrV4GFoPh15H8DKwoJl9wHkCLeod1HxLWi4wepR027Byo8e4jUbX/huXkFUcs
gxkfqUWuZqxJpFI2CjwapVDu65kmkNM/Aqj+HJdxFW6gjT10bZevkK/kQF5+4nYb80L54yy9JjzS
pK0nMJ90y7EpEUSCe98rBuBiZ65GNeoFd+Zp8UnSljdcjC6GTl3tMAIiPi6BfZEymTyjE+fyObyI
71O3KAWJTKgATiDjCIPI0ETJ8124ryo6NEHOz8H4X2TjKXwdwUZQWQjHjmDkEj4eJRLZ0/6padL+
lzuWY7UI3BpPVJD1IESLoc+ZfAjVWRvawXnAW3uuo+r4JpMaRBKRiLXo1OivN7rDxDlOLMtWNcLm
9BSABTrzbqFPZRWgs+eZkbbIvy2IIfE7rgXAK1UxVpUS0H9OnuyVneLzP1JSRyXG+rYkb6L/LmIx
A/hQgqSQjVYCvWlg83tQyI+KybVAqPlO6DPIfLufsZNNSXBpU7NtoliV9bRf8Yvgi+SUNGV7xvBU
zKEO9XWn4ruGKvt+UPvsj5mmxWOJPtIbyWavYCsMfwMSpvUGIQZNz+shfGwqUdVs1JAwEt7Vy/oa
ntmO7QnzZlttwRicFs19DWrdEmJuuZo3dtQpvRD9hDQJczPbddjDeMUErVxvlw8nN8yljFNu4O9e
r72itwDKBK1MkuTqk4hSDt1SI2QhT8iGVLEvgDxJNuwZYqsOg3Qkr/SfviHS1YcWTLyRbQFJ4uPG
c2OY6RyN4XlqP0kwLkzacVJDavxk86PtelhTVzgw+smYBfBuSlYGN+M/fjLBP8V1QmwsNx+wKoIj
n2c8bzIBHueg4ExzYGAqTZVsRWTIjJNebHFi/g3RyjiW0L0Pyr7iJalvxUU/ZKiU3Pc7u6Y4zdlM
poZq2eG7sBeW+VMHAb4XvssuP4JTz3Sp446+ODJENUMLqe3LoUQDZB7jr0xmNlufQWKNwnuEDtpp
hVKrt8fJ1i88caSRbowbK2LNG4BSaPm7M9LjeSW3jG8fW2Wb6UsvUcaA2SRAIk5cm1bqFvngocj3
5wSl4fmHGsW9FbUO57/KUt/pfQjED+V/0VweOuV6+hPgcWEC3TjCYTSLcC3dKh/1QPcy+2iyND6i
3lUr7p9n7bJtmIJSJVUQGQhF7DTthwaqlFwAjHM/i2C40GuTmB5DgQc1I5EtNygK0pEot/dhIK99
izz8JehFO9i6AokKCJYoRt71T9adW7+05aiY6ovr6coPTgmLr6uil40ilX5G7KwHDV+x7D5Axspy
kJff8D0mhrw892j5jDCrtblEmVhCzhpiWqSTx4lDR8HDGZ3DcklUwRHoSZ+yUmclwWHOu+zwe88X
Ien9yHFD45raHLkPNP8+FoiGMM/C5DnQtF7EpP4OLP13t/h1vlBQuy2h6Zj6ETnaeZqoR0xC1Nc8
i4b1KSzqzDTmfYolXm1CCy8OiiOCbGDML7CDPw+TeuhKZOq+7TI/CselPXviDrw/3AiV6CKEb5Fp
mlQ75JOXrGM3Y8PyFXFZyVfnQ09PurBXkL36xLSdfxOtgh+DaVGxw3FCuy+kdMBCxHXFpx8Sjct/
ynBnLVaaIg+J497B75mAKWfqMeEex4WcDC/hWun/0ArW8qoikASpI/H94huvGg9LoumzohM0z6d0
uEcYGYQ17DT/0fuarwRPpCf4wSLqExgET561VsgSfMLZi+/qrJpnT0kE4rgbIWTxmowSn4v8v+dX
yE5JCd4neQQmgmw6zqBj7soEgURf66cOJ5a7r2WaR54SWBtKMLBcNdwqvzNIZOaaOCVXwLapJbRQ
28xTwqkQ5iIQW9RTn/dzl2xHYnM0t0YwdhTYDM2gICg4pDH6vWE20WDD7MkKl27zq73DZqAy3HIc
mOYWUgjWx7tvvx1/GI70gVcywVIK1DTeoYzaNxtWWAf63PLqGeVahucs/w4e0xO8qxCBaFaG5j6f
JW98JPGks+c6HQz48nodflu1AGM3bIQd3OU0Vs2c25E7eDiNCWXUTxg35eFsNnxnMEzoN0Bff7Tc
t/7sBz9DgHrZvxFYRakudONso+8wapTcPCVzqLD/wTZ/PrZkJydzQrufpp6OWXzwefvBagXlfPbG
QVRCvlivsRMzwDwfxHZb4jd3E9CrQLAsFfzL0JZTCffLICoJeTiT6UvFMZ0RexX3b6p2pZ1wEpkF
Rh9qqGTJwhqrj5BaXYgaj4EWz/EqEQimxUpDrGSKvttPzFgYL4gQC96jt6dY8Y90vc/VK9wbQwdj
y5qyFoFoz3DghvidI7E62WrWprkcE7cslrkc/0f1AMoivhz8YJKVd6WKaEyNlG89ctu76mJdMukc
fK/ACRUJN/KJzNfUgY5Bq8el8tndwqw9iBJehy+AEqvicNR3HVCpFZpFtY2hZwMP+tgBDr9WAUzh
m0D36/GtH3NaT6PRgk0Nr/KYWAoM9hKscz9gD34r/3N+7SNV8Ul+QTSu644ZVkWVIQpVjwsekKDM
zkNI9Z2HlaTYbnnqeRmKmejtBl5rRUKsiXWjR3w8GiU37TkQZbRJT9Kw055mLe85ixOUDaXecSwp
qGUjF5jbQ6ttM2xncDGfK+xwzi6XKitJVx1lzDhN5gDa+REqeEWjipwtTpZ55hNnjENnHjaH3tX+
zHWNAmo3hBEG4g0RZuA1c5r65KvIaHiE0MnYyB+H2GkDAqhAjVH3dctJTC7NW58Gkkv9PD0RLC5i
4q5MPxUXvnr2FmQg9w30VKGyXy3bgXoJp6KSFCd+TVKnJq6+xjBn0oyTWSusuBFQue/jDqQWTHf4
zUxZfk8uRpvzmS21GlMRcZJnLm5/EcrX5fTYPs/2YIe7vzvcovmxsggbutHxSFuf7iDAn1FFyLl2
5OPnY1iM4JT2x+pzBDCqZ7dm/gXFUNgGHhnJyVMQCNS2KAbXxu7ZQhxm3SVf94P0cOHGdmo961W0
Soi7UQ1VyirQFgCmESNZ9LjbZy0znt7tl42yTBM2omXgsSEuebJLKA7lle6gIDgiNsARC6PDo6bY
vOKFEliI1Zs/4JHbXgCdfZV6zEMJ1UmUehpcnoYRdtA9I8+Qf3A4/MIE9PazMoNDJQdOdUxW+OML
RKsorGbndsnB2dc7Fx1JPMDy2QX/yBHf/lEfzF9fSHUAe8WP4jSiwclHfN2+fJbonFD6A8R9dwXR
s+olYJD+S6rd86IdZBBzgUdawDBjDpTKvUpu9G+3Bxcd5C7crdDIUIEtdddg8EOR1nbTCSSub4Sx
FR68CmgbJNXSuPoIL/GqCRyLyVsEanPNv+C/Cnm1Xdi0jW6MNQxrQRLmS16juEonoD4dWYuMWWAk
lvFTVeSO3Einp+04ar/S9Qy1aQ0OaX7YW3sRCESZ9ek4GIxxYNpQiiQntDrkV0ng18Q4xehXM66m
4atXw1QqkZmpBc8tAqVwdkBkkumKL4/sG/7wvdYq+9CFRtT+yOGaH/XsFZ6dDqyBHu2DhqtM/40K
2plXfdRt61xWL9nkMCMcxHJw0nyP5oD7Ixq5KphG88t+u+xHi1gwY1QBFa6zXWNgEFDEnN4CCe/0
5pAivqXCRgUuCiue36YRAQKD/d6BGb3aWy9/XfPLrO5bs6OQY5RWOJkDW92Mpe+FTRT1+UkGg/+U
Rm+ol2i/wSOkWpojStgcctRHqSWJmQLFJS61GJxD0BgHrumZivDeOh1+anhw1gJIgEPea+84d1a7
IJ3NWBxF9cBHlHnDdkBGwV7D5lFT4YEPp2DjxlUWhwF8XJiG3D54illAMwmPWhHyHesau3ZQMay7
FIn4DQrTyUG97QYHYIwGBeJ4sqAPodlLqnQs8jprQyBqfWgbt29IkK7soEBSNh+jrNxlQh6Xn4WH
AFdsAuS5kQmgXKrYRSRp3TRVapSQ6xwoZ4QDpcXg+6AonXSe9F/ZQ1tPwdPSvrgyWJAWKhPridVz
07G7olQSRlOFkVRraWn43L/8S5LhhromSoLhG/8T9kAkRw68COOsqHj7xlsPpxNvkY8MVbUWSK4i
mG2+NhAPCdGk+pb2kRSEacKbDo7Rivl2xTnftHv+i4tjypozGLGs/7t+XRUg6z1C7FcG1df9mnEL
c4yXMT6P6zp2fC5Fm0q4ZadwNqcPIAO5TKyFFlJ6UuKxcOORze2Dnf77X0uoWIaHU4F4fTJc4HK/
dy80pLxxHbCYF0r6ncifp4jmm+q3gOfLcDKchiNTZwuwWCtDGitU3NThxx4Pm/pzKeEIaS7wAbI0
Rx6nZPD5RQybt0CgS4PasTZCYrqq45cQQqnwhsqnLuZQ0IuTyxVSb2Yh0gpa6BPc9/bDk5qVca4+
4UwLkimIrby03S1LLr+0KT7fglmHZ6GEzvdQYmOl8mftPkVnGIIPGoSLuTGmDCJ6q3nV3fnvKrmm
2ibu/DTrOoadrV6BXok+iKLsgKBdnIRdAS15zjO7dCAuFk22o1UqrNei7dszs2jweoIK5hId8X/p
7Yl+4Ll5k6GVMyqWugd3zMjG1qFiJNncLySksQDB5gmD1rpRSQMpsapWBiJcEIyo+dymXomCw76H
AP1PMTvwAF5F828Aze07VV9DhPYh8C+y3Sly2j5LbFjsbPcCpEW6kDcZZDmNCqJstE1Tq01TlKaX
yZNoMHIzua6OhkeEA0CaDl7FBDIFOEFpeIeBkjkKAAMYDq6of92AVs6pJ931quQM3AVTOIQf6pjl
CtCazUzB4P6iTwMScSRinro5w0JpFDF6+C/2C/kzQhrWNSoGlG45kU/OLZT41zBmg7PMsD43+851
T6D/f3ttnKt5yF/liEbCnjXIEsdvbuf6fYetBW/PqrpqBZO81EJ8sO8uEqwhGzavI6pedWNrC/bG
emupSF/4XpJm9DK1FuWiWJ0PV+YtBNPBDAqy3H1LTj0UNQqADJQQxyshZIDqRsVe5BDzo9UUNVNi
wrpRsEAe/PKjjDY5pDFr2FrHVH/YNtC3FcPMHuFI25Co5fxI39rNc+Rvaz6gXIm46yGMLtYaWOxX
dKZ7LBP/3utFRP5eOI9APyedEzx0JjNH13wh9S7NBIb/1z8s9a/yycrZ6L72Fju91m9BPcjyhVEw
5w8qqCl4TZKWGQoykuDeUUn/Gx7fZ0Ol+Ib4rAaXwY5V/YG7fu62Cb6ee6o5psIKpivJ0AzoYjr0
E3w6QSF9aXzndz3UAi0W/AOvEhfmW8FLUydBEiLr8aq0vcpYHsQDvxJClKT1DoAqJrcRGoR/79g9
Je4TNOWEZwpL0Fp1Ot/OAKqHLYGxmn22UwU2IJXLZyaMEqOwkJvZr43+lHlRIAKS1nBqF2iptwZ4
Od+gx2l7XZmQfoMd1JHvunnitK9rekrl3EU1X4CZNMLc+WEQ6SApzFm6h1msJovGL0LmEe2piHWU
zhsJdG/XXwsexx2/77/s/axgrcz0RB1HnhT/5FF0VC3EGtXYJnZDkcC3rAhwptKUOTA1kqRmU9Xn
IjVAfKY+Na1VBEbEXOLd1cshfSuWx8A/jICuk2QEm1ZRpPHLY6xQmu7hWF4F+RUfVatSOTBGxje4
46xumZYihNmoYzTZucivdc3YKtNnF1auzE9KnxHcrhJ9HIo/KTXPC/9cbS3lpRb/SKG497zL9fHj
op3bY8LP5SbQUt5wVhPkIxHgIZvCyEkkvTFW4OXYP71HJUQlUh91H7VMTK8wwwW16hsutqTsR7bz
SLxGEiyV9r2XDB9JN48q97Abkk9MVRMVtF3A/wINKSgIn3uWuEjPX9M/kxxuqQXs6mp+XKO1behw
TZC+ZtoC8TA8wUqLeM8Gh3vReLpA42PSMQUfg/3NzWGrcFLn8DRwxgUzDH3AafoxfZDsBL99ikvY
Vdz9agSGpzXPgtIDfCmx5Y+4NVHfImQHulQtFBwwky54T7R6FPvKaxhRXB4DzJahlDatRtdYuHQk
xU37XOIBW+BSnVeNYiLCU523nvRW7Oe3om9EitP2A0O3FNd3OWlg2hbIyOJ0MysgHzK/8jk5X89r
sOXBd/9PxwVIqNmTZ1xczWZ98iKDaI5d6bqE6QYijSSs/F7jLFNvTqp9uEHrN+8i/S1yOtflJSrY
/6M07XRSvn2tNj4EY4OohTXjUv/YIN2yXAN2aNIqIJtorOAu23bqIRweT7XRLLCWBAv3FwIVGumI
WjoE+8BlSMkwb5OV15u22YisTGBm31gxCEbHrZh3SLRh5PYIL3fiG9uW7Gzrl3k7gi3vvDLUkbXk
DEHySoem5HD1msT59K8hLcp0FFhiPnjVH1YdG9VOTBnjSjHiKx38oJTrgWUU9z17jFwnU+Pp3QWQ
UqiRx5LLrUjON/DbJSuvWDQ+MasKHri4Oig3HKR+Rjup3Ds8BkgOR+v3itbFQr+EfprCtTmJqgkr
BttLNukXwFxRrNwGO78g1xHgM5uHaOl2lkp2zwqr4/bKzYzV/AHghkVLKdhxm0JbTiNToV0F2k/Z
oXz18P+7SB4yyQWXNKGnnaWEFO2fy/OVxktkzckduicjwFCSrCJVzFiIbkOkZIKgRk/8uouA8DbU
84PwvWzD97ZPNfhYZWBXvxMDtYP4APsR+9Tdz8KfIk8naOIya2SyPMStx2ZnozC3rX9jfyBd8+lO
ifjI0qF6AoqRAu+b9WCvllEuxeDfeNjHsFOsHjo5aG83eJvmOGiE8iGSRRlQbtRXbsOvlh/agUEj
w/iRm80dodP1mXuITmYM/ho8u8M2EpmC64yoxoDqW/zd3oDUU7cb3dn+yKv2CawcwmBmrTWWJFp9
1/qBeoCvqb2eCFLCP12l2dAgI++O16dOt7GfUR/0fjW+4lN535027KRtIju6n7CCc8r6qTuZT8iJ
AIqadjCkUgrmNX79K6XynB1MaP2bVALpXHZG5M0gAJDPxw9La9GSvNNjLdXMnlQtZZiJ04IZWaPg
t6A1iGysNBQbOOLOl0m9v17q5x0GZWR4QTK2UtJU2H/49Lt8ySFpyrsspd0ZtT6Ah0QR8Zzyrqjp
3WZIGKj1gSoQZC0HFnHRUH7SyLXhrzK7JAIWkTDMwaDg2f4HgMXW9fJHgizGzwUO8PYFfaaBBWzQ
Pm0lmhFlYqkZC7vKgk2njgJDn/0ZauwW1TX8FGSJqghMJYwwzhsZJ81HBHcaV9mGmWOHmg5nkxZe
MeLhJJwOUxQoz1z0Z9lH5KdGYOWuYfGL7z4Cm3c0pU7Mmw2IRRvT5If6yEpD9bn+O7+LYUwFzHia
wtPtN4x1tqIUiEpS6XuoJVN9PeNqFKbZbWDXlpx049zMT70wFbRZhQKoHL8EOZxYIDCYTqutmjq9
uE7bfd9acNQ0XRjP5Ust/LjQkVTNmXztmouY7P23DCPdtH+92K42aGrvf6N6lXr17vWrNN9rU+vL
GJp0MZLd3xOxzQbq9Xr3ttos4QfQFrDeVO8B7ybXfX3dX0lpugd+ZC6tTxAE8IoEkS0T6am26HKd
owltxGmklw7tkzCY1Zq8OwdJnjq/9WyzFjXdEPeeZQ7reLdd3pso0s0wNe2dIeq3KWxfd4JVQpPu
DtTVkRVO9MJ0efh3rtG0acmO6zzsQvKCLK1S4VtTt8fss77/xOhCfhcVfvPwM+pI72g1y6ayWW2v
pg7yxgZOCaDMdiTuQ80RIu6AshyIwzyuLLuMX/h9fISnpqFzN26I0eyFrpVrAtDoyNDl+BW0Vyrp
oWuPPtOTc6t3hvBRLqbNeVj11t/RSWgwPSdq48ZGs5X3tzcHGrzxJ2tc98YRBfKKqHRLgDG1ItLS
gyatzLD4obV/qo4cqJmCaDN4obEt4jLxynKCxdihUCqfQKxreYgx1lH2Cc7dNhM96uYizuEY3Vkz
qoWb44Uwd6ZZxNlB7/jb//BUahx7EG6YZJYHOltB0YF/1uOTXkg/CxEjaHe5XjVC2IsHUX4hV5Up
QDOtFAVplyECZ7VJPwdAFyjLUOcqRzhFNd4KZeKYpdf+1TrjxbI56Qpq2FZys7rZxz/kFX0wA9vX
p2j+FLAX2sYkr02GqRxo25Ge1L3R239AyUg+cPY2aezaKtxtNW8wP6+A7YjBLvYNEVzVEBWAtpl4
SrmfEx6efx4UGSnrm5PM9e/F4Oa3O4bdLPOMs3mPak+xgx12FlX/OkOs5gpFbfGhIZ4VQmWPGSmv
f1vSYewt6j8Bz0YTZQg5JDpr3O7m3ZpbuCrduuBY/oIc4NhDUxJM54GpvUt9UR6LQg6aFn+EYJiR
WaMjkzwhW3w2Mvq+kJ0ohSHlVjXVTVhOgFYSc+jwKZ+1DezhFmE6enECni+Av2fL3TzrTJyCetIq
dHqTpz30eWoiSxIGLU+QkWTpWgUxTaWZ4OX5ZnQ17TWpj9REcmFtHSoMVQYMpQa0xzG18s3qSAjF
jcF1tN3PrARBcnPCNAlAN5K/P/OnscLZWDU8i5YcNbmtn7b54knhUBWiN3Ie9j8DZ0ndUPk1wpNM
W4hWMDYtaE1QKF2K7DW5Os4Bq+XJ8HyaWjaEVdG1VoW8ek4ee6bF55PbKZ11KBkp0yU6p3dVLEgP
+CFA8RuSy1qXjbFz4wjHvmz/0dWCoXjhF/NYHgl+DW8MJ1F652mWG2WYq3O40xgmEDt6LiWRBQy0
fDiYMF5swSKKglQHAEzhH14TFMoZOuo8997FzJOftvEYOVAqFpY3aK+E5Vm+iu3/Xx7aeTZdh4lS
dKINAflTG3WAz0jJ0stKdIzDi9ZRZSPnnX4/rRMREkymzckXknl3kQrGmZ90RqfFUKYHA61RRm5b
Mmot4tHFYI6ov+YgNi3d5h/F/1je6Q5qVN8Gl15ymSad2BDNOnCJ4WenMvAioZQoODCJuX5mppV/
z2wdaMceyz8/Ikv38rVFqpROeurGiJTshQQX6Gy3bUdAsrAuynXSxtJv8bewevD0tzGTZtgo3qqw
RtNpE3wIPZ8QSyVoBxKw7mnC90OVsN35QmoVih+jKEMkFV3hGoabXyojkUWKu1wGnDyfb9Tv6E/G
D0nJkA9pH7TKySgLTze/JrSKJdQLABedEaK5DKs6Rf1Q/kCi607mQQ0H29li6zwvb5CW5ZWN4Xu/
K6JfUc9E41gfJeOx/X05aSuobTrV61WgIFgK0YHrV0aytit/3BM33nfp7atd9jc09fbOW0l+qGyU
zZfoip/JOHLDaVpBOpSQFl8Spnu7mLCGGL6Ylhi3YX/Xgt+L7n+EJp3FNYaY4N43U8mc91QQO2vy
ATYbRqybff6Bx5QBHo8eFJkeg8kf8MSzZ60EbJnBitZzjfmFGeZVcUr8NUJlRz88eTJ3ld1WUa7+
IrjBpZhzsy4WiQ3Pp9Qu8DUoKepBDQ+LGR1xO4C2xRcmYfPMAIVe7e2iKnIXgYpE/Goybm2mSQ6L
4buiOoNWAh/w608bJD5k/SDJ0npLNAH7F2zgrTKfc+aVjkbx8gh2OmaF4VnEsja/YAhO0xmsgP0n
SxBf/9E4Y9qnfYzbh8WQMQJSafOe09g+1piS2UtSfR7QZdNeh1ciUkEqjjnnpQaxCAAU+z/V4eZN
Klce01VELqHS6T2Y9xEK//22seqtjksb25sUWiUYuCHJvejed2hbsS0VS0oXfiuZigL4FS9aWjw2
/D2Xky/lC1NLV0JnjOiubPGiyYTRwJ3t6Rnyo48ibsd5vGRHAv9YZlm9iBlvUGZbSLwiXzw5GHxT
4z6aVCTqY3+TPdQfiDcuOm/0mFfaVxdNYx7VSJvCuDX+E+Qqvmcg17wG+Z4UbL7ej8TfZNmiaHLm
BYssBdimXArRtuA6spD9Ju5eiQ8hmxP8k48A9C0NavhlooW51A6aoPWidFT0q1C5tkX/wHbC4FXQ
9kL4QxkfnxhL2yv0jnDvpAU6dJEfRALxCkS6iVa99ncgHHcE3kEKPfQDQlrotqbIZOiiEQ4Ecc9K
52H9Guyhk+gV6R+vjETgHhar5yB0hSNVsmz9WEzad7kxa0Xe06hPTfXeIICJLLjRImDHSqv8Gp4F
4G2ajChMb07DtrF7cetPg6rGIjqBfjVpuJwA52TnrQJnsJorgqISe1ld0HIyh0qQSm11+dl1uAyG
zsSDQJepol+kZtgRYx/x6EsmjerpmCDxVp5fOX8zs3OE5qLRp89DtDmjAoYq2GAPr7dQ+5/U9rMB
fkYSbbRlVleu0oMyZznCT/5VgKCjZoIKtY1732JQbdZNktoRlWAQo0T7kdreFY8ltCMzTRqq+Ce9
KPHtj5EBdyf/MO1oRMRpEj3N5TpmJwFCFTKU1DBBorUxr/7ls/o8V2EX9rjJVozFNRrKzg9RQHHx
xfeVYz0d9hOptMgzXGn1yzn+8WWSn9N63RgsdqbxLEZUe7HysN3Bxn8RIP0BaAFKWGow8wdCWMWm
AqUOqBf7+JK/GW6KfKosJCBQVIUU/yS6mYtx33U8FEJAHXIAb6l4E0Ou8xA7I2xdf1xdyQ71bJ34
ePiKfTMFQYnIUU95+VUZQq6fgTZK7RvpwxkL02F2tGS9oGBBewDr2orf/isJVakiGqgQDUCc5X7y
5cTppCp5cKRctcyIMig+WDLDNnGNuxbg4Cju76IBsW3WHqjQQIz2RWw/ljg31VatHRsYyA71hF5H
5IgZfYiDzLQgY4PgSUXuXSANLQT2hX7mCjbNUrqQ1DcC3wDDLdfq8mQcQbvF+lnqGuqK6Y4/JX+/
P8klcHxNkIzr1u0ss/wTy5ymZBNsNuTdCMJM3ujBhU9kWPR9nin1HdEnv2CKWNGzSh0UEzIneLzo
GYvhqvfM5zs7BIyXwTwDh5n5EXyCdcJPp/nGRIjTLq+GaI6JWYJ9UDQF+rM0kMixDVAHVMOfbTQV
EK6BaW5kO5tvoPeulRudJBs1Cw0BMAVawyJ7mZ7VFDjfcI76+SO6vfDlLTaM12paE7D5YWpx0gd+
2GU//JJPlIUfTQsF/hett9kXNMkNTVysUuUrbfkrAPF8F+VUPvgAM8C4xX31ofyrwTbI1qi9XKbc
hNohv7lohtxSajbeXg4ezCfW1fTX0zaCnlRIONSh8oYNVA95P156ZRCaru05xWs0dqbMwZ5FTCAJ
U0D2fu1fAVTc29CJyShp8bffQcFVow4cdGQ7qVvSYiHQR/m4I9x5VsqVp89PMrEszXvssSHTfGTX
ImUgR3uZhcZsEib4JOwz50TKDzvhDG9Hc4dzYUL2dMg6+ECB8jzB+Xt6K7nmpLLZeVGBvq7/O+eR
BLg/bjIUKWdXQqpX9ItqgopYxEmO+52yscdKg6m0qvhnKYjfp8vaNgIHXcVXo3TaPgYCS6OlO3ch
jUIJblcjmjY4ntVfLfpKNiGs3o3aCxz9c7hyNv1RXlJCvc0TKn5DO1LZQhypKL4M7t2d4lJY7nOi
hrhrZwJz0uPKGTr8O2hQUUako7QAqrJ5wSIktsExj/JfbsYpzDY5TYqBfEUzKCzTmWFvhkVp+7MS
6uK8H8pW9tQh4B5fWq09qeV2KTaU9d9Sp2flBzEs7m25Yet/A9LrIHYHpb3C8nTkEHjcbKZ1BHK3
XnqMLyARuuhPwEsh7cMT4twBj7xlMGshzsTbMUgl9wDnw5l4Jiuzb8tlQtwTXjC0GyCX0Zu2D1yD
PqQOsb2kfozzkJ7blVG/q/UGa4hBwowBlAgrDv+ctXk/zptVZ2nM3cvp2JThGSZntBzQXlEZ/yiI
zeicXLei98y0IM+vns9Tp5XU8IvVJBz7bfplLImm2SlGQi75GKhFl8DTqqxRjI5kfh9+IVk+1DcY
FKhCajPDnxAEYo0kCskbLS7EqfPBM/+QYJ5MHddJ0SzIv0i79cFCDfdr7Pm6ZQzjo5+qedlQ0fMC
nqFaq1K4aEfFwrTpVy+7GQ6vsw43OHnOA65ibStiC6jIHB+Z4jcnWRbJPZZK3lnhAcCQCIk0wDGD
yIJL7o/dgso4R7gBG5BcWZSc5ROzT3pBQ9PsABaW5nP2X2WoxHskTLN3EBaUE4MANbmozrBNE6+l
l53234ZHqEiA4Lbn5bYZWjpLc6yZ5q+x3yE5kksrGHkx+UkqSVh6ZytNFfS/Ug0Hyo6G6R7VuU1H
NRiJkyJ8N7qxiVo/taJoTo4PrvaU2yFxU5l3TxOPj9IEf+juqLq1taGBVtCYkqz2bCgFHXXWzbCD
I5uk/NWfGqxEczjctgSZ4Frtm0aoCO0Ok1qPOaYLYSEyPFCSdCN5Lwm1FRQJ2A/xXpzJRm+gNJQ1
tZhfzAepOXQC5rbu1Mpk6gYXo11LDtAsTS8mvL4iWNobKbrWy2fNGUqItsyXp2q/JOrFnB+Rd3nU
psGpd+Mctfz49pPPsyy33zS/39A5zoN0CDB10X+8MrN0wciwrICNJ3mulwz8fExjGNDjJKvgkl9d
54eG6t4xmLzKnZAgatyh8Yu/Dvza5GthIsr8zZ/W1CCaXLdT0SFarcPqLaZfbWrUr3VwgydSYFc2
2w5iRLWwKvhLyJcqTwyFmCMRQ/AEuK+F3pd9kG11OkfM+4/J33Fy89V/t4xYz/nFwHo3IUw304rB
a3b3eaSaPPQyFBwyo+vRCKDRDFZV+RcJ/eqoPxjvEoo+/YjuQRQNyOyp0UNV9bdcP2T215qzAVYC
kozscuwEn2xLTaveZAm1dMqpwx+vOVwD2ZLArcf31imA++04hDIovVxc1Mhzoho5TX195/QNy3CS
FOtWxFEj1z/JtA32ZK1cyhWIB9SFydWVa+Rl1qq/KYrE1nGNGFtZNUawTcd+n3ixFaj9CR2CIGz5
tKybj3F5p3ktXVuq0U6M1MxEb1zJRIf4qZLMdeSVxOtGRdbfLKbHygPXCUchKZz9L5TfLpn+UhtY
X3l/8f7Zuj8fMAsJiL/Y6PUxD6lcIqrJDC/rLDK9CikzPPjauJLrlWEPdj2C1io9a0a4h3G8mP7O
6QMFoDVfU2NVkyz9lQZ/ec6nE5FHt55z0AyVYLV0f6kpXnwG0A+rPFlpVJrm3gohAyJBGZozUG2s
Fs9eGo0mv3vZlxpoUg5f1WC8u2B9TTdnaxHrNXsgLMMYrM1CdzlclWEHioNBFJIXwMWe5nS70qB2
3I/0Q6mjY7331jtBb/pDOnM87uol1X0gGTRCNsE3Gr233OMnC8A464NO5S2UsebMv/xnj7w7N/eD
eX6FfNi2HbwtDebCpzf35FFq27hITBxqSLSUan4XSS75g4sCBdW8CL7MIAic82w+YkEVeKTvsns7
KWbtQlF10XJFlgRfZ/cmwqJXK+70SGIRH2XnYS362uQNe/eBco2ZGKiTBsRlmKx1uHc8Bvto5Wdg
6BtFxLsEm2K0fE1Le5Sgul4FK0Yune22rnLrBs2oADkewdZ/nnpdtvIke9FF7jeHeIlRIBMOw5KK
0h0nhF5amaowmqJ/hrB0rtqs60fTo9JMXJALAanokhIfnhqgGKdq0tMMvTKA9H2g3keEqvgniPcT
WX9cDLX+wEDtrWCY0nTs61GM0ENZLQYA/WsY+DWPb8E4zOixREvoJmNafpplodl8WhC6kOj2I+Q9
vmXA1PUfMDgRr856CXIYbFqhZYXiiw8BZn7woHU0Lwyyr7IPusqKojDnWIZAglbPXGugzeUzNI9D
HtfaP1TjEggkQiVDYExqhUgV9pHhHaoEr8vpI7X6FhKVHtAq4BY4h7kFuDs4j0m6t3si7rl1SnHP
OGpqyVePc3hXcHOpCeCixkNNbW3NwJjjsrOlsoT1hHl+BSmkyhmx2/OL3/wt2+rYAVD8ZkMpSn9d
DdlbKfutxopVnE/6nZI0t88UuoYVcvBSf4kkjZhHkLBfhWIOqwbEtSQpPHr4mjE/j2zXvWRBI+d9
q24SEbq8TjZnNwUp8WWFqwr5cjd+PbqYL1lTimCjfwlRp+04esQLONRyNykP0ccKFno+z+4J3KKg
KTYnorj8o20R7l1BaXvd2T/5ircFEcwrSzaH+MOm2/TjCI8Pxkr+QLjWe+NaouGyPDENc8JhQUI/
qe6j2RCsIiEuIoX/UL+lVevSo7RGNf6LkcI4nQxf2myi8T0VaKb9yGZhnH4WaLA6WGSqS/asUq8L
DJmOKIOYrD5vRWXjFO5MQS9F2F0Koqebjc4PRXfGYDg2VzBvNyHFcniuzYX16Q1OIK45Rl9DJoh3
wvbvEZRXd2iVh+OcBOdAAFtpga9xkeXJNPzs6IOAM6YTEuwNDuDAG5y9jwH3XTipuuy3MghgQGRE
4vefy/p3taCe9wCx4ZMpKB5Q2mId2s0d2uGUh6jAchCgBj9xVbte0I8+HhNsDpyEPZ15YSOd/P1v
Hyq3rOhyxB4KANNY+anaopvoz3n80swMwtIVQyS67TqZPSrHguxyLEEUwo38uPxrvYLLqfOsQsy8
DLK861ZOWYQ6W4zqAD+E1h84//LxkZgRY6m7xATaJWL3346WdqRfWP1Vy1diuN7J+xtJ6dNhkp0t
UBwJ6CHO8MCv9nrU/2z86RVL53fst+slCQfEDw81oTWbBqfmNFOISqZfX4a/NojbjKdXXi1qxVhr
Apq0BuD5J0EGQEeRDJiWtTGHDOfPBroiMc7uVYqTZ3+qzJlRq1Dgr28OFVgBayvPKNWpCPW2md2r
ESAJWdJ2WFq05mw79PdVgPAOPUoFTDqrQWzRE19hK+lI92/jPnq+lwa2jzXr1a8RZZdpptl0sTKf
Szk5FSD21d+qubcJohqhyzTaIKNHlQF5r8ar5PIS1VUTZFshc/zBvP1eQgETGtY01izUD2JlcnnK
xlPtCRshPF4Qz1wyXafDNOdjN1fcqvXWvnvipg7N31zcohlJ3uGxyxa9Ekap94aRQbIMXf+l2JRB
kAYaMvv2/YoIwCNOq2spqopSXD/QIVMGzohf/VXm+NompRDx5hvoJjwxhdZcy9Hzk4zvKMM8CWos
hCd6Vmq7o59GnY6KbY7Ste70mMJGML7R9aKtFxbFFM5Gja+aU6CpqKpbkPVHW6DhuVKG6n5kRdMa
woOmwGw9va3YjhH2bFSUCzD4ZNAYAiHcGK1n/Mes8qZzirOTT2qBmf4eIqUFNVmsIzHpf6EY17m0
rrU52JOOo0GtzhxuN5mD2Y9DSMzZbdGjT8sIAiXXFiHgjlTENuGz2pdHtRtZRswOwkXdQyZoReyU
oki0CsqXlR/kzPkFGFAfJMpVHvTYqS2D4ZcPtQUJQVWSyiWpV8U4whJQAduKvfGzFcYjSvu++9zB
ape7Qg0o4ux3Q1RUsjnv//6uQ9uVmIc2pq13u5XvJDanHZKCoJTv/cRqpWF/2PuZAmBenvu6c4lU
rZiZBD2PWaVnFqhSDBK2L/0wAdRXLBxsJPSOAMKZBZD0P8B8V7Ogi7n7eemHvsnY2VX2QNTAx1ZU
518SbSxlGG7pCMaw1NpnMO89reqHwqxzwxCmxENkyiQNkS/ezb3jyYa7CPIraOWEoKi7MwnzBPOu
XPVNJ/uvRDOT4Wud8gAioMKz9vPWbmtaGw9m0yd2A+K7i7ImoX1SPjkUwvw80sIMBwyDpXWmlErM
RNJ06m5Z7FvpkNxY9vb4vypf/eYSaz45BT+7yQIytHNvXgSw3aKAtlWV3erUYVeBqHNddcguuiC5
6WS4RGm67q4VDKpPYXN5E0DaecDo0g3d1g/pxgDGapMdJgrah8Fu7X6hSJwHzj7q+HYv6L9Qo3pT
2XT+7QNIW8OnKEeNAcAFVhk+4Xuqa/4lbfFHhRsuI/OeUSLoeZrcK09Um36sAH1Hnv582TbiKyf2
GLze4uXaqrkXCtzvpW8Y8opYcHqSUB/vsV7G/0QUt1MY5lWbvI7YRbQ7wBmfIhCCek0ybyw51E54
0U5afJNbR0uHUF/ZfNsiJ9saaUXb+OXUr8CSsVN2jI5KqGYAnkwZ1QQAi4qrJezBBiE23HLSZT9n
DgCrShu2ngi8/4ZHsBKm0PwPiBHNNxunglPk1TfFXrNHMsTqVVoxNX0ltKQ4qBwFi7mAOLIIEKkV
tm6hXCcn1dLEMQnxe0XGNUmTcFgSB0Hnu1aidH2wesI+TJq56Eh4LYXypu1SyHK/WsQfG+btOzXG
ulGR9PdLFx7L5xIWkCFjHJGBvIo1nX4CeK741bb0VhC9dSdDt+1FzuZibIFvlBRl2OWQ/h1jLfy5
mncF/+jhXWaLhQAnSjicE7vpepP6LrZUXdmaz2Urk9j7xtHCq5Odj/kyDEh2xL12bAwH7a/eYsjd
RFEMhju/T9hjVhdp+ubwM5CO+HgGRM+Nl/u2vvgnRs2svjnODCiZ+NmSK11BMpUscgv22pD4R5sc
5IwqoUUfYZ/odUI+Vts3stRSvVxIbXC0+zLKK9atRFq4hJe0axk4eMsdZokZnCpogZmOQD8fUSED
gOR8mNyTp3u/i67+31PMYMmc9KE6WepvMUm7KloYL7V3y0WCbT9OOrDPUGi6ItcopA1MEy50JIXB
gnMLPpItUcdutfcOtDZdOTNMINBCazf9CinrCu1BPOVJ1BPa0PxLVJ50uMET0qQ+7ntTzriD3dcf
ITtY3zAJZnxUBfbUW85hDdIND4h81tXKTlQZu4cY4vce0FI/ncqAGUQshnGGX84gPKF8CIX98Uak
5qQJ0VNGp/M91iLR/uIlWYFLQAiA/8wRVf7e/DHHSIAtUvKDxrqQyOXbGipIXx7Z/1ryKlT0c2o3
ydDG6dmWaBmqRQPBbYJ/jNVP5Ps8gkL4vFp+HlmAD9y6lriXipEOP7bO3GitoDQbRgoyQvZz7AMO
EA8jGu1JQRBwkZHdenw7Eycjbc4dGAlKZhHf+zapnB0+Vcg4vkyyy4OKFZjRGy3ccvoRlLdAOLfy
CY+px0AP+iOKWJ5wbHYdr5pdBbc16Jz7ykgau0KXyq1FrEVS4oVLdMuuA3vc4FST0D0h1gRPFtuc
SkQjc8tqiCw+lIsy2eXZXSOq0P29rTv40e7GdH/Yy8WVRYoEqcsCSMqZeu51wQoeBOAQouMOYgDZ
Br4voCIKBxVcgKto+R+mNcSpqoR9Z9RINVxZ5NaZEDFhxZGwq0g3EtUAWoow4aNyiEEN57lmBTON
dqWcg0rYYtNxakRHbAYzMdOkDdl194E+kMJz4OT15Gh6vzLAs0aGZNov8ynQNvaFoW11rhMrN2q9
j8Gk01FN6H4zmWGt2vjQiStTSl+Y2BQyasm58IMVBZCF994OuweUufQjUQ7XXsOM5EQLbLUtoSKW
bVtBck50U5YwcEXEMiEnk4WHC2FwvKBQSxWvs5BsgTIgkc4VfwfyVuh3tpyYAkeR8tqn8eJf7MuE
PMusaKln2Okm1h0reAn5c5LghPX1xl917NDOl93SsfGVX1J0pAosQ4QnsKoSsbzNuXBZxEYBhY0L
NHJaw0yEmcA6eGO44hit4b+WqHfN3d0aWaU2HbpbhVhWJjdKgPYN4wM7GlZiKscYXHcMKOgtAj/y
p/iF2wrEDWZDDkAGU+GkZiDTqnvG2Dxj7ruTnobPSofv49qDaDQooU2Rdnia6Y/igm4NCiOevSHo
s/127+B3UMJsteNVBBt3BYuXHuTeOtzx9nzzoj1mOEWW/F+Pml9OITsv/cOQuXzUYaHnMVlOFiiU
c+g5bXQ3ZVvESkXfZnS7FUGbzIbK9K110B8RHWoK40DHwNTNl16LQfhqCrNQWkDAtjZnEb64miZ1
lqaZeYfAaTJg7snyK1DEx1PGhDMK+q6gG8tBbVcTcgiaihvQt7sapZGiQ8pXb2F0Z1n3ZXSLhga8
4AtPZhzaWopakF3ZAUwqykDc3DQQqyRYzIpy4OjCuqCijwOmfFI56c3i0foVJ5o8P+HEMR5lfm7d
apHgdw6zx4uNn9LALmRBLaPe+CZUBc2yVXF6Dp799beZ3zTlN55261WRaWxNoYmREnc5m49xJmSa
svs8vkfy+JZpFKmf+CypRbThUCfTSweVmnA8g9x3MjrRCEfe2bFuOgQxNB/wHrf5GhObeMpPT/lV
a98D1umuqg5x7IxMJA92Gvzsa/+KwtM/7O24bpt66UDeMKTYEV8fwLgbuqBQMadt3Xk8m0ROFatJ
IjUAkqaraEILQZQryJBZTmd23USyIOaZmHQ2RuDGwWDOM1ZyGhqKUpdmFIg3jhz9IN5VERgURhQJ
uBnR7yMMVjpqozGydeTFIWm7DHJRYdhu5R4AP6A+pWNbG42P1duvYULgtB7vB2atKhC3rEDF8rbL
c+m+70YD7CalkBvbrcZJccY5g5IvhamUew2EJLg2sPWG3m23P7UrRNch7tW3fQMFsDKWfbp+O00d
Kg2O98P8T7T2x0pNC53+G5eMtJQeGO1ZQP/wFHXFWsbEvXHsLT6AfnCPcStIAC604YV2lgSeeNBR
jCRn8X18nW0qFsEaLseRBMhqRLNXkuHWJ066CRSuGSQ/CrC5jsDvbbOceka3fipNUoJawg4WK34w
26itEdd3xDwZjb59Y0Sh8HsdDGQZMRnARBAMREMa8BkxiLW7hQL8+we/jsskx0qm0H1uTkgj/ixR
hJt05B6SpJQj5lzMTPUVWC2d/fGBqMURn7K56g3CQBfLEZ53eRGbzNDRE3/zHQO8emKPxEkBaTbt
c6OPWN+XATROqEu0YKOrn0P3XnKDbQJ2f557OXf28dafbfGCIjOEMLakwHMHfKoT14oTGWoVwP0f
lTIiRiQBJwuLMcxLhYiqDHiwkbFHsQLNX99ry3apZwx6yQBv+fZllWSDqMHdvWqtRq+8Gqer/Lmb
SonwqfYRDEoxDCZENttQa9dLMyDeulHju3OeSSLwVMFWsy6ldPJueDpzfqPGz8q+r44nrbl3stgn
BFteHmb8iGMvHPo6uw9Hh5t+vTztzmLVBVgxAAICqhxrncHLlfkmgrhdGejb2ijqeNGL3wd5j+SA
5YdYmgPcZPkBg5/saPKG8XrWu02tQp/KLqo0lB6PiYbFdXo2ysJAOuBIhjSn1phEAkPovXnDqV5m
HQnh8/Nb6rtdYgRNgjrsSXlGglamZVqzJS1qmqG5xVte7EfX/ikTBZNkzJEQjWjF9DkbGBGB5zOb
lK8FIRj3cjNr6lj1u0vijvSpmaj/bdhVBy2FhQN3C8g0xe150Q978gyHXf9nFto+RxTuo5bOjnp1
+RHWxWunDmBZk3FpDkzQiUa3y+SvbrIl9dj4cjG/doQybiHR8MLct+Z+foPxoFPCQcDuU1DJ876Z
4q7gBqShEub3WyOTerKuZK9k1Q72BM5wn9q7/i+pZ5Vh4jCJc3J65xpG69OmBQCVNgzhjuRBAL8Y
+E+ZAFBpBQRY0UAvLI6oY4AGRml2TR7GmAx4C/2s9HNskLLCh48VEN7vdpKxZSI27c1Ry9oODkJo
SB11survX9U7z6BYeoBUNMSLcpe0gWyCTOFxW/r3d3PhBw/Y4NXYWIs2YjmtiLshr06Olpw2j0vN
DPIRWMfjDb+ChMxEmUnjFEGBYugPmEMnRk5giPFCyTBGmRZtwEvXWYrgU1HV4CCGbZVMilMg73L4
BKgBcoQ5Lxtfs+LZAMQ9WnssvIY4skcqYBYUKX0yL9xUi6tKpm14NIrJgF6Bn2Qf4phS/DJhBQG/
yCnQDa0ns8LMlTiJCRP3C0XNlbL9qheKW99Nn94OZZq+PCeyztE0kv4gHyxrUZpr5oqXtb7CysJo
BOJ8aoemst2acYl25TErQKS1qcVkJx8hgTNuZsRF3b73+Mp4A2oxuJHnmntmbcZzwD/BvpCJ4Rwv
LSTLnlxATy2HiBX8mnJlUo3Yrs1PTVA15C+aH8RLN3g66UutKOTxwixrNqSDxRpq7/tg/fN7uevi
e3X0dXVv9V8AXhoN5gI8HinofCYleB/Z2oIfdjbU93QEirydmpYl7rXHenKxbAyQsEc7UyebnRna
Eout09m4yurossYLeY+pBnYV5VbSGbrqotYZ+7jMXTdwVa5uvgJQwPwNMAdCW7L6M6+obmMwKgw7
hRdlwHPw/T0ws5xLkwV2hk13Od2SiWgzqcr2uSSiOjpsrJObFrz1u1fCfVuHrEVw1daLkE4MDZKn
rLWo5e25dlQ8FY0+FwLu8UzPJBADD9ZTVp3XD4vrYKMfz3TgL0fsDutTqRLckQ0WVItwL61MCv4o
C33k8VZuzf5S+0q9CqnelgcQRITscThJpyCIT41R2jVhRaYXWMF2Po0IsXVhxXEA5QTg7SvgTjAI
rS9FX1XwQbueSBjq7jgkcRYUAJXEumn6Djq4wSP/MuYT4TPqy274zM9Rb7/BMI5H8Ge38OD3FzYs
wPeUOHIs/6RInX9Y9GAFzvPOhU60HXkEhN4JW7sRoEP7KFtkXmfjzDzv+b1UFKbWtpmh27ZhJI3d
qWY975V3Of6RdG0lu9r8eMM6blUB08KwYd4QkDARMu9fcq0q5v7f3MrnB8yHQQ2W2GkEgwtGuI7M
t3mNw1fl1hAOnwYKwrpxvlvM5KrEd+G9uWDPnM5ngbo03yQloWF1g//ak2KT2l1THN0dAfABRt4t
oqu+LgwMTk4ObavqKZj5S1IDBooB90IoHNyCOyq9ULfNhtS8ZGkC58UPpINsoRJLXoINLZJz4mYd
26UqkXk29TcF55/Dl1+xNgVxgppp3WWLbuL/Ykp3sUAl8HimiSJA0DG/B0PkSuGSkWd4cmU+MvMb
KaTcqnPcY2Lfe9ZD2+Tm3W9YCJKw83kK2yhzMD1rzxaFla9W/IYImnCuwhGAsQ3daJrtNltvtSC4
apFFPOdyCIsqxD5aCSnktp5DlQLf6dQ6aizFUHGsoaqtrU+x4T+s11CMSU03jnKjdeA3mBSu5l19
+zvl6jjO4sALl5o/tWHdiTixd6rMKUwag4J2gaXKphCefG4FaDDDcgTO0bhvwBVRryf/PoYb0gEz
/qHZys4J+iHnLOS2DqWH75sBPF8uZxlwhMzkUtZDB/Il5tZ3u9uRth/UhFF9lItrO0lAgDzeoij/
WMcr0GACRhm+BoXq7mMEc3FkNT67nIloq/9FbLBthQG+zEsidvkT4zxEex00Q3h16+YWu7DdoBgK
KioPwxq1FzcmmaVfbPAHDzzctT103MUMVOFuMsw/w+YhW3qDB8pntFmyPoRrRdwIDxy9XZto8Ny2
fz58DQXQWtlo1VBo9drz7Yat1HgfT/6FD0V79XlFIUMvr1LU/cqX3pSOlmOJwkijNw0A6hYIp8JR
10tYnSgcf9WWg2bNAS3pXH43swvd4NEJSl7PjGHR3VAlXRSIEHzPNcXP8QKZHjuohju/Nsq0hDUe
q6dQEHZ4MzoSnDPjSG5qYFwRfRc2qsiCPaQFLSCo0rLi81wTJMtq7NwsVJL+JmHZlKzvPiERqUCp
AkISM32bfLUk7yPBf9RHa0jTEmxA0CRiggSX82rHFsx6UmQmG8XFGyrQyYAgxSTyKitqlIP14hdI
B8qDFmUX29Ws8LkjregGRgUd7wdsTpATsIE8ZtwLs2ER0SuBDDWXMQhUpaBGGS3R3qYI2qPc+S98
1dqiejStb7hE9FcHAV07RfHn8+E48NsgpTsy3urIozHpo0c2ZxZQxyrvme0Ahr4VmAB/KlAAHsa8
fdrEcPajRx0ovnouPalk2hftAJo1EJKpdLtlvKCO9j+2v033wqVYzhOOaa0lyGIzCzk8qEz6fK1d
Sl+bBaFd28rcwkZy0nBF09xFhpij6zpqk1SoQhJ8uO7C9VHQAIAB3diTsm/0JCLCydK3Gsm2CCXJ
OjNvQSo50zOuyNECyLpPOS442tnL40m/eVxbw8lv3BDDB6RYyKVSJi+DgwRus4tq6zYBCt4RgFo/
sPTK8HePfvnVXr19Y0nhLrUvvaV13O3W04QwiBaR28tg07GEt6CQChptLCezVOhSIgMpwWWYSZhM
NdtxMBbbjF7pTk2U4yKWr6fW29fftE74AG0kPQz+vI5P9PaFXSzLibiarLsVnGSx6gTQXUaGC2aM
RQ4+XmYWquD8h8jcYRyVkERCch9RmOQBwEUjrxd5mM0QDYiuuTTKyH8gjg/gqHfl0OXUrF9N5gcx
EVNPP3dk7zMX8v2rdxUZq2JM3U8AnovONOUqtWN3JJriUMgb1dml0SEnXqYQUP4lMEpDJdqgF2Hv
lDBa5ubp2tRmMPKZpP2NehTUVE/tAHQ9Gt8cakJRNTf25/QVSulrwIyRyQgC6rQ+mLANwSHF36lB
0UAplpF6RYpC0a3k2RbhN/A4adWip3++1H5F0JF2mCQXugu3PwzJa8/AvZ116iYb4RNnnpUzJICC
Qn9MIO93WDCnWNM/LEzCHkRJ/hXzoQc/+9pjGJX07JhkdTR3CIsVHFjl4F6Nl6QCaLocBk/7hN5G
DQbpq2rUg984Hqpu943q1UL4fwPs+KhrPo8kAPu6Z5rec662vFSS+4GPY68ROAqlvjmNCveUYdqW
Ykp8lFi2XgyBx5Z1WDubMXICdPhCPNxEoIt3lfaBA63IV5WFtjfDlC00PhpPOhspUlShbDG2Rbl2
nRjD0cDH0+7NOts5+lXECVqgtEjEn3rNNb9u5gyeUGfcS5GA7kU4kB5w8KojWWF4C98hMfNxQtXp
KdpQpXdVgwYdExzMaN4kFXGnePpBQR+eu192gpq5OZr93r7bGlPTkCdj4LyytNC69W8sK20U7kSI
1+TQCoK0Hj6rRG6A0/ErECWKNcdRN9mCMuEhQvmXG8gnE8w9QN7PZYnOYOJBXJf/zF2Qj8cLZ6WH
nsNZjzUWa0M2QUP1tmqEJAPF8dPkzmpkW27f7Fj5NwQzy8hZWHACJS4Kd4bQKYIlFGfm3RUjaRV+
KVsrK7Lwf/ZfeGeDIBGVc+PR02sRb8AdxduCZKiMwuhOoojV1Rj+4ht/7kZdSPkabXGe7GnsFASK
IRwcYVV1t0BH97U+A3n+aWZjb3DxxD7/6kNZijp7aXBMx8Ot28hoAMs3uVTiaOyiFZ6DWPa2m7sV
JAthAN9J7TRl7q4XfQVatajfJMYZN6KqN4u2MuhZr5smZITTPUk5wpaDuv2pOxc7EXjx2QZxJ85B
QYfP1qHjqCDPfUvO2r1O6vOpLb+0D2S8KQ2VIAEqZ4+2kt/9qQUtg8lmomgIDfKG5FaUwuKrc8KO
stZZlTv6dtjin8KXLdwl/bnW+setXTtgfoR38KqbbenO3C84zk+e3cvRtokFXbwYK1449I82Hcjp
cPwG1UcPslo8zS9dBy0NhRXNqmzMdjZ1FXM3T+q3dhDzy1uDFFeK9kg3rAv6DphiyzZXHwmYAgRY
bvlb5i1C/oNsUb7lR5C73ftmo+m0H81GvnmdEtH7x3TlwLrgChV7Xn6VP4uq7UBpZHE1zA2H3RCw
qDnPq02m8BcCs+Ysp0ADseUlJcUdKJ5sUU07KJ+DvK0lkGQVBbo/KWgPoysmX13WCseL0IoYtRQ9
TL+G8dqvV8kh2j0q/ejPBBWn3p4qHNAYPhfQyhAc/3ajmKgXBM6dM/0g/jlVTpnoZhuyHcTaYlW2
HR786z42rIgQt4U7t3cb325sqsWSD/NvYvskM3InRy0iodAyUkdSilH6m6BtF1WVMI/bcykvHCNG
bNLJCFItX1PBY0gT+YkdshgspL+OvtZMyMSGBTQ86ORL73LvzK9Dmlt887n//uuDba8jrQOOzFvA
NbMPKDOQyuGADLQsjMlcMQwaM8iFm1n8rOWVCBYuxGc6WppGvGcY4KfZVbDWM8PClUDBmClpUmJk
uddWxh0r2KUPDsHYxr2bH22/9abpkeCahWoN/+Im6ZLiDI8DRTs3X/mWcGE0ivEdrak/SxJp+SBG
VehDE368Cw4Q3dTofUZlu89l+o33NrHgk5W+5Uh+qcqk4B+epiYGdTTW3k45YwJPWUmzh/A2CRPO
3EBB68EjesJYdJqU6LSkecnEPP7dwDtN/yRNDdKXsEF4wFd7my/EFNBS6D3KKa9PEgR/7T3gMpH4
79WuZ+KFyOODlF0oiWcUWk2+hrG+GvB0nKK2LgWx7lnZyinUXM0Jq3Plejda0E+YEkPdwe5j3IKc
m0efQNwBn7uNQCPq28Us1wz+SKUj1ZCuv86Mdl/LfQ+6zmHHUN5b/cIb6LXn4I6j1fmbzAUKvWpK
/vFJwqauBgFXIwKmP7nHIafOduVjrScC5/gSEBrWklD0W1fczEjUnXGA2gmXcohKTC1l16qcZpla
wEd6+dffLMC1eFctPdPjud3cG0KE25us60OMHGaKp5NNFp89D2ikckbXbr6F/R214uQkpDtke2Wr
ATTbCJK0BGoLsR95O5BkpuFyH1AFNSoi79MIqwWvEcXnoU7VlHfdavxu4ikvhaXhEeUqGwZbyAc1
Z0D3Q24cMz0M74FlXg8tRcAEzMvkfh+j9AVzmPWeZNnBRifvYzjJ2WI/JaEEYNkW1HQUcr0PIhVv
GxkNeap9XUJlS5mhM0Y9CrPDM06PIJ2ESTGFdfkeASqxn2NmOc/o+oPPtUmb+5glwlJQwepseGO9
iUg+JDO/0vKVL7MPCMtJhtPazHHbzQgARK7FY3Hadl8OfZdq1+IA9dOFCC0m9/219GWBmqVtwtJh
trq8SLgnVRXpkP2xJpQ0rJfPTi6gmt/ikVfzJXWikdvdkbJD3jmJNQR2kqfKXNqkOKWm9gczIfFP
K2860QNtgLTYr65CGK9l6YxAonkkfdvz9JoLjJGTgEC/p2cTaj9mhbDVrhzWGsY4chogaip3magB
lgyTylSJ8OfDL/5fCZ+Pmde0W1NP8emIArTse59JLEco/24kk490lTKCbv/EzdhGmk4l5OMH3eBO
LZMBd3gKjhPiWMb9+mDfK6QEz+tfR6vkbfB9tnuEyFNiwUcLqP8tMip8DMv5aaOObDxA4+0zu6a3
Fs6vle6l7VLKOrDoNbHlNS7aFp7w5I7w/L4KWf8v2xEMGtmnaJPI16TG+JvTfr2t2F9VJQXe7dNn
YXSuh0sT+d+SIDt8wDSMKP78UzXoE7G14wD5Q83aLXLk2G7MYVuEpkJvt2s5uWsiVB4q9zNXoptH
PWeAipBPfkppRW4gU7VrWM6nj6gDh3s4V8Ourmb0ERmN3dVoTRuQIiMIKBh57jfmQCt2NaJCbI4l
bWdNLV33rSb5Ha8qGRU+iE2R+BmuDcAIUm3prnuu8VLuOsjEwQEyw5Hgfs65WRNledPNEfgkN6GN
LeF1KZRY30UYmXqdheBEEblFcRTIktMRnfwKgoaILH6F4pmvfouYUUvLz0+sNZ3hjquXZNMC9vWq
1DfsFcC8qqIDk8LJbn5TYj04geX/rDbvdWQ45enJG2wrmoD5EYI5Z3m/1jOMzLeFheh3VpJ4SMat
p8+PCsVRUFAGduMTCHFXLo28PRVJIsaeD1/MmbeRQAWNNg8aecQoVqjX8lTRjSv/ADR79Xbm92KV
LDQeNP1DrWUokW9JCqXmJb0YF+t+wFlFGeyk3G+czIKgeFKMvBZRfjfaWlPfLCEH2KZ9dcnkhD01
k+9p1i2nKH3CN9JYah8GieTC0GqGq1S+u4e3m9zh13AGQQOMvroq0UKq1vsV+XsScGaH3iUc5qux
ck5/ErJKTMzNJspHY5vqjy5M1kIDw4eSp0u+bWmIvaH1koQtNDPv5ovUyB3OAeY9BrsXeXSL39P0
bAl6zqJzgOL/n2XylzuH16lcZEAdLlVMqYL9/25Y0y4wYlhGQiuRXiJKD9f0JEb5yrAPZiAYsJWD
vv9AwXVjerIrK/rJcyE7TE+X1Drnyno5aCpFRVZKz3Dta565q/PMQr45PbKgqeF4GzkS/cuYZ2Im
APFinfmBwcwyWHtJPedvF2SCsftNXeKLge/KIu8fhUWeZujxyMxHFWUu4F8TACq28q6LuexMiAMa
nSBSwNQdqyWEbAr+z/ANe7Q6zNx08xFfcq2WruSPIsCaPl7IxrvS0/A+KEWeYowIVbY/bok7uNkW
FzpLA+e95f/hucuJjYJwYtPh70KkCnLSCw5i4OYauaiU51QW2Hj3lLlNNRmZxGP9OKSRGt6grfmD
8EHhJXGQehZ9NM3pzFnQCfH2R4gmqy7MAf05I4cIbQa7gnItKm8bTL5s0u3peZavAKo3jYCjVkKG
TgZ3WZqAyWe/Av+e9/ktmuJP6jR4D4zHtthPqbyPF6V3uoJJmD7iQAe7pVCNzgeJcWOHMN7OZynG
+NhkViaI97kh4yRRO+oxLFh26XFCqbFt3l9dW/1A68yA0ZB73BotVOO6i0QSgTKm/FFvgE8v4vw3
pWeKgoPO2Cgs/AqOzvUxmRmAVTaihsGXMVjYIaDaCV/4JsuRi41CqMKO9KexshVcunvEftWiNhBF
rRgf8aT55e3EJ8dJKiszjgHIsur1Gb52ljRl/SOEoGn9O8FBQkcK9kufF5ywPXwh+rpoDnhj0OQQ
cLbKvXzhYLYuZopG1yuCU1s+vRzVzi9nMSdPuF54rtyJaWnQKbxLO27kFV4T5YuZ2pWjI+du6V6F
BWi4p0kabYLdBD99e4qYNS2EfTcIFIcY4i2mlcTXDWlEpQJYj+UsLyoeRjNdzT/SJmOFMuYUd+J3
+cW5qoPuQ8QL+J9wu57FAVN4YJJdcRSsLfZFLAFHoHoWy4G9ZGs5kNdberTcSOVcEvTX52FFDgWC
4axinx4eUWysyK7jp6OJ5HgXozPsZAYexSRjxeZAC5GhskAAA1FA74ftO3bGPyJBQCra32RfAazq
Tg6lI90lnsbNEqsMQZfNEJORoJtOngja6aQYHxy41/ijGcaXcGqZbsKkLpOc5hc32QXWAeXsKSA4
OtHXuOCD6tGYJ9e3knQ++364opB5mfiL905S9Ku3+7KT0YrN0ZC+zhSt1ujzJq2hCw0YUaiZj8zA
CKw8GU5JFSNlbX4632am+uUJX0gzVD5Wy8gdvtzOSBfn8D4q7z2HUaFWuxb1xvEziS2eb6XTFGEX
HbyU184CTr3ZJTqaBs1GjNK8knuc/bI8XduMISnB4vKZ0yH3pXbmJg7+rukFAOJEoHmD2iaySxdy
Oce7VCtCImpRR6O6P4TDim4JQabFpvOVnGk6SnPD6oZ5JTggivwtO0cWVPWVbI/GplOEqHHcoWbM
GuDmKhNEOiYjRNcRj/nJCqQ8Gc8OKqonTIbrrynRmTjFzvNoTkFoKcHbu1KaknKcDOubKyP/YMbJ
NPw0caqRQ6GkyNO2m2WY1lNRKv2gVf36FxOd0/uWtrT2cANhNSRZGr3d9hDozVIH6yOS2Q89cpYk
kqHj0954BDgteF4XhD95/juXTYy+EYuxa5y24gFn7yRoZHLMuynp3PVrtvSJHvvY91ZOk/6crc3p
xdNgAC39vN/7p2TOM0w3BBpyjT8oz2YBYoiACLJkqnD6Aj5Csg9ZTuKHm8mniIMrYqpicKWBxst3
f9jD/jE9wBznyk+j1CddkKEtobgZeOuHTseeYu5hMaKVp4iaP9X0/AhKFZecPMA0EwHAHV8fBfWh
wNHDm0pmURoyYTs4+Ct+mgrudpb0JGLf1ZT1I2MKs5BnXe22C9qIPKOXpwoI5UlbumOoWNtkPBwd
K5jhtWrbWTO8H55u2ZX+gmAnjUFyFedFqBE8OFD1FD7dHmrpijGJ6Knu6gG0w1xR9VTjkX9ktwX8
p9izt9mvpNmgMkojA9OOdys98GtOMuwjydwjcYav0yi4j0rdtiJEzq8KiXppCoxUWEzoDmDZ7fEw
vK9+jfHqLKKCwPKXQ4N04pTte5edEpCS8LYf6i7sB8gIb/xpeGR6aGFKkdv2LvSgsN7kj765a+OL
o+UUGe1f3NpNmEMTaDS0b/cVPHmps01KhkTC8wY0xrE8fOiV6nSM0XXoNI01ytzS7g3LH2fDpGxx
7Bt0o6zI3pTDRsPbNlA0wShbLJAunewr898BLRWmvMBm+3fJqVPcyMUsiJEoHldUPoTFP8WoKF8z
Os0OdIWldTgI6XMH/mhymtfjTWqgsvCFlnRjwdWGmSCtrWd2o+0ngx8Ta3XvxlFeOZ7mjWFxaa5o
pCQM/XGizsz4rTuom+Fzo8Qk4slWltSA9V/hdNvCtZWryJbZ6xmKFxsSDcI8xzCKtTiPvaISRats
ZEN6n6DFtcQqWe6CGDGY6pWzJyI+WskUBWY0wXxQU195Hl7Pejy64ydGUqZ6zpfPsnzycd0tvQYA
ANE2/v9LkFlKl8Tx7JPsnYjtClqQBFYUHIwo40xruSk+yHpygiz2s9eUFE+V/ftQI9TBoibS2cmr
eaIncrI23NVeRlIbaYJUUy/IxZg5XyNEzlMPWUufZzG73jdeqXECxHYdGvbGsRJZw/f4gXWqyAKI
RJfIMYsJLZuISUmDU8f6OTIlvtzqS762ar0CuAwnggkVQB10NRN6dD/wKSfzFFAgncm2EQWiTtFZ
LNRMX0+kqqbcdkrASYCpeON0bdGbQtuNTTUmG30zRXJ0LvYmb2tyZD9x578OrTBJVDK1jWalHeUJ
ZQywEaaosVMobVVKCZoLo7/RPxTml71mjrnexAXB8YViOjsZBSidUE7cDePPjlnVov4ilXcJaEbQ
8Im4W+2UVnI82DXY6twlIQU4aaq+NuE5Qh1BtwIGLqz8RpbHVsoFEvQV5uW0N8vrAh89VPKQtPTc
C667V/93g2vg8ZpuL1Pa411VlJ9mchyvMdOB7A5pObb1G7smtNrJzDC9CgBge9wF9dQaaOtQBPwZ
BL7aQgtEZMtrwxqWlQC3wiwM9NZRb1osbpCKzK9Mcwz55WhvvLKwIYrNgwfU41PT2fAglMQFlCwJ
fT0n4KYiwC/6JHlm59cfs9jGG/87N6wdyztOEGZtutLzuJH0c1k4A87RziDAJO7XyE50m32RmxB8
wBurrdUlhy+SBR1dIwnIFqF/9EvI6FhTpcRGuvLDt2uvcrV/AdK/cl41vTCl3mQMoUgnofdrm3Un
fkordZxwhcstLtCKWXZ4IVv/be7+Sav39Yyojm9RqE2LQZtuCcsHf3Ag9wA6IQoBuuxp5+oPzm4d
ZZbng5J9j1FdtNp1HC2u69mJDopNfu6UsFLAORItrIyjJfxu5xsWZ39MDgeKjYTM53hL89RqqtCz
lGQfA39f66AdmJwhoaJUhscvqV5ZrH30du3fQWofbjChMDEeXngtx5EnJ5mW16VPwCtCkJW44+Us
/OAMm0cMGZgFb66HWtEO5fTIQgShKmJifs7TvujsHi8oqsn5r0L9Fm3Fg2ZsCR+SCQqSZh+wRiVK
7M7Apix2uV/G9jaQdLsbQCWjQtHC7hUrE9hDtfAIlP8hqhEs3rJzY5vx7g1ghi8H5UONlcZWS0Hz
odB9JWdlOf3Sm8Dtiua25EB9A7LZxKmVmVhO6iMRJSHgbg3VaYxk3fBADb4lHdNrqaDAS4PjcPHY
E+6oh/4Xr7KsXhFsYF47h52/I17hwpWBbFnYXoTjfoaDEhXA5cQ+xXmLHwtm9OYQr79R1Q3yRrjD
n6fV/V/mSWQAcYVzOqmNVIAnPdNe6UbwlcuE2n9AvMqDVMPNbhnfi9FtZbrFE6wlDFDGRwKSO/KG
CNZiLoEn9l5BYrbC21YKeqMA69o9C8thV1rLcbCLD712uHkxe+yGiTgGLV5NZwBlnurLz9EysR0b
U/Vmi9ezJ8/ctHeECMt5/0uFCuz8CkedE/UYGylZzRulym95GJ14nGGpKfNrPVAPpmpftuuzF4VK
gCACvQX37wRbe4PRLFyava9hw7lNApUTDFzTkPrfu46BqXFvehQ7pFTw81pCekcVAg/l4Ah2EflM
srcXNSt1ApWbQlTUsqwuutIsVRZL4olJV2eU46zwbdfNStvTNUC/NhXxdmKhwzW2XvbXRS4RQnsl
Xgnxs8sThVNi6k5V3p6djQKNKqZjgiW//qaUC0fZDSpp5cF+7/GU1auDwZ6ZAt42pcvBhyx1Y9Me
IC4uSpZZOkfhzoPpmFJIEkHVaOpQNjiT/fP/TheXYRMrm1HRjRab9h4dS/g0UtDScfQKC7+VvaO8
AuBCb/c8m16l1oYIW4DmhrNiaDSOVfKvwjVuJYQS0Yjwqnnye9E249qeuvmUavvsKXnrkQU3vOcf
/TzZnoKCvkujz7EkZ2knzu+y5z+BweYvJRGI2VKVaIcagj9M4uZ1ygM09+Ae5mT8S8oZ1guX/j7m
qR/YH+BvY8uUntRXFgbVeIW1n6EHwrOY4DNKIMPNXxva+rPE0YZHwRsFMnrt01JqHYK2xn9W5Fkt
xuE3qmUQ0MFiAVUzLZubFnNrZ5Z1Kb77arSsfzJPcOYL+jfJa+pxC5t17h0n1y9ev3D/e2fpuTyD
/8JkAFpjpW92RrSbseGXhNxNDHXWjTquGW9VTaZV2WEZe62biZfUy11PAC3RBNKjgHHKhdLohrqq
btdfa/AldDh8sa3QUGJA0nYkCp3CjBvTqBorK7zTIz7dJYfnVi+NXo5lRx1GhZFrY5fkzPI69qei
Xw8rXLswnp2YqQ5uIiyWXCUT8OMHmkFhLqkelkSehwNn6mOgFyyuKxARnJi9OHhKwuctW5XNx15e
PQT2TxZY+sshe3+hsCoNI21L7vm5aaVbk1ALsBQqH2b5vCxsbMij5+dSdzFFD7d/DeG0GZh6Xhvc
7P6pBaASa+54DtQl5lNm2ZNNo3F8WaAjf0osMKa9MUFo6LAHR3JoXkr/T+LRjEFVjCoNkMZikgLZ
3ByZFN4D1SuscTWUybAlUY9CodE97Eg/PXwKxCxoARwZZSgpJtd1MtzxdbpXOGjhzo4pbHUOEUzg
DrLYsV0D+ddF9N7YdNpiwCtQai9yoDaR6rkwuK9pNV9c4nSlP3A2E89o41LdyVWcNaHQ2K8Aer9Q
PKGW1L/o7RxV45rbsDOCL8Oh8UYaBTb5E4UWYXZa4afLWy+R7HtwTyZtgoGwM9RzMLHkz1m3EMiL
vN0gT8D40GJ4aiR+pr8uEn5GLLHXNFYsp95qd6ZFd72p964ZttPKbPvZj1LdiuqDCOuK4B2cK+BK
OxFVId7rg0I/AP+RywsLumE2cZu/Aldp0XUvDm6irmGFEt7mjaTCjIgLEuMvOB8kQ7S+T3QuKMuC
DUDVBHii7/EvZHQkRQh8xn4WDrWKrZ9nTyOPVfxTi9EAZjF50UvB1PSDzaMEJJgoitO+htvh/gVe
nZaeqUvI84vsotb93Cht9PlR6Oy3Q9Pcy5lmcNW1tukK4qi/pMyudLgy0yo8tncmwxyE0KgwGR/3
D104+LX8R967fVS2Ne0KxzS2n0cIhFRD6ul4ew2EtjcaTQopjpFI9zJ3k/m0wa/JNfWkmrdbx2Wi
jauU4ew/usO4WncHpLANCCkE9nrRd1rbeIfA97XjF7dkIQHiQxZ64DZuSyj3bLrjMNp3Gv3eS3F3
4iVbJIC4PND+jVYAzzV12NJzPVk7TpjuWFbX0Pq0QIzEp/EQF6rlomcoOJ/Gwb7TKjPws/jD/9KY
wYnAWtrMQA2sC3hsJz3Hb+vxOhvTPq54xHWfQ7PXNsYa47l33twSMQSn0YhmOmbasECFrtB/+9Fh
iZeD+umatthYqhFd1DsCWe3TGmo7F0toUr+M/TUEUDOJZxBSaTIuBykIJyilgbsZO34pc2MYg7ht
8OaifRy9tN7I4UtTKgWj6kx5hEHt7+cg1ElaNqa/buUC2YWTjEYWMmOinSW1/Rf7s3yYgdWLBhfa
Bez1YKK3d0fx36Lnt+EitZU3egXZPv85Jsk0PN7Y83+qBJWeen02dQ0W6piAMX4+o4rVB0vgmRsJ
gF4CjYM0S5YVRVQqZMuCYMK+2Oq6AlqGYnMq0FhHirmF7zEnYZZdgs/9i6M7gQ8+/7bNDboVrQt9
I+QnSfBM0CkvpW4JRZaNHllKNs18YtQFrW0E59BfqppYZuZTHYPWG6KC56Mc7g+F20uKQsslPjts
O/fb/9sU7o8qc+q2uEdrUgjWA/7P5OxeNrAboIW36JR5Ea327dVdxl7tGsLby3ssslCIyP8MPT/J
Zoiif9CyE3TJITLSo2n4gs8WCfCma9+Dy91khl4thInbCCVdWavzzAT6rdwUjgP3HQd7LLn5meZE
wLJSOxFFc6YmbR7QMPCf2bVFnMiaKlz2hEtQCW6tN/QLbuCb24KuNr0xtAQWC0aVdTaUTxQFTmDz
oLiGO/uQ9rPoJunjD+zcEbSdi8bAEogEQDsHsaFloN9HyHBmOZX/Hybl86q4B/TDFUK0f74p822n
NLyw3/g=
`protect end_protected
