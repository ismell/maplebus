`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y3vQYJGoi3blgkeLg879oEdoe1iB1+/mlgPLGvrwhHjuziZvWcfMDQFZS5sjqzLt31/gRDV5HTMM
ldRRpb3CDQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIFkgaVIz/lIyn+ihhBfHj42UOgxqtW1+iPBc/E70csKfvykrX4u1seWzaBPfEuarRV5vi8m/M7P
AU7E3JXglfI5x99BDc+HGZchCRYDHkjgA6esCvNlhVE9XHv8eRQgqZTj863FbU8ayruVEcFz4r2O
LHmdpZwWOp5MfhSm3hM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kFLRSb+px7e2wwv0x+CJxmHcwTssJsTFcxLC2a+8paaRd1PBHKA4Gacci9U+MJctxdW5ViL2k5mi
Vik8BsiJHVMyXnWtozpPERCdP57gSsT+P/oawRTWgr6GhjloTipzMsZy4PPb1Ta9wF9W+boGqanG
/QZGJoJl8IQlujJn++DXQ11vhAvInrWNuDu2sK+4sOuXx4Vj5zicpumadaDJefD+H8fa/nkgjSm9
pvmrORhPDdOsoLbbZN6Pal7jiqSmO+WL3xMhYfwpXe4nkSYEIo70rwjYPq10pGY3veB+OVCxVvqL
NB7wUs9YQeRJYuHH+9DZW2csOrt3elW1u3o6ww==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a1/FnVKqm/JQCzg4Xfmv8syNjE+66CsHGs+bi56hN5aYZnuO+bLwIfU9rOkFY1ITNF2HCBe+uD/b
mFugEJCYjTAKc2kioI21ZeAAvgLK+JwSJF8iJX+vS35/JzfHfFEAqRVM+v32B1RhWTzYCyXMkYy5
FFqSnRbA58jKB2xivLk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Wv9V94CAS9tEczd7Vd7LCj4v7RZvLlPgjHz6rIlOXQ+PzRUxuzRzx5D3Jtg8gN2SdapVssKTXLue
+LUwzZ42sXQodXJHB1tTHr62RO+lhxGGn66XEqAU1v47f5nog0L3bebjPOX4eq9+7y8WKLpXYzjJ
mTe8DMdjQl0HmBbJ+GnBk0oqNzwYHrol1IdAh4mb40/mpu9e5GZbasd9OOCdrVoijfC7qhc56KXV
LOhSTfL74ysBmCRb7G/ROSf2sqht0eS+HA/JAcAaK3Q/Rkp1dhSnW+nDKbv9Q5/V/HZ69YhtDpXU
K0tEysZOg0pygcQBo7iEHIdsE+IjkqmMKbVqbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
OD77meUxaM1WFcBluioChjnE6mbJRNDWbUEhdAtPgx8U4aBD5w28Z640FE5E3YcYP7T/kBeojGda
oiAtPYw22AuavPb7NjhkegcOb/7FUrEa7a1km1c6ZfpcFMnvpUi6BHF6HaVmB3BEu47Kcc2ECkG6
5RhyWiM6xdyDxdzPHkcI1I39du4kZReUqWJbTHx7QPdoZ58vZLr1SOG0wZdN2BAZaWIZEPGbb5CA
YI6LqPEAuyMqb18/9eaMWcdakbrWuDPs363pfEfRUYlyqcHDO3dtGTwA2JbAO8mueIGKG7hIyQzP
a0PJJdmGCVixLzZdbTmXkZSFTrQ2dj17pZTu1PjYgYpHTzbMdRXDgHd5QFkEaVvrn2bKIBeKRrNs
0n60M7wHjJoYMW6u0vGmKlIYH0EKw5XG5Lb767JqUWQGVdYHB0Jw1iA046Zv9BBbPpXxT+Ghnj5A
626eJjqDDXmuRzBBbLco36gOIj1wJO5FMCwtX92YI/3beFS5y9HdYA6ESfI2gGqo5x86U1Z7Z2EP
iQSHNHP86CmYXn6RxyJqpCwtSbzoEuTSQ6TD9+MW8V2SngICz7J5jduvYCSAKaiyh8y6uparEaS9
gw5Fcc5qjHBvvVFV8uy9Evmc8BvN1RfhRQN0YFTOHQlzVl4iuTu6KGcAHSWVGpCZMiNSc9Yjo/42
n+ZDiUGrAYcvkH4tUJRmBieP7dG7TKn2QqvPXs9oGugdD4ltqBDCEXW6Tz4sbiB8QYMMjgoxZ2jQ
KlIrL7JtcabE43EWDU7+ykoDAPwQmMHhUnQm4xpMmRXLnnijBXy7LJUBeEH6snRn0QhWFLzJ7ok6
d73+mTH3ec5zuYinjxGlpN6kFV3lZiG86DhLafJiH5x/Fp+sFKw3szFNmwVm0p2CAQIcM2oeveSR
u9zZtT/lRdIC7T9kSYjlohx/e3RENIDOtAzQFGtPlPZ/VpyEzaikNUPyHhIEh5kD49pYrmLGFxvd
OTESCe4DpeSGHwU2egVyN9Hq0P77t76md+v1qylZk6+tEaTHNh13cl0ZDX1HjbkjrFN+SI+8ZPcQ
10795166QCMCIoGnpByzobIFBLIUmb0nPuqLoJxO25pxx1aVwcocxDIFvjhuOCvwQ1qJVqX74kVq
t2DPHDvDjfRpEgyYCXdEu0UM9JcZZfFijk8ZTKMPvyvQloa9JvPWfEb7fmgIg2+OLf61F1fFI7PH
/TmYJjgilW+Q8SB0ole8GQ35jUc//ZksmfGRqR/ghmef51SnMFbzAusS6/LPvWF1cSI/pAeqJ8Z5
+eHBX2mf6234v58JYRvTLAjdQb2tV/KFsozDYi71XRsYh2lEGiwV7AsaS1y2r/GxJQSx6Ho+QWr4
q7V/+2wbW2UeGaqgauZPh9U2gVSL+kMLDC5z8DYnt06JKjxESDvUChD5iRqfdhOKG+vwumSfp9gc
KGI5NkwTjQ9XQ1pVW/MFo+HqQaX49xZl2TH6RdNqzbhfjgFyNtlnSuNBrAzjK5lEffGcVy5JNeQt
QjEy5e76SmfZzOB+4QWeFlpE+rzTq7E2X46GWyAbZVNe7hbKr9VVFz+dQPFRcWCPBBw6ZktvXt4n
tlUJB5VtFwe7k9Y3xrol9bjQJPYHLnM9dnrBzPc69nYIOMpjMVp0sDvFwetKKjiO0mcNKa+39j7g
pO0d+lBl+/NENZYm1159/dZWM0yAdVy6Os2LJ7wv0o1SWrXr8GNxd8Ap5ebM4JU0G+88WyA5kCBD
iuE0lfbg7s1Nc6Y2b+euLk8sc+dENMyWoOtN1Idburah5hWnALZP6CrCGqCvdNdaawSqbYfqavhY
2+kxQqdavvIGxDtbrIuythOzqs00FNfyFb73XCRQs6Lfe9QGzXl0yyCGY2bzyP1va9kDP/zMsfbl
uAYqkQLdoIC/iyMvNCzkc8X9vbYqSrtB2e5/hySKB7BvWXFiqUNIp98A1mjk9EF0iCHzCi+hdV6H
UzVA5+m1gm6b0G0ERgYL5vi6RpODjRDaYXp4l8RtFihiZ6XtWMzu9toqlb3et8oO+kgPqq6FGtSi
lK6mFBgFbGpmFPS3Yzg7FvcoDrJFLGwL8j5TdmHSwFki0mlbJxuoWjSXtHKaCQk8Tj3fG2q7g3RQ
Si6SjwAk75+iWwEYKtihKZ0ujzu3RSmNoPfzFmNcFPsgvX96VFJyk6lGvt8PDjJPEO08ld7Nr/yY
MZt0iqpbgU3IaOrN7gAi9t+RsUh1ngmp+8LkxyTW4szzTES93CzleTpLHC3OQn14SKKQ3uEeWqeT
Yk5w8p3qJpqbg9TIDWXk1sqfAGd/xAgwVbRGDYNJBr6M9rdxpBhFqvbRqLcrSY8MVe1EFEUYlzfO
dhvxhirvurwILlDEmzDoI2/hIFDgHSoLz8S8o3MnE0HLTZEfEE9hXbITJsqgt+O1ao/EVg+hRj2W
hx2x8dy0uH0nMk71SL0qNaInnPb9VQz+DzHgjIsWIkiHJJaqJKQOLEfvW7aT8xL+XOreS90ql8Vc
BR+AdD596ndTrS5T5qtAQMWEJOROHOWrfYwg7vQCHQooySFRw5awLKMaxO1XJ3qHaCTw4ArLuxVw
ojG52JrIbepm/W2i9iQZmITE9uUcizE9FWqTVPXcm9CbP3Zs4G9TxvSzFiQvJZSWH4RoGmfeo+Ec
P3thkx2CWy59u+F72Ncu3uwbTF3JsQRPfc09LAeLrLN6pBBz7+xGN8Nhinzyl5wTO4suqT2xuO0/
VVmvwOVSQhUffLcyTSPQRn1CvFfEx61jFm+XjFSfdMVb8snKKADP2Kuj6RTXdsA2ha9Sfw7Syy8u
5qPSU8XZADRb8ATxz9gDA+EozGIRRSGLKKOusutkjYGl2hdh7O/5e62ZUCv5mawETbCgRmzveW+f
mLRdsH59TRcyqcXhM/upHn55oy2rLbWcvPC8VyENHqBM7yLVaRYXASAMXteL4WSygtSND60XWZAG
ag7mlMueL5pP6SxK/E1YWJILmJBQsCDsFVvehfc+mdJ7+Vzf8bCOeDmv+3T9GFDOo3bjLjJvSMnf
dY4G69LH6RfVGRGZTYi1HFeNOAdAbW9aoOpu7xjDPXdSvwIuTJnc5o952eXJlpiz4RGruSvPcZei
RTDSpUJRA3/JeVad3PYXN0OmIYFhNeaN38J+8QcttCrXQF9WHVe0pni981dBV/LKn196eDbVeouB
GDZ0uog0XOCUeY5hcEyrHjdP5kQIZop3Z3RwonKpaJz0vYuHTDTnDj1V55nwVqFR6AguMpXt3GNG
0zzR+MnUF8TqchZPfdWmQD5MBdoEBiwKyj3O8gRvMxuhSTgCLw7n+doBXINpcn7PC0vHqsAK6I7z
YAV1lQwkm8ulLtIWUQ8oVqyec1pdfMpEcNil3l98uPoqRGDhl/rRq396WrxdReVq33IG13uYmgb6
9GElpnKTImy9xf3TRsX9RwVvGfbA732RVEr3BoiuWO3XimtltaEzzMeOS9TyKc6P5kXAlzJnE+B+
1VuRUaRGauvn/B9f3JI0sRWHBkzJamqNPk3hyvrFDf2fNHN+b23trTCoOdArkhMfsc78DSCA6YWg
1bg7B805iAH4nUEwWi541i0Zy0mpmX0TKsYYnMcb9xgxRmiqsSYotOgpeVivl3gjX5Vh7bNZ+2gr
ilFDTtQHsg4cBD5Tx/L22UaefxEpWTgxEjSyVk+Cc3okZnf0CPuYNRTbQ8QLoO37GotLjqobIWnS
FQaQvb/vXpttafHeL++Tu0bwZ+8cpPXacS1kgKqxBKwnIIG26dLp8HiHNwNh7JJvr5DlsYVFRwaW
EfUs8PNjkcWlW+q7UcEFMYxO77uxTi7/T2J9MFA1KBNv2vwgsQiaTs2Y1V+Rz4EMY8eFh3D5SF/s
nyReCWoqdOZY5D6G+DMsdntOPo+LEHwXqCGYPs8rb+Dtrd3fCGP2+CKyMHfP1hlJShfqch9Buhw1
A6Psic1A4zZw9oXd5LpTJZ2ygUtraGFoC/2qOC/fzSijQXOvvQ0SzH74HioV9eo33UXaYIocT18U
9RcvpgpCrXa/IVtrBYfywCEu/TBSRaCZ7UYx33YMtgB07VFyG97H6tmYG/UQUzrikDgMz1+fiaJ3
mx9Ng6aXKe4/+HktmR92ao8QFDrebuTCuqmV7RFtnmYjyxz721PgsZO2OjyixvPT0NKSJ/cRAQ0q
WHd7JTk+CBrQnhlZZslGs4vLCby110j7uIBVLg+/XH4V0XPodjivWUmZrsZMVTSMNjOGvXOm/5QL
enYIihC/sBzbTxAXJCV6hdyIVEOXqfOZNoPf3AQXCdjCJEZo+GYyM7wsmKIfFi93m30EU/1nbddI
hxGXMt4m/qBckrP06s4GUFzh6Tkq0N2Q3utY4eQTCgj+LSrBcDroJEL5fiHCLamqkipmrjw3OTQH
ksTIEwer/BzRPX8O406gBnm+5L1rwI39ZRVjNhBmMkUsPTq6xuKkbnsa1TRudd/ZWGzm4FIT2dRs
kLAt1Fe9bNqQW/vfu6hodxPohHflQmV7TN0/M4sBTzHpAI8BkTNAKnx4QsFjLCU/h2VN78Os4fj5
gndtB+JlbYiqOqymsE5GPNTSDmO+2055rUE1UVPjk+dJeKSzjtuexcWlsSKcj0Db9JJsQLGs5dQD
FGfMzH+WKOKm+iHDv1OJRSQnnrqd/VR886ubSowhyBcHPv8EI4V09rpTcFx21qIVKVGRMn6V63Me
Y4XUwJoOD8uDyx8rQaPeaYfJ7UDa6Ynu+6mPcoftpph3b54zNYmLeHld7zyu+9xXpl3t4lX1cTlv
OE7BHfs92gf8L5SVfcS/ypx5wpNQUZIQdI052IqCSk0KUz5ClmkZj5lhQ7R5Cnx3x0BmDBePDqtp
lj6HpvaLJSsxm8f9pPcd7/Iy/v/JED9EqLuS8NDWnD+xJhqZpznVihdZbvWDZH1seVEV9RYcadtA
sLenfiTZOHRxB9qQ6niXEbzPhqh++9gebaKzi6PGoVfF/3cEd62zpnWpa6UFCe6Wln4hM3zakLoV
gNGg6yn4MTR7rmy/GAmutPEhKoq2UBzeWncJEn+Ut2RAlSS5FL1tg2ry2zbjPFEZx3mC1JPyctry
uaS+0A4B5E2QpRqp6js0bnrHVl3SE+N1wQ2XoGFH9HzGzB7Pn1Wn74rajqqhwRizpd2zaoKujUr+
nfxLiAnpgpbEYi5kKWXAcoUWI2PbaeM0d5WpYLFrQhtkgaf7D4klio55R82M+KMJj86gqWeCij8B
XXC/RfDtZj2oEWAAOhPs2cbNd9sliQDObYo2JLQSl9cuSpq22IkJEh3YmfV2WHa55h4Fd/x8tOG2
G/seozcU6rgPUGQ+5i8+yXQTzwuhiVljgeXy4t6IoS9siN6Gu5CFk4+xDpUIJuk72WAo1BgG+1os
CAPSD3KkTR4kTMbIuBFYLUeB2kTfq1c6l7bcZA1I278rAjC5U4SPdBGD1hdRRRIyGymCHzCi48jV
aJvQykCEDqW7ZoHU+wuu+Ea5ONu2fRS/ob5HxHwYqrhtNBHiqHu6u6jg53RCdfL57EmJGfvXbhBp
nM3wooOnHLa1OBWHNx16dqM5+bkQ9JeSsD3YclzuXEEWYF9f9cRu7dtmfk/V0W7KYGJ9wguX54C1
i6CPhZ3EuVm3uwkKOmuoYB6IhpgcQzo5T5DUuQX5YnhgOBdMVSoVQxVqN+y7UUqZNUFls6FRyVe7
etWphBZb5himM3JM4RjpikR3aLBJCUHrj90Cl6cqou1JeNOtxTlvTowSN7HfZvvW23nkRiDcLvye
WcHt334CgagtIus6hWL/WX68kRSQR2VDXcl+Gn2v0YzyKeLzz+U+nXRPmCS1qVw15DaCtGvLnrum
9xEadyfJ+7dOV3HddZsIWuUuvkCg1nG5ZM4lqepD0EVUze5DljVfRHPto1M/wZRnlZ5t9Jdc1yez
T8nX3WCIEPd2eZco+6qE5xgXqVKp8C3CB6cDfotNbOaeLsm9a0NP3UdtBwNee5PXS9eWm25+WpKT
8bX2ng+WUmrc51zbwKasIC3dS3i7b+S2sk1GFQwmR3OmUQqvDTx4993nrH1MW8BCjHjd2Q8v41CJ
46BT+6i6Scr0Zg6EDiU4uE7KT1TomFPrdexKM6UgowMJteh/NEzFRm6MVwK6LJBstJRJr1BMXMFo
p3S9KWPrPlO3QKgnt2PW2i/aBw7d9IeaejJ1PC0odC65yZ7kGn24+EcYvK9kKC8/mVCtJpKWoFuB
NYKSq/gMkD7SYJ+NVLrDFZuPfVaD0ufJ4hf1y8UbIrl1VO9ICtpvH/gsArE9TUI+C+PfpwCfowPB
/38D957HznrWgSheww96biwxudOtI7fly66iTEOVb8zuHg9UMJfK3YWj9bN1WwKBve7S1qN+0jdr
3kI5YRYtdbaUR9IEIQX4A0iRffN6dAECqA+vXBmaJignz4ACfeIiJ1FQHh9gPihIaM0aJ88hDVSl
kalMTHhQoHMX0w6M0DDpEpWApb3WLRJaD4QEX4w8RZlP7xR1MnfDC/BVJeZ+0PtpawTxLm29n1Q/
Yg4BgzuHgDbQseCwUoE2+rOyDAWzaj18R8kBwy37h8U792bsoaHMEYpOFM60qck+DpxqvuxtGv5Y
/lr9nwlhKAq4mtKrJC/sPan/aUWaXEgYpVWZrrMnyNFFsMFqrhrYIe3JXFO3BMdCed/pXWuKYOHG
K8xe219/14aEZcZz1ON15Sj3XkrFJUpcHRuM6yeK7MLO8Hrs+kvHTmFGwwojEunbIcc6k67KANW6
f2Wj45h1N4OxjeJb2CLXYXBpqIn4FYLu46MDd2JGtNToXHfE6cAGU0KxVbSizjGKASv1IjacCADW
kq1fwuvNVl2Kw5hkR+MwLgDeruJvZOPmhQ992EsgYmtyPKpCzAFw/oWB/PudrFcp2FRicDnUeZ9/
LS8AauM7Qo9Q1+aB5Y2KHUVDIDyOfRGHWqKeA6ONfrmK53iJ6lrVM4t9g0eUpHsOh/1FPQqJa+l7
jbvSHPsljPt6uz0DLIStr2+61mDIss5+CrBK+YAmk2XklE3JDxuSduit2FjagYEWvLVdy70js/QB
80ZuUpPCttkhyxJ3A7bMWVVfmUqby5oThSInR5AD9GOM83ig6/s5Dk3uzzBwTwB7CA6LVn1EEZWB
OTGErTam6IDkHV7ygI4gQXrsBlD6HxRXfBZIh/4xk8DTS3KV86JkJ86ewh6p6qMojTO9dD1OooiX
t6nW8ahJmbJG9/ptFIdCywz8wmIMdJQyA1hdeRC8L41XLoq27vOqCgOj/H7rpIBpt2JWBBFi148O
9iGjI48KjDTzZ7B2W19oMpKesPZs3iwmOAVbrOGR74hUdUVWUgb3Bf39lH+pkos1+1/BL3FG3RxP
E2iCKhFgLKBnUTTRkG3zJ7Chf4zu6oC6N71A0cXmI2jRBHs4olzX2J7nXF6VolzkR7Q0G/fGvWK1
7wv0M0gekvdV3DgVFcbGwMwpFdjYqVqQMUayxkGN6PyLiTDyWBDJHEuMHixmaH1L5S2IcRUdLmXz
q0DWPhb6wpEMni8K7wP+PggNz5kohZpvZoSwt0XigBzFc89WnWigfprCZwqu8tiKg1L3om/lvjG2
iVRjySaDqU4llGRD/ZspNr4cH9U4AS8SHjvwPJPQ8bESdelTXFUfMB2xhF4Glu+EGfYT2EB2O/nx
yjTkiJ6NzRoDcXfMJ7i1w7taumjpkrmvbKdnWQIX1RkOW/A3SIy19uCIJe37Exn/PNVM98ZJLuPM
T1F+L2cpoqO71qs4+QsWpCUcjGx+zglkIwZwjQPHrf/u1vIXUK5FgHWWH+DE4agrbKXdXSKlA/JO
7zofqKzsCSsSa8XO4/AwvSbmfFcTC19qzc7u/cSGZlpSNElWMO2oX1Ued8sZlnrdiZVa/JoraTMT
xVEbyT81mfbuhABANLCh0MAxPCi3NlhjiQfU5wEmTcxN9edZZPpHTMs6CAlfV4AnWE6Y5r1GJ4Ks
WCI/PO4Gz883kKqXxCceSWl8Zk8KjfrS3H6atbW0zTIYUpB81jhJhISstGEZSrPW+a2wRmF1LMSs
llWhFTrwl2tayyBAuXAoXTY3YRPQNYFZUyY8Ps1dMkNL80+aAW3errN1fpcPJwE+qd8v5CwMh0YH
4a4vHddUhIw7Ty6jxDaSalEFEM422/YDbuPdB4L5SbIHQ1r+KmVt6jy7VwADoj+UCdGfkxIFQB8P
QeE1b1VPPqY4f/EKQ9mBoOyhF8PXjq8fzHgwCS1BLHBtPYrVt9s4rixfZCnBt6P0s9WBvJNtBpCv
iHxv6EYEbTaviyzTwrKTyPp6PAeS45N4C2st/TzVbdyejQUOrsNqmtKbtT+jakKGdyWynRYXcNOp
mWK+xjCPSq3/LT6QRYPVHxy8PjKdJ1PrM1GOYmKI+upkWCSAzNibdS7Ic0dUgu7G5ZISulFYpNfA
MC/pzwsJW1/K6RKiX3mmJTRxcvhI/+ArbfnyyrLaGB8/tQ9FYkvvvIJYTTUHt+g8zH/7IZegl64/
Jn/7Yh2uFjlQPqvzD++nWF2wXeGcjoF+t06L2fXNvI0Glrp9/SFwnYtPnWqRAcsKkN3IkeYS/rMb
h/hpY1GimovQ0h6np5tlu7/BLNx8Povpk3pSqq7VPTrpmDFsFmMnAh0AMW6el3AE1j8u2ZkkCi2P
Ruz0/uvTHgMg49WzfNcz2FeveIcPQLERZ2dVrgyImQzoxFLTzu6N0tz49BdXIRyOCpsglv3NSy83
OvHQ8NJyAYlXOtch+8vTkQ3wVQEg6g4TuEz9ECGBaoeHnGO6K8Hkz6KNEnHcSWeby/hksDUxU6yA
GAXkpswm1p71Hawj/f44MFGuDCqeHr/hEOhFFratlrRns2TSpXjUGkpe1ouDnr8cz9QOwn7lIHwI
HgfXyk/0H9P9vfqNTdxeknW679GfK4sJCy6uKqHKfqkwPG4UpOBfOmv9IWqPeAGbCXjsJvMO9uzq
cK4g5dMVzoqooPA9vEF55/GoNWbmiVQ8sNjtBps+xTv0SqalZhXDJnRT4t0naN6WgS3Vb1yxbd89
V9I5HmxVI5JfMLvh2jZw47FaAFRBa4Broe77RZqho9icaACia32b+FWQEJ8tetTnZBXXjkbQguc/
zcpHvuqLbLe0rGfeAkr0PzYne1stsAFS7Z47DYGKGLDNrBAoJ4STi5+I1KUXsRd4t/wcL5znF9Vu
NNqEZVh5oI3qc3QxzlRP8aZ49AbO8gwaGKtYejND5OcnLNSVFUPjKU8ijGblw6npgPij8AnRX5li
J9yt5DRmkY9w1Aqok5jxLFxUqCXp28f08YwrPMFAFEqG9rX2Znum2QWNhgZ0XLs+glPBHDsTbC1l
RxBMAGUGVAZnq2p/v44ivCg+5SJm3fx4tub7QmEnzV+zEdmjpiuPXQpE+IAvFfhUaN1VORFRpe6a
Nn6NnGgtImQNAx/FqP21PqR95D8s0Bv/Cq4/mSUMkY+Q7qVt5riHspdEShO+1Sw+0Bl8yCrYBvsJ
LSvfG7Gy5NUYt3oL8ePP5cNhpTouSpA1iRDUpSoENn29lM8Swtsanx0eilOMf/ZVNO4ckUqRTDIK
2KpoPjBSKkZ74z6hZS6mDNUMfEQCttfP5YfkJd01AiDAUTlOLErTRPVK5SAOHBuGhyzVyXRUi7FL
8wxy3vWX637zzxTWeON16fTpvRve8nk8qD+M1AcpM/ybvWVPCS9hXVgxlxzfjoXzByeQEtw2wir4
Xs8hD/XjuNZcXy0FqK/N/3mK2nqyaYk3Y91qss4n9736d37CSs5lpcP2KdE69BqvSVCbrwUmHZdB
Xeo42466LB0Q5ANecKtkHPFiBCrZUX4WqplizyNB1JA6x9SeggwiSqAcp6gedO5sl4H5ku2GlFm/
/JOnqj/MVi9TEaDz1CiTSkWE6QyJoebu8S4U9FeaZNB8l5Afk8wy6NoVuUYdcly7q98zEk4qOiNv
VtBBrSfNBjDynfMQY1cJ3wXya+RBXonr4WqDQVl7rOtxtjvPvYpdorYwO7N9bH17EFRRuAZELQHF
ojIf/szFddTReG/ngym3jD4BSUkUijS5sUAPPp2niJBNyfD0ixRGNWemvVPyQ+WKNTHsdwUEs453
jPsI5TxB65T8bcRUMUqJniodu/bah75mmxyC5pYehyMnvthcFQVmIvwMm3p3bMmE0fDg7Nca0YbS
Ldk7aIt/HC72o42YpYcFdIJZsAKCyYwRE2sNdYVXDX2MX6RxS+J5zVYNkVBZEn5AV25xJcKY/AhT
g1zZCbS1S183WZeCHk0tVcIetmI9rfirBvUssRmpiUjtnZGHMwcFr3YGk8Ir+yerBNl9zA2ql3a0
g8V67zZ0l9qRbiyiy/vv8p1vw8NmACQRfdXf5utgih7QkTNoI3rJOLg5g5+spj41Szcjd+G39OF6
3VXyEAW4PD6QH9V0FqO1owNkrsUsiHpqloS3hCOutWnJ6oMQjmIsfP6o4fn3Ysb4+GtJRvFvWsAY
Lx39KebO8NloEuFbhYxoMFZtLPVV3KFQIHEzla858YrUhWsplwrqtSHnDE1G0zLRQ5CZXHtnLOFz
dySDAxTGuUJwju2syGywif0JfO/TI+7jo1ZVFFeNlqMJ3u6/APTWp/IrVm5biY41oMRx7lCQXXoF
gBpEfr0WkPUn75UVR/9ANzyEqCtFvO6TdBRjWXt9cdz+xq/QrjjYNv3vUeGab9Fzj7+JJdENPdKD
EwGcHFbqd5ruY56dDTFfx2rpS3HzG3eNczWRG4c1C2Sw4vCKwXB6d4i2VYlmyiwQSQsCn40reJ7C
cVFKtfecLC2NMzVca6NcDPwxDwCMCQBF6BpdfDTeFPZSUJ+xIYEm/RYArc172KSsnLOuUee8L5Rv
yji3TdVJgVfoM96wg2OuD9GVj0C07qRIh3iQegwXV/KiMaq+25iKo2IQATuPV6pndYKMSxBb4FXr
gTathq/gEyYa25/HcELEcRmYPQ9L7hpQs2v+jvkz4sdhxa/CbPdOBKbkuvCJ+VUMijDres19Kh9P
kX5d/NwD2oVtWCBYfmLXst/c1T2lT9Bl+JNxmQXaHdmjLADfa7v8P4ytp6ZRC8RFUlBDoz0OHFO7
Px4M6ZZlmIGr/TftR6VrjoAExZaZXvqzDuCZbjbwK08b20UrHaogY+dnixNuA21PMQLrF1/JQtms
qxh1Mcjt+D2nUAjCrRVDWZvyecMwJxQlonwR7xdNupuJiWqmfjBTnv3XGG5mZLYdQc0qbnWoHFOY
6R5ZeUbxWWNC5q1/q8JmPCvWVbtP/cJWPynckgbprZNjCB3x7kqplT79NZI7uJ4HPSwrEJzxddVk
/b8d+021ZF+CULqHR+yfQuzV+GIelpTAPvvBdBQUG54tXVu34eH6Bdtns8NJrlNn/VhoZG6dWiCp
/8LkRjKZqu35pzsTr+HsQl85LirAIyceurdKa+5xhH2KpE+oPGX6AeDZ
`protect end_protected
