`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qOipVmY3fn0qNeJcBgG1sNHjIJOb4KstB81rnTtb8GNEMjlu+MPGjXbHiFsd7tiwTZIAB5lnmiSJ
hkKu2/ksag==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mGhRFBwllporpLxI60+dRp/4eGRGHBGy3DIcDt6ess1EfQNt39yaEmH3/epnLkz2L6N+WBDQj0dN
oOfOwEB0+WQJt6J1aAx6KHxqG89t+e/knjk21TuIBuV0M8CBHOC7jZojSH91xue39VWSzezWI4Vk
j6ix3IW3HNCbVDBeo3U=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XqbYI4GvYTVvdPof8LLtoyIUzAkdShzKP4ayR4CfhZYnWI91PJbQZOFsgIfX6A3BYMlkaivrvJiq
YvAOH7CuQOI/YhtdyHXMKcOAJKrw0f5UDX2HWbrH8UCv2EeYjG4V0RAGXESUJ+myJ16w4G00+JNb
v/RwgNHqqiHbguLSuARpf0vFVGScEb4WyrpgVT0NrqAtcBcmsTmXUC6CQqFFN6BvzDCreGQ0ktTQ
dEWG9gkL3GIiHaF8fXkkxCgiShjAYq1l2R53CvS2Yxvvzh/Ho1VtEEM3cAJnO2bRJKD3zYF2c8S/
LQY2uCH6190IFW5CsgO9IuvI24DnaT/56aYHXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
keYOERLKRipzOBB2uWzVpHyCDtBAuP1QXo8eS2ad1WXCfAaV7Rh53wnMq4g4cdIneM1VJogRYc7n
4kuvPEeCWT2XjsoJR8WeWZwkkQ/Sdy8Ne1984QxR6E0W58tT6AVA4EJIyFyNN39PfgsvfYIsNplb
76PRpomFk19FAVAU46M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aM/cTcRyKOUDxBTfQxqpzOnnTVFSI4bzG70fvzamupKuPyIi3W+LLR1JwEW6OqIVEnQr0MScTes/
17LlIwNY5MP0NmQJl5RtOaAZQJ4auyDcvhC+mDQn0tsqiuUB4AcF+1wGYxgwVY9p4IGAzXx9vaRD
8UOguvI61/vR59Z9pMhjo8cMXes3QBPww/cGA+HgIG0jnlQZ+UmIUsPJKwOvqbYIqQ37vTVtVX6S
PtvL0auT1SGCP8+Y2HXBCWOARJ22MNriWrBi+HSR5WCTJp8D4S8LJyN26t9S/LuD8hneZO0EsASm
W8WTOco12jpzuPoFpAXJFrDmuFd2+iPU0Eekwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
PzWnawgXRBY43rTD01QMUX3ONSElj0BrrBdOK+wstylcq+EYFPfFjMffIR5wO8P/f7BcdRgcowk8
l/75ot6e+g41rkeZRFv1pRPLXnD5KrZknYweJ24moFgAxoutVPbZz6jCoBc54n/+VAg7HY82R3yA
eCUd1Glp9IbdnbKfLUU/xXELXzcT0Kqbsb5qGFxb/Ml7jUwZ7xS1ZwUqpX2vZdrFKIpdN4w1V20z
D90/YtbJiH7Fld73+2axzX+ZFTmM8Yj5kg3emgOSacN4bAtFk0LG5yVr9CYlm6wjNY5STgje3QT5
TYxrNyNTc/Yoskiw77XqG9xtCsV4Q4gMLMi69pO13fkNS6VqgUW1i/lUjli/dLadmks1zZtpQSjS
0KKcf4cy5tBqlDAQ0SEz5Zckzlq+hAH/2QqkzyVfl7ssQJxYDaTei8GKJlqb/MNnkZR9PyAd3E2x
H0Su+tD2xRjHCrXrGyeRxmUFAJk4O74FwvZ7Xh0aVY4+mEZOxeUURdVJSg2FU0r4ZRMm9yTYZHvq
l1pUH/69M95YDJrj43fxIudLBZlXU61CtMQwUau2kQj7qg0gkb+ROpCzDzxVF4K5OY2uwmY03pX0
yJbefQS4Ysx7L9ncTYpjeKANPvGuGsvNianpG+Gi+m9gvdUeCC8l/nBygIX7CKAa9P1qv/ixGDyk
pYo3A/FZlAzTFqi86RxQwr7ZrF6bYbExumxM/6iLNg/AJlpvPKDoIp9WKIQtaU0tEViwhJNikQtD
Ste3DWHnED7rGQCe9kzGqDbUKlBRiZG7J54i/7AWUAisqRgYXRKwWZpZ+r5RQWzhJUwL+KeQi2Tk
ZZVhW14q5ho7rS0wHEn4naO2Z8cMMkmUrnMSHvQl+UPr1OhGtEUTREoPh0p6OpfJU6+ieZKZI3lN
vEoMnlyVdaTZpmn8JlEMJXSWi0TWyqgF40rmCju6W4gL2MDQSzhwoS7WFEyoVhMFBAazZKIWsVoO
n+jdNLUg8svGqrIVOxn+1oICjZPDZkReqnBRrj28jfsM7FmZMu9xfY2FQRMbZclU0rjQtiGTNDaj
2Jwk95GWz63ysx66wPNx/7r9oh05NnRkLFpfu1PPhUKT3Rf+CDIFIxBbDeN01uRsGqk9xKErAAhX
jBqixtnx+dwAuw5ptrKt29ON0BKac5sL+s3oupVogtVZPRTCx3vE6EbDAs996ssIJUBt6pJuiyCF
kZ/Rr+kL/kxk08s0L+EtONRWdNVQqyHLIPZEWBImzI7tUHJmdOG7SAe75bvb6F99nQ3+v58IkvMV
bgdKOoxYtQQIfVaseopLmfIqzFbnTjOTouirR1ubO82Z5rSH/CXJQSs+t0nZEk3SKOHabE6XK0Mj
5YobPWQneo1OctVP+NUxKyVyqSd/cF0TmpdQKqUucXzGqmNELy/TBMTplALZKDihXTQaULQ8XYG2
KfAFPidxoEoNIsCr2wq64cTLPIFh0CbH8utsFs4FpDLKm0ToNzd6MR9AmCapBFn201J+QheSBgun
1AKvMm8uTYzJCQLmZzfaQ3PtEwOG16nG0usFgn2xOqvGZxIWK499MHgWIXJMvLsXC2u5LqWBvrDh
srE0Oh3G57q586r2a8q0C/R5vxaIk31nc9JFHBj1o2NUL0UHHEJWni7s+xUZdBVKAkCpgs1/gBAl
q1hsgcZo8MBup7SX5+LrHylqmfLepoO8xib77eGuGBSQXfB5KKTOeq8wr5gKB4z/Fa98FNWTxZ8d
A0Rxajn6xDf3+VRZPG+wdq682jqqM6F1GWG6hJ8OD3ylSpXXEAVtFgqE3dsvhqQVbtRgEyD55i8z
VD9xirPlutn0MyWYBSbLdNyoKq1JbyCtwg7hcOUjudIH6NpbSukYgIRTe2jVRbNQGCKHBigblpXp
WTq4rSTFGlPgFsIw0FZ64zCm0Z8GcCKK/1PrchqYfffTT7xxtZ83wgX7d2F6ARq6sTRt9B/tdd3Z
jqEntCSxY2xa0YZLMU0ZcumTaWCqfWFthhLcW3godpMX3n6s9fTRNzolsYJNkXNt9dg+Km18kyh+
0FONeRT+EkHXVHANAQOEIVoyybSZvoAkkXLmcdKKtjMG9BCdHdPB0EPRsbwspaEoA7ZaxcYWSvU6
EtpK/1mFH5bDK4rHU900ohDO6xckmfUTb5TdJJGI7gct3PKFwt2kDYoCAofHk8asWsZRtNo5HPVb
rz1BVD5L+htIZSUDyLAhBHpiKuDi4zfUILRwQkZAkOLB/cjwjlhh95cFzPTeP6A2waR4guXeoWra
8Ptl/6aJlxMQy4d+wzuWKR7aa3u//fC/nN75AoDQJzavGZjd1owObelBYa1EbVy5sK6BWlAjym+W
6CqG48EPjQZKoRmgeiWRPbNCBiMAY54fSpUCakNtvjWZ8LaXgBG00FCLsNUc0FVDp8UQS8ifNAK1
9Mq+qOBYM32Lh3/8sd9R/SygLCY+qzndwBNyxGhtDUQiVPIbNdM2BWievUVQl/1lnvrkgVzIqfHj
hbkHj2vsqFj9p4V6wHjCcIPKgFz8rCWj4vfQ6kGBkfuLkl+Y62sMbeo/EtNBmFwiHcRQiGCVNZ5z
3yWj2jo2TE44ZDuTQHNKdMIHOr5M9fln6X3u20vehUfyg50IRbHm+bF3JYrGXzmlGmMSTRX43GdX
y4p7J93m5j5KHltyoxc/rDBM+6k5oxFh342n+RobAwD5sf10wftxFLX8dlDLbWzbROX274u8K1w4
fQWAlVi6idhYxRoUAoOfjxbhHNJ0PmivUiLcdQqEHHiBtC/B/3slcX4xB/JeiKb0As6/gIk+94zA
u4usq3KmLmrFtmrcOeCJ7mAdRJoQYi2TfbpkkXUcpHzfoubQCdxCVH5mJmH73hWZpamruBgcbE11
bjjZ8VgdWc1q0kmEmTLicvfxwUV/sSr01l0mjw+dUkEBj31GD1CSmMepuQQW3ZgBIc/9gP6/S+SV
RTqRV9eoAcDNO1gdkkOhR6FHWn1oOxltJpuC48BY+SEGj5dU7vf626vFEIyZqoi6nvhDK4VJeFrd
JrJqjtMW2+Bz8a2ReA9YXN0F35XBhsX73v6h61fjYprb4PGlKw3dm8kLIvKjFLa+kOD1z02o1YVI
2A2f9cNEbnwr8K6pJU7vkqtVL3LNw07vCh8Hg9R/Ue/YYKh0pbw72KtX3b7W8mCGP9M8IM3K3CZu
heUjAajEJ6JQHUS4Ggf5ieG2ZypwBzbS2PIk3QkFJnxx0Eh+7DE/vxhsIXZ9I+Znr0o8OgWKmjpx
REQRPXc/Y8JXgZ39i3JPK+zRoT4/LiQptcwByDpfKfxqEiK2e+n1RjVsQBzcQ1Pe0/2M/J3lM7p1
qlUHdTCX+a3ajfR29cWIb/9A5gABTW4AnnrTy68ki4um1VO++h/egY+gZt7aGKc81VvLtezSyEBO
wUu4DBrRq2vGB8tnU7x83Y7wOnRoIr+2/4AXJH5wIUJagtgYNW+qcVKbq7IjrmZYIzL1Hom4MQck
o5/issewkAZIVnBGB3hafRmyVWdrhmAjfJHzg6W1g27E9XKVXmDqyQ6oYgrq1wqmuI5kpBcZRYQM
ZLMdjBhOXkGmJTiXJj+nPxGX5mQMwnGocBvw9tZ9qYea8R8hxN8UZ5bT7MZlh9MeLvSnyO5NLyGS
iA7l/IKyUizW5lUSQ0fZ8AQmQelwkJDkoyXDAeQsQwTYITYGqsRMHRm0hwa4jf9zQcNdZw8L76wf
7j0/2p3NCXX/WhzB/oTkHkOQEAamKihV7rEAINXNe2ZZii6y1afM6x08vxjuy0fruxitVg/B9mv+
RQKlTwd7V5ChFXGQ5SWMC+MMALHhvq/oO4D+33o1rFIW4Uvv5X/wB6UDAi3TER/pmFr+Dtsy0skL
/uGT2IUCCwEd93FURvw30Pbg88kncvX3bhUFRKF3SPB3gIY6UPzb+tUp2rpBUxNJqqV4zIw1rcqI
rT1EPyc0tXi/quv5IOveij1eDMzpXx6y5tD2QfSg2lpyHQmo3uKJ9CZtNSlGT2v974mvVOMfXiyn
kK2cUWdg+c9ZPFB1eQrVg3LMk8SE+qmhVtH5FvrXk0/48rlCYXRd1qXGI2OSbsym0zuN9OITRZ9W
1i27QnHN2FJBs+HmS2QRjKOxXcw0nXElqO5reesC8SZPJzac1TOxuvkmvbZQNInYayyZcLRjaokr
AqHCPIbcR94xiHCyjQ/0B3gni5IvU0gM/fmRSqXDLkvghksEwAIXbaJSvTd9PFoNcMT8qJB9TH1U
mTyT/IwZYcU2ruFhbEw09bzYQ41GawJXCR5egQa+NTggtbdjeMy0bCdTivqnt79UtJZpBUoWK8qA
ZnXcJMv80CXleV+RsW89u1DYeClfBOYqnBSeg9wppyX0iLcWYCxxkPfoWZv0Iw1ehWYENycn7W6e
5PwK9Z+gOFR6wqIoh3xjy/IGsEhCJn7wFpfIbyzifQBM6rrmKoc6UumSVa3ROxL5U7GhWhvdkyHH
7RaN/fZ6qSzkE++U98aMRAXd0u2MhpE9Bi4yTFjlL270SE2wxx2FpjBxhIIxmxfSPOsVOKNpGnhd
CHsnFhxWDOqOPYzHKbV2uIpb0OFM4vcQsM03lnemQFsocmOaLtGAKvwfVksFWQqCe566VLKF4/Ta
lCrNKIAMb4/vhAaVF5ATA6ao7CMXzXp0BA2xuXl7YFivtGDETp5lg5NE95R8BJzSqKHfRlwC3R41
jG6UTJ0muttMnzGX2kT0/gZkg4vaEr4AJtrUd0mRL1Q3H/zcjWEpvYCpEC4VnPlWG+X1QUpAm7oi
ra4dYqyNlATyn6A8gS6eHoyLXiQt03HBgCCXReuZQkTdIee5FyzEpsHYkWINSY3CcdgzzVHoepvC
SOlAhYZhrR1NMpOgvgBuWA1Za2ydPnM7eSuidGLPt1C3i5V07OKXQjDDMZu55EnCZGaeXaU8y7Y4
Hge8tgCoeNMAbIycWLSxpSHbu6lhYLsbqbcNHNFeXFL5+ud/ZSCwUhher7FZy/qQdKvhVMsUg/up
jrSeE5E0KU+KxuWpPTTI4nnYz0gAKNGBGH0Bzbo/Iv48GvX6Lnm7w5Sz4FjCWR+cONfHe1DG/Bof
n3zp4AAHl5y5klFD2F9wbxMjwzYavJb71soMG2f6P7SgDY+tqIFS7/9+JXjzIXbyJ1Fk4dEUNPTi
ePT5PM7FSGUui1wtLoXx+xpE7/fmrEjKhHgdwbN9NZ3W8j4ZqctjZ3CiHIDAZuA9nWC0293SmKPh
uTTY4R9bNzTRgDP1SMO/32TzJCi+sN1yCSf8pe3r0+meuo2Ri9Fx7huBpWnFTW3b8S2hI9VQDYoR
FtmC/NjpxygX84mM0Gt94A3eD3Dcl3rXC+B1CvyUpkK/LlnGADvBqNEjNmzAbmlvl3KE6UppjQvY
pJXbdCqebZjSYs8o5HB/RfgTC2CfehHx76dMjach736dxwsqM6MCjmRR0R5lIvahcKh8i5IFtrEq
MGvM+5O3W1UBkr8oZYOW/o7bjFSNVeeWUOPRZo2ddXdk1Qhesgud7id+5uxuvc1+uJYesu5OZm90
ZKJ00llxGqq7lrPgsR/WZ4bxtjl2Qo+SlMyZAvquB0sbrqItCVgDhkak6cZpUaVaK5t72ltN/AMg
ipAaUvpovkxHXdNrWCuFfG0X5jBw8GO7HNmdjm/CIfkn3BzDZ6outGPE1mYsMY3jQJgaoEXMsqx2
Lugg/1ILn3BldQCEB1utdrvVurSRa8klTYpCSf1NuLSCZ/8439nhnMo7tFRGPJmQhvs+gCsgC865
/8W3Lj8/dOYkr9ThRQrJqf5bvrsNkXr4eA92tB3Z5OWeYdyThXpUID+G+F/efIalKcjs9t8t0vnx
MOKPrnI4sekg9La+io/WYVK521CLuNbpxOF5qW9NI51NC9Nh/OzMswxPszQuXTLZEEZsOumbTKC7
uE25QaWJxl+wQYYTq4/9LOdb9TPajQ40enUaQuFLkyrW8PcvOvYmnmb/kWFryysWq1bxLuHNkAnk
lgGUX8h/Vl7Nf0D0Jso3jHiCSeowtHq6fbFg2MsCBNuJpiAyVnLi02EVTGOv98VU+tCAxCQGgdkT
OfxqjWtxVmkR+t0WA52XRM2xUd822ZkufH5qYzr/DKKrq3VsRyGNJ3OCjGungDlX+7ugbBBh+3nE
JbLa6AJi04OUXU4inxtyxNv/xJBYMWH3ozBQMyEWQAnK2BVBw5KCMydVn6vNrfh0eykDHHrVEkcD
jjoe2V+6DByLFN9rlJrnjeekO2M2GvLq6+KMTnl1Pq91KmnMiB27Vu9KDU2eKh7aPRaTScPfp9l9
5vzr2t8m/k8uc1fo6ndcrfKyBcQyffJW74zRcMlgk3hOgnbWQPIn0HPrhh/CcrnjM7jwFWNxRI+d
NkPQs5vEzFS75Xxy7U3ndwAlS4ijgjr+Wdejj61AIZr2J+E49plzAzwdrxkvrE0FKRRMGK74MR/Z
EcktgNP45gUlaABjhIm/51lIL/4TPA/6D7eIqD4TAVgn16xM9E6oG9IUf/qlj9JiDYlvE5M6IiZb
LrZvBGOmrFzJLIRYEorbGJM2sshaKQy6sPENQHjMxdSDry62YjAUhjyARwHu5ygR0Ohs+QmAt4xs
kNA991fLRj2PX6Bj7T9QyMccsprw/lju51Qsy9KvfC9XyR15ndpfKYBovSWUmW2/LOiPT5Vv0GDr
4RM5QQBaXtA7WpoCbo4N3QqA536ICyWV3l/6kFAuhOPjwqjaPtWZtaDxnKRHAvhI6W8et+9Hkx5j
U5AebmXCt3fXNPVaZfYtdzMcJB7QScwfs4atGumxpOcg1/S6hDhvInodki45ig1mS14exxysgeOp
mfmspQwHC/ikNUC6GfoOiOZLMnfMZ9NBRKeENZ9lPlY5OczBa0kAadX5jvU509+C5iuszWlWqiII
PlcmWSXg0BtzAMCEsS5//qQ+K6lNfLYt7s7ynBxIGM5iZJ1Eqy+BHlKAVwW00MWjaX9dYs+UCpaq
f8JAV/O2Uq79ZVvsnUL2yTGrFjeuIBoCpuyLer7J/u5mrnDT9odoWIm357x9pjZyWFhCxBjPphjz
J94m5o5d8L2invMMX507cj+w6s5Qo3U0lfcrHv8sB8i9BPngAOdh0+AMZ9fRMbjEL5eLhkk3FEar
f3tmr0/MugTwHFpki0144zBWmg5/+zc4RbZdaiIAT2+2BsLKDVy/EYnKPTmTt/0w/JDHzUCJxjDC
D7/jkglDuf3SMjWt9fHbuwPaZD9OfGvXInVYxp2bGJdiA8R6OYfFYmM73oyPNZh8WchOPFO//d9E
qsjb401FmZNN8zWUfIvaS9Oe1Bs/0ZiPzYCe0zwKQccQ/3UZDXTfLZiUcOv1Djx17Igbp92XYmYC
SJoorSk1xmh0ddzGgLfPA9sOpDjaauAB/IlhNQV6AgKKJ1dzw+2cVu0AICU8f3ikrWDynBMTPt3R
QadKe89/utjvaCrlx8lxceJRscFIpu2HbNQ/TzLFPheTowJ1VXIf3/EHsQF2rP0PzxjEeBSXI8OB
0gUj2gMB51te/4QrqT000+pXvCY//kGb6QhJpZVqsj/sUeWJLUyiH0T/dXunpcZe74Wef3yQh8RB
9VQuzQcEBThVl9bkkB7KIME+LIoHgzrPtfApYKpODv+xoneer3S018gFTVTu7UfEfCFfGqfevpqO
fuNmMMRroJV4htQdAC77kd9qdxXRXgbamssRvd90aJBJWzuREReewSZADJ1k6pqJ4PzQ7V4KCSoI
SatU3hHewu1n4SkH9dqYqB4SrH4QTLO1beGvs4ALHuIKzV/kMxegHqd/6ZkHu0joSQ29angnZLOB
qh9xWM6igDB3OoI8K7HKG3dy39aHdoIATVwlfLLQonLgKdvOY7jjPxp+I2o2dvAKokPz4o2lBmvm
JVx3/xhzdbzxQJS9BNAVO2LzrbaqxKQ+DVDKOj/spAXgFvU+T9cwPU9WIcRBpIpmjfBURPhHyKZu
t74/3cTHD1QqmzqPQxntnnWTUzccisDTvDONYcR61Hp5x9ITseZm1y4t396q/um0xlxwRSzqa5jU
NX9WWdfFOWHz0LbrotfXpLLVjpxp/YD2N07XuQ5lljSULnD3lZ/MWJCazWkYhMjtFri/Z7atU+nb
s1UnY/b1Mg4od5XmBH1KE8dZd/jowevPhgk3D8mKqDgg6KZj941k5OYcaONctHyMhFY/ALKa2/rf
0cVqL2kEcFz3MU97UbIJlNXr1fyO6bd4YcpBWC/WamoCPDnt8v3FDfixg0ybs6Ed1zoxWE8rhkor
1PwamSELsJs6mfk6M2BG9LJDixGD3n7RfPlq75KlUeYOBh0troC44apEAL+js5LQMK4m2cVWb5AW
hHKfa/vSCZYIV5IVeZCFFc+m0KTpRVFACLa8noUPG/Hdq0+sTL7+oaEpBXi9iJIH82toNYkbt2MQ
EgR49MJSw0Zi8KpzCWG7tlS61+ZtKIfUrkDwBzWbTtmubQ/plIDil1s/LrGiWWLH+0pNQhp0zRSR
1SbFlL2Y0EW2G2aK8jSnM8DvPx9T9OX+HiRUsZ2BZeniaWYR/wbnHTVXXSxh/d8ub4jQbgUnyGdR
RaWOfeX+u+GlIlKlZtlT4mnjWteG7F7ai9hpeCbs9DyGcyZhnoLGl/bwK66O8OjJzWNZfu2Tlc83
RYaFi9OJRfA7TCktcBbUSIOzh2ap1KbQoYqAuNhdp7ttW+aUHG5mnVdCTaRfxUQtzAcxwGW4VKE7
zK7khsdNHMGScL8cEwBcxaBbSEO10Qq9N3WN+PsZhQsnkDDdBG3iJk1v06e4TbY4tlZbHnkJWbwH
Pi8QQiNGu58jX0hsUO4E9O9/llwpUgiYA3F6juLemwfk12TN4Lst1/o4Nsa1Eo2+qeW/HtKYHBbR
7liQp5HBr1m1LROMHL/4y5dJZRxc1iPRzKh9pfTwD9J3kMEt5fmJoEXypA5MvrvjO1RNxbfdZ2Bp
1XTPBWoIEp3ovjS9HT1Ozg3UHX08GrU07bLx2xsWbjzTkmmH5W9f54jUouqHtQPLwdkP65gyANNr
9ujDq5nUYln8C4w0QiU1wxSwNAqhn1i7lBU4zn1Dn4JVKkMAyNNfuw2or6fXvK0Cvm83mVpClVrZ
TCkm9H89K7Oxk7ehvQZCWBldYteUt8JCRXbTVBOvu6EN4EIx8ACRaQbBuJLjcUrE9zD2coBOaTDP
cn1zdIORGwm4v1owom5uK8NpeXGMVZERk0rO6hiehFRuPr0rvjzpuHeH/WpYxeQ0hHLwjEzQe5DV
AEHXj69g5aIv610GyUhbyZLOts61WaXSwpoPke9RVAK3iWAvWl+9cxUZwwo3LuHd6DQ+n1NYh3Ge
ccP1V3d6bnvq+hpB1hCjHtrvvtecIArz2YdzSLIp9QO+VLr8t8suc8KTVGB8ddj1DKL3MGSkgy0j
2tMK1VP+Jmc25aCUyokkusE5fA2ZlqyFJTuAoUbXbyMMjOkQ4LNYxAM9GP2qa8J78lf4ger71nqT
Q1m7JogZtsc8WHV3GmkGm6Z3FYlJyCtthma+nuqKiQZJthWyMYaQJ/EoyZ1NaZaQkJpwf0Qy/VlD
z+MEtNw6u0WCoWLpqMwpnaBPRYZWI2ncUQ879bofB7OUCuA+LeZQjSvgMB2GOLwa7Aw7y78AlTUb
WnPFRPmR/0UVWXvgxsATkcsjqf8KOZyrRMhJKTbmGh4e7BkNdjftPbyTAo8HBT279pyvcdZtGbn+
4oYV+mYILWi4iVLzdKiAnMoLMPGj3v/Lo66ttKoaIpQ41vvAP3DPFvSOq1FldCfSIBs9rIjsejXL
oZq97Jp1HBtmzUBLOwDof3dJqsPzz5La71RptMl7KOBEkoCKOZXVLGVpSpKd7ZrRAkRxBzKX3+ed
EI75pu4h5eKQg8MLNaAzvoBFqoalkvhPLzqGoQL5bWxCL4jgSslxGByBWkOpldZgLVv87/xXcU4o
YQeXf7yOc7WRWbEjdfuRbKh2vB/NthC8uihEM5mY+FtGl1RgY/Ral55rOWwJKyvWAMX/xAXtdLKJ
9oi931PeTwkN7INRfPei8oi2U9iZ1fsQxdpLy1ddSvoFkYfn+RKAdBaCBTLJBtbCDfyWWZwXv6Rn
UUuxI4/RHMXZHu3M/4CYT+M2/3KKcd2o18U8VUX7szSOpQQUZgjUvLnH/q5RzqvYMaVSaj8Uvu3s
yjeygVFay+0gnAcCwsDGnaiHeiCI+b6pIN9YqyVnmmqMMIvtTEb/ehHoOUZbaLpsqUlZl5I/6q9F
bUQNbEphNsHGBKR29m/X9FPu9aG6YNiw7ds2AiGtRsjl8dvZBmcmt1XjvlZ8SCpskNGONDEbMHpt
I91V4ULoyH5zPxc/Y8X75HJyQ/82EFh9vO+M4wG+BKfB6pOnvVd8LWEvdBSBsWPm5pi0gYEAQtpd
yDrV4h7sCI4E06T4RvK8Xtf97Djko2cOOjs/y6MjpitF/DrJy/f89OaZfJkY5n8iE2Cnv4x/k69g
eq2yFVen0sKSS+OCZenyFlQ/GzkEcDb6Vd09GkouWALC0D/X8e0d3eoSbwXqcQ05D9qj1v3u9vZ/
QWYPiZXIyXRM1B2shcOYWxIjFjN8glneW0AUePQbmISP6KJP42jK7264WoSUdEyAYFSY4wjuR1SU
N3VW+0EV3MMsP5PkpmNSR6sbn4dzQdnuuko6nxX02NreeBqe0XL98evY3Du5P0a5N8vUoQhyW25k
OQAMSkAgZM1TdP5Y9OnAHaxJfkVKXqKvHtZWK4kLY9Uv5ilMauDON0nInsqR565OcULQYUyyrcff
LtLRj8cPp8/Gh57aclfmiCk2/AzexGvXD2xXblfLtukVOTy1ttgsV28qLiYyNIRX3x6313FRPKFG
tLY5nw7vZ4AeiNNZjof/MVTSz6iy7uZ16Sz2m3Ow2w4dvzwVA3L9BczOkECecG3xX7pHqYBllCVo
SczF7BsRDZdbjukjqpOhd2A5rBjyGkulH10XiYkFWL9InHyppP9B6UubtRRlk++G+Tm0wDjKPCQH
RFeWM97oqjsXPkLEDZa9os9b7rdYFszq42TEjRsYx3FUIcxIkUu0wnGf+stWUq0IJr/sb0dCmWsn
1crSP0+cLG6NVNNvNgkRtz28SOpQgCwCSqTg5xY+UoFvCWjQqDEGiR9MQksm9KfPGP4YrWxS0BYV
Bddxl+FReYYETM/1Ahit7TnKm7Mwi9n9CuqJHyDkn6samL1sibxO4aLbOBEhNOPaWyGEjkWN7kAF
ecWCgq++0mH2NDfpizDWaa1L37CrJhQLKRuxg0iUxhsevgYjNE+SiVFE1Ipnx7LIe55IVwyKjd9i
4dxuWP34TNYQMkdWDHn1DkzhM7AwD7LhzV6z+su7qyBBzpC7FVpRkL3M9OCsfwzyy5mQ5tZg5/bf
/9+fEzSkkyHyVQkUNBSUsGd6pZMYGy58/bv72P8qE3XqzJP9VGxfxliRFwnLwjLhU0QA8h5vOz3U
YpgeXhidFLJqMZfPylok5PLl9kV3fVJxxPGDJeHwfEHG5q3nlpblpzCdXWozKiDry/1lgV7xPW7l
G4+a543Np/bgeGpOHAr5VD9DeIfqRu+jvvA7MxdLJh+hDDWWvJTMmyvqvT1lOoTpcJ2IK4863+kj
/rZqWb7Zy0QDXPbpcOr5PLEN9oBOCJ1SQ+S2/CwlW7pnXneze4sAMFah4IY+qSCvcp4yvxF1wjMR
dYZZuEm1gq3YkjR1+bNE/hsFFauVBI4X/e7Lfm/p3XnYWaIU6OXL6ftjmyNgtEwwkMvjLiN5KDV7
Zp0hNidpKNmarHp3qgqJVoe67qW0mW/Zn8SP6F4IYlqZ1vmGOs3+Q/m8qIvQapkacLcI6R+yRAY+
gEqWjCYdtz0oq0FZqRNCFtxQXqyDST1ZSlVqIUmiA/mTxcOik2GXzAhgn/5ksb/AGuK2Erdeirjh
cOyvctP0lbQZ4Guw2+hZPZSCi+zNjmhU6hEPYzhvFlzYMqgkA8RaJnOUUVvnSsElQHS+92at2G1G
TTXx2yIZaYA/IkyuCVfILAnlJwSVuapPJMdlEGmrjGwsFV5X2O0sPPgQLKv4RmoYib2gwWdUix4l
SoWP0w5hDoLmGtDL9ILjPz3aGcuQ4NhNBOd+yHAkWwsDMHCUlsoTA5zjSiW47MD6Q/vsYY7Z0V9R
6pW8LqGVA1SlBnJypCyjqN0N6Pa3iJviKPCGmXtd10YT5wxziUCVXDRSmY6/Pc7ZrCcgOXt3aM/9
xtCoXhGShrStO5WbBZXnRk+Sp8l28Raae70jD86WdFXHT1NNuOTZGFAT6l1IF4crXmjRMQOgUHDx
C01khYrcpU7d2T6PzgCGTTUmzl5U24BadOTwdh6L/n6BaMDSW3GpLhqUFTbx4bon5EiXKYcoY1hM
S33o9yQfZQno5zvaz6zelCgoKONDMcKPnuZ+1f+G7plUaKLuCfh2fhfY64i7wqCyuorB3SiULNWg
miBl4kKPSaeXgyJ+pvaVwKuMQUv3HDcUPgjYppBqlspNoYFwuQhhrLWdKhmMiTqVjFLuVuONBrfd
n+bc8eF46aUqT/fi/EpnzeFUrlcG/UhgO638SFDcU7dLANmKBccZFStUYayd4NeV4KD8W2cdNUY4
oPbIv9YC9T94qYsoaoc1X9Eb7UIw4INELzCSBPtq+a1n3QDMGHRBJFiD4oB+r4XB+HJErlpB3u8m
kvBFIUZFIrP9CbOf5yy217j+SVmxJ5xF4JKtSwtaoIxmllif7Zp/RPeiSySAoJ5oIDKb4dU3lzOY
29yO9Kq+5vtqluv+rCNY8Wwo/GFCPSh+FPzURemNYusHLOXZmBfDpjd49sP0LLuDwxZOJL1fIMNl
Y+gy6JUR5odeN9byRk2tdfVzfQ2kqSxIH1UIsT6HwD35JWNQdUXXRBmdNaLTap+3/ozcgs8MNYA+
WkUnR/ZBY87G6eoVfXgVUak7vqJFMKxKb30J3E1uzk0vgj11U/TPYT4WsnPcYXsXlwHENZKU3cNE
hEo3SYRQstTBnnBBI0bN1FJ3J59PH5j3ycv8dtHTPAk/N6siPGP//UMqPMyAdPG2yt/CTxeTlN5W
QmtSH4JEq5M0XWGtVJHsGHZDUt/jW+xL6d2GcNx0HYmE4VG97xszkMVxS7bp+URUXL04Ayds4KoB
kWUvCikGvLl4ORKXlCOfPYWKOFu73DhxkrMVVEVTRu8fNlYLEYnPd/SZcvVbiDBtxZjhXqQM5x5x
JJsb81FZdHe2Y2a4W7dDULzxJmRUCgC156y9gnQ0P8MWFh0032n+kXAPMivHY+1v29IR7igmh6xp
tuEI+D4NJHetJQNy9hLppQrf+AbPTRx1gbAD0KvLietGBHtiJVoTNUa5yTWzwxi3TWUzGcU5CFbx
a84CAvkxjPxAG8Aj5VUUTygAUfe8N4tNVq6SCDGCnkPC5KuJ7GJvtW2eo6K4xRCOrFDGQ3VT93Z3
60gobCiMfkeOv25i2VbptESHrM9p74onAE4Sk5tUnFKqU5PwZj3J7GJ65RrrjiyfshlHZbvnihqW
6dEZ4qlEhYghoDk4LwSR/fadkHvsBQmOUjVHaxySj8wzY3toYS9sUOUDosKGyRq/HxEWHeKYoQn4
1jKENPTNqt7VMdK2EywnDBBP+Txrh6y79tCh8A5ElIdWxzIykX2FqA44d4+4M7OrjdA8PLEA9ieb
EE0jXa6hwFuz6oEH3OW3Qh3+uZY8VyVtMvnybsO0XmLRWua4PgJUHAiHjkmv3wFR1eb96ckOrVW7
TucolEggUx3pWsIPpJywQN1GdPcXyVs1dEi/PzFIi4kMoB52K2rV2Ks2k1brdEYR2gIf7wTDJwto
nfICRxrRZY1PE8uZGe5F68s/jQ+/YInNdhRW5O0jnCSMRvQS8/OmvzRHiAazSz8zpnOM3JsDCS66
aAkwDEPrgve/t0kBCTct8Cz1WsCdOSN8woSpc45rNYgoh4ZTXzR/gu3Kev61EZeI5porwkGRjgpD
OYVn8l3trxIdfqYCypf3tq+vM0b1rFeKsepfBKILdmQxHAHlAbeMzRHZXG7zn9z36EunSjjJyi0d
IhZrpTYVMhY6dcJQV+Baervsh0U3ULV5X0GUzlodGKv1Dm8ZLCd7R77z1BlFMf+t8o/7EgPhO/sG
5LucTCPxrqAkbhLnAmdjQQH9XjOWdePgVCIP4qq0YGmYJ2xEQzL/qV7RyeRAMXz56sXM9ohhbdIJ
AeYNUJaunBWIR83uwsjL6tcCnaJG/SRQ3Sezdbo7a9N74Xn0wLk1V6YwB07jEjgLqHwmDJPiazvA
mIGy2kOEdZQV7887pcRCimH+sYygv2puAOZZhSo2O57R/9yAD+ILaWrdQGR/YPaFInWSV/llCi39
4ksBF6ScK5FKK6jbkDD2J1W7VdOkFitY/otvCmKRb/ssS2KUoUxIW/CQRxmWtB8hpDQ8jr8YSCqt
MUBb9CVQwUoOtEzJZKMGzmKLs92+QDLgUD/Wm0CAmFYogzYiYlQ3UW6ZUw40pNFh0SxleobosIql
EKeb/ecWHdjnVDsEbb7VVZAsilOriKW5D8Dp7H75gdCExvsUsdpkVzCz5v/s2/sQxrR+DG1rpYwE
2VSukKkR0LUsoB6OJB+vmPu516FQTMXyS+pCHFo6RIrIO9nqREqDxDpQddFDD8OayITHTrVC0TBA
2R9ALGIeW6wGh10vN8g/XFEkkBHhvmMOxYvBeXhrAlBPKr+oADqDvDnjP11AbFTL/niC0YRKKsh1
WWbpgRmNaerN5OeIo96Z/SSbYCBjgKL0I74WH4GJ2v69koIX+K8ct1QjHny2zMcfJZonwZlMaQXR
zlcaJQg63Gpyqdlc3BdWhH3bGB5TaI1gQ3dc2iSm/Dj0GrziMQDU3lHaEJINHUTFwfmsdHd6uc71
uReYbhI9L1AhZf8f8jgv3EF9D+w+DI6pQMb+HaxDqnF6m9/M864wkyZCXzZViIhpWp2T7IeCECfH
taSHBauq8ZHAxi+/7VkKXY3NTADT4kwls3RXfXJDHF9XRAhdEECrtuUJ74BZacPt/UCcoZtw81tg
V3SoH0zmlfi7iHEgAflCcVaglCcQIZm0jQP0dyGj9JG4rA3ge5Cb30BToJZvFRP9Yv3y5ygrY3tE
R9TL8Cb5zr2/wCTpm74T0SAaGVU5kg9iR4xHms80drJVbeRUUTSecE+HxYfjy5RH/G3d3Or5rOVQ
d1H4YMjNNHdH/+q+BF8l8tSAktSP6Pqzd9tgEGFPI0YXa1jGCDeT7kJi1aR+zkBWD90njKafyxIg
9G7xOl0AZkI+OTbxbCV8c6ylI5Oum1PeW9/GOYUVS9X+Fx/ncMxM99kouwlt5RM4RUY2SO8BTTRm
4QtlUpELKY993xvG63U8WrOwiKoX/TrppLbx87hvnKu7lFq5XnosKldbGnEjtazn1zXHYTpfaZmw
sJ3iTDvuy2MSdjYvZcnyM/W/g0HpI/zrtpZJb9uhWbssMFh9QPq05b5bSeUoBnzoYaIZWGkpnzgC
shm3bkx/AOFIOia5wJ4HldVxsABTvM9XsNnvDvisYB4M1MLgtw5UEY+vv2c+l9DB9ziqyzYMkuSt
q6H237dCm2d8PjfUENVs3U2VNV0SuxxYAs+4pn7Nk6aJG9gvrbjYa65M66M38qS+zez9eIbizMBR
29AxbG+oc9xO7DFKay8AEDNiL/rEZXmC7engL5Fs1jzJyj368JBX/pUlnyQyfFDdRzo5mhg/GndC
EiQlSzyvisvLUfuOxtFQITJywIe3E9gJGzc+gjQsGP7wu+hFgl97T3Dsi0pLxiMonI4IPPFA+G77
1L1ASFz5HM7hL+MrqALWtm/y/WSUQWx9jI1NgXHb40OGkvKsaDoNsZQUZjfN5H35PeVmOKJjxzA/
1U1pOnmBOxxZpPEkYaxo4XZNk+fSZ7wbIO1PhD4guPZFfH66YY630iQM7HMLDE6btTAFrybPvvtr
2Bw7d8JtGoryQ8xVoFYKoOsfb1Q1gEIvDCnGP8lPfFBKG7/51ZsETBKNX1Nt9kWHQZ3hbkdHXzEP
Zzh3KSyAPvyTYdPFCTRqwtbaZhpRlPNKaINykHQe0LB2r0+6rhQMODSzEaqE2JqG6fofGbeIrKYs
c2eLI5ATxburOAmkOjoj+kWN3fsnTkxP8UIY3ZRheZlgbyb/R/k1WMZuL+HaowA7OliRqBSpxG9P
d8rzYg0kQ4cocSsh/tsJoOrkpaTtEwvPlstIuEYsRLfUkPh3ycuS/z1QDaeyOS5z72/Dow1DgCAo
FUgOXXbz8V1WEjdho9LWCCjNW7WfCDA81c3Sjgw4h4DOgftSc+FqiNYirW6GMljd851Ca/G/4vK7
Ii0Cp4yAsnnPItK9yAQsKjQZwWsuTOZDPcL3IlNk+j5+Ov7Ba/NY5ub3DTdznZ9o+hOTcz6+tM0Y
EjUE/pDSs1LzC0uJc4vvVOoKAfkiXVCks3MpvEyx9NmarKKgjw6/DqR/buqwQtkkariG+rRI4+wT
hdn6wwfokIDssO62Ss5f
`protect end_protected
