`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L7QXUHa+EKO3d9U1lByc/MlIKaA8hoGuMRU7SK0bjih0q4L0bhKN9mLV6juvon/DsSBgTbASQDzp
XjUIABdnsA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bVntC3V5hTnRNy5jl2xsvCSeeJuoGDgwLuLST+wn8IdrQ/NwFZizL/B3TlZDAisWeOVE7NtE712E
g/7YbbYPGFyDsJ33ap0iYxiSCmVrIMH6N1pRLiUQSa8deQqYXi6ZLcSynx4/VhXRXOjw1GIuaWP4
7bM1niXwXkEu6VQdTt4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m5P5oF8fWoOo2eqmes8S1kI3tnhVTxoj2C7SHK/+x0f3aNHd44dJElPtQNe8++stgziqASN/TLwv
qoIpiAEDfJKsHZ1leHdcRfuAUeqRI2cjhWS7pRHVGfFSvKKxkDxhaUfv0Zq+yQaKcuEAoFRaXw6b
xmB+5pgUmQtuEHvhjg9k2N7thmtgPsqW2Op4FW+rnowp37Auj8WXN/W3ylviLvkH0EXE+VtweEak
PmFCe9+hT4kG5xbj3UvnaB6HwpcHRSP1iWLkX/k3w80Ofx/gTGgbyCtUv8x1XW7aptfSwAaijd5b
AyjIAx+iwew75VN/VW3g09bZeuGeXy66zQ4A2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jM5h8bfBeppi5YZJSfABjcI9yI1ktEfvRORzdvd9oTHH0f/cou3dzwit+DcXDs6MZf7DDfhKMh2B
IGtchv6rXvRZ6M2wv1bskIAF8VCKmXrnFfYr5mRque5wmkwBYVg0WXCF1cEe+w3Fx/EQsEXd4NNy
upLu3LkUWcnh+iqHNx4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Be5+tuEiORBtxrRPAVW2gLIVJB8wW11O71rfRRnUk7uIzPg7SgInlX44eSrJwTbOxlxlEHBLpLwN
hMG89KzDC0Jk7g572fHVoZszRBV7zEt5MCNzLsL+nqIgdnKnvp0w9Cm1n4qrDk/vX7M75o+ekwb3
juklEkpM3BS50n1nfMxG4qiSpwbcCAigxZYjSX+3RC5mAtvUDTCn28WbtUgr+BFpzhYbpuu+eIzn
DuY8CAlEhGR905rSl/P8xTB2QF2DKCJATFSSQBRrFoRW1kqRlnH1E2m8aow6k7QKpdjLStGomr4L
ufRHA2eb126wPMn/r4l+csMwLmzGVqmGXUSNhw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20912)
`protect data_block
sbRX1ypEr7ivndxuCOsz/Ev8BIPUjp8BluEeylB5RDgNrzN0Bu9f/SpfDzdQ7P3yrG+PtlJfIwcg
6UUMHogUHy2/uLSs843RvfaTZsi0ILpvKoMzG712FK7s4SVuQfLICsqRCjWpIGZDuVWjyxwZgS6V
vZeuPA5JOVT0gPkORuT4OPzKdwM1vu+n1ese87YsHp/Q2tAHWtpf2EhI7IXSnUShzjmo9quFFm+o
pmdiQevKRQ1DLGdV3L5/MROXI34U6AQXSU9gj2xX6eirLVaJsrQacJblxYzlG0Rm3FcIltueau9j
7ABtQDNgtw3e1zT1odMUxQGST73UGnuCPaXX6XqYPn6PmfrSBhMcGYZixRveCqkc4DAc4CLfcb06
eDiUXCn6RVQrBaxKAF+9lDs81XCgu3WStuJdjxI8p6Ey73PmxVjii+u1mQBlZiJQCFJeHvg43ylA
qucDljeh92ImjR1JrgRld1TnRPPXr2iB++gxBaJ5HsQWO5PWY4MOiHVUQttV74A9GYEZ2Vhg5nPt
qCB/e500JFqtY4lBq+S6N12iGTbqnWzOiRV0CtlN8YR87xyo9uR4WeXYMvlYEf4kmgSsAUZOiqvF
XkHUU5p5LvsltYt7JhYjLynhb1ugjmFQhvARXEvjnVbZqVu41X3ElDMMFgWs/4xZmJlxk8PwWUup
RjuKChzTYYyZavPpwaA7i89evtqRA8eGdSZHNDHKLZGshrIVJlPnkl6h32U775s7J5C6VxlvHTXZ
v0Xb7xQ/pn1B4JsEjwzUgj6hKCLJT6c21cfA1a5kcS4W7xmbd3ZGHia7RRBoaRMwysSaVs04tgQX
i2wXDCKfxcpk4nui4FhXKytaIrLvf3irxwvDLg6DEtTFmSMLjE4vqY8Imut5EvncNCGj6XAyzlEK
rZFaOSJEdQWo1q+dch6LLxSKjdg37fkUqUrwF546KtpMdR5x11feEk7fT6vIG3uWuW/YGX2wCJRI
KWByxtxsv6wSwxEApskA91g9o3LriZictIbOdtyuvnL/jR4EY7yfz+hkQKKSl2DUoYKaosIcmcGm
1WpkOz19qUoZWotk9aKFEPoENWgCLm3Yoz7cBfGYu/tOzipKZDbsi6WGIdJPwnZEqGgt8KAkOj+A
JTE/peYaMV/sx19g+ZmLOi3doAXycyFej0ql+xpNnxsgVoipHWNDqVkjn6YDHbCR2iQH5tQiLDB6
Bq93CxejMZUbFv4kyHR0lk/yfNDm1di5pHwiE49PgFfLerLexLBGDG9sCAci0g2W90i/KwKiiCCU
7aCqkEBlpiCQFTqbwrt4rW2hhTuVTEzotTMbwCOH3aY68Of0iNEu3JyBoQ821EdqLeHSqul9ZRAq
dnJNkUZd4SDOK1xlu2Z6ZrjxndDmrfTiYVlOwLtdpPUZ3eop2fkussndB/1vAAc/UzI39hg3TNuR
ozlvqzTP6h2ds8Tl9ocutPQeMcAACxRnXOUbIMjRpO7+h8Uv9DDu/+/2pAtHNh6GFbR1Msx1EM6c
p2/fF5J+g+TZN4WcWUd1uAKACSxv2uZk3e3RXLC1v0RS4955Un3pgj2xRqeCX0nPMxrjdtTzyAna
b0ZMySfYUBEKmklWVX2Cdb9GQgBjcUvjKjhYkHhi5f6m9QK56iKa2cYhgDElxFSw9F3D6mj+Bk06
pdM9pl4Jgy2wOunJcXHKIdo2zodzed5vHu9iimQxhwzCmvmHG4EOh5F/QY+r0j0kNDLoLV0GG7/Q
mIOWl+eHnkfRUP+kdkNGseluWi12mxkpKgHt0lWN4ksZdzajE5g3XGVKrcqPEyTt8l96JWdVv8rP
Tre4sb6i1f2w1NuMrpZuuAOCz/BamZBF5hpY4GxYuFmlKMAq61Ny3wgJiDVr4JdDfU1OPiP1iUy8
JbfYn7o0gYQB5pkbs8/DrS9ne0Q7N/JI3Uk/mtfXW2aVl+rwkghXV+W247ePZMWry2YdwgemtfeE
wIxAUGJcj7V45Laezyn06aywx3Vi59C8RJIUYJ0zfgyIpFuUMWIr25C6bDzNZrWjbAzcfCSTDeQL
OZg+AxfTO3/uIDmJhUS5QKiCNhsRgIsI7iOtHe7yUBx0U5aunfLTQQMekMC8RK7MCi4jt2i3WNPE
MxjEBOj3Tx8Y6aBIyZH0lUbT89/37KbmlBAP2XhDeDw6Uk4dZrPY9WbIFw1/x7WtTL2mVOQlvz4G
KLAmYO6IuWJGr+AktN3d8l7fc1QbyzCVES2nLMQmklcne9GWVTsG5DyuCJk6TKKAlEItKM/U1AmZ
Pm+iyieFemD8RWRMfaiN3CG1BOrTluiEfy0SQjuNqa3cUupZskrnDIGhBtzoH7ayr6UkrZlNd/yA
oiAiP8MRledqwjT5bIOezu12nesjs1sc7Ce/8oTHefZrpb8dO4cisaF8o4JD9D6qL8V/eTTOsEmT
HpwZFCTdz0QFxlIlHcjyiP8NahpU7b7LqG5bxi/rBaMuWWkdn/n36/52ITXuJXQQJxxop97jFnWV
u+iFRTM6JIFc1LAaKPzVmzoXhIGsRlMK068S8VQXwqWUeVs4uSi81Z2mB/+FTg+WvWORL1NXJZk6
5HiBINXuPgvvv6Ki+h3eR68gzK+IqL1Z6JXhwQb2OmBJhwK4xKyn1KrRP6R3wXdv2oPcMzanXAmZ
odJVeRalAcNikKCu4J9CfdqWrR/TXzN3aFCpVTCZ9jhKS5H1eWre9hamkKPB+SfuewDkdKg6yykS
+noZaES9yJA000n8DboA4wLgWGD0FC+G2whsgmRd5s+ULzmbaUh173i+d/UgJ9jf2f3C4SddmIuI
Uql9YEKE92tHOm4JMV1V2FParpavaV5CYLQCbcCklEqBoRaa6FQHvti8/HWzsOjLGX+SMYWkXIXg
ZpxhRL4kP3iS5lIX9jdki4OW1WJuV1hmgbI6xysngp0PTr5MZtPKDd1rwJNQfrixRJ/CHMS/msgz
ILjhOiWFGLQ/80aODSC2bVuTNGxYPrVSV8u9YRdXlafQzl2CTiHI4s14tm1DqMIVuj4aY0gBQxEY
Mfyd0l7AoOsoUOhFBNEJvNYAa/Izvfc035vvyl3Wmy+SJQOxK2LewDnA5Qo5LsQ6/F843RPuYKSc
jKcC4/M7QszouqLAtoaFZHcI1Q2XmW9pzmBo2svqOs26/vhO+ifmKD5YyLGIkvY/CyXaza6DxmJ5
Bv1lWIBJmyfPnU/8vy9G5tMgHdDeIj3rccxfGCVVh5TVq8nd+/odY0X7LV17wMEdsTDa7HydeMoG
m8+t8lLSFTWdOHzCSVvT5GMGZtpuYM125uwS8TlLC4nmQN0YQND+85T/VwNAtCgVgSj794AMOmQ5
16oRbnBIy0M3oxC3m8SoKFM8cO8QTi6WcPvgslIGy/i2KAjWKNUXmSiS0ySvqOdDeVnwa/GT1id9
o7crhw64GbEw4CB7bTzyLNPhuhMasf6f4S9RWqlR2RBpq/ns2N/3r2Ta+m37pUY81ju+cCah3TrH
fSYzWm9Edu0wVwKCQKmewXI/J/HrfOXxT6Whb+uCH8zlAfbKX0xr3ZkSoZA/gzxaQ+R9qs1HOuPq
4SZTarPdntJHKpMhBY3LrMye2LN5buQem+i7agKoUCCDlZZ5xIDvU2PaDLP9zmGC03qUroupN4Nj
eKoVRc9RSafFZOelVVaPaA5TsXuir/845hUI1C1pYw7ARtOnDlOip066C3i0bGdRiKBrlDvwtRm6
a2EsIn2PJjhtb+56FNnz/hAEC0QRurY1rFCxhHH2kzT1elY+zAgMFAIu3siwUNeH2Nh/KdF7rzzG
QE6oLxHP7UpNJ25D90BPIJo6uTuRAnq7stgCyga3WmaujfO+TlZNqsHFaXkdGWTqoTG+JS/5RZVT
MBWIopLDJMDB57avtqGrPpL6jWRMhct2z2Eh4gLjVR8vqsLdFr5PGRVOwYJtZIbYdqFu+TBzUIpf
b8fQQn295P8W33blDZCosV5cd036ToBMaCslDg50rxOP3KnNTdqciN/PIwcLAgQcVHGjHargK0wR
j37j3HnBMNVva0S60e0R5keApZLm8BpCSr1OLqnoFl32rhMPFXoI/513jp1sCPx6/rmnXJnFEwSI
lpK6XVNqYPxaD8wpHyD6qtByW6GOYPZN8gwgq6VOvOH/ej8lO765pdPSQRt+8QcE2LrCa1/Y/lsx
2iKAIuLtCdch1W3qb0oWl5kcEaGGkEU53QjLIs8093FJH3VthOYXcc8VQpv4rzP89YiGjpbKbmb6
bmcQwwhV3UiXC29TJ3beVYe/omngqCyMMevJwzQ+YkcE9LbrXlIa0icww29/ZmcO6OwhmKqTKFi8
lL7Msc5ReIuyFwb/jOfbzj9THlwtuRP/3i7N2YDQTcuZa+8bWCWDSwMmXQ7YpP6A9yDf+rjk9Nh/
S59D3/q0plKCbmLj3HFJF9gPPtUgDrzALhQmtDcQ/8GCurVb8TyKq5PVepVj3riB18LPtstF86b3
qgEsimmNTIWk49o2S1Fb0Pu6IZL4dEaBYlXqCs8+w2p+9cI5T5F56ysBMtk61p/dPu0K/OzNFrEe
EPHVSyW0AWk7mQTohnG59hfeRpA82N8QmnciIAv/47JtfP8HVtB5oRgQwe9Zd279ZivJtPZSBIA/
W4Gq1/JPDQPNGVbheC2nS771GR/1gbfmwR9K2u99Bn7nIGvawrHFx28wTTHEQ2sEqoYrp+mDWElF
nZJUJo4jU3vIN16ZWiKkcbSUKZi67mO3mCFxhzrrNqVh7Wn4STqgvDeY0HWMahFVhOiyZ15Xn6Zv
+UIj9FK+i34e6/Nm0fUJgCIPMmc2HXzqo4yJ7E0RcQlLFxFB2Ozbr2ZcF07kmyNzXJ2kKJH5/2ZG
yw1RiZrRzQuZtNiGilfoL16sLRKao6AjVDpSL1ywL46noSBJp4DGvvhsVRM0cUl+HXyf76hOi6Sh
7eOtRT+A4dZoNsZjENmf1bUB15YKIEN9yoFvEtUu7hTuw6gwCw6idT20707e9UCuffenNsUzvbGh
HgsOfuHJZpw+cWH/7MCXuXg59ivrNp2h8OA87DfV1bimGjP3msmrwTKgS+W6FkHoxLYvFQHNflbB
FXlFbfZ+IvRDQFhzuu5IpXeh0QSwrFooe6N9awEUKoUJjxXLZSbFWu13Ek8iF4eGIYYTZOjf/9/9
Z4SyxPcJha0p6XZAG/vVKWXc8gOt9fXp6/nL7zLSg+UxFtzT801GfZ/zrPkEp6c+esRPzncPDv9b
h3NXjFDUtm0OEBuDHPEtRAsVCet2MLAccaLUMYO8hR2pe/HdPVFrBqvRP0idpJdyZYp8F4Y5hbvH
2nUdft6kPzfXaHrnNb+/hQ42MbtvDlpiRf8USb952OiS8Crp2r6CMxBhdqJir1ExQSqpc6Ih+9W2
/bzilRSSTV0EPbx55Acn561zRZFIagwlsT3z6fg+8nvTbFqYUWdh+aVZCe9unf1T2s1SZnS5wQxC
jGXlB/Te0d0s0kWnx+MEY+2KyYF/L8Ij6GFEsd+mCg18Gm6WXQu9/KE1f1Fe1q3byOtCnF0Wh4nA
rpGyr8n94af4V1ifxJAW2cy/X0M/jwXH/7MsbIZFSKTn0nwsGTLi355zghO6P6VgIuc0jqUY2vL6
iMte0QI1waPMV0uz/BPWvoe8/l2q90JZmMjriPT9N1eaEKtkvZXgAD2Qn55X2zygWZ7I5JpqOjMS
MqjCsUJb4/H4CiOgvF1B6sTw6tbAMyloSUUBbc9pw1vD1wZj/JGQZuQ1s3AvhRw4KI4kqQ8cxq6K
Hj9k4vxbZUPmKuexRx9PGGtn/Pd79SMb1iZJG/TS8pg+iXzhN9prp2k1YvTSNSKRkVs97Uiy0zNX
T7c59nnbCpxhGLCV31uiGelP4c/zB1dTAZtMwSmJnXZeCV7csHoErbzrseidjnUgxqydcwR7/6CX
sTV7yzJ3uf90tgmxcWiJa4/Fzj6zbQDAgcx4wQKnYfxNZ/fUzH+Bxh0HiQmYBdKl3u9dbatudUE8
a5p0hAE515Nzhy+ud+sHC77LrToKpSCfyxutIkgU/M9ZzU8HFGlqR30SVbAsPLVAv0Gdt0ywMD1g
47s5y9xkYEoCGWlIWYXtQmA3MjPGhWDcyP5OQ4Dmn7QsnkzrQaDF4tKeVP6w0Kvd2r+/ekoTzwNz
WcTTUzvBT+4KEbxibiKEwaHRaBMPC9T9F6uei4U3rqw2BU4fqNrCt9rGsmLFbE1SrORuOSesw59T
xigYEFDvyV8Nd0b1HEVMd88wthKxNzxfQid6yao/viacJ7f0M4AE1dpbS8Y9k88bF85HWeCYy0JJ
zOy0gWy+jMXQJr/djN109HbplDi1gQ4dTSFvKrCi9V1g80ZJoIANcsIKZNqeJVWVsrtIbUmiZaGb
Z51qOy/uS+NUVbVqmWEaD2ouLr1VFc3rtNU8oLzq8jdICp6DKRFspScdnXEaM+IzkC2aclDA0Dsw
k3VRqbCkWHTIpnnGuifQmgqikWrdOZ62hp3/BclkPhg2RNMiVClKTi320g+9nSBjLIPu9Je8czLO
8j4SpVp9vQ3F1ssHlLF1EojxF111E2njKETvuRdBbH1Oo8x110Yv81vTQ8JtXSYi9bmR/EMmVdv6
XOIBDPhZy/VLSrZPTFkNq2i2ub9bbgE4zUsGyHrRAoz/7ds8/39cKrPHDDqRjifznU81yUfYFsUd
p8OuV4zx3cu7P48QJU7666M+Gbdenr9Txh6yN0KCA8+p7nGv/u7FlOWseAGu8iJDKCW2SioOAu5h
yk1y+kippqQNLS3KS2l8cjH6311nAMZlVhCoED5DtjLEGfmv/JIva7OXVTWAzzyZ1LgIlltU1sHc
c/TXBFDgf2O3uiUxou9Ry6Dygzcnzqn8XEjDd/ZapPFez9/5i4RtVTrGZHw6H4YtWUWPIoRGgl7A
RxgN3VUtMno1lIYoYWqtt7aZ7W2dy4I9fkRHNxeGIkl1QO2LnMB3I0MHI59qyuBB6DMHgbQ2/gRs
N8IN6CYI440/U1Ch3IPTueXyjRq5rPrlUnPML24cV0Oxoqm/0Vq43EvuLudVu1wzO4tg64GgdRVq
mBrXgWlJXdY3WqJDS2M2Kzp44X6V2oh4mayMe2vcGczB/sbsE+YG9frllGen33wfGVrrjaTdD67J
9jMrbAvkv3jOlk1M5yMoJpwzWoSGDAMSS1TcM8blri/7fQ0euEkRK1RXEzteFP0XcuUaoL6+cTqh
2103FynQti1YGH68guqh13SmFkBVg9YZMEt0x3W+/8D9Ldm7myK5TgD4twfrMxPFRXQ5bhY9H+iB
tBT64cRLj2jOZw5i2v7fmUsZwf18d8jOaILySrfuvD7mQ9uK4VVAcc3oqDB2Tw3lBVGWTr2mi4+F
bEuiYeB1w/zh52+KM8bws31qaJm7KVZ74soCloARg9IzHPYa+K8vi/d0xkyjKjhsAtT6o4C4p0X8
Enzq2NG0JXr2Qy3CJerkBycDR6t0BirSNvQpotw1L5kOJe41Et9psfJ7Bsmz/J4dA2ohSOrnVKBU
G1iZ5BlxM4aXNmiIlJmpWpAQCOI8pBxbvlIDYO1xjgAlQphNhjH692RVzAJKTvvxGSNbeRtE2TMw
YzooctDf9djl6lDtWvfM9wtzOVX56q6t53H5trbGl/tVBysZWxjqmQUwETR47mlMm65KoMadYKuc
A5rnHeVkZB22fneCc90EDUWnHt2mSnKAW4OUhfo3FrCokx5Jt8VrIEAUrVKHS/7czFkan+TUNQqt
Vs7y1ZRZVCCptcBFzEG914X/YmubOnHfwGke4Z77Uzn1LqEyzyh5+82Ez59zMneQpmI9Ss7O5yyg
REbNI5T9EcAxjPn+4QCJxUOEf3PwDtQR7VUjZhjlfXFhVxH8KKF68abWBddYgj0C71wHl/rjGRnM
L0zyCz1W/FDYwDUOibrcXsI3G0bPD8zExV79o8i3ZWVV1ZPTerKRWeuFFULWEBuFvsRwhiCl6M0C
y3KWcuqPeReYVNqNv+TuRwbo4FP4CD5gnpTgR0nh+d/v7TrAoY1PkbVg8o3kXeHlpzqtA3k92ypq
1NHMv1UE2GeUpE2Xc9MFxd6oGQnIsngcuYgI1dP7gM+ErUIcSE5g9VzKfV50LcLjWVikfcb2NTJa
6ezMlhj7U2ZR3cEhwM+S2kTn46MPbydvwKbIS4iGdIlNU1NB131yCydxemL+ubaTJWY2iv9cGbOq
kJdPAbLF8+toPTKt0Y8OE7kS7qYERFbtodfh0f328kUw/CqJvYtJZziBWo3MjITqPMmoxE8rXnz5
MI3XtxVQUFaZI41kjLW5C9H+eRbyWUYDp3sNAJHQOzC2jKd0tOLqh9CVrhn8f+KDIXRNcISAWv/W
9qKPmKjpClxy0MK72qrmbgvP/wyHdgQyR5XOpTnwCJZo0D/V128+lWcVqJBufCO7lnBRDrK2BiQh
xjKY3s1zl2sfpT0lbtqjXoEhR4RUj3GSp4b9tBEk8HzwLDmxjKio6T83nvqDNPTgPHtXD6f+s/IL
vNN36qyhNznbzSDmPnkRKxOaVv0c5/4bqABZDOQectb5cO+yXIawQFbSJT/C6+lEB6gUteGOvVhf
KWFQ4pn+ZaCygFhibTg9eRDprfSHY+U8U4NCcs8D360RzdMA8JWjeGkxZoe8S/qjMQzdFXH2J8Ip
7r8pJPJi1jl15QzSkBI7lVLlKWhcp7ixmWD/y8rgtVkIOXm0Rn7bJTC3PkLZicaJd2Jw8AXUQZEM
YQy2ktyOBSf68efnTvkoRj0HGnfleHlLG7eCcxVleojlcotpF1Q0Q8OPVKk9gnBnp4mrOe7Wa9UD
9iVpuiesvzsIpMe9u/A88KAgZeMPkENW9pm2TdiOtt/b6kS/bP4j2bF5RMJk52fxJIHkyoTzC7Xk
umii4VPAJ9WvN++y5cvlTN1jWLcEUkXpmX73GI+FXsy0wyoyUSkCqDAxq+bakG7CDixsH0qHbx9O
P5KsNKDCizTwU/3dGtBo+2jtbqAZTNGqvFRnikz5hW44bXFdcrAfoCwYMSO5FFbJBloPb76/Bx8e
IQLFE2Ia4ErUHSl94OHOGdS6gB5RWvAWDE3zly2480yFGjBq5Nm8VCDoI1HYS+W6QX5QlpvzxQ5k
zkVIHMqyWQT7sNl0+N++QSM7KJSSaguX1MCUH0je0ebjkOQ8k15oa+DKwcjffZvdr3Pq7ysTDCN1
GaN+ZcTOtfixVTu24QWh8xIkp4GAB16zsVZgWyMXDwgTPw4LSMGTUmoouGGw2gZ2KnOY6RqPebM/
/blSf4pQsS4+tyeMQ58AvdDmtjqJ4dMNHDCJcsiF5UGa0+wQ8CRQ5uQDbW6F2rhqo3RhbXe1jU9J
WHga83gsAvuVcrz1/w59AMB7/Wl0WheCwOkdbo0LhLIBvs+uBtHOS0q84QmoDdsaj58Xno7gFal4
al4tGEwolpvzJdtfaVN+FU5vav42Xuv4FnWJbZMakeXrEz5L23doqVtyMWQnwx4BfL8R9b/T4iLZ
yqq/GcddnORdGwZ9FxB65TcoU+HVM4R96V2xSznofA9f5JgRSxEapEixJhnfGbSCNASVyRjc40Ph
9KO2TJQ7mBeoe2/zMn2a9sWqdZE+ZZJATvPFCi0irsRvNGTUQwJgzu1kv79cZPr0WAXi8lgLSlFY
sb2iUzMGom3ett7HEMh1uKI4v61dGtChFGtaicKBpLLNHdWrX1OtAqoE7QQOWDkkSRozn9gUb4AE
ObDLriLrpYwW72Y0juvgGn3tEIIu6MWFYksFofXTc/nlcTxoWDTEUh3MN/BPWRD5EN5lSJybfIPn
J2Wtj6//UrESuRw6wya/j5leP+vu624zMmgpX+CHxtMxVON8EnyZUzseHUdfyYzzGGWvCh1zjqCT
HQmPw/n5C6qcCqOGz4EBYLKUgGc6S/M1HxGUuMqQk5ROvK1FHsprSaowJyIOJ9maL1VKwtg1g6nA
sFlOiDKovIDvXg8NKqnUBzm3EgjUWA/vBzdKlBani5HPphnO/pP7NRVVorB1VK90yEyOX8Kk50dJ
wThlzbE0umnEwWv639g0ZG8IK/OUTCg+fvjsGjcf3CpOvYTTC5eo5CR8rgXw6mbJoDq+VPiZbY7I
rGGNwVPh6P/r1Rs63a2uiTXXpt7hrhUCMS2vNL9yhxTpQPi81EV3bB5zMb9cxpZkm8RegBoLPaB/
teY4EbWp+oh8A+azGfteaAZsLgS9EdTTrOT3YtIZ/75j663KODQleyIvVVuRno/lCypAFdxuwBuR
Vi/6nNLqISItkXioXHe4Tplo7w1c+RRG+07vAKwnYkXCc5sgO0dx/ZsGfS6eDQ1E+HusV7yXy37q
nJbdYYKi2DaG/DgQPt3InB7gXTYbJO/OHS7UJqisXr8rLVK8kHtkvRzMszH+/KQKnVB8xKmwJBOQ
3NVB8EyNCzQVb1HT/Wq48uTas90HCZROR4VAyAoeH9HrK0fhuHDvYm03QuSVbSw8WqxJEKaKrugu
nM5rBEEULB9kNDvSbu584muV9bg31ykqsfeyq4aC/J8oYA3t1NC3oC2lHtjvEBLsQ4rPZkFlYKza
S1Bnd9ixsXgL2IPXzcbEK6EVWYJ75WhMwKbt2YqyqI6IvqGcjt7HybwrUEmq3GEaJlJ+etFCdhul
K/NQHl03xI+COeG7EYB4bibxyDIRzzPIz8w7iNNc+k0uEHgVwQxdnlapxDkSOB1WPR6V/0hx3pM3
RnHeSkMB8fqUPa6gGJiDxyTvxx+ASJ+56a1l5dmqsySEvsNdnQ3egyVnFGmKqfC84erzlG2wdnb5
n3axMolTSlbJhPc/FrC2ReiQIdYmXofqTe0Gis46OTzcqAcH+ZXAd3azpQfGXf2uuK2CZzhYZtSS
pg+imaoGmNDfsmWxSrMIFHiD74f8QUL4QKKl0cGm8TyFHbaBm5XqNkESVLI06ozAAm1vttI+X8ee
r44HtpKTxtF87We33VhJ4t1Mt4nidE8T0UVlaNe0MTA0G7GMbNtnQsRBwmOcImRCl3Rr19CXdbn5
N+/0/yFxEJ16k4UGkWvGeVjKypAIz55L891+1zXDi84UEr4IOSxJjddXaGoKgi/uWSta4N3nX/bG
hpXD7/dKENpWK9u/dvLTMkQgSEI4AS9nus9QAqhz4eTS6Qa3q0tuxyfcL/emgHjAmi7exBjNig8o
PsWaMKyxCnNH8Z7jdgSmOhpQDIDLW/XoOZep/MO8PNGTvgy/vD6mC+YPIXjT7t/p4GLlQ9j+pCdq
nKFEJ39iFx8YwQtKWOE7Vm0elTsJvXXDprc6XwJjlJ+8vdtVlC+3JT7SeoMo9vG4xA7s4FZ/ODXI
BYBatIcmPMlP1/rixsaay08TG02hw6Zf53bI8jRRcUcAoOkrscOtsSae5cwsyvpkz28JzktuXT77
UeUmOoM0Uy3Zfv7I51FHbkZmOJEM1gXoDqqHV2vsqOBUmRXqU7m9+NoS0q6nhQLXQfDurQj3MozA
BjteJfcMphuMV+wOUgosePcFU9CcR++mbujqaDSGNysbXqzm4NwrKjbVpncQL4b6jLSS04gUd77I
f9HkWSAlwSiyquwiZtQZ0koiyLDo4hAYzqxEK8U2vvAoA9vMIl/JImhNjJnF712BImuj2KHzoZCL
7Tzzo8YWC/IKpRV0JK6h543ltkHVieCqAN48gavTOLUo9MHBSmiJrFR2MZHH9qhCod+V+4xDijn4
Fk2kKyYAVbaOe/ttc2glTfT7rNIOwTfRlKe+GzpSwmQYGFLw+PTTAorSj35Eotp8sJrCWO8lhidU
5eWPsNoQfztXJ3agwqS3kSYf/A/2Lkhdtq3oij3Stgjd8imYF6Dl+UzXD3e+KaPPfaCw8P7oluRN
rXIKJENZqZO6WsOjxR7Eo0YZrq7Y98jGjGkyhjZ5qcaaF4KUPSsS3n+n5odUbjNoRhw08BPZ1aaQ
GfqbUskxLWCfTe+1uV5aijIglGNe0DYp6SaXL/WLdtLToLPkUQFTOgOyQabfRAm9A5gmj7vEW0co
RodXCL8AnXDIytg0jzhm94007QGOkeH03ARNozdEoVqO3nRLCiecSB2hr6/7spXvF+A6UC1iakz0
5wR7sisiti/zvtOmWRqyXXprDFAJxmPO9UH3VijlbL8JBDc9T0CnHz5LR9Q0TE6DsSFmM0oAA4a9
8DMNz85NJt7gfpUg0UziCtWuQrqsl/5AF5xdB00m+vOnEnJlkJV+dVzldtEXe/STzTatmJe8Kqpx
sEK82uVnhEgqT1uqpEzoVN+k9sWgyCI++m6t46wGcHLVaTVbWcvtz+RZCH4s6iNAzp2GMHtMpSsw
rgo6o9wmCiyYDzzn31S/UXlSSoqaeHwiAmmqcd4ANtPloOhOV7wNaIxwKcrYlDC6UMCjclWI7K4T
sKg0gFLpFQaHS+w3pUUxq68R093t888PeeeuxPXLNXemnRFVh2s5Ms3O+vEEDcRg6SXO3NrVi1zK
XwC3Z5tARYlxDyNvLQPD/uJINNTcREgYhSX9fe5vGCVUG4gLDmWgCrgdklRY0/2cs2EMklsZtAxm
Kx8JFie9fxrHKEBaZ8AMmvuofyWcBTvmb+O/ldNacyyn30nScTaCpFUyJxt9qz97kg54EVXb1B+j
Q0doubS+41ESHFsuDCLkEfXU6jvHIDouQ43j9ZEejWvkJT5yt18+HLwC5YyQMB1WBorRU+0To+R8
cY3dAGlDMZoi8QDHqSlVCSI/mDOr5QYDhN1EmxoPy8xRaJpL+y/YaGkr5/k1Inb6G9dnDHMCXqEW
ki90msitR/96TOYxdF4yLeUOL6Ce7oCHIOgpv4FNL1QKx1tFqD1jbFWoO8wbD5GC+9nmFcnPLEzR
cdkZ3uZBjXD2dvtG3SW7w7Zb5fAMgs+q4OU0lf+rAEgn/Kx9+uS/GjyXwhn09rPp7iJAXtjJf5Pc
JjLFT/O2geXyKaoJdbzHp1emaFUaNtLC3f6LHFp6KX8N4eHETpuj/71smfBsP32O30cWgSrxPOEB
mTbr+MlDhCI09l8ukvV1HS7nhkKfPZn/pMrO280f34OSn3N8VGZyQ8zpMaNu92vyuv3Jt9262MYn
QybCfb9FLEeL9pHgGSq4rovUytr0JYGmWTQPbulWjrmgq0c7XDJ2lt5o2dRe3FIWFtC4GzPHoY2k
8j21edvS9ZGcBA0i91tSi7xsmSz5ROwukh/zRftR3W9F78uak9EKvAjTdLDcx7yDenXd/vtuuvd1
yKe0DmcTLIkUPX7sJQfYI5eQAn/PW/+cB3NoHx9Ou5yrRgL4Rq1KZprCWnrmRV+ylO7MwcTRgMSw
uSzSa1m4K3Pot19hnMaAeep6XVA/i5MyqmL3+dwDW8VsuJ5O7ZnQGIgMs8+Uk7SVL6n5N69ufnQ9
2pDWXn8Gf1lyyZLTqhAgY3HyzyPVW+BXvNymogI+NtPN1ZlFuVJxAajkgzj4Y2TJM5wC3hvcympv
GbC3aLpa+nxYo0QykpDtdrAIVWoD0i7DkHtDuFpKIgqZN5BiFnZMEJlKNVl+fZBCdSuKUDk/Smwq
8HVXxmWQ1rMQuww+CCW/nn1aW7CRQBJ6jrOhmaZp5RoOyQHINmIhRFg4BSYmuqyt+LWQODA4xHFQ
cexwRnyFVfauVsOb0sdUVEiEk17xS5fZThWJjAbvBrV/egGdpaVQvGdH0Jfkv5zJwSFWWlHbLT1/
cHwoIOl+Vmby5XvY7MuE3k7lz3Z0QdgkmHuKpyaS6h592Z50N3mE7SZFiQs3mLWC/Jm7CTMZJBe0
9oBYKpJWSsflwv3I59rU2MkP+XUruECdWamwdw4MWACscNEnOjmPiCv/XQ+HHNT8lAsijfrNl6a4
9eGgTpcE6/QDEqbnPIQLZV4QaRezj4eHSFhDXKeryxP4QLWEibHOP/aC5sSCtIlm5/pDiyMrJISJ
jproHgXab6nsRQoA5fQ84FoLt74Lz0cSpt6xPnwXlHgN+6WCV8lX92UuuBVDkb8zJkHBXt0mssCy
2DSo/Ns9E0gGered7Fbq13osofPIJ0QupA5QOtirTZDH+GgZx6Anbhg2mu7lD0Zl+GK1la9q5dVc
YH7CB5guhBLJQ6koO0hGZc7g9F981TgDF74Mt11/XwORSm1UhQ+UyYH88epG2kqbCCF+4Y3BT75+
e0KQBaKl4vr4HcPxwCYVLOJO6BO+1iM2x3VHEYHRr7UeiWg1flA6FvhvGmsN/CRKWsMK3zeIvQfO
Igt+1rl3WNCopcHicME2Ya4q5s5Z2/PN5muXYeyisg2RL/m/UtnZqncQrpTyvis28HM3O5kFjXiu
X+Dp7FGntpz0qtXoZIQZ26kgP0fycSgQBbj+EoXEouccZHLa7GmNd0BEizXmrI9vZOHx8LzLRKmB
/wz83QBwOmAe+a+NZlmAmML6Gb9zsLTFaDq0LgP+kEP80UvdbtHcgwyODhjTX8vWEh8qlmK59g/0
QSecu+8xei453wcZgM+xvW1+ec9T9o6oIM/+wu2RezGbevdM/39JzKFqHIZ7y72BMOrWJS1/EqsV
jVhXZpMjS16G74GJUL35lnNAhQ/e8Om6TeIUNJ4DnIUBSWL6xpuEV7KLaP0jX1Rw69cNYx67Dn8x
3mn1gGx3cc9E2uGSq9mslLkyukK+sEC/71mwEIG9XOf5l05AnqaUhFMfY/m6MaFR78cemlZjglEc
rrEZU69UdITuJ/AINe0xVh0MtVi+44lHXJZ8EsmsXhmyAk9nHzx3xcE5tJNkaQe4Q6UIZUB662vi
GCc5GbHzNxLoGSzehUPYgZX5fNTPJ3n3nqbtMej7r0hTQ2apDAW1fFOOcvGwISXEdFeKtX5F78bB
JUduUGUGgDEtSweWb6q98bvcTLqcf0my+oLWSpsC51xpz5ijcv92gI5lye+TO6T+KleRAt9xn9i5
0iP6wPrqgrf4bMN+qzqj2+ZK6RoTw2eheIv78GfjG37GGKqk+2Z+32/a+plnalj8+R75MG6mHGkd
MqbAvpl0nfXDts/PRb3wbkArilngbNjkAvX9mLtnWBcpr4wKj6OGv6TYbAsBp+ojXti/7/wsPYL5
0yKOBTKj2YaNs4mnh9knIvV+wZxNWhCy7BbbCg7ynqRTdWpXHfVhU9YHEEdeOwCAWkFD+YeCQG5Q
OrbAQkO5wkntZREGYo/TPMdk2SUot+zwvolnhjTQw+THS/1oPltQkV3kWLQMEIz5wYRvYOic2xw6
FaHs43sXuQXqvwfmtqopI1sa4Bb0OFEPZalwD3aA/nRfzgESt++oD8qYg7yRtWBEWSIGGl5Iw3Dm
GfWwgXLdgjyIMrh/ZYvw/qSP8QtN7LmCVpT9ogX6pZEQm55f4oT6xRa83pdiXe1tq0n2cqRgR00H
c+X5lJQX7L9cTrC6D22nGMNplvTpFaTYnEjJHMVPL7uPXqbFh+Suyl5MWk6HDdneGS8hLdai+vqb
I9EAw0SMmF46hbf9Ym22Hg11ec6eiMFmNt762fGWtt0I72ypzGeeluD6b4Kxx4pmlD3SEXZAVz7e
3QlMVSxzdc75Dv5htM5weLvTWpNApE9/SxvQ7Zq7uAVSC3vUILrBmZPieBpdUeqMXnNsynOKY1Wf
2FzMdpWhOWACaAVj94M9pDiEqesf4LgnTHyLHlHO6MCrJioU6KaiOnMcT8kaYgcXAQDMh2p/s0II
nxIGIbY4K3qe1pvNY0qJzu/Y0IWiXa2VnGRbprZoy4a0lMBwi3hBbl52CBlZ3/tRhMpQP4F/oUnn
NbV5GQlHC07jfo4pizwKi0lTO9Hv5aqaKSw1hqQzk820rO13kiz7MZKnhq0n0F1B0tfF0cFZjZb1
UjMDsf3iO6Ye3nOA0ej3rtN0qCmnVwblcv3bwSKxWhvw9V8fV5lG3PMyKNXtUjCChOK5sfa0/BAb
WBI69UIX2caQoNBmqAYzEgxjod3cpWdZi/ao6cQ7vhLOQk5x9xZ0L7dxVppfSrnaJvwEaKKH5NLi
goFbg3nd5rO+9A7fn6uxwHYfMU3zOjqMbbYwe2PWqn2loTnMde1NMM1vQm3iiPTtm5j+NttUD9Ot
B+y/zv6t1XpPSIAt8VqIM+3JDMH/b3Yd4ztC46Iq2rwsZCaOij0yCdt0oLaWMaSKGLvllPEh6A6s
THYgao5uJzDZz1vpj8zM8yybaq2qdLFg80bv1OIanFUe6ietihr2vdSYHbGb9ld83EWPiX5tQuYC
RiZSrKjSvQXHMFrIrJNW56XbyC4i5iwBKzE1rPrMrnZUViawDGUybvA6zPhfIKcAcJq0u52QTG7v
TLsi1xelcrG+8e5NfxXsJaVbpKjILS/avPPxTYJkMchzG+BTKN632A/vCCpkSuaMynZm7SUarAu5
5v7YNHSpXdw0ccJ/U3N8Jw/HDG/rvmb7SptpsAMATasUfVkHLEg29l1VU6CblbTfuknnJmtJ0xTa
0t+CsTsMTQgYikdlbTyfBm7OCR7jAmEgFld6FmFgRXkDeh1Dw1uR6PO3FCrnbmwMTWVoG8A62MYO
VsY7r44mDHhpp5jxKqAXQcoN6HpigozgdFgbBEJX/HPZ9HTzX8EGBaqH7UFOcb3YGht36ubbocu/
j84lsL7mD4XA1ce6JevS/mTsR/qOZCX5emNKz+i8NE7EXdQdG24nU2yqEC/FZ8PMWLVINycjWq5v
F0JajDmYdLN+o3X0S7EUpnoSqW9Y2OVDL8afdhaJk9JqsKO6kWDSnQ2RJ1lFKsaeMlbBom9wa4T8
+ij6BwDRWc9xDR2YpSyLfBQiJVKjU4+3cDWCN3DjE7kcr2da8E9sF51X4N8T8+pypIHUZMXFp647
kNC+4SIBhzF/8hXvOZHpJylwuXAK0RbUZB5Ewv6knFMbZfumKyZDsBe33oG8oW3ex8HIjgoBimKu
QLvqWrDwNjcTI7lMo0YNR8kIJXM9wgYY89upKIu4MexBS1sb+rI4Jqk3JzMg/eg6VQkl8KaY80U1
wu/AXIfSwkeYP9f/GR21yR+u9Np5tfc1PQVDRAx5I0wqPwWnA1zCiBRMra5KO5ZA9hiwClt0AKlk
6ICxwwbCSOxK04mMjVzbjSHfEl1fd7OGivTzf7XNwtXtpyUKsEOfOVnQTwJ3DV/Oil9/43920ReT
lfmMDmxEenB5Wv9IfNQ4rxAnlvSuJjgEQ4CsBPBsXlZ5R7YOHautmNRXvnqeLpkZif2zO+Qe3k4O
RUXxFfsTBUFoUmV4UZ6e8c5aT9xkXBoMIkMDymaZnhpQZXCLEeyNeJ+8FAmL2n0odNrOL0Ob3jg0
PIH7RKbrR/EOFuqXn+mGXbFSUk27AG5vd6DXBSF1bPCoVyoVbvJZO09hrIxMztYu6oNTLz/30zs4
QtHKdRiwcM/2HI8K3epMRZkNsiq0HTQXZhgXw6SetgTQJLqx4HcJGszTl4oMiBeIQIZBE0XUg3l+
Cl1TPFrbsSuaAO4SqhAV2lp6dl3T3WG82NIJpS4+xeOrAlXlgEWkn4lWUjRIdXBXZ6XQCPblViJT
XrkBfk1pwtM9N0y/TAytzzKq2ImfTZvpHiofC6Nh3WBwSSJEI91BxE6yF53hO/1yzuKEs9i/puTi
uLcLbG9/Im8VD3+heJZFq6aDH/8+3e0jbw1n8lz32y3U8NMGpaEZ0aK30+IzidBRbUi1ORJR7REu
34BpUx+iE0JKGEQtBx3F9D5W2jSXZOZE7Ww71jFkoTlF1GXDlELVIRYFAuqerYjfnygQzBLxC3Bn
PCro9rcrgkjareN4JMTBY4BJyQa0CU7Ttu/E0aSZMMz2B2JMPzJbjlPJH8Ls7W+cZonPE8AtK9+8
Nx40rQG5HhoM/gyfJyGKsrNVX8JcZ5qJYphc+SkyvI+yaiNzPX11MfxfsinFOcoIgAyS5XRk1dXh
Hil3IzIpQCLXdSeaB9b7JCWs3meD0ur9owFz90djpn92BDFFIGiRyUhaHG3/y/XbPmHsRzAEML1o
rSM8Onfl1E9s9c9lvKIxjjRJG7RHC2wCjKgpsqH4aR/qvSnp8KPJ5iK/a8dmOkWWaLrm7UEkBkGl
+sRG3kRbKGHVlpRjYpG/l07lVTexP7fVe2e5jfQ4Ng4jAaLmHyPlLLvXA+kHZXJ2JF25DMIPDIJh
+9HEnmBCZ5isHgy5ajx0h9EXZRKMhM87iIuDBQ+ykbV742+xkroivUJ8HQS9I6o8x8vUpqFKTQ3P
3h4zzbgcS5YCTSlwsSY83DA7eAZ3t+McCyrU5extde0nsM3HeUiQz4eJZkYP3KnZL0rJnxPQhjzx
bktb0RlrNYCnCKtE71CIRXIVLDLqB1L2+lcK1X7KJbprh6yf44ou2Ow6/bP+ugu2hGrffJbExFbj
21SbpB1y/Ay0cndmoeT7USs7a3WMvUFOUnOFh42YLSQS72zHLmGYMfPAAh5sp51DMhgYiT3EiQgs
Yhh2EnYohUw2ajMtn8PJGuGHjx+9AIGdKcDppsRcWUrX3yT/oN4gIGIe6zncGd/TcFTtwjn53E+N
7AK3SNGQXvoUx+Wkt31cfdW1bleL1ZzEN3vGhV+otPgHvdSxziU/u6B7gefb/Sh1y4rmmTgCCKcT
1V26UX/+rxYsp9sD1G06XuseTFiVIBz8lFkNZBjzPXMkjLyI+tHjY9iQWyYcxSUgfrGP7xroFjX5
6e4uQFS0xqWw/e4Xvad7J4iflvL+o2BJ6iH90Tq+EgU04djHYXiBzk14Sbw7E6Hv3ij/fkDyACtx
H+MbspE3f0WFHBiZLml70W1arNB7rZ9Y6gzbB6FqOhh0v4SabKxfoJq88ePLUuw5u5TaJhMw4tV7
zmQmlXnPIN+suzthBp6xvUTp7pNlXrILPwqU1ZLQv+MSVXHRl7pZhHr2GK+yhr0FEofrofpp4wLM
5c4vAmRKeHSZneVxlEOK05RaVgt41XSoJe6Add6IuUgD7gzCojdycOY0mJiyFArnYCnehl3kuiPa
plu4mbhODvyWk5+o0RpnU7oASTVeBZ7MJ+oMLP1SrMo4cI2gUg2Whc0NQkPaTTmI0RlYfdHGlw/Z
UPaQnB6tmKxgFqQo46zz2gEGP/YbA5dr4AvZwbOxkK2cAoPdPUV877kQ8lvzPtmgc713o0F3TOWD
Mgpsq5sp7xfpq6EfWwf2ZeK6xy7AAJEZSS1QeW9/R7rLO362i4sLuVQ1NpO6hcd8bzRPyVcxlX3x
2zuwh94uOXuAr824MnMC4UuOOqv2LnkguJ8Ce7fC3KQsAtko6NvF8TKeBXTDPomAq2sLYU6o3e2y
QXEmk9rxiCyUF+PORaILjv/nKOGA77fQ12FoJGHfYFeqgOQo/Q331QGtFs8g8J6LuibxBt+m5Jon
RJAruV4gagLGex1f/A4+btosVAOznGaH5yl1vXptPtugFlnUecROp2huLFFQnRyBh/zJzIMT+wWX
S+fmK15AJtMSalJL32+FQp8gpk0w41p5kY8mmzh+gt2iLt+ZBvOMDMUkm7X8HS9MSa64yOfj6WGT
bMEXHDPU0CZojLPRUnT8wAOLs0GnKE5s2w+Yrfh6upCWnBR3aNRUU8D94P4fMlUYUGZhiAPPAbUf
MmbldWN16ufowuYnmr3Pc3lrOHNj6TICWSVMeGjaKozYcvtGyCs0I+uFeGu6ORJ0KPHLfWJFZIQN
WBRv/8HeSfMo0GDj9Ok0odqhIycMso6HM44hOTWZZawwvp5ZTcIakZDcYJCEuL85Rrlq3ghoOh6i
7p4iqdxPGplq9vLG68KxqQKHEI8Qj0NZu6Lx0EUHNTqFPTwnm1xKaYY+QOhm+pggPQtXOnXjc5j+
RjDWoVu5ltVjEap9fcJlhR5RzyVch+NzsiC5K+G+Nu7P8+gHCrP2iAfKng+xhkV1qvwY3h7K/uwV
d1nlw3Bwl8bnP3GOtkO4dVit5T08j9fSWsE+RPhVsmrt0CuXVtywMztrrvE9mZ6QNJlLxkB3Zbn+
UmIq6pb0zZq/Ei4lxZuGkxa6SiVE85YGUdjuwJLQAaiKHx3QcdJEprRIWiv+kacaKCsZDUNdqyE5
/7X671NTSEEi2cGA4skzEWLJBELAQPz7m8o+Fe8kuNhiLeGmT1zRAQ+AQBUR7xFveSQrxZiQT+UB
CP1XAc4q/pcNZrFeqPOTk4/Mqbi+LwzLQrJWFdT33tUFKXZNzKZBiHfBZM4GJMZs0FJ/yvTILI2A
ilpYYJX8QnxzNfD2WDeN3FM5084rcIN9m8MYCoIs6QDYgy1L0/QO2SuiHz00rd8yP/MWiQtrXq2T
Sb41wBufc0C6UokmS7Yu8nlh/J6Wrkr3dCRGXkk4oFTv0vIFaM+7CUrSMf9dysWdAUduCn9088qU
sc4Sjjm2lquhP3+BkfIQQjb16AmypmZa1q+6hssXk8T0AfZBTnsEagLjOEs1GBhno86uwXjIkNGh
Q+5SM3HdAR7Ig+mrfWc8HqHlqaFim29rt6YcRRQX9tEuecsj5eR4iVh/W62rKPmRzPZwzBT+xP0Q
JgP+chp4XWBGBDPXedyMg/PKHZxbbDwbRd8f7bul4J0tQNdvPmdOca9fWVRjQs6BT2viNifdUxtz
4Zm0FgPEjayEU8CQ8mut9esUz1rohVKoPogG+Jm1Qav+ibny8jT7w955jWaDkN7FQMXHG2V/gy3d
ea1AjvZnirTKN0M8Q5WtS1Q3zG+txOTrYIROF06WpHrA7QOyOaeFaq3SQK2aGOvR0+sfLtJiLiNy
yCSosfBPw4w5fTCCAKkGc+TIZnIE7qOL4HTNa+89ypjw0gdKiWQgCROp+jIdFcnJ7wwPRZ+COi4b
JnXwxsrMS9Gwe0nOX+X7s/UfKrrWwqBB16/ob0y+VGjsntjyX+g9YZHJCdtRRC+Rc5fTmk+PhXTr
nNx52aI6SKrPoX5v71VBgNcLlS92KUiHbyiUqwWm4uBIn2afT2MTsAbnKUhUn3wq/L+a3dWP1TSh
zVoqgv1pLCrQLEqxdBTL8jWR/r8O3SO6fRfOUDuqncBp3wC68H7qCcxOB7nRGh3s770Wfjasxrcq
Xijv2M6TKVOMNMV3sLv7hNisNADyzVvyzkXSBcUbj8U6z1yOZnw9XwShwuHDMGNgJMNUY/4EOoKK
vrDjnse3wUI5zmz6Cw+zLTnQeJYAPO6w7fe+E2V/y+KYitfRQa3vIbv93ONhGbJyX9UdqxaFuvGa
j8hfhhNlSu8Ap322RW8uCBkURyA9ogx24IoXXWZeKulxono3JOB5JUctat/Il5Xrikd1bncDhN/w
9cZGP7Tkmh1iSE739uLA5o67RIbvmXA9dqt1rWSryjN4BVbWgm+Wu/4picibcZqPDNl+MdpC6rcG
jND55lTgcTD91jVQeVNNMCx/3CGcC06TJfxWSzFaecXZ8fI/dvmpeKamY6minyWsRpP8ToIqlcjo
PllxMIpDLnr0QMpu5k01uRMFGRhhwW81VK5lF4981paMF5Fr8NMLLCya3k+jCqjRDa6ncXamOeQR
UnJg9p/wfOt5klG9fn/H6d7ImIwnRJhO6MjXq0ZmV5EcolVINkoZkcmEDT3zieZIiwYCwaQPqa/4
rnFf1GxVxMuVW/xB1KoDl8nC2SBgLRGi3s9FmQysnyP+PMH2V/KPcvHG/p3/Ah8QhAOzwRIIPyjw
04RSaLUEGkRcrK2Z3cKrbwA1EevILt88NJprwMB0P9EGvebt+/QaGjN1qewEFFM+Lu2ZB2QoRCdW
9VvwfJh7L+cgzWK6LLqdH1hyQ0VbcIW/MM74xjZ7KuRvlE4lHln05C+UIuu3aV/RL4TDHQxoK+vg
1dWt/ziYQJOvLh0+bGgZBc7Y8fbY8vR04wIoaRqQoZmh6p0J5I2/+chE5BlBbejzp3iqNMj1GZBr
/n+Fn5BSxdWFdcJqmAV6wVT1a9aW57uqTlTCClWEECMSzs4Z/KDxwwf8JaYRye0lKUB+2R9izf6n
4ggVMgrtFmBlzqvY16FFQ1OV8IxB1eYz/4QRbKpI9n0t1TRPlMJa/IskADW4+1yRMOqmqj4e6AYb
Ufp81bCB0kltCMQQze3u/h0Y+czscauErxCcBWG1orndSkDM/lpheCWDaQ4J5F8ynHtI0gYUd4x0
qu+jOf3L6pRlz13Tho0QKbtlDEIPXFc5mZbCLPjAzuXEV54A1N+5quW7ysaPbZJ8xGtLeP58eORF
zGgVNapMX8s2F6JVSZ1AM1ev4cRUsFIedj4e9OgDXaO4agnyr11C50sgqtXeGn3EmSqAF3do3LcT
su+sjuel8UZV2fuTCs0/97t6z5dsFIILp7DEsLMy54X0MYl9KJdWIlqnJIMrm2EQnH9TogP/yKGu
GjHSf6vdYDPmhf2DgLiAKNkvTzSIiIAYknYhBI8aiwgIvuvawfDmo7Ak3MPoQgJAiu79PwSriguS
dg62GNsCeA+yPuoyNrxcO6Gb+QdnP72CtOGXVhQL/kllUyPu6hfhVdo+urQ0q9ISsIwE1ZxrraqL
teesyhvTJMmJI0CGFkndXV2+BlwsMb5MEUwnyEQF7rs4Y2zBKi9LzSY5yvpZlWqFSi1gvTWD9yXb
kn8oejDKynroLTL5GzpAsE2AAg2jXn2Fv3O1TjNsYv8VAZVnibehC+Q9Oln9r5xu6/woSLhcvXrW
JZMOF3CkLgmVHVFthZ7KF9bsQCF6QDBEDK5K9PGuRy4iw6e3jDIH9soIpPh8La9Ed7AM6EY2aSrR
xuPZtEqp9OIkOQUyvsIoZPpbl8LfWxFiO6qA0WOVC3cjLziwWAr+11vuUvQCD9IV5S7xUapBEkbf
Z8vorbEzX3L4YnPbpr5SPR0MeECwTtRcuAqibs0U+GPxlZNa3Ye3SG3YXmx/T+P97DKM/3kjeCRe
q0DCI5NHc0iVWi8knpByH4k0EBHL0e2O+DQSFpuq5UVJ79z/8Xyl3ZCrEFk8b3DKsAfWaXaozKVT
w95Vv14C0A49Fb6YsxlXhf5JP/eWog//7Z4iOiQEPGv5OmuolRV7NUSAR1Rznk/lsSxvNy9I/Zlp
obeDI9qS34/cwN0VZuw1y11ZzVefBYRRPRiv/q0rum0dhpwjbRZz+oka0J0jtmWz9j0NKpvGUO03
G6XhpsHAHAiwL0ZWPNHCzGk+HHsVhdHGKVfdqoBgjj27ZKCpD5IqyBTurvkW1fFfRelrlpJKV3Tz
p9rUHbjiro16TbTMIUuLaR1gdFtiRhWB6CIaBdwH+XdTWXQ1scNpImRheyFCxLzIbBf5wPrZoAXx
LAOXkLfLGFuQFqmYBcWDWhQL1u7MQkpgigTQ1M0BZJmEZEQeBqnxse7qFXh22xoaOmVYq/Np8LgO
vWQOgkeDAoBNIAPLNQSbxCWgxMMq6W0YdQYq2MIxemTf97NOJNe4iIQcTI9YF/L/Ma0gz6QRDLFd
sEvZ1bIgWJzSJ5mqUWT9XD1uxuZPKL+XcPI9eGaahyfdgBA9CQdA10gqhvU07FoAEOcTCvc+lCc7
gd4O6xXfxAK2WgQ6wmh6eSdjc8+uurDMK9zBMlCg+CRCI2pR/1pa2jR+ToHDnTLFgVTibEwk8CWP
OhXP6lGGtw72kBc3Qv/FO275Qy360NKle+9vyztshJaIma4NQ9L2JhtM75airb8kMLhwJHnFkifK
VkkRaM7QkLUzigVyVPde4ympBRVkUaizAP/Ios66wGHXC1Hza09ahvQbbDGXoAjCDni/hNXCeK0y
G1q65jDDf9RAYq/PqOxXOfhCbC7M2Lxiaf9U9sUVgPYljvZ13Nbnuoz/mR5nLVTdtR94cfcbv+Lk
l6OOjIVDKmqv/bvMHnLFA+xlljxh8aWEYUgWWv9mZQcUPKWWUGJiHALr5RbSMDCjT3q5s5Ufox6m
3zvQ1rFwxvdxbpJSUN03IbDaqv0yVmholsOsRJGtbqY08ddhEVP0rD+Lyt3YXLjyvjH/dlEgM1jM
2pgYS2Xl1qqRlWX5yQquq1ngBYeUoC2GRds0tI6YlX6qsjRQ4rboHbL0TF+hJPpOgvosoPpdPGTv
0ma+SX772a/uRL+hyhgxcOAJgyOW7v7DLE14k43XXfPHYjY/ba0vXcUJWdIvEzxacKYBKLmvtd0X
+CayGwHBjkF1LDArYoyCrikwzbliZ61po01ppmAItbLk8wW4yNoybcp64jgUF6LkIuGfFMP9vwlJ
3JHjESbaeSg3Feo3FnOpJytZcBJ9wXp7QFed4IjLmCqE5Cv0VqbLkU5+SMPrC2+JWNG5omuQ55SF
pJY6usr9Q7Yv4rQVsCZ5ozxKuUM+MEI06roO7SvJtisXx+ZpTANHeS6SkpqoPH1iz6c+bxHKDo5u
nNDas+pOMkrv8UDxy9DELZnD4lLsv/HQ2N2T4TfY1XqyiKA/I0oZ5p+576sb0K+sN1DO2FTc+U01
SRQD4xqdir3uRIGd/U7JJUCzdN3g2tLS1o2myEg/awBg08sccRGzzMzM8hAW4bjofihDOBo66M8u
4rP+1rKEIHdSgJMvznHPcUu+K6pandyLWsKaUcg8lwhBOv7AdUc3RJo3Bzz7cRzCCa9CwyOmhmB5
Gxi2UH+CuJAXo6jgwsrPBCTWmnKAzuyLbBYomp0Dr3SHUKT7rDVINLyrZZxJWe2k3pSbCOHVZjpW
yN9WZsr+jlAHnF2Uauowen/D27AMJHFpjn8piP8OXQl3zt+6qwU6IANFgLCuICIjhqiNxtfaML3h
VQfdPEFnVYZGLalX3j5gl5+byjx8+hcBXCZ8EH8170ue0NjwePDQ7N9vqiAFrb2YXO8OQqVtDu0G
D6Q3tzgw8Ga0ath8UUOHSuaBAggprDElFFv+H+TCZgZ5AWjjJchcwIbyOPz/c4PTEZ9ZAFM8MFi7
exhl8LliRBW3fLBjcmDI4d6vb2bsLjK95kVefkSCy6b5niUIjvvOdUxSS3l9YtcVUloWEIBlpjmB
zW89pJfTGBFtQKBv+n8ggUecGQnNplYTHnMeCOxkAOg7eLW5P6GoWlk5abkARKjJ15VaH47W7EIC
480tYfaejB6DNOaQDx/IeWcyI6bdzJoWguQzshbcS/Nknlp6UU/UR/8PCK6z1Ns4GljhS47kvmmJ
o4dCFiNFevGUL433XOdHzadrUyxyLoFTVhLWyvHotULLGOaiiYGhWSgpuWpUqxU7D7UPg2JSWe8J
LyKSmaZXlY4+pcQH8FhQffpeHu8nkywFju9VrK3QXaznx7OHdnbsDPFxlI5dwz3p1nCkQdspJWFK
PoMXlTrc/Vm39IvGLTXY3ASClEYLDuizHKEE0bh1zNePABeq/lDv1W17QD/tPOiL5nQ3ib41f1t8
eVqa6Qqx+VMMB6XrWxdsRhptXeCbhfQA9wUEQUMsLSkZLnaTA7H+54U7uWZP3lqBfj1ytaO6naSL
6d7meA89s6gvZyLuPl6FcEuPZwD4y5IYlbdQtBqo8BPVBA72qfPyX3/6CNnqwVvJ1dRhFe/DboIy
us7y8+RqR8+mR7j0N/+iQE1gsZWp3XrliENopUyZ/n3mGy7fadyDy2cBig3e/0e25PJkTCaqOp4L
r9flTNJG+hiEVNdZTSl/B4HCZez8/9oEbQH912vWfXN9jpqdlZzSmXnootPrTmlslcEeVBaPqXRj
BQalV91a8awcyVwKn6+UUbS6WwRX9ZprRcEXKxfhJgQ+PAb6cS7N+KBn7UDB/6T230ywpMgL+JBS
mK/R9G0ixXOfg+k93Q27rcJXPf/bEJAiNEVglNqNVM4FswKNq+Yi97L/HzCrptAN9m1ISWy+qk0h
E3EFPglRKKSD1alMQFqPblh3AmmbFs1Y8jaVFzA9tQNqfxnTXC5NqfllvOD7pbQtIBQXCkNMSBIv
gcp2/gRpUBMscuUmAFa0Xxcn/9QOCvDd+wXMkqCYVACU9YHUOAaT36br1pTkd4Si479FV+DK3NJr
n8NwCHdlmPxIIYNYbwKBQpj7s6Q1xWDBtvtPTZr/RXtZocyHHs7IEHsVMb3WuiKnui0TqSiwbkQZ
6MT5LjExhKnx+bImcdKFEO2HhtprEUErl/4n5Tgd5IpUHdgWo4s7POhrwvZ+8j6+coHEicqeKLby
EJncbzliydmbA/r28wmQilcWkDqhSaNKeTaWXKDlbCUMGar2U7cQMQ9IG63RuxPuS4ZnfZ+5PLm4
AVQimv6Tj5qIbOc7uCEnXXBuzNFudj0Td8OlZIrlUt1K+jdyYlN8AvYPuAma5gozMmf9zQDoJYkG
FV5qhOyQnVl62ZWAMBeaYlb1WcYnscMgfJ59THhu/UIcqmN+kevwDS/ITT5tTcrw6qA8jlFL3qNt
+FpN0TFvhs/8q2Fk6E02lJRz9rAwZPdD+hUZO21loxAFck/bltJHiKWh7hmTqI1qXjPxn0BXI5WO
LevIvttoZ9E4VN1lsJDybxTmH6Zd/7qTvk7e68mmFyHs4PnrzIPpJ2J75kjONrIAjG14hhQO9kfa
DS8YdJb6OWpkQ9aQGX5j+Bn4co41Wfo2zvpg5fU/kEPrY1iTXAquN7Eb6JgfTa5PUJOJuji8L3Z2
ja0gIfY69s4fkHmJKLssTkO4dRGgTBgOz0iZnVVj83mWPZw49Bk8P9MgcOiIFNlcLkXpqK6lvhIC
o6rcY7sWMaTKyFVqIF7wblhg2DtE6/mYR+dSxeRDsh+iEpPVQmqldst+UiM7PFRxGgeMEp+Vn0Yv
1XYIkJzAMTYXHM3g/hFHDTA4lDzTJ4GL1VqKO3CuqbnfLs4XbaZPtmpgiKAIllsMKUb3F6s+AvgR
xggPghRTt1dQW3GmZyFbT8DCH/Awr04MyEIQravrZRGlf7sL+aDHuI2+p8MmBPTqIo7UYt1/H6B0
JbTqTaELZuy6uE2IppiNBfiGCA5jWDmDU3e+rJJwC1H4GEVX2qqCiOBlaYG7DTH41YU6XXmBJ38v
X/m+Qngh7dylaq6rVsuk34GyNCI8h3MficBgFbNl1qoktd1eudBMUMDEpUg8lritrdVvySUZYCCq
XA11muNcSWJeggTGawSNnfopHy6fFeZo2pWxju6xI6Kbf5WExR6M92vp5jchPD9+sAhcub7bgYlv
bZpFhoJjxnmO4nbJW5sXX9w/45KCIZSoteuUFrGY3KE+iA0fMGQX5CS1eEYB70gZww7WFAr/Lo5e
Eanl9U4q+IwcRsh79jeExCtnOJpa1BjmXW0VhR4LQlFAaw5WgLy0a1X99C7c+H8UY7p8sKZbbXo4
gDKNrR3FGBmDrp1Khb+eX4do4GZ/UwJ8tL4bZqherqFmJSd2rC1UpqGzoT+2KUmboa/9/y1a4vY/
d426dwJ1dPrAbHtFjKUxlAclNOkod7wKk8/AJtCpw04Q1YAQQsncShbdkXFIYxH+COy3LMPz62yd
7HlXaSd5oEHDY4tRrrAsLIoRriqMjzke97yyHVbaBt4Dvjv2fNZr7l4hEMN13TMe1miQSl2bPyN7
Kyr8kKwOFNQ2P/+wSz0TqA3416j00Q8lNqphStD0voKPCU6lud2kpCopPfNQJKRS6sUe85JwDi2S
NTfo74gn6iKlo2m6fmDpRHn+LzrK7hTz2Fjky9N7YDIwvKZor1145pcjagAYhzPEJ+V0h3qfPFvA
wsQrcFBSn+6IxpmOKCeeu1t+2g72z72BkgxHN/v7ZUha9wKKA+4R6/KpPp1V+JfIWpSUibjQxZ8o
zKjPtoKxVR8Ne35IHiivJ3NKWfaUKK3qyRSqad9cEIqEqo6LLgiRJKQK9oXqnkAWv9G1CKD6WKoz
zEq1oy9A/LNq5w1z1r6YROcynvM16bTE9txm1uDdRdOqL7NwZNXYpUy5lzggV4Ac7Zk9FxEG4iqR
YjRWK6qmE4uhTxYYqLb+/pd1MDFBYa9Ua+RqKnLfkR40Lxcl4VjjEn6qB3eoUDXXjRvHhOgIvcos
LZa1yDG3XDVUY20qWvhLyvrhFWz5f4B9GdPepZq+wB1VREOMsIvq9JKQCx6f8RzfFoc=
`protect end_protected
