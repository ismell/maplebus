`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DrFNe3y2P5nP7Rx95qyoQtV577JZ6mHlWcJpkpgDuMk1tMBHYOxfAvMPjf6auNpYR8gPabRS6cnK
jRny4T5vWw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IxQn8drvE7Sb9/3BUJVMQoZBd8cj4z9U1TZMSETxI02fgVKYupGpiEh+LiYhMW3es0I1ffs6McuE
bs7kk2EOtcuTfwPsa4Wu3OOcvxHHeC98yBqddgvOLVJoAEb5RNiGoYqws9c3o1iqC3JCd5sYhWwU
LB7ySr6E8tZPaq82yHw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UC27eDrtTOjJIFtKeyx8ADcLMtfAT4mJdO9dhuxbE9av5VWQotisvd42RGIAgggOPeCblnuSjCFN
MxJcsj0Ym5C2pXnWD8k45HFBUtM1CZYllaNawVznaxCoU9cbI/F/quA9dytfQ6E3nYD7NRUiQeXI
qNLRVlKOd3sHDl4Ml8BUzkUxkau+CLIMqPeItwxQ3t7N51OKF7jRvSKtsM42GZNwvj8StkQqJPGy
f05noKhb6G5GDYG/WWfCFpt3qATC3nfEMt61wsILal4ZZQnpwZN9UWH8SrVihRpVT0MA2gdJUbVX
9rjCb9QcTD0k1vglSUdT7+KsLKo6kCJgvn2v/A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iqIbH529vk+Zbr4o+0lOrJs0Ntf6Ib2MR0xJbZnnBLs3D+25tJbl1QpWtBcK9/Y2IAVXAleMTcjs
fxnkiRTPlx6HRCqglrfz+Vz0phKv5uAumD4xiUGt4yaxyu2wRfEx1rMjicoNaeBeKJNOOrM9a9FV
tnb/+g4KQpZTMCq7fVs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hK4UEFPXCgC7q4kNPisRaOqK53obm3ze8ng6fW4VvFqUMJP5MFWxSphzH/GYPeOeKkZBMmwyzQMN
47e7HNlOFny1piZcPvqRo22Qje54G7VKf8g4sBoKB6RwAZcCt47fKr2fP6BimKj7lZ8jjoAMqczT
V55bVQ34EHRLyi4l9r3Q2wQBGK4UQoKHoiSiCQoY2ZpDaDap/GKR7pdAqwAGcIS59GXn9NtJTQyZ
aLEkmd3ecgBvcYG/Im6ZmTT7EkS3zPDAAyygUTx3LO/s2tO4zMX2OySkUFOMbQZ8wzRO0TJ8aEkg
fSuuEquk4K9hgaUcIr+/UeW6VcPEOH9JB+BOtg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
mBVw3xJ/cTlKJIeI2d/aQKXOIw2ew8K6jdLMNJadPGPriaNdkZPjrGbWctKKO5x+hl11eZzH0d7o
csL3S+obGbzyDKjtH64QK28sn8vRMlrPI6Iq+8LOhyXxE8Q3ZT3kJNrrct/JxsAdGlMtIDzjwcAx
BHe0Fp6FoJZZWEO3JVA98nn0ydJrFn2p+MxU+Wk7Ja9V7xGGNzv2Lockm5AaoL4N7zwrLnqqREVY
2j0Uv/Du4YWX8WAVY9jC7y4oQMvJVTeyaDN8dJIxDXMPm92yK2HB9Oku88kA5e9V1DYmyRldV2Yt
2I29LXI6uhG5uwxbvUdqllm2P5CxKhpyKpipJDPgYra3CRUw/sJdgqJUSR4Bln5Gnf1r2bVVUagT
UJvkhodkcJmRyfaMmHnMzD3QmjdLaLEKmNUF/eHaHFKtlFFr7v1O0kXIqFrhoX0fZ6MAD3g5VP2F
lXa7VBx6isbyhfPTjaN+bGKSe+cwgyBhgVYBK/hOnMbDSxg/SsDn4TIPqV5Hteyhf+nkT0hg2t2u
Fg/Elubtrs9WQmaQFvhs6Zu/9rAAyV9M9e7BhuBT/0v7GDQscHZOhjwr+JmRwD2MdjyoFoC2OhR2
A8Ib/W62GtVw67lkqh2Wps0F5uSPm5smxw+BnbdFANnwkEizeFEgcwOlGuCeHcmS831uHlwCqugx
KoXn3Xcx+5a3piZNdRb3vKkPwhSiKWfRKFF+NdXAPrR5wsngoT/4YnV3vK7KDYIpe01aD/YhzXPr
KxiiaN91nKMDFi13LCAkbeQyshTFzICVwR0n62kRtQ2cmW53s8X5VpMQpdV32LuocCJFxlz1NPDC
YW380BAGENDBmOMiQjynRbib38mUo7RCuIwNIuGN8Tv1InoDR7/4PK6gi6mZKEdtRm0ltR9ZLRec
pgUZW0u12BsGqEK8KP4s1Xhzk+3VGoPkGvMHUMPVSlPT2dFPkxktG+ofYZqdxbn03hx7/h14xWZs
t3aYbtKrzE5sGxxWBJXel0LZwcxFME6WAOJQu5wDuMZYp8CZVioQT+MLm9A0+f5KqgT0OY4a0R0O
K/q03WQIlj4aYUlGXPs9GSh8vt6n1x53nyKmfNxQahIBVaaeShNWt0UFMsDxjjaFpIqSFGB0SWz3
Zp7sWW66O6jUJI81joaoKzszKttpjtwp751gId+O1ewTpSiBV0MqU5+gCCI9a3QP9Rp+/frXF+Xc
BY8OSd7dqKp52qCXYo3wEY07p64hf79FQ8pEHWrjLuwBZmHCqmxF+r/y2gMC+o1wXqETzh57aAlQ
yDuHCLh1h5dR7FC7Bi10wiKH1DnrZ064sAqL5cglr5xIiqOZ5YmtSHVryTqnk2rOmH4ILieSFwd2
l6nUkKgZavqF5gGoXRMgKIGotBOZqA5fiFFewuSQdXCE0pQ7YmIXFXIcA+3I6LFSizSyxC82A12w
h6MY16bLQmJpk8QhtCIEiba/or0qkL4lqxrqC6PP86SHJoRpSAexC1vX7d5EIYDAanISCMZj+/bX
2kOxUr7oigcM3BtoT0WKTW78zaNu+R3yFJcxugKGpUG0xmBnrKVx8DCQ6vCV9FZdchoQ1VRg8vzQ
1ma0Q0vPA81LCMWjMPevBr4jvb6V1EWr75GtrVQjQXxe/UWBT54R6YYEug3MiiGyai6Dw756gmYW
wBbJceyLyksnZ4wCg7Av4UgpCKwc25PpuYYpYRDP8RZ2Cpy4TifEdGzzTY3X1v0LwOeKYlckACu2
QnvUZ+tsFJOQFIRKg8blaBZRhHrqljONq4OiE1arWFiYJmylVGsm9w0VmkV8A1Z6bPe4+e37qVnx
SKiUK8iFxjGQyUWHpR0wlJzrfVPm7IwIA95F40WInyHXIei0KFxtX1dh1E73tI1OLvz/SPnD8VWC
nkziaS1ABbvoOVlFF5lFHFBosAN411sLMBjaJvkgp4ONZVbdq6H7JoadEtDfeK8LeVtxkkep6IKY
VANVecXAxkM/6Bw4ofMa09O7XCKBAnRnA76Uis/hBOdKd0/k8ciQWff1OkIEFF6H7lVS8sQ1+VNh
dbUJlfFYFCLoCr/I7EZpfZ8B+ivk0OgyvTszkEO+vvxVUCmUCbWYhMYdsiYRuyGpjWrg/6GHPvHw
HDARpVPLJ68vGFUFFMnV7PaiGIxEb+lyF00jZkREnhwmyQM9zyeghVZYC3/DjX9UTH37cPGkWlxh
TK/I2Ub/Cyu+5l+QMWtHPOQBVwUEZQMylTlYMYA1FAmc48Z+imO5XgE8ioGb9FzDsBr7wyLgV5dy
vtp+j0q00rNOjeDAvkALEUlhXEVLFhCbmQ37BYVN4sm+PF69tmh9oSxRqyE2SBcK8nONc1XXhMfe
L7kTvEvwLIQfbfheyWsyFGeuv3hJKnXB5f//mpdI/j9HGv1/tR3GAHxPF46X69O4ayd7k3/HT4Tm
E5qKNT0oxDyvhErvlja+gmN7os99D1XrgxWCgoK4BHOPrBWKHwBAldHMgBIh592BOA/7z1keCM8D
ZoSbK4G/Ia93z11IiVC+He3zMl06tdOckPt+dCVqePgnsdy1JtY6ayzouRk42+aPdJI8ym0iaMcZ
z1V5bBfpkSHrgEgdDf/U1fyFCFwMtenlw/2xkU/q/6gHRCN/MN2uXuOO4W2Ad92RJHmg5sAYar6m
QWt27QrZWc3wDTulwOMlJgyxhAhWEl/uClpTj5vMCTW1L19Z+AsRVKM1MVG42YDP63GH9d0vt3H5
XKV1ga4tUtJo3J+vfpGGjVwx16icUwKm/EHcIs+oQQ5oN8MsgbJw0ct8QttJEFACRUqFbA8aR7zd
exBHF6Rgpl1xMQQ0CdoXSd4+3ZILJnwF7hhktor4K2rUpqGIUWqH4P8pQviW6eE+QwzjMmLr/zUF
dbW4FN1F/3xMzwosCbO9gfLoP+mwC031/ytplUgWHi+UNFAtaIJy+Ar5EZu6rRuPeRy7PlCb8kIn
mPiqa7TUZKIZvRLjJvU8sB5uQvnCYm7E39/mkGZELL/P52+B7hZU93LSYAd4qgRnip6iJVXjAira
sQJEOvJzonxFGgwg/0pURnFpL7z+MmRVWKbrDWguf4gMk3tfvARu/UJOPOL8JJji6h07tMLufLAC
FoYE0iHPaxCR2LMyfpOGgR9WtQIvTh/OVH0fbass9yHi4EswtZMuiDBRy8KNP8sotmTSOePPal2u
6RLidgNcPWA52IWLSvjhMhgSdTeiY7c2tvDpmecR2FlFf1xLLh4TmrqEehOy79ry9utenZF9ph5h
lpxijrOXzBfJ8sVOEwu4N19TrWv5APdVTjqltMb7VZRzOiw9Y77babkTdSnWZ35Rmv1MMxg6DI6f
tEPJ6KGdGmeITHdtkP6bLvPPKsxKADFiGQG1zonfjvO/utnNeMpQRFtPXqfq0OZdpZtgsfvsLth+
fSj3O99iQGpYiH5Xm8VV2R20oM34mM+Rn7JHucw2ZaLN9S3rhQlT0b6zLPEvKFZ2PbVdHTpqXxiT
PBN7IcSipjtmp9q6IDcADOo0tRIsC+LCXRCgpXA/PyLrZWKHiFbJEEDaor0ws9avkjSpRtkq8dlx
L9+K5Yj3k0r3JfeXBUpEPxyYvpeky0ceYEZMBZIf5GyMwWcB04G2MdqcLjTYPFut+HCKMs6RqMmp
Rzp9ThsZbvLrFI9FLUbOEWXA3s9dbB237ExK+OyLGraqsRII928YHNppCnW3aj7II4Cjkp2m/Lh4
ZjeL8yGZ6ZX5M9wktRYUyCNAxaWxQThzBdjFWbBOYkmP/eyeuz1XgSIOZfjZLTAk3xkoBpYiDpx/
urzKCE/ZEBYhLmsdDjoOEWeansX2tyNjebFX78aHCUNGMXrGjnnp++ndK3PTTKQHKhSdF1aKYoBx
7Dm6RyRZsGas3iyjLdjYKoDGLmIQ9eOPZLu7CJOIb0HImafawtvB+HlsRY13eBe0f0jhdk8SXBD6
UyH3c4TaBtEA4qEICx5zm7EWJ0xG4oX8bmCxpIolgB1ErpusqxF+jUsBps8fGSxcgse/1lgS0aYP
2RpXRzUa8IBMa29pgYi0tyhDCGYzXXu0EHA6rQ5orKl34E0uysN0fVBZcRg7FO/qbB0GME+upTeJ
sY6HjEblURxMzRaSmqBfypGy4kPVVbLveRW5juO8MM63zDTUWn8veNDK+2o9GYKu1/EH2Ytwg4oX
8GTrnJw6Mq5Udj4XdDpu6r8z6XK6GdHthGUzhxUdzA1ySuELgAosxtJp0OtYcgGUjkoYDc3xQJ0N
vJIkFHV4p5RaU1g/yMk8MDkx/lap2yk1Bx/Oh9sOgLzPq6h4tSoSTRnKUKj3QPHLFzC9+EDX7IAz
8J+GvmTUgtaU1nEI+bJxtwqXhnqHyE2e4PVaVgeAzSHr5nS+RoPlbcGj2V6gw6BlasY6sRuQ+sdP
45YB9vqiKLHADV6I4Bm9mZC2Mco+AonqqWfgVqij/JFJbbZjq543Ok99A8SiMPvKTQny6ha7pd3E
gSlZ2fkAq7HIm1hRmcHlLJpGswqfquN2ISOtg7Q0djUbNuF2JS5lc8uNIYU7kNSFfYZxxcWAUBBB
mRluywu5YT27HchXbOXs6UJB/VcmtOd77pyWIaT42PFYFRb2ox6KvRPV0dhKdL9YjpcGNRpGA4X0
q6aH03XCzEM+lWMEhzm8MaLrCKw/qGH8sX2BViT4FtEI+WP4B43eunWOYB1vjV/jMzRKWIx9z8Hc
xaPxxFcZJK2JT85Bs/zXLKTu4D3BjW72NEZxeYZpvFtcYXXV0v6yrw1BaPtMP1YTvykaHNaGSNxV
vgBmve/N0xgeoOTYrrbrLABMur/rPcXBr1Vrpp7g2oFtpHsPg6BL258G5fm7YzM4Hst2vyY6pAs8
ZneHub+k3FNRItHL7CcHEmjt4sGRZgKU4PRuQ5RjkyB6T1n7JGFCTzELNpQmKKO7677JZO306vjS
HXK6GEw/giZl9obHqoo/kXZ54elkOrQ4HzYnAWXJELcQh0gHk3qFyQf1A3RkY46Lj5W6NTOHszRP
loKBZ+irpbLjKMyTE7uZQLQj7aoV9Tgk6qzp8BavpvoklxBodijrZvc6/ahLxqTBMB49I7FLJfN/
+aL3ex/4ADjvcsA7lxQTpxHHBnmQkr+eEdGj6kgRBjPKSDdi6Xh939l7z+RRJZNFLj+v5mfnPaWL
nksNXNzRPmlHDJxiO4tMEkmWsHffSzqQNaIaXiqM479AN/hLsOtKNK/d7ow+wnY1g/aDfCMt+nfE
H6g+gNxQ1Y9Dy2iSOjTpnVA7vvFfUUCvDrTsLJ5cJNj6m6g4kftcPcSpXEJCTSUccH5BsESulexA
VFr6JDoFk7KZ0t9+VqsDboE54HslTX8gdNEMt5gs+//AA/8zeNONGtkV65v8aFhqUe8C238FsQO9
dMFFZE66De1nkDwtxLnAEVtwpt5loQZBGZpDJWWDeoNFFZ387/Dg3vBrVFoYMnrvff+8T942ICGe
4IV0rRy7VxZHUB07REoMQCQP9Bl3hh5wDtjIpqBEcR5JKml7bOgbRKKIaDtUvT7uyL/0L1XnwYTd
eJisQgJYl2y/Ge+2KQtvpBcLIezzRsdOZmqDB3bHFiYrg8/YBBwtodUx+3jwNN0WWftPkbEt5zGz
pUO/o+layBaLlAHX962DOXwXBh/3R0Z2OGven0PX91WMR0g1Vkm0pdwkz6vpOC/XTb9QbQeL3HNo
wbtFLjYw8HdZCS3zHnRURQpElNyXjKtnUA0y5VhNh4pH4oZ/tB0jifj8wv90t7xaA+1s3kfYOKGY
GHt1wm1ed4nm46UxcCD7IVchvGx9En5jlpPdbcJBincLs8BBA11yxcNzx61XxHHR9cDeOjLuq/OQ
XGvn84/eyb6N4CQ2GpiwLhqhAgTOYAbXVU7wvU7xEb5M+DfSAtzp/0h0RsHlwMh4JvZ3Ib3Kpt0d
osb/Og/yiIcbK+LG6nnXuBfCFK1ynQBBINUHqnD9D5iDglMx4SaqKtzWmWkRs2P5aF8INHkNhw82
FOa/OswYb7XvPrCpP5BfScyf/WY0mB7gdjkgaz//xH9lu6VAzClsy9HX0H8hmMAQwuUufrdfT9LI
gO5C6dyFad4d7SbUl4rZwxM85xvB+wXSglP0FIpXF5nnlWMn8IQA57q56GlZc5he3eQDZNMXeOII
qvL/RfS6k6hnhA778Yg3eBXn53U611D5PXF8qzgQAHOVRyFkqS9CeEaW/vDo5GLhvhOPn3LFtgIv
mosqO6f2EUxwNaRe3imVYshVmXNDASaLBAO/wZVfTLkLy8pPzN7ZYuQ9M9v4uliMnv+zP50auHbT
tx1Pt8pUz3nR5m4sIxNSDKLvJjEoS4GvdecIQeq1Y4W3+zUKa41CU11XWXddBbOo0h5W445tNrc1
KU2u3iMMX7fwO+BGELAOZGGw4FszWN0bLYYpY6SJUvPO2tqz0n06uPcjDbli0Lu9vCpwkCLr//xk
vr1fSK5qp5Rn8M9/+trWz2P6X7nc/euMAGIDktXRRh75OskbjSH9usHeex6fcHrNXV9xwXO+bCuy
V63vyfZ/PBulCQfY0i+9d8o7RWdZCvb3BDBcyUxr/goyuDyWMQ7JuBlWpk+tTmjoYMsHNMOfPn52
GD0C8ixjbhwj1AvsHe4R1X9Ba8KH9tPgNXD7IBitenLQUTUQD5HetuMrEZ3t25nWkqGDtycQTEVN
OJ11im/CHjYpBfG9EPV/IfESrWFlRuas
`protect end_protected
