`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dyILawmwGQGZDshK9S3HVDgrSwUXT05tSn5ITcYw+qwXE+4CrGOq8xbVwSvnRZENpO4OzRp6EHXi
PfB1Euv1xg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HgIT/ngeSihqgRJg1VNwSlPB50chggUJQ2QTlvivNihdQY2HpQ2MjhkvbG8+LdSbh+H6knY3GYBw
vME7JcszbgHVrKupBJHQ/nhQWtAgvqGB75DPHb7nW2rGhCrlKgI5LUzpvkHDFvp3sUMJTO8EBc/g
y9tCU3aGuNPmoW/s3ZQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eSsClp+UQlXlPRbk3/c9zIEuaJzSsXYAOp+6j4FaJKFBVavMrz0lOYeXkqm3vbWfXKvjZ+94cSJZ
9TDsUvjDMKZXHwFAzwK7nhOuXuTH+9d58FhOD5eiVNh+fK9CcgBjyukEFmzHscjyruXtnkLTXsuT
oijpJmjuN70xBn9+2BV5irkU/OuKWDWlMB2RfgaHapnxSyo7zRVxxis49ukpuLNJ1s7ji77L/dTE
mTrjcY5HXt4vDeB7oS5i+fEe2a6LfcqvEqSmt8XCWDroZ/bkupJ72Pr2eCByTkKXOQpIsYHF8tAr
tk7zknMoCXuaTXBLhBUxs2NpN9M5JjwR4Z7XRg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NKEjLZYiJaqqJwb18oJboUejfSUhI+6vzir2f5HId9W1ziOyN9LZR++H42q6BiYK2U428nLl5Lky
4TLGC9M0JZ0xEDxJ9SKHUJw2Gl/Zu5LEFsCCJZg+i8VSJAyK4PAVmrnAmI8EYKR3vznPP4B3bUlv
reDyy+qk1hRxNWOJInk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ONTtN+n3/ERcBK1z2CmF6C7QoGfPZH1LcV7U8HP1kejEhHEyxDRl/n2mwutGMCSU8evlK2qZJZi+
7T5De2aIA8zfIHudu6wFZ2AIjayHKK1aSg/b6QPhGTXJKd4Z8eEYnoMvtKYHxd9MsBJAEQREQU5h
+teTx+TPlHpYJcXT9IehrikiRdS+M5CDb4Q8TsD4pP8KQ8SDZQ2J0W0HqcXoL8lD8SmfanXdNfxu
Q+zoQAU5Lk3LEvylNsCshNmPvidYUoMpp4FZFXMTMCm0LNfPskPP1cj9a84KHC0HR/TsCCrEisVQ
XBAv1zV2H94s6E9WOcmk66JGszufyVHAWJaaHQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21824)
`protect data_block
6LFSsers+VcL6egmrABxNRjB0HEtDqTi5R2mViMNUn4FK38Yr2IpKupfUiNI2CIOY8Wce0JeGLnm
ckeskYHhbc/tGquZaAHF53F6gDhcVrof0Th680/oLFkgmsb/OdXcccxbn17mluXCBhB0a2UkBiKB
aPRkTWt28XQQCsu5B0wdgf35lji6gRJvEEHAinVjG5Z/+w/5chdJ/vpcbC8i7FcGX6dDaJX7Tlov
24Clu32jl7KIj2s0f1M79IWCLBcMng8z5+dqXMT6ckP8c4LQwk1bBHN/Q/knCOqMob9iXT2qVaii
RZg9y29/MGWcC9GznElcHO30/5Q149IBFzFn2qAfrGXhU5EhSvmzSiW0KpKYzc3oe1nKqUfq6Wbp
vZxnlpFX4B5Grqgn/jAUH0c7nslKUHVElLLRRaFa8u63oW2AtoTgC4zj7CMi0hPkMWLYBYjGrSRL
xf7yEB17n0kqel23UGR7++NG4PhKPFMicVY+Gmfi9OqrJfc8ZbebeG7/QlzzszknmrsTfNPPuI/J
WpadpWVZE7mBgObOQcGoI9178SN8rinp4FYhQFt5wf9ouLiOryLOOf46rm0/267ysnGFCOfpdBBc
ft8Y4SqJrfvDhNkfFCXV5uu8nOuiFfAkWf9D0QZcYRat3BzbH3OztUeieV8jiPJ50D31F9LumCz0
zgEFcgW+aoEVy4fNu4n7j1vFQOyy5DdyI/W3Ny8YWQoasxDO/hLd64n0GHZQVVDilydJtDX7GkPm
MjIXSkzde47MxbeozgvPUDQPR5tZXntXvxyoo9GIjLREV0e0TdzpTWcd0fVOukcrZ2ta15us+L0P
Tjd9SD+nzgRj+7Ru2+Hp7Nk1PMbDFKVFw3OS2cINa3V/fXNcnLrQEVfx6jeKi7vn2M06bNbZ/VKv
UuB20V8TM2f+bZDwotA7Ndf79eBa50uc1iaH2KvS1+P25WYchl0eftG7WzSqQz/0lmA7Y2ZX+3WF
TZEokt+tCDiQZdnN2HYVyZ9lNlui1P1QY1vgITFRlvhyL17NW0QaSOl/mwxno6KQYeOrFgiugoI2
kznySSGGlESE0/tY2rg+82mpk89AzPADK/hNysnXE3/3wIiShs45qRz+OoTx75YOsrYCXRe6ACZd
rPeRyJAEJsqnMtCdqEOMdpufCH1kBBaX++oiiAhkR0LI69UPafvKmXIRk4MhOqlxi2jaFKVyEe+s
17ohuQZmCHl090PWKox3HbX3Vp1RljWAA5XDgnfNebZeymJpvQ/6mL1Dy9Lf2PF7/lwyL2G1Ml+h
gPE099HwpA/VqrbkW8XyJ6lpt0VFuClckCpj1ZsF5p61p6exrMnD1/5bbjpyczQT5SSqiVTVI2Mh
WIIsTBh37yn+h0hMtida0LnyB9hm5L8+v85MyLMBHqZiFP1fcpuJpNoHJWDWtnhpcHXOXcuLjwUR
4IyXPlLig20v/ijL+G4stJ0WVH9UGTpXyJUSSxP3WnDU7/zCeEymzGMDUk/26+cwOlAqz6lazlbw
cozkSB/+sIzObdNvx62trCl++b1YZsS1gA6RKwKeSvUZQF1ItksaP9jmO1BvYBY6rj6ILEh3Vv01
g0n5219TVzqECs0F3r0wcuyNw0EfD597dUvqp8SSDft9Ak5po+x6G6lBq+Xxt6yfkyc/spolb/zy
xt3Vv0SMPPVrBhWz+Idy3eTuqUWHRJpp+i7VVE/8LE0Q/KDRn9VKsANSpK37e7QPsfiGXQAfydsi
m4McKLjGOkJks8SoPwhvAkpcgNE38SPau2d2YKHpnfqcE4c1znjzNqLXgK77Lv1vOO2RceaKWbMU
XZtLf1KqHmj98Sj4TB1F2jWPVgmXIHF4PrsguaCBfR49KfeqeBKVVl5yz5rp4a0iaNwyahce+42W
ZSrHpe2VMh4sKZJ1k9Wa0r1LW/mpb4tiRFeKQHu4bsHQM1eRksOs4vVe4KF7Y1uPMGmWOg3j9FHh
ez3/RwArWZnTtkZMhD3ojYuPlsuHVqZKwWiKrbq0/1wQO9OwuOb2WbXLpzG5wwvqnUykE0vCbYLb
csbr8EoYbKVZPjL/a2ckZw5sYWIgl4dbudGmoP+rSq1GiKOLp1rr4jLRiXU77wjNUVJR5OdNPsz9
LLYikWK004Qi6+Kmpbxr9f20XuN2TRUrtwwbv0hH+5C7trgmpVI4A58ZS/2b713Y6+6ctL3nX/Db
nbLHUDCpE9NLHcnhKDlGutNPLugt1V0h78gd9XXkZ1fasIwjYBR3zPjo1vA+Z9Ug5NFpQ/PZGV8k
r63ZundjefB8JAF28S0Z12lawKQbgxT+W3/cSHFJYMgjGaWMqnUrnSgvrAyAefzU1x4YrNg+PyUD
NHLlQTFwFk/ndaGj0AR4+CQXs/FNSh5G8Qx8aiWgPUEmhCbK99cdHO75G5woR/kntKtPRhglg6wI
M/t7JmG7EvIkyfbyJc1HrU2C6ZaVbNObbYMDjG7bna0uT/6/EUY7WhiP9lkYwKMSFLxlfVaWnP7p
eel5T34Ib0gD9rBHIuVThiFbJDD0RcLRxgW8ocZRtoh/fI9jdT7Ow5lFkkLKpfQ3aWP4LUKT4stO
F7W8S8dcRMGmqNNorLfEIXs/kqqXDCP1gdkrv//EKNJwt9SoHrbORWUQ65J/Tfwo34jwzl1+YF19
TBjD8nebIVGlfBnJkFtzMj2fynT8NQ55PildvXHsSOMzYPEBZXrVk67DP+mnv/LYlSoCjNZ0cAUz
Py1FroTqIoiZv31GkOKEZuy9iNhkBqoXSgK5E1NP1sQv/KaflTh2k+pKUxxeWDpgAQbCh1cS7ZWZ
yV+8XIKItpf0C2eQT0CPpd52yMg7/owkoaa4/9xToSxfjzda0qQ/w5v6zWrE/pCTdohVTjroQyjK
AEHRDz9Iq8CnnAsK0Tbev/Y5tHjsWg/q/4IPNrNIG+c8qQZ4QcDje1N/cSghFfNMjIon5IXh6dZe
L3k3RhxQWsHD1Qaq/u9jxVG4hlkDge+xJPrxK+srHB268R9YJ8q6D8pHhrB4jn3ck192qcEd4Ic8
+7OIUepiSVC+bxKng1UIlr9fVotDE8UMvcS1SQKfGsCCnc8HJENLH92G9HzGFE3eJ+N/dGyoD6KE
d82FDWQQpCZmC+v7qKXMCXE2hUxOpzVofkfLhvfnsuax5WDP+/IMkONLbx1fq2TTrLDJyzbejmGy
vY4IB0E9RYQwRtiSfETI4WSMYAbiPzQNfKALKwsSBEVUSVAuIZWGL4aSoPJeDaWbUH9CUYAm1kWj
RKSaMRLWvm9OKJoAlbt7VwHxe/Ke/1S6jtZdaaWLoukxjTMszl998K+DgbaCAqLJIpqRFhEgdkjI
c/PDEECpEE8OEQEJ8ULHGA+pEXLshtuI2jBHGtSZwDyshM/pB7kIol1Xozlz8Hrp0u8SpPs3R8FT
bptXSMrQRqvoGUra9/XcV89iaC/tEA3EeGb+1QulBPylvNFNqLVOXIDtwmcQAn864dltloJEFncd
GyQonIDUYVOq9ufuxS55GptwUHo/Qzhn8hYhrOWrk82ZbBKmDlRz9POgFv6CGDu8Ld+JIxOUSa1W
/ex/mWEXlnY+rZnCGHbZG6XW8484U+ryCAYEVGyBTBGfjcINmjL3C4aWjLPE9cQpGxgNZwHWa5zV
Gq5JRsQxrumDfYFaSpqEfSPW0EzbhddUzY9ebTjAHbcbFhFvgKlltTX5QLRHF4sGPrPXsTHySKxs
IMwal9p5aDpb8sSZChNY/F/Ce/C1GPy7YSxN5oPV63i3UvxIpYLs90+bTx0Dkx3pWTmRM+pa8f+l
kQ73QQ1IMg1AAk2ept16AUf/sP33c9h2HNLFrc+zNl9CuCccZv7nRJ9MrkzlYOvs7R6f071sbKm7
C9FgdhvgZsIn5HJWVSog6p338VLgYM2/Q97Xy1gNRn3vhXZ/ApJODsO4VhHU5jQztLlSkAQ0Q2WC
rp0zmEiXGo09qxkDW87/rQh5KcD5/voURz0ZAbZp7qOn4lnBicrGMkV75hXv0Cgc9eGUdRMzTDRk
qu8JGVuWLk7EbrxT7eH8qw/S30fVnEhm947QdlmAkQL9ZwfTvjGHEU1ia1/3tA3R7rZFJvCQ2gFg
HqQ6hz7dvkbe3i9YFroJ+AthQUjytY44DMl73TWo0YiW7b1m9pAwldxzBtCt+cv9uSUNNUu74kqI
5+JKCNaPye3g6t+KKZo1NDj3VXtudlw0cOjp9frx95IAewf6bEVsTuiN+Umr7dnWTzDjo6rvl3gg
uSiIo34CJUzBZX8gcpADKN0D0EExDbDyZ4z2ve11rwGM+hYb7t4fEH1jm74TyxGcQQ3Fn2JCZ4UV
m4KetWI4R94z/ctOw3co6Dy0h5iEaw5wcnukp3krpcfh1kqt/D76gOtxacLPZ3I6nYtI6+9SLsF0
rcq4tjLfecvLDjH6uc3vJ7nEbUZB9PGnUBb0blYgRWcEEIx2abbrYkHloRTZACvwkXaTmnvxftOu
1sbXMx7yQs2GMkvigvxBdTSppdwBcohvGKm5Nfm4FSxJGWAOuhEfvXLGCgi9bIYmvx+SuAM4V5Cm
RvnewSnnZcfpv8CTGE1IJKaGpLpje4T8I2n3vNbelEyPhNOxnomTzhxb4GgvqYI2GDlH1qkz3DNE
KzFShO8kU2vYqjHYcwybHMA+vXnI9Vx8VIi+6lGRYe4EqOO/CM+le4z9B4Z5UB5cPRUBkj4n9ZhB
K7Sc00nELdt/8ntbkE9YwLRHQ5IVCuX9ZJdPedgkhJQrqrDm7XvVuT+YqkQm62Lp6ei/5ICGC66Y
N6z56uSAJWgTd8lfx2wPY9vHXLftp5oJE94mxaNoTkoEkOB5KaJxf9yJgdMRcIWASJAIal9ELxD/
KHyd/KGwwzACQiCr348jjAKQIr3dqquJzz0mni12tCFYvS6mpNhmelWo5E0LuCHfZxk44wjHpBFf
JVMLMmAV7NLy+geUJ+PZ/INOjzOd9uE62DOQVRmnf1yqOGlxscIKlrYpfncSvHnc807R5JM4yZad
XG2y+ylIeub5PuC8zMFF/PoKiErrERQZZA7Ol/XyDezAqmFVvb3f5uE+KykSbzgHiFmICwqrNOn8
lQF0Bg+zUE4fbxBxQ/X4SDjnExs0gvxitfvz1AGBE0Ou1wXxlMTLX4JT/c+9ZfAyqM0yhzZGIjwB
d82KpbVmvPx18b0dhi2B05DFED12E8AObYeml4encFcFBlyqCnA/TuH59uqYkEEdm3bBvmCh/cTE
4bnGZ+S3D5+GyYygzx/B3uuOV1upu/BOk4s5XajOhNIBUISa7D6J8wbINLCpbZBHqICeOQCFA2QE
vgrVqrbfLexdj4LVFC4oxkUy3hHp5DXyorF0AC2k5iyRg8Ca1YIqm0fuICuB4e/SUdpcpjQe46bH
xrOTwNijVZnU3mWzstStoE7RFSAluQMr7Vy+nATpghF9VW663gJYEKyalOzY3aOIuDxk8hKtdL+C
DnH01j3C4JPGTGxo7FTPpe+lFDIJ/wvfrAJJL30S51c/Kzc30X0YXDGujr4/4ZuZoBN1T7VGT/lK
XsVlo9fdmXg4n64A23q4rSd+hm9qAQrKxrtIdtm88Nc793QcJ2Al54try11irfuxJFkyOck4FsUn
cTRl5AFO1lC2DQGvCc/O9KMkULxgFQDmXeIfYjmjvrY9a5POZVs0GMl8reKxHAW1R6Ajmpuge+fz
xqFPdqfcSlQyWeklVvyFi4w0F4lAwbIuB5pwaeSGg00bLQMns/QWXj54MUd+/PHvXRYbF0tPXG/P
1mT3B3tQtgSSRVJSey4tcSsBp2pEbN3UjRHlAfKJQs/Ib/lCNk5fBmWQn10G0mSDWFy7H59aFBZ4
HyoygbFX9D1tbScIMKtrFP41cN3iTWTrsLh0rnvT58hsq1WfCuj5jWVe0DhzJWtvX2hxlmDWrvLl
UDD8iAAYMo4InIkKpxHIOas4Gfvwj4ogIodTtf0qXJpW9ufWH10dbOFL/E9syiuRyQ2cznYCHX9S
wRmpsze6R+zS4vZx9kRGbRNtK95uIIelmekMup8xmyDvltQEmSF3stjMQnjd0HvbanVTFwdJxnfh
3wBTt7CTeVZ1y23EtydxkqQsKWme+te4Vj6pPYaM4/z7WFBDBMai6nxoSE1b+iLlt/CgqSS/LUfU
+5+y7t2Qrk8IZaH3GUaopxH1TT03JpgepHSvrUwLUlmjyoj5xGvYWt3XKzABd37oQ9ihbuXV5ve7
t5iHiKsHc+WmQNB3XNwqBwHuKciu5AxQn5u2zZMd5eWtEy9m9e4Ec/Ib1bOOq5B7ratdo4a6zX+C
3nj9/p+9Mv/y+MPyTrI1h3qj7FuZmTqgLxylRZaZOoVkfSmrTglR1bRR109MwR6R1C/t3l5RxL3E
pC3K9usB4bNrWElX+Ccvs/w67h/VPmEBi6i1SfiYQEE2dIjeEEDCaUXCtPttHmG0EYHPWVHGtoR/
kYH2mQRNUBIccNy9wpghll8xhMedIrPelnwUSV7aDaTVEnLuewkMykEHnhwUg5bo0WBSNYmEc6Ne
ccPc3fs2DLO8nfyf0wO0LZBtF6hbTJVN9fmMfJdW9tM59kVysfNNgBuUQsQi9r+P2CVteXAKhnPM
R4CKIczK+FSzeFwoB8NlAYJt6o/M7O3Wskpg9RJnzmpfd1c2vorvV3NSVXtR3uJ+LiNezm4BU6HM
RjGUb/f5eratJ6K+tZH/nynQsRu+7azQIWZ47evSJqEWO0aNUv2mMFx6QvZvZRry0+hLJA9NyFnr
vU27X4GdV8V4Kxwkx/YLMyFXjOgMUb9YZp1Shf2FyczSWnTyUxXRUkeG0aZZz4PxhAvHqdGqWfHw
xfsP31KrPME85eZMJROVPnVZ7pM6ZQrDnPJYbXprHfwppTYJkxP+GAu4E3foO+rYRUluJIDIes6o
x74k7acLaBjamgUrPqBTh5JABKRPH4wcwFmZ0dgxQf0EZA7X6iNI67qyIcWShkuJg/ACxvQ6v7Gi
4tB+hhWgvcnP7IVBGlBxSTpSwf7qe2UAJ9rUqXy6hg8fHUK/Ii2kii1Q66kSbTzb9EKydyHTE3CJ
LxCzXhPMh9O6+qbGX0ktOVy221hakXTaP2LAxfwFFaoP54aUyyEHqaPtLaKr7+sUdBpDzl1EURUa
67oPASqf3A4VzG3K29fHidRsJePzmEPJRehndMsStNEiiN7UxTOjlBvBs8UAZ8kgfiXsJDXvNXIe
Ep9I0mX/EISHSeDJ5A6yVg1Om+xOJGTKHiGmbJeFVIUDwkc40l8TyKgYcCgeCly/m1wtIZYdcAxO
qW2pE9SHrljvYrhg1BqhS1MAPu4S7oElmxhRHBCN4zk8JnUNaO8mcFOhHxr+wy9HI9bqNBO4Ckdu
ZEailD/91CtUPa5E4eAjmkMVkGEIQBfpOhafei5HKN6M6Rw7nMn8XNXZOmdUJY5BLjMhaL75kTqm
TIYUgaa3nWGzPDwg1PKqKXgSutxbJ6wnryJjYYVfMnGSucf1euzIoqO0Kp3vCPgBTDEtDJqvQtxZ
KMSn3C1T3IbyoClF7X0gcyzSUIgmdn4+fU3WVhzOhkvLqOTJZF99hc9/X0R/DblEGDcFfNh+z6Zr
53D4ggxFv4VotrG8CdXP2O+w0msdMOkD6v18rfLyy16WwicH2JGSZAHPKypr6O/OQGwK820ePmun
N7JNwf0HbmMq0uCqKTNoohgAj+rYkXtKWhWMlNadNOS5vmjfNpnfJLJoRFBBwFLyAMuIvoT8bsig
8WVSWSZIwlv0drBjAK36nNPz3R2OZoLvE7GcR9KP9icDBjE4pTk/NsSoIgoJ1w3OGPZ8CLCqquHT
yIFfTDVsKtpofGtoUl1mkQhuaMW9cXiutV8D34WxqQStxGokYZW73UBGITEytefsdLzxwX9A5O5Z
WlMZDzDCWJ3WBuRVyMAYws1+jOD0/xPj9O76XH3IWJyVSTaq9kedQyMeqeB65CIDGTWqQXUy9CbA
XnHHPnytPYPn5n9nymCh/Y6A9863WsR4sJ54lCi1NVRp23ogtmvFQobpDzwUCiaY60yfQIufUhvQ
cKlcLsniBpXf7WrLbqmvfwBTSb8pD5vUu3QHVt0bv6P+u1QwskUIIEVROs7Eklhif6xuvQpstZD4
hurPouTQfXEWhLVgma2CKdIDxJ69Z5zaucMZG4Z021ChWzxpBzUH7uZVwcU1DPSJXH2vlC1zczMF
MMCgvF01pFBZ7j+jLIJnyZlaeZM5WZsh/o+p7+xSOamHL8Gl6RDlHyVE6XtPCWf1q+ubFDZoxVFh
SszxCfAv0dTpscQvDLqk9Fg2tgwL9iZDZ/wSlnr+7CovQqYgjuX9+r6mqnQZqIdmMPXbMG6w1pHs
bDu9KFLaHm/He0uAuOaDfWJkrrh9+G7fMSKIipyxUHlmK/9xwZyXH27NEcKOcZjzGz7AsKLh2hXo
DB68KRymQgx6XQWBVwwc1eftypa8L95T10X8bjxTKjJwSnSae+AO7UpIgBXD5Ma0FFaMQ7EyBCzV
5/NPehGvLZ1HWn7m2+wn6OHcgRF8Ju16Q/AGVz8S1sHxqrWiBQG1aX6FTH8GZbZmLCYp/ktXCuBI
ivK8oQAwP8slWeu0CmRtfQHcORU5SpYoJtFB31xVNj0RztZ7cAzdWcT1wgjJ1NnjfOLEAduJlXlc
9JfFKrhwmh6GsKe8k9pGtjfupX42q/dE0waJGZ4BHmxpRnxyby0T0LYvixtahRHQoPcTmV1wGGvd
uW+gjlA76IMHYNpLa1qpxrhve6YBzXwZ/fZoAUrH+nPU1dQvR+uPGa0umywkM0BdjJS1Y2cSDcIm
TjVj/fQQ2Z9RDYYCYlLnFsTSssMj2wHuFLaJUKOeXz6PXuZispAEGQgoqn3jl/iQZsJA2DDUVMHZ
DO9G58zKWcGj6XR3mnrH4H7/tpdiXu0MkPcaZRkErQ+ExThw7fiJq/20JSzrvpt4LH53K6epEfwf
P34M3ZhngBPsi0BYZWnvfkxlEjgBkeE9lf3OJhH6ZF0Qo9mia1oYoRIEefWMgO/pt+mBevDWb0It
PLbGe0SmEawzfESF2PqBK72GGKj3N5n89+gbWqKoOA0vOW1IzXETiE4Oa3rlEGW1WjgvrfkpXStf
/QGO4uFS8eLxRJCpGP4g5zw73YhqJ0D8PSZMpNN4XJDdi7wwFteLbL44/zHTM31VrJRxCIVC+dk4
S1pY0C9ZanAoHMUpGyxxVghMMFCRrhpy8ut6cc1WfEptUWR7imL/7nlo8RgvRRZpQ7B633a+WipO
apKynDO/JO6LFiJYH7AUSi9z60hwqk8riB7PGyVcUZdtLfPXJngUaU+AtcW4Wg6ZVWzcSeQKZDOk
QBoggDdWCU3Km2BBE3KKbKJbFr8O6ccZFwHHVoohHVU2V89WImZZM6sSDQUbZhMVE0N5+mbksc5u
oDfjUVXPZRKAN+5Gh916Stdlcxm06rJxOlbJfGvUVexWUt6445jxATF3GGVtuywvgqF2HtzyYFwA
wE2P/6etvd3nh+CfZaMUlrZQ8Q5iHG1hIpS45wZVkwBdC4fXXOWg0/VOXY89eqsNuwYLgoQL9RWK
WdB74t1OglR8NAfzWs2MOcmlSmoRaAIpaKQF7c1d1vKw27R+VjvDJ5aKwfYgIeu1atq7pzcdyhii
yASMOykMwsP04FXNPnF4A+aUC5gLjM7028zXIS8fQo5R1cFUvTQrIIsmYVK3tgr5Xz6NAf3p5lJh
0QqApubaXCDKl/LKL8Oj56Fy++WM1cfoYobM4TpcpUUTmSnxdZqownW//Ecx3jcQp5KpL8WZgQWt
Q/1hCMrYfim66r3ZxjuPaGkDobJpKNiSsCm/pIPqddu9FEElDbPpA5FFG+JmBp+8sifW8K1aYMVw
bY12ugryA/Zi6D4Dbj0eeWUXHQKA1UEA7tVVTOxDPnjRTT/sVrRCqLn7tr+N30fHHE6/yYEHYLzs
yLh6a3ET1jfuEmWSyXbMpvG87ShRw/zOFjSh+pQD97rCHpwHjlwms0TZh3VhjiukLIhVWHASfuZz
6DHA1ie97W9+Wxv80CY2DpAbYKD51oalWm6xHuVY3qS5fOWBUFn3HAR2GlJ2QVtfXGm3wZNSQDZz
P/AYCLI3k4ofLYE2WVl0RfnXDYCA2+UgtGuTzIrtAK6erp22HzvjWtjCaUmyW7Zxa6nIRT2b8lUf
SlCzbT00rSBSN4AmohtJorEVowLR9glmP5WUM0dWBtFNNpcTNwUq/0C75uJsXi3kWLEeU7epYsYp
+cDLdpMf2+Pr7w71hlYRh9xtST/fySHajdNVGwZNjdhLzrssxYcNMX9XUUz40h4uduvFaKUy88C6
FM93M1KdgDm9t9d8F7T0D2v3Y9RMGdiOSS1SVWbbEOQ8hLaybmhxbjWtNhlN4QDn+j30SqwtzGpK
UNv7ZZsxLgqyG/Ypdzdkgu5UGSEwfZs9ECrIhP16DdZ+S4dm+Ih77PEHRHhxWA2IqgNjVasfE1/n
VUdkMYeb6tpp/C3Rf2mioqIMZzfcczXSP65Nh4a7iqXFiTHd6JBDRCusYGetBFjA8+ojWMOmSZA2
bPDGLUlEqPtUUycYI4juaBmXtmRtJ+UWmbELU8wIrBPuH2VurHSGScqn0NPEyAiRQMKhQXnWtPPK
YgmKTnwrL350pL04kGJ7DOJrVozifj8u4LnzUvXNBBUvIcf28b+CtIhXuFPm6MT8N7G7ZqidafzK
ZDXr2/K5dBcdGL+EUeK5+DFSQL4DsmuEx9aD4qtbawP46K+08WaQbQxQQmb6J+S3KvZjmjoenEVG
7rB6TRiSOC7yIo/w5ZQ6ozYHi/P0xQkaKWnv7LGsngGfd5m6TciRY477x+mfhfMsWY9q11XuYNtJ
VeqoU+93xS76nWH39p7RaatLTvj0HSMiO6fjfg5IWLFK50LQH/LXW30bAjmHMeNd1Wf+5YYmxc1D
VVyuAbfrlYu06rqGWhhUbWDjQPSYuuY5OX1mQLkC6yDi746514DZPJCJJA5Pp6ylMEAhji9fDTHl
+6HsmGwxyZP2OCYiiQBCWFCWfkBDavcjvxPG8cQ0DoN6bwyFJycmy4xtDMJISLjgHB6Ql9IAkRuy
8qwo9OgdmcGj776K7t1k+SJ5FXbyBToavoLP898qd3q6HSDN71F5fBUSQAI12RYNTFp3Gp86UkM0
lG2QcF8aEYipmuFEi2aZv17NzDFPUkgc4v4LMyQnJnrsZTbetB+/LSQj9WB58NNrbAKJquhNNJRJ
+vZD2fDTOJNIN8GchwLBaSpnNZsnXPMEDUaH0zVJHpb2C9jGxoIpCKKLG27VojxduR0aectIFPHi
c85ET+z4QC47b0nsPZJ5DjhXTnZbP3UJ1FSabedzpVYMznWUU5xNQARtlJy+puh8Sl1jbekYhWJg
YM0VJV18MunMYcJQoV5L43Dj3kdNV6mtd62QNyPy+tD2Sq0x9Bl9+28tWmkdE/RUYFX3UTq2PeVL
NNCKc96agDZbnGP9H/NUyWBilqT8MdEDex45wHwdbv22NsTKdv8W/sJa/6sJ6pI4J/ClUKDo+2VE
FutNZpz1c2yiv6miSfUCluJoV1ywOOFZ2ECP8mMGIBkFEbn4GAV5r8uqnZUsWR5KTBxcQ0S5Fojv
Ro+fKC5h27JTL3TEwZDs7BJIjIKPGOJgraOm/wQONVryKWOIYJQbw7vVF6rQL/L8K5El+ERMz+tM
WS0ARRRKlOG6pSEslFQBKZV3L0IHUn1RYwAyW8t6vVmYc+kwwstdJbtDiM8yDsG6yPSEMIor4tis
EBgNeUXSfD/oUru+7bXWsNrm79+6t25teO4QRGMaPiKUBIi5/0+GG3DXa0FanH+VNVl4vEotbaFV
CgdmwthNkqrll4XRvuw1xPVnNTFiLzTOpEU0oL7ZXjgFqhf3ibpi3Au2LsaZgQcJ1V5C5wntIc+9
ZUunJR4GVZGbl2NkWW6S14gkXSJrZTbFMWeUzEMN/pZFNG9KWI5L1Ni3qEA162sOJCDrefPWTmWx
GgwmIiOxBaOEKIu3Bu4R+dBwFyy4MXvmJAh84qfMKqHrAJ/oFjR1FmCZrDawLvyu6lraIsomzufp
H/qZHgUVVeS1sONTtpvykx0ZFx4N+1Ga7x+UwCLPhtRzKVdR02u1WZMN3Svj1dUvGtEfVrbmI2DB
oWQL+5D/Ij5ucgaq+tPXcgPFHZYTWCHiQC5BDxrjp0xb1F+0zxr46FrGKuEcLLP1j4heQfQCQOV5
igbQCPAKhu9XhGjXlt2sT8bpY2KGHfaTovM5L0WtNmdcf3XZw/hgiYz/lKtg9iAqHjbmvxa19WZS
00kxHEWHr1/vzP+iB4zrA2WNrHnPq3cagdc/YNZPZ8Ve8/Lui/Ske6albV4lRwfqwDHCaoEE+ykj
E8hEqDkp/yHf080TeenbTPDD4Tfj08hCl0qmX6a654pJl0zi261KxGMzMWRUs8EQJNLlel8OY49E
+OhayI1RpLBOYH2Shpq6ZPiztkhookGhG5t959U/6x8Lv1WmC6zBDPoY4Em24rU7i/OYVB6rK2fi
8wlm4d/gX4H6aW1wa5H/MoLAQt+4iNa515d4WmuMiZfNt7n8hGb/Df3YfBcWqvLjhQIGN+KXM5FP
70Q1A/TedAxpKAESnF4+RHcjZ5ghVxkIAz55NtHTM2MkkIhBbEsKVjOst4oPxb0FaVrUK5EthBzg
aVpaiP/UHA++A+kwDyA+hjnNJlEZBUrvPgnhbEgjisj//jkB276Kagd28A8rHlWkltTkFWmvt/7M
T4ZwLZc5ARjAqHV25deiXveWzHM0a5e7Y1CczIrrMrXn6QtSxesNu52pbl4wvs0oAXwreeYqeRlf
0TnUC+dWoeCRixPQqxlQhAL8zsJZ2vS2x+VmY+5RwV+3+VwSqykO2pZ/ydbjEL0FlJ57nyuc8WKW
pc8fwvY2qkb84Ct9Sf4zW7hDCfLRe1SXhsPWpStPyiNMOYvU+P9mGlZImaFYXyBrOfUCM2FWtD8t
Bc9/jIOOPeMEGtvuauAJHrdyR8JXgWWEviIayYfayZYwi2AsS1dmhadRQGX1TmH3z6wzQud7swNV
wAd/01+jfsUZzbHmBVnhePL0U+xHMae9uw9PmHb9bfkwVJGtkb94l5LbFWXrYwjrBhlmsYQZu5BE
ZXdXP/adFdtx243mQSZhhT7297nuTHWvWVQo20W1dEynvrNGyPr2KITRLPuKMoBCERRYLx47xlQA
6ZFoF8Ot/zZhtxhWYj+itgyojBEV3BHVXPf5daDdFzzyS+HUOQ8EccRQvOWSwEjDreIwQv1d69S+
RhcSZH/3x0gOwcTRxKD+BovW2iRSwXf3rTRzzFk0ygJ+J5n17GB3unwaPzaOCWbt3q3BuqGD0Wl3
QnnMepbuk+AqbvRPD+T4cGr2tRpOAqaOLGUolD1JjjiF8YLlCnXT5MXZRexzetcLojixuL6bA3i3
VyXR+7eipWfJ2vJadjTHzLi+UeHJzZ/ZgwN4E7X/+YDlYMT6FocMltePc23jt5ToOQNvrYrB9M6k
aGUfFeHh0Epwjn6rzh5Zveadf2LS1vYKPaJNS+KsF8zwiZHBTa/ufiQnBJ8Xihwbu9H/XKiCJmWc
JF9Kp3/g8BH6w0rRJmSErCB6aA0G6TNoi96mLXUPhBOBJLNjqc7gEho+nbEaYUdGknf5IlmJ83m4
xm9EnM0VwZlQqUN4Ntyi14oU2a0A/wwggcmZIlaWIYDe27Hyv0h0b5keFy6T76UsW7/hq66pAXCB
NM1aFFUX+iR0nYaAFyXqQw5e23+OiI534EzrI9qbR2EjYbjeJ6eG/5GGbsPFPrUpNiFRqmfey837
5AUqWOnLDpP4lwJHsqHLyqblwFgplo2NCGJiqv0C7k/xAOb9K0EWM+8GeyFWOfxpo5frdol+0/yO
U/I6YYXstTVrQ50UVcC1zP5sOuLuC9TnY0n2AQ39ZKAK8ZKxro7cVE9+RmosQTKOWEV0LZdS0GuA
62RDTz7MfkQWXGa3ffUeFgBf0tVDwnsdiGhIFRVtHjz34/MZhZNKUNKa6Oc5ybbM7DkrGMtzfY/v
HglqWrNyTHAeHcY7XzEmGxQLRH11v6FWqx1RCxeyNx4rqnpU+MJ2w6Ia9XZ6zo2WXzHmfmX1Rg+e
ZlX/lFUlX7KplXCzhNvub0L0c5vPoK29hjI4KqMqYuMyGd97NymCjEWKVjbY67bpKdAYIB7gcbrV
bQm1uT7piFkOBvSEmkKT8ppuL4+qFj2zfcetMIHF4YGWY0sei5snFg46s1cIUHbLuW4TInFDN6gy
QJriwym/98sZVjW3JUlUUdm67phQCKDNDdCtnmZdyW5OunpuFWi2v7WrNSdN+B3M26UQtJDsk+Ar
FudsXmrtBcS5qgAf6BY1fAKAkDb8WIrec80cVfeuCbuEcinnw9aMf6kPu2R3/ZqNQOtr2Oyg1Pw+
liDD5L7I5Pza7UYLA3Pk201WvOxhVAqzLox28OjsdbRIz12u773TDdynkch2pk+WWSd/vOE3KXlR
mPJHnyAlFlyPKWoIF+Cs331oQnJ9jmNDsCpEGSCUIZLx0KCP1qDTYM5hzv8cU6oN0brWnZW0yc5e
0irYclicVH6vEviw/xavi/n15Tu+oDYrewkqGGxXspYVXlsPfUQwaaKVWYLSmL4PBl+gxy7hSNVK
0QhZaICh4hZ8KIAm2h8qLBnx+XYvNziJVrOkRGtZBvU1QVvZIX4AjvviFIvWrOko/wFH9rda/Fts
WuHS5AVLiu/mQ1DnTXTPQB3WEZY/bBtsAFQ/Wg390QdmTnefw9dPXzn1EiwvexPAhJEwjreOD0UG
WrEa/BbCrYNwcudPtykq4SuvE/unz+WLamMgIRtL3FXO63D3E/AQCfLc250+vhOIuzRdQLPE9ayQ
+NpK/hSkdMJIeoiKk6Mne7DOaABsabonXSxdteQznK9wHcNvZbjqvkfOl0DWG2DBcIdjyQEbtszw
0ZFQLXNWOfU2CoQQG1Cphzf6skFdqM8wNJXbYS/u/+d0XVgT1LCfR6mWcDYelQ+5LQyR//xais9r
zmAVWzaNYY0gMUIItrgvWG3IS9Q5l5Q2IxvanRP2NJSB8qJ9TFR6nja6Hj3W6hbJpearoMroTpvR
b7sI6HcAl8GpmTCP9YLH+CuGVJn0561CO5zgO2IiOK0hVSAjl65WYowNZpNmFIwaxqeJcWcbX+vH
KXfpp1pMmpVP3QsjVFum9WA0PcCzPJ0jFFvwUiSX7/6mTO4YJ1b6M1qzeCIAtcShtoq34todwhTV
lChlM/MUydfsCt360LTLojqJsRWiHzCDkLx+ENZZ4VCSu7urJDCsWTeJnApMBvFjJ2o86c8kmuOi
dU95HHZSNrRHeegtivpgA4qRDBhasygGtfu28QtGl5OWZHfaD8wbBq9HJdiCKMejmAzltfaUUQ0f
1jVwqIDinK98wwpuWNkJSS/MrqMzffUBdFbskW9VIK+GJKqrQb+ZbFMbJsUWvuymiuePFJM3B+iG
9r+KOi1T05jJO3IhvlT1uP4TgNSWkwHZ2DJmdczGnl4Xb5Mxrz0Q6jbYV1hRbPNyV5K3nUDEhvH2
nkxifjuJ/s4P4aQ9iEJlvp9mE8yI7VOE6v1/yyzHOOuMFbOoRtpeHcUZRzrCM58QMDWHy4uzMBFq
54UJUvdXeHqcSqGH+5Bbnwtv+eTny/dYiOAXFvN+NG4/CW9cJhBU07M1H+BB0TyV0b3Mv2x26Syo
A2QlXXHBqAuTVy1XDvLauO2sHVG73xJTVmtmHsnWOH/yIdTWcrweq5pfcZ1+dCpWNjb7bDJRG9Oc
Ewsgx6vOKgApGDtnRek/Id0MPWsQBxpnMYRD6SOv6UTug9i3VyyYfQY3H7t3ymgIxu/W87HJBjxG
io4I2CrVQgliPbnX4BASQTjcj6zEz2QqTkv5Hmk+EAMm4vvir/Gwk55tqVApqDRWbFRbU8Xx5NqQ
Iq533IsRyY3ig4yxlbLilTDNJEVU9SSoDd77cLsocOJiYu8jxuUZj6so19qsheRKS2JbfWrYlztd
HTH+0/vz9JPuuvvk8JcqV06Vri0q1jUXdWmuHqUgPttHQt8x6wE7NDTSHigev9FELDkptOmtLrml
KMsaKl0d/v70EeGWl4j5pP6s+PWaiQTSmhFFMf0CoDIr1q2EDolxc+6nCvm619t52Se6cIBzfBmo
ht3SAg9pDEht0xGagi+GtxnMzlDlBqXx4+y2ciZ38FVtqbWOn8drQAqFujPMzb0OaBzg0VFLJDI/
AlHB5uc+iG/oPAImAJc1KHDtjhPogH31UArmsTWt6fd+665G0rPSM8pASMDC1iVQJ4t9MN670sEn
ZnAueWM7bgbd25nuub6S26Less+pBQVwVPoxj3Gsy0Uan2tzW3MPR7IRHEW5yP0Rb5RZ91Kffg8T
iH+qHNcZkEc5JS5xiLVuv4fE38Z0oND6L1E5qfrxZ1UE0GMZADYdPDZx9lmF1fVYEsUtmWO1+dy8
BBWAmFFV5AQmdNtuoWogFzh+TTlbmR0kEvkbox0HE7oo+8VNuhF74gxn1Ea3/yTVJVpAGwmF8hiK
IuEbSJGq1HnlI4JMwwQ6digebOAii2xQxSHqu2sCVQ/09yMxoUS4m9NjGyWT3d9JDJLPgEL2tRen
o9szRKsU1GS2ooqX9En92BC3dGb0Wx4yirMNYbut3aWUYSzxrsvwTZyfM5DHJvZSK9EsYjnbokKk
LFtgQlTL+W0x/kswEb11olZz8AOO69DcAWEDd6efO8SxrPsnVFsVhjnzEwA3tKW761DpfuF74sMT
jnA/FYX6lAl6+/iSft0CagDBisOQA+HRo0z9zKcW3+DLgou4586UHbGxT3k/puoF4W3N6E0FJOo/
SdQzDwbvaxtpkbqa1vY9MrE5+zLrkg3bWCq1Vnwe4EDpmzwTJb4flTh4ZYZZtFbSgzGExdC4EwTH
oCg2jGrH+vvJEcfX7JxOVFovTNS81hFwD3qnwilJ/jWeUwcffWMyutReEN1oNCJcXejUomIskbhw
LP4zUXSjEI1EQw/PSsxpE8zkpVK8nLTJvv+DFsPddG64RRRL6uycH6mYbf/0LsaKvpQENNbRM9SA
UXl12aiClxxudf10FED2t61u4SE1oYFL39aJOO8WQv0NkBH/tnNSEm+Q7wo3Lv9lv0NR/MZDhJgw
rAg7RZVGQcVd+vvHW44Jw38jtlKw9JR/z2z4y+y1+Y/lVyTBIY60DsxSwH0EPLg+HjmGIZy58s8X
JRDWoLfmyHnXeZ/XHSRrlask8LfXytGiuYbHtEE6W9s/HyQCj3R7tRuFLxH90m4P0X8cjsGCpeYX
ToMw+3//iy2b+qQ2q6uHkzUcWrVPjlhksx4RCqOP83fUR+Xm5vIQA0OhxQ3tJJsvfanqLkW1bUT1
1QI+O37h1JZQPojJWD1LIQUSx8mTE4AMNzv7fP3/YAgiWheWyVEZzxXP3vrkU/w4Qm+Re8UjBTrp
0Z7WiJhzsrULH00LxhXDRyrmI3q25UZDxTxfCQsKDxsV9aacnY/lvofk5j4KIA9GcZhoGPYZIWHx
8+6mFyc9kVhYkKVjtY/QVl21OVkcTpj9BehIXGmOvH+Qo8Q8MdV/tgxoXTZHJ7r3ugEz38dtZOkj
H0hpSN841K1MYU3vmtjoiNG3XKCeFcBW6pVOGweWlRcDMtVm4F7HQeSKzPSiUfnhJHKthRgZCko5
g5cihkGOyW/ewDpi2OI147eUXj8sy5V54jFujQG8H2C3h21MA8TssQW7EbDCG1SFt+J+rmEqUMoL
T2cCUOXEjGKj0yAPLhCn9iupFUKEuM2ofA6AayhR6RxvNs9epOETdkddpUWo8+rXwzI8bZ6Rdrf0
MjSfFdN9HDfyLYUV1l6KjX1R2eUoBIvW5u9v/THViWW6hOnDzT0BnrKfA0SFeHxnFu8R6zuiO2Vu
5UvzC6QXpJ+pvBiCGuh74Q6ohOP7YPX+2kBgh3C0+kw4e7sj0TLKueVw3jwz+g4JPsIIJWYRyoEI
oG0keq6lhHQgJ8OsGQ9riHyn7I8CPvN6mNwt7pPgPpNUYpuP4cwT4oa4eMx/B0acctEcjHHWZs75
Ajz+C0QlcwsJLqnoeXWW3W7maAgBGonGRIfdP/cjNoItQmkA+eQNclDaIIl4fx0ouyPAOhFVuDNe
SZorhvvA5r4BSWubOE4h9gOCH5LsT7AlhBw1nqfe/MhTD73sKilhJizt1ZZPmbiub3MbnaGlQHs3
1olhMtFx+lgGkLseqd3+3Pvj9TK0TSnRQSRFWqg37alUjaq4ENwKfQrghGVnyM723DZwB+2GmccE
7LgG+g9mBwHzquU8IyR0qG8XOqDq3XhHgSffygf/ymBoMbXP5mqpe2ICTuMnm6RT6O1NROD6ujV2
mHcHfqBHOWc3WfaQtIGQZdq2hwpP+AhZij1kx4aC0qd+cJuj0ooGmvF1dPNYc8x9U7N0J85TgnLm
OetgpQvWpmpir1LA+iGxszpN9zXW/0m1HJfCvoYSqQPCMxXwBoQl9FRK7lqdPEaNe4e/lPLqiVuP
Vz3E51lNvGZWFhWcD9IqjYpT2moPq3cwk90lfKoS2e9rvBSjAnMxYIvBhrcDiuJgsiolE+iQ08A+
n98tGymaVmyN87PRTZlSg/k+3Sl4FFmoponmIzAggau31aIbk6M7juZs3fOFHRv5d9OkeehpozK5
9FYJzGytg7igoDe3SNqe20mXNiPl+DpKyyXBZoRvKcJFjB2STWHMHonutpQO4SbK+btLEx53b5EW
aQl/33GdidN6TJp2SBJnNa1CSDZG47cvQgZGtPZZhYpwLjq0iznTv5mUfOGGmp7Rqt73kleMERnU
zvXFgvZCx0DynIjmnitV+4xrut27CGxyq1hKeiWEkNR1QUHe1HglTRjXpzjAsz5/q+TS+VB6JT0P
jgnNjAuR8af3ng7G14n6/1WQiwD1ncyEyecr1XKdi0JXjGGYiPynJnYyOwO2aNUu7DTxIM7t2N/a
TB2awrL4u/AZMHIWIRNDCswgDdO/qla6r2xuvHasQ7c4jTg4u7oVgkZTZGnSNd2qa7TQ2QUY9F81
+DWCQP0OTEV/HtUESmkFaazQuWaeyiVibNw0oOB6rM0fwbaOLSwUAzMyNjBTwasD3DovgJd+i86K
UDqU1rurfrrdEPC0ekeIV6qEEmKWzQ0xeNBpCWEpkObm+GkkL+ME9usfr9LpRTDPNuAAUePxqFL6
fxyjWU4BHqYbU8wgTlaPG9AV3YqmTYJNIUYlUPKkH9RR5GnqMmOeZbePsw6pFO0aAcadNFg2yMh3
hgNK8w8NSYS5n0VNDIRlBpgzayaEIB7p6ZnccivtZD5NRn8dgIFBao+0bRXENLnRn81+R35DGZGR
z6+D+qcUFE92/RFiS5ainiIFMTDEVJBIcZqBJz0VM4hrXZE7fbry0OOlaCo7H9csdBTd8vlO4wuk
I+VVaeEbBExr3fLWaFgi7BJzEHFKROVoaWZah9i8gdrbHiqwMgn4NK+ff2GNdiYDgf1yDz58OjuR
3YDHWMlvnMJ4EdTAHS6duDx/VZaRBNtt5cGJRKVH/FpnPwV6AElEwgI5E7/qaDX8XEzl5kjXq9tw
wwISYcTtG+fuGf7SIh00/p9jZ66onh2enL4TLd6BuCd9icdPEeHgeaPRRfQqiY68y5K74phIUa+P
+7CG1tzTI+ANmWHPza6MsIAmtfWiOy+ibR0uVMs4Iz8Nd9o+cMZt1nhKnFrk59dLZy1b9ics0M8J
JRe8A6tT4zRd52ybpEX/MapvJKLjPiHcqwsrMndw1Ozg5OGLpDgix8v/4QoM3LvYS5Z38Tqs3ig4
JNqR7TvRTcaCLTSYtlCo27mwYTgKn//S+6w2w3wO2XfTLswLxyNwSAShAExHJ0FpeXsibvzHFy9s
OXwni9ohqnezj1LBhfdBPKboON0seuLLxV0kW0QOz5tU6k55ghgy2d9lCyN1Yiqta3O40QP6xI1o
+xuQVYurDL4j47FuoIq30ZQ/OCh7OmK32kX6yVZ3SHn2+tzVIKykj+mMgQYiezQnvPSiHhEIV6E7
yVAQ9Gzn8ld2owbDE/wwL9vpL5UV4KZMP6JnMbt9wDgQthS9NN+GcHEShhRbHlDoCf6H4oPw8t1W
iMOFFwqPxgLlvh27aQuaksny+ZvcxBQEAUwqyfFSfVrr4OK/1qXom1Yhzz6ODnl1BtPvPYBjaT4z
9S4PJOWouSJbNy6+oj/a0b44sNvDPV68vtaam9UAFvk8mjNXLIernYGKoJjdXyZXIICwmXt4HUMk
ceoAuLT2vFrtGSiB2fZM3XNzJh7NWAZyF+Wpl28IWGHoFdCYSU3sLduq/5BqQnOx5lOoRP3sTsHv
Ndyy38NML0AE/wDYOfF2ggzir5kT5wQ8AW2Kh+6wFbZF9e3lzMUnKXbH5G8Qh+oEogDdnLQpJAkl
vyAW82ZDmzm/x8VbKos3yjsnK17rNQBrUqQAYsQ2ZCjZobkprZkAWPy0myIu0HuBkqBssWZE42il
1iKMsOa49ZSlkPuV1oUke9jVtYgKTMgHDveVThy+GmLDC1NIKslyCpuP8ivA7io+DD/mbBQsAXtv
rCOCjUb7QlcrrrHZrdae1GOj54wOmJsCDTT9KWAUMbB1fEvVGbCHt3s+0k8+yxCyrEjegmxCwuCw
iyb8jLnT312pCj2afm9iqybGYRmcIp1kREHGVkv3TmqWTAE3TmgPraQbHHtDAA3XqXsCbe7GClR5
nv5GQ0gHKQ5JIEcdIMNPCuuIneJf0xZbxTzxHfnsItQgWCvfeDPERiNhagf/wuFlK4j5aUI0/gnZ
xKx4oqoXAlast0x9g57pJ3olPZT36IiYAfCulmrKptdlJysIldbrPAFVT1zybIDw3qoNa2LKPjBe
JJcUdqYajKi4tz7MC0sOIlBFpxBTL/2EyutQ8rh1LD8bC2xpRJSoKmjfD7kzRPxomIQPT+wRFIkm
vDp8e/AEqQqvOJnZety7iKB8zfUI3oGE/Y7+d9260LzIXBBd9BmE2G3Glo3k7SKh4fI65IYPseR1
PDpqU2gePFC+SXr6pmHIss3rPJUOBpuZMNVaWFu6Oe7Hgj5Bko5WiaNUgNKw9zr0yS8ZOGY9WhvF
Z1KOKRqx06ZNrO1mQMKCBeI2ZAFUJ82vudJ+KSShVza2DLM4hfccS98sWFOpXTobcl+iVKX4NJCa
CHVPIPWSDvoTa4GefvbkEeUGpBjc5jHR4a4d5jDt/e8Yll/kXEEVF3CU+x87F6w+DD8Ng/c3vFAy
EafZzgZchSt5stk8EDnLPjZIhwRZeoXXLzPHuz30cSU0/G9f2+swVb/9FVRLoaztq4jdc5IMGAtd
qZwbrDZE2j/LdRhyaExlfn2+duwsvbU4N6maTteppBy+I5yGBVPxtB7LSD1LlDFNwqgjTttHIfWM
RtfVCPalnH++IUf33tGXZ2eFLsxYpgZbIQd3B5jdWZZuuU1gdt4Tjtvka9D5C6T6OlptyfY0oPH3
Cf25qGM2dAfJXezMUBdl6lwZVmTALn7i2XMy8vIyDQUAPywL1tPbDzzVfvEp7B23Poc2kd0BGiHy
FeuRnPyB9YNJ5rHnoK/IUZsmlUovcYOm/qtqiccMIMjm068+itUMTvBF7GKfmPv4bnW1JOnwJmPf
00Y/E9xTGIkC5lw3x7ptNFA6DOYmAFX24HHKQFU6NxsILC5zs4MoxcOk2FdpwhyXFt2gIfUx5nMD
Fwjt9bGE1v9gX6RII62nfftiGt78qWw0LSLLbIm85WDi+E6E6oyP+uh2XhfWNxwzP0+PW1HTb073
jBtAPVnRz6OTXSGsvoJ+IKGVrt7o7e1MAhjajbixk9uiJn1NULm9puK33gIiLAyhwOd7fDDRdPUP
ttnHJJz4jvr7T47y8TGzH5hMct75lygd/RBDXHAiRNhIFsP1uW8qg9cR/WaYtMmBNaSpGGJsjvJv
PLMLEPnKCHxHAKCGO0jengKbVFaM8WpAo8AaXgdQux/cvScTTWVHGXR88yGErefm0aYcMgQUptDx
2dB05JGujxiAGU4wT0KH7dFgtxEFT/7MxFn3k8ZBc1HqB2PQfy2t7a4/uo7hJgXVvjfn4FqfZ67i
OwVEtJT5B76wgDAf43COEyG2Tq6ikNWZk4HfWSHtLS2arYzbNYKRYNMIGwUDev1P1iklS7Rsh2OP
1qJLGpemYrOWqH59nwJ6Vt1WtBQLah1cwTT0MyREM/JP7MsEWanOhCqy/JCF+GU1hy5DhfCK7qqb
IbEoEkzIsYBaKxxXryQjjvVrm2GfznJQotLuwDUtqsD3DrDdck69uq3/HmIBB3M3M3ZGAdbVGN8u
5/1hh7RGR+SJT5YIYxFQxPG+YDziCIea2WmcZ6voh3tnesjPOxBwmE1gdt/8xwm5lGtHjpTXWQXy
/YNQHcM6PAt1oKMDjVrPYpyrMLpi78S/FdiVknOv4BpmUBI3jQxycPs9wiZN2eERaw2nO2pgvy26
AJUPzEM5GIb8N70Rt0ku3n9X/e95I1gtfXvnVRlxpSvLTQIjmNGXGJsebtwms2EccuaRWlwHynKT
wcDbKVHIdH2EGnUD/C2vHT3ehJzyT1e5C9rOm1cO7Uido6MKNASh02As3p7N02N02VtIHrAFDjxH
woTmigisKxWJmaIWqnwEw/9ig4LDIVyITki7dOjBiWuxNEOGxoyiUV2b/XWpNIsTzz9bKQF/lsUo
ao6AgMhSMbEzVURNGui7xOSIWPUwIQ6elCuirULcHVtjllVnt1LnmdkvHCDI71OQXIoUeDEZOXhy
OqDc7RvRlR3wTkcHdgmn/2qrgyyFoh9U+DfFgE9SuxjIcLlvumDMGpABOvXd0lpnw27s+zNXXMGz
vHP/I7NAY/ainodPtLUOuP753uH0KOY14ftZP10pTyO9z1zhR5UEk9aiW+Hm31Wwle9YyfZstTyh
LiohRpnU6DqbrDOfvUUbgI3vnXMQU0snDIYJHbXwiV7fhtbgo6ipiatTEL8l0Eg+VVhRQ5/srmWQ
J8OPbESzN10Pmgx2xx4/UYfWypIKDXZxbT3Tg10ftjNr4dcAQ8EUyxgJxHaLuCHSwD6Aibcm2vxX
AQTAEAa4jO39Ca4Pqs2mEonBkZppWnzYyEDJOhFoNqzjXbd2K+EGbiUcgvjSgoHoNlWHnRWfB6Or
rFxu57rvnqdLu8SkyoDG65BvMocEdHI/P1w9+FH7+K/W9G5ruSSV6zXxLXb0dgM7dsqzbgsCY9o8
uJkBkco06ls8hlvzJ0DNtVTtotmc3TXOxibVt5rDC3r58plDNx6dZOX4mWvPIruhv0Xj5jL+yvEy
V2335n8TjIt5WqoWT9f2wx8H8DcIkEiEvpmTskHXj4wtsEycN/px8E2t/BZ0yRJdV0zCPWEfy06t
6PR2vSORwtJHJWRFUG5/K6svkMMdlfhr+l/KE4pmjbDtksEiIokuk0fsPoSIsLbBId0PnV3rGOVw
9NQiQuxsW2pdj3xEPP3P27oIQ0v3Cvjn8y7zWzTNI2i5/gcveZRQ2BY1YAWlNBE+B2X2Gk85BppH
zk7Xutnr39pGyyWWxcEVf51CJnVUK1qblkbBsGQuzIEmzPbccsBVJleKiBFh212hx61vAkw6uK1I
BTOvZqvUpA7AZp5FubbAkzwvMpvSzFUtb6iNeBCjqojCGPngyCItKzkn/EddPTPYDQkhTlAjFX8t
/GkK8chp0kLU9zuwwAvlCbqiw7bjY+zHMguDYLtUvobbKoIIEilPg3+mR7/UNUEzvPRbwz0Fb1ig
60W7b6qm8f6uyNF5NfAdx9TlboQMB9fF+7L6gxvYer2p8N8HnLsnTI0qA58YqN2x/uhdli+tiXE6
/7HmqrmuHYvVKqCwliQju3zHN6dQrxlfc3Xz3wLxdkd3FgGNRMuDv7MJYzH9xwF22Np4bs8Vh+pt
F4k2X2Vp8WT0/l8J6Zx7nKdYZK9JwOnuoxroGbLqBY3jQNZHCDjGpYapgfld8REDTpl/FJGyy72J
usQBvm6ZP6SQTGXcyI3NItxYShx5NC/67uSWM3GdcknbcoAcbgLfzRPU6nnqcz3QBWyXuP8/Ti2p
pk/P8D8zB6ZF9Ge8FCxTF3NmjXhGCYKMovtPYnKGa2wUZqYv/c3zDtpZcPnoqyUtd//0rNpiEetR
G4gpFaWsWULPZeKQyC+5NPavTn8fIaLBI4T+7elM5obJCcDks1cfbHoFdupH28WPo8JrBH+IgeOc
B2UcYVhGGgHgguMr+iU+NxEJXMtRCfpf8zpFuj+CQ1+wOW+F2YjArkpa8MfDI9X8wZ6r7z9P3S/D
SCj3qZpCEfCZ1fWubA7Rpm1wRkM/pQrCe2b5yMN8mw+2YYMpKNgV6HQkAcJ7jrCiGnFy2PwMiCmB
kVMno1nqfrnIDajYooNYhBbbJ2jnufMjeQia4hfWPxVjioxltQd7gxhCO2nh2TcmRXOap4WrFYZK
stNTQm095vJeoVBJTE+GpqIvUVP6hJlfwmiOASMZon+SsmVjun4VBERmIzrHrxwqRsjHOYS64cW/
LhZAdg5rx3s98qjN+5tAdVY7kj8AkwWMWxzWDY2yyHNo4WoEUOLmSXtYZdpWgmIOVWoiYVd81JQ0
CYYE7vt6+P6g0egeosYiYDhSPgwyi1siTIfd4CyVO6hNTstDIlRCKkfdhSj9fAEWFAYfayZPUURT
4A6UWLayXu9ixtRL54nn0b/stYIqg1zQtCrhazRCcxxs0yWLG/oRRItQN1IEKidyVcaOfiiFEllc
WC/qkn+3laCRcz0BsfrIIsip8EyV33TjLOriah/6z3llgyrwS5Nxs9EYUY9t0wvcc/hw4JEZNxtp
3eB4LfXfipHKz2mrBXmR1fayElE7SAClkcZ/wp/n76bCf3pdBRr5WwwNUSbjrrd9DKQYYKDXj3i2
Tlbyi8sd6TJdlB9hK/vKQkUqbd2zf3MEdPoV8LcBGDGVqiMyuwPyUVWDsDjaY/IQ8FEyBUTs2eRn
JhG8K7oGSXk1oR6RfZyQY7OELezOCnivQpTukkuMDhhd4fl2gW1Y0KWxxR+H5CdvJ38bZMCdHnJy
3qlqVz13rACUhvuo7lb1H100YgieXvDM1EWiCBmy15E2idCg+NIsn54bLozVVm+4VeGh3Efr/Zl1
mKDwdketSdxjtQskR3yN6eYW9rJFND6qdzelC3vDqkOZo/2xT4FSmGKrVu++e5kaCUR8Vo1G4xGL
+YjH9MPeohsdYbU83GE0wuKYyQukqHXNQiGnM4e8oOpmDk5dw8+FeoHyVpi1gaHJoSa3OjLC9OqB
Zc47MS2/PtDqXqAFMzzQn7Y4phl/SaDAZiZORKOYJu8G0D9nR+qRWB8ZCCn22i6LBKx/wx9UQIzx
u2Vugxbl6+ooPsH+fesMI8dPpP4tQhJrx5ZQusdQH/rp0A+11ZIrxRcwnukmEgbKFZviev8Vn90E
OrG8Tll6Tu0Rg3KET3tpRNSIn4aoeN9BJo5jygYgBbwRaY77wqS0k0neOb0Ct8ZT941u0+mxzIFB
keVBBVY0I5kopJnVTF44mtt9aFqC1hPb/O9dS9PAH3DVWur0gy2sr9wRb561LoU1n36PwQXuOHrm
UWF+jYZkFSGKBc8M7gJgyVyxUdta0yWSCcZrtAA8FZ6SgheA3nXbeUbcjr0ca3U5+mcGw2sOdDiE
PBcU/2WCnhF3V0NFyetXUCNje8n4XNBuAW2BIXzxbh9RUUQbtQXycdbKFg8iHvsO9vFNk6c1DR0K
u/ezmqQDdt51vp1+F+4w9ImoZ5dwzg6HHDOJHFoijNbp9/A1zr3loeObffi8DBCvTqq4ojg3F1q7
sg7DC3eNtagnp2/OfGFc66EGsF5FR56oCglKe9bWZubU0BNj4cJPGweT/7asH9tDFyxzux5Zf0g2
afW0R36NKQCrn/6WNQG7FcDOrZwbrXlUqxqH2rtgILojeCyxObFBd0ooXTfZRdNl067NerjQhPet
AQaD1X5zHhOY/p3EFhx5wOwX6HiX/osyyW5+DypErVR15On5u3KZTlyjaYb0n2yz+gq+VfbEifRF
8Q3VtlFRHtm8bVrNjNLAn2lr1SPgS81E4iUr+DydlZtPHQdKruDaOOql8vHEpPsK5CN+zVNZv0Gs
WyJQi4H9jPj58aNyPzf4Myk2nSiRZujK9ZDMMCPm74TaQZ3/mDBSB21RPmZ7sVMO8Jj/Usw2LzXH
6/2vt3T2FkPg77+DRgWV9zv/jq9DOPDfvOI8tpeH94LwnU0VXyFYZyJ+3WOlkFgwbdJpO9ZcrBgu
U7S2pi7jIAWWWtpB69n5ozUi5cxxPVrsbwypZFD410zBw5HGrzLIhvGFNI7ER59JWwG5PTKs9MzI
siGnRJjfSrNu4UtEILueGwbSsvQxDRvayiZyDXrGTknsg8wvRad30ae520o/0Pgg+Sjx/SYe7up0
W7zGUQlqLQVzwG60cP7I4lTkhSjT3lo5FAm3R9MljiEZKEtj/jPVqIwfp0lk5vHB2lNlyn7KIXQL
fI6eEh/Z74llYjP96oAOHDtygeyLuF7XVQkfOwyG2UZh5FU/NvMmHrz4MmXgxQmrfwHjiA2spWKb
DcWT3j/MtnePCD5sr8+QKnTN5hW9xvP5illuipbQrP+mxnctK9t9p+ahLFCYrs0M0+qvM/dIBm1L
zhI7Gu/MAR4ZdRI/uRM5lFHb0biYfPgY+qVBxUA06DWZTzY99KelKGuKugFo2RgCuYjnGUujRKN/
WKyRStAbBKTM7ABQfntEJYrGl38UD1tDr7770HFvf8saW9/RfosBw2tqWIFsamTLgc2LjyfljXgh
3DRrBAmeJWqG1bvwz8ozz2TQPpk03Sxn/6oRgOYfkbdvJ5yZNlQMiSGmbln5/DYdhlNTGDXuTsf3
6Y9VHE10h2hzMttFXxI+ezr3t9Cfwui+rKhB4HWCzA+f5smFailOPE+gJZAUFFusQE3PShdyta+Z
GZoP53Vt2I1sFdrK8UoqqzUq5iNs4GdVoUkmQ2f3YszcuJy3dRBWEjxOkvRSOO/029Luh7ThX4b9
4qsnCTygK3tKjOYm2PPVAATysH0QE+f7KKkiWSiChLB8Dvp6QDdJ6Mc5ZnHddv0QlIKM5MWNvJjy
hOurqz0SuGxfA8kwCQGWOPdcFL0NXKkncDTXeND8zyi2TkDxQwESydtoS6ZKt6ObX6byLvDH+sbl
bj4xjGEopPJeaBfVbVu1zVyzThHCHWmE9pOe38mOKVJ7RC3VeKV2Uh+T1/iJB5VJ36x8ICWzqvdy
QPPODfel9MgalIXOaomuPMKZrOz6PF6N01+RaWsV4e/aU0DOdVftjHJsEhw2XgnLx938glz3jKDH
YgFBivUgZRuUZm1qP/mFukJSjWFpLSxrVuMnFbOd6oZ7krkl5tXTJ+a7fX7IWlZSFipjtSaYbXE8
AEpdixPqYU8RfJV4oy5omNI92w7e+pz6Fd5Y/xooG/WaWtVU3uZOjMPYNVlE+UbEmHMCADcyKFCU
SB2eRN1MlDMEVZ1rXPpJc3JlCZSYy5ibUXsWrmUgyysmgVfOt1NL1uru1iJduD3cPUJMQzCHTBM7
zPfunmv04ToECeZCNrkf9tScwKDCcOZh9Puds3uR8WwDWKhB65LN1219wjHhBLP7qd+3oNDeUluK
1/ACfJZNcyI7S/tyWHXfCodLX9TMOIgIlmfAenTWOy7SxsGNS6mfQ+5rK7sU8+yNS9ElmKOIjCrM
zywdbnsKGByN2e86Jlx5pZZgQJT8DKKF0+hr4Dk067GZDGIpZNe8iPlFKzYMPSlNxuDKXc+U3Hs4
tKgrnU7RNUYjhzlMNb96TL9glpmxIvHYqEivaY7qNY0/i3tsPSBprXzdr5O1dRx/pUxHkki5Gqi+
OJuW5xE4vfkgPJ5xUlJiKDDElsYUU60FnyZA5Y4cBgCLj+3GNopfE6qPDTh0S2IPRfMNIPy5UlpE
ZoyMmFGxsKSMGOcB60vJs8sYN+h8qzhFweBOuYN04mEH/7PREztqNrCgu0oPHZnIqkrE8UxC1zDy
ETT9hs+czXEhuu+pKqMuLET+D/Q28AFNfnJCElUTpeZRkF5LiaYFQzIKgaBybGWzWnQpMN9SGFb2
rMKQTg7MPsOaTY9K+ztmn2OHuerjziVkbLO6rTMLffHs3NF032B8ui9aE38Ci//73AFWUOCndQE/
lLeAO7/LyKiXcpdC7C1IvqUy25nHVy3VDazVK/t9UM2QdAIn3n4A8eYV8KKgGTIfp+T2PfRVPJi9
VInceHFsoSipVdVUrpV4Eda6D2B2/QXYDIiRnYgpzz3ARjz81R+7xBYMo/pfC02oddqpqTAX3ZHL
e9k7VD8+3HxTYY/4APuA5siTDBtUJsxWV4UtMwudzGfOkEPKtnCLjqpE/7O0U22qCdxsdvGUKh4r
soRuqQLPpXO2OvXcj6cj0zpgSrB4QR4HtVG3Hln3f/mO2rDVPd+jQBDwsfWnbE6qR1qcSfhGcbAH
ElIqLOxeyOXqToVc2+tYS8m00HlkcIlGgRL+6oxIGKafYtYEa0+5VIhzWsGX3eui81hMflfPL6mA
Bc/iQgLcCUaaJATEjusT7dS7N15QNPt7vJJcEzo3ipJ+jcc8knmTXn9xoY4h9+q5+J0J5j6bTxvK
vfKelm1GqSklRfMLI5WPJJzdN3VtVlq1uxWTpLSk8BBHSSwaO5tCHcmpRKPkKZ7uXUN1JDv+qlGW
KEXHC43qXNTTfqpYt0CgSe4xVJKbqcgeodwsECqR0VL3a0nvAP09BKL5c6Ms3ecd84z4p9UsZovp
fAnFUz4/3k1c532K+8WAv2u2m+y1Pk3kowWMbYM8GuZVIB3G2dmjNKOHZaD0YBLDsigMpeCLTzBT
RVax8heofH8C9UreS8UESwGXD/tiPUkhbSRBryEwWd5+PKOdIPrLqxPrcvi7WsigF+KG96h9oBOk
MeBj9AoVlcTtoScEly8gBaHTDJKywRjHBmVuk4LjJgfYJ8dx5i0dL8JvBpcfRKs3o5jO/Kpx8shp
ooERzJdXt/uPHsr/b+GknOoHeU84ukXlaEYNpysMDVzsoLQHwQZ4viT5naQTgONy3K0=
`protect end_protected
