`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L8H38Pn5e+65ZnMCPrgePq372lx5QboRhoemdcS8kzXm3WxhEUO4tSa2P/S4rld5sGInB1EDi4BC
mUYJhaWatA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YCgZI3vLQn3JXWTnPUPW749ljnkBIShBSx7VlBLDLuJKIQcDFoTqIIK9sRuKRCNw8yOawhQEgaD7
Cr3Bm7UDRo7f+Hc+zkxV626L4tuu7+0Xs86Vg2gCbuIWRqH9nAGGgTiSFvU895Qx9MT7u/sVJ5CN
3KOe+zT1EfwRIC7tGxM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HPHzt+lwYO8YO6ONuv8Lm/QQwSgKPk6gIRjSaOLRR30MiWLnY63NjzuQk8b5EzuxCH53czJDh7/6
t+eZjQ/fHnD3Z7CvNdQnXdRsve2+qT7PxrAfpFghWHkk4VKh2OdBy+sti6m8EK82BFJqOVqbmlFO
pFJ6GlM5mRRsjsCYyqjgLfulfGNMMLBVd/UhBJhRj1mgiHTM+IjYJ6mZ0x8iBWaF4auUS0vW8dkD
8gVOMzK4t8MD2NUFp/YtRdr6uJqlX69e6uKdCFWHo8H6AZ4M1V90B1BDr7D9dxxJKuCiPvV/mmVL
IHnUshgpq02c2L7zSjuXJseWAdSAzxObqgeapw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1seO8D1TglRAZwDExL1q9tv44rCD8oyQiE2di29aSVb/lPmpyltiwxraF0YFxFYpJoxUb/8eM6BI
DAzjTRT/7qqXzC2+tPQQnDQsI/INhfZb0mKldM+JnW0yyVcexTk0hB/0lhGHjZUvpim4YXIShAGc
Miur5wRO4grMIg6LXU0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ltrmPHNy0YITlTbIso3YWorJhJLaMzmLqQZB0I8DyBZLr9si2To/bRkTyexOEJjV7l2AQoZaR5YK
PU5ebh/JgAlxw1Fai+rGxLhu49Ejvt+96SvUHJksQXU72CvlZly3afoTJAxrDvDTDA/sgO3zOIJc
qSkMuVNgxnueJZMhCCgEuUYWhTVM7VeXV7q6nhh1K+gpBYuElpfrKwjLVPZiskxaIStImZGI97ch
KNlIX+M0TEOW15zVA5J4Nboad4XU+SufaHZ2AyhrVA9JYlyZhCS2H+9PNouGFxy0BGlzAR3h63oP
4B403UvgysCyTKigiABXaWIB9C2wODNpfJ5D1A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8000)
`protect data_block
oqBwFI643hiaANpquatYQIE5hYd8VrLdva4XEAGTFddOKwOdgKICSn90S3UMUK1SfsgEd5Q21s6W
2W5Ls666D6+Hs3lGU7iZqCc59ZmzPKGNAf1MEribo/iNmwRBRAziPz1x2eoxxWpVfvheSQdagvL0
w15N8RYkfYfdYhl9/FN3tWo18Kaj2F3+bMPWEhL14wgJi3dFKgXDLLYsYGBjfjkggDrzQfJXoAib
wDUz37bL1Hh24FBfrHjzRZyaTC10o5EXx3Ulv7pTMckamxmC4+VFK4KDg5TRNieQjy/gUcVUThlc
6WFE8MDXrpOOH+B8i3GGDW1kZc7bMYTu4W1vdst49lUz3MaAzZwNT7hfKIHfUL5mXzSBrdhdWaQu
IWZ3qMVOsKY+Ba0KYWotzmmXLnIP+PxDQxN8DXwkq3tyLkXWbzWQDQuwXM7lG6aqLRoSXROngVqA
vEH21JjZatJ7j4PF+d+CvA4RWqOwj5QG0WTryyi7eXL2VLvVJeEEO2qAnf9vrv9wpxGDbFjLkJYo
xrKbGP/yLmws8hB5/YqOUJCUw10azLcet511oQmHI5MrEf8BqQZdlDh7oemKu8yNtDKwE7wmqHba
Y17QsTCRnXI42aCGcZF90xPb2rMzZd0Lw0ru3RhAThsVY6lh5ECTBlz/hwIUhKe7VSUsZ0v21ihu
XmoduNlGbWwWxRTydHO3krL8m66q0yFTx5AQ+O86GDDRdWDErvsIjFztxnIOb8EC1ShtUB9mpXas
uZIqMUYH7MH+MoUcOTStKFgAye5Wa5xd4/dhxlGEuvXmDvybOOdxqGYpGEqHYAraFtBI+O3J9BpZ
J70a34oMWNXa7FynNGCklCwYSWAby9KqIcP5isz6eD09N4HA5hY09CMvhP5FsRWPDoD2VFRwlpxw
EZ3dXGBh80IlicHJCJtbi4kehI0V4JlCgqLBSNqP7LFB9u6krgfdQDp/vpgKk7UcQdT2y1+NW2sz
1ly1EHXydGTsBlrTQSszbvfCNo7EZe5xyyAO5o8jNbOWkxuj8sHfr4cjM5cvM9cpSjnLGVBvqxTC
xVDg7DOp5Tlc2WoYFKmDwBcWAZUCrlMx7xTXNFFgtF7CN5syKZq3nU+gysc0U5kUVPEWHQcyL6H/
BTdt4Bou2tfkBX4QIQlCg84jhCx4QCNawJ2mVP0GWKkl4JZwv5lDTIhW9EcB684k7bNPkx0gViiO
6fDUg4cYcOuK4zHO8CpJnWS2hpLqJkM6YYGl5pYVymeUK1Uu04+1MKpmSVKMUBISYuXKIFSFErA/
kTNnvHEK8pvvIW/8lF+g9qA8RjAPVouI14e4pH4ZOoo356zqON+VCrKZwC9zH1l+kF2+Y/O8IzNP
OjnwOv8TjEjYfB1wE7+CHzAjrl9xy5y+Wj/dBTLt8ciu6vn+LKz6UQOcHCDnZSZd4/AzPPoqLKq1
iaGQD5xj77q/wCx3htkdVNxj3r5740GLgSbVOoyquDS45AfwyfY3c/r+R78OH/EO5P8k0fJN+sAm
YqmATIJ+O6QQD515EcYi8+1tLjj28ZTxXoYc6CMIbo/7OgHxUkh5h9WoAyn6Y3FjKUU1QYsoG9Gk
4BKFpleUyu0QpDxtWeFxFp5DxIRA35VARQKViFgIWgrGRqi1NcW32+0QDzpfPdHpQ3lzpSJey3ke
xOuAf7tTe9fVlZlcjLHWzVz2Q6JY5CMRijT5dKSLLbuVqWjrM/6LHDv9eSauqd30Z7ZVwKC2hl9a
jnAr34br8MBzs92RyrjEjvh/0IyVtXJUAPXm/zsdYF8u8AXaDWii6VIZLhDEsbOXbDIIxL3hXoLT
mALF9O2QbojJyhiuquG1z/bpaFQSHbU8cUJWUqAzpvAYDIqOAhJbXtq0Y6oUZzFKVBCUG0a9bQOK
+YHELONoWPUiNCZJxE3Up/8Hs5cgIuWeRP5sckjdMWM6ZFaGZOR5/5VKFG6JKifVgL0qgNBAmUDA
DKWM5bTOfjIPAvj30ejgKHhR4luNzNXvviqWefmj8yzI40NvW0iZocO8NT4gClbeHs4oXNNc4LfE
fALvcFKvdOsmnzLVQVySvh571RxSWvXxvbPLyEoUQgFA9gjG8ZKy4+YXHBDPb/Lw0EqUi30SiKce
TzkoxV/x5T9el27dWLGGRGANQt8hiSigSb4KuKG8Z01S8rLBexgLYoDBQ66UGv1JIKO+1KBxxzET
cpjzhUxoG5CpN/atv1Yer6BOKoupU/vRucVB8sOl3YqOgo47ZFCDKMTNQqu5jB8y2rCWdmajAaVN
pm/nZktPAqUALDJtNySliY2hc9Zyz3gsNMDfOHtN8PSRu0pO5JLkOHoByUO4F8Kh865IygrgExqw
72lhZOv+hFhTn04x1D+uawwKHW4Rnxgz+2zh5LJjNqfVjNPtiJz8PnZtj+DgBC0NH4aq3jIvZvC3
FiT1c4+q7aRCJsWsxePVHK/MnzF9v5iLraDPXhUUFEZL8dQJuW5TJNAz/hpSbeE5cmrJiWDGuflF
5oWrA88bg/daBzIpdanud7vYQROwsuyYRT4+2w2l3xCuVj7KgIPkl6Z3WMksbIt0Rl4k5JieD7zC
cOaQ4lGRQs1vNTstTuLL/33j0UDaYD9/d3zCkWvrdUAYWC8MshO2Hi2fjY3nGg1WnIm3eMzzv4bm
r9wMgPZbVOq6bFdNg2UHz74W38NkEo9NfSlhHA2034zupRrr9weWOnrUYyi8nezGwIAadElLnu9s
Nh5GwXP311vAIsFh/Wb/DK/dTPHsYxS7hg7B6Ic4e3OHB00izD9OAfJN4w2riIZIgwuPa9F8Dnpe
U9gBMvMv6z6Z65RJQG+CkBaMEgV2aJdXKRIAK762ZWxM8AQL2Xb2XzP/D38/qjobi3xZAN+Z9LNy
Vxu66UeEGhBU5myTI6L+DxwXQ7THYZ9EYz8Y7egdYWJ81362Jv6ZL7ttBUkG0aCuSzGrj5mPDvhG
WIS10aNWXazSmewa9upolvPjftaOVSPKaaD56JGkPuzVIhe5dVtUVk39z62Ac468Pt1aozPNKccH
vDE5zvJWCZyNCJiwpRc737AHj9CKnBK8xTSTDuZ8w+MvypG8cum180VKpl5IN9OqoDZjbM0HY8R9
AJZW9jyvYyfHA2UkrdAk1wyX0zz1igsF1pPgd9iVa05pLkR0Ecf2xyrLhUZBZsqYXki1xab/Lg87
Qc6iSamKmm437yjh40PTv5jkVGzqpf0fPl+GRfQvgnmAqCvpH7ke8EIeMuR/NOHp6IBLwEE2Ij3b
PfOcUqHZwLWfcdqVWtbRF1j6UrEAYttk22RRnZn6NfTb653HTWrbLPWt1DJgqu3HAxXdHRlnd9ui
v+cc9tvqkTyK3WvwWh7DUwXRp7d2AWe4mOFW00ISv8gxUssEOk5R+SjqgBkDjJf3GXejOJhOu9iY
OEB9TUVGl6OcBvgaVMpzjoQOErfvzuZ3UYtkHZBUUkJ4VAREkvgcdRwfkjIokr8HcLAUzlwy/FWH
JMtaY8YgPdkqhhhMTGh2nw8z09fID0eu7f5k8x2WX34SyRvG1HvK7rExvBT/w5UyydC2n8hSbkTF
p8+Z0ap7F4XSPn5bRJ4nl2zTW4/PvzC/WjukVUDcphdo411M/XlQBpUAEgI6toYPmk4l5zA5ypaU
bW7pXKIJz8jfWnzDkvaAYYH7/HcX1kidIwDAC16GyB6HXUQr5m8/nzB2P28qBlVonUW+zNRCAGEp
9LMzRcD53wakAZK1jWHP8FF1/44PKiyJ5AO6qK2tAhrbeFYXg9LA2W1f44TFsvWX9opZYU43HLev
OuU5k8fL/MFO0bRJjEbpCScQ74IG9gZe0QCa5jBp3nBPbjnBGHJ9dJfZ4ZnGZZVT3zUGWn7ddcip
+CsbygCzUSdnWe5oknjcW/ukI81PlC2rMcDkfCfwiusSi2a8mi6wPwkvZ5MpG6RUsSG828voSTSL
4TfmbSZH28l6mkm4liZwPgEm1F8C+2APYqCCOhETiRdFff7IZTwtAnb6gjwjVTeF8NERU8L8PLIl
2TuADABuBDTJC93rgw2s5c0rJOw5jcqGqUcGlDZmzlOQqK56/fbCqTAPB5KRthkrXeHEj5dOkYNP
Lo5hX77MBewvyLPn1b3YkmRjCL9nsS4i8EvQlWOmNQsZKt8F9G0CogamHoRS8JMptx7XLPD2onhn
rNTeeFo7/YNIbc45/P76F0rLEgZPsFia+cm8uySpGc6h036NX2beThRVnG2uEBzBxHBLeX4Daj8N
SSaza+hmnzcRtsuU+Y1ratZnsZC43qzfBz5jLNywEGmIguQin6kbHQranbf4fRa000B/VBEOVNJP
v+xXv+4CPOvC20GWxV1rXl2C1gL/C9Apn3A8y6mvZWxFMhOA4sCpRgcuM308qdi1yNfXbqY2Z7BY
qrfbQht6q3vXVt71rT3AXx0KYx4R6biUqCnwQjdtlRLeHUuJOwxPFP04cH9/6dOa7qIt+U1+dO4i
rGIC23wo+ZUMdbXjUalN8nyfMByRNj5Ypu3HDY/alt3kkVrsZwPLAmr0PMXAdYL3x5/9HqD9ul0u
ileHYcRCkgREhbtDeoUJYp92+wAYd5Gh0U+Q7F71YhC9/sMh65OTb6kOmioQhJap78BS2kQmPKFO
0zQh90d/oomctwdmNmBJaWBynyilcvSDv+r/9pGwplgmyzcAZwFmg8dUDuIUzRapBrwjPNgeoVPP
xlEf3kBYDBS6D0B6gB6b/cfBjFszIAW76lk2aS7jNi+4Zm+kaappz55JCNPPcbC/uZ6SaX5C5Elw
gihsjIxWDabCj1O3pOV1Th9NPa65I3vuEdkJ6I7f1lFq+hKmM7EjN5FXGyv83NjxO1KStdY2/MZy
CECeOg8ZY4X/oXoOP9IC85HZu146BL7vT0UqoBRDdRqLyxLA4hUeVtLx9FkwQRkQz2wUHsIGXks3
J/icL9KwUe2wifv6ONxT5rb7bHHak52PtINQoi7PnCnlVFXZCIghuOjw2P4DsN7zsoWzNqbuddlk
9LKPCtUO3aNJYDkV9b3HoxCNNkNHVbMku5Q9NaZ0X928XGdkh9CYg8UBJVFfCygYm1ppVZyYG59d
uqnKxUG8J1m3VyVj3mCGM2K20Ip1N4EUlfTGhASPHd47PnZc9FXNISzo/PZXGyAQAJbyCQnPC8FJ
kdbY+QHtos8OM/NKLig52mkfOdmnGSlyM7i8mwsJ8HTGqIF6hKIetR54Qk8WGYXlPzjC9WzzG+Jg
tFicNLc9jt4/7v1vn4eP+94VeFB52bjg88NYDZJTNTpPyQEdl00fNILRp4TTrnvBIyyug+ICiX2a
J2NDvTfk7jIlbg1VIbroGA8nVFv64MW+ZT38PiYvjYF1K/rT9lGI+9I5dvcmZWnC75QoRqPSy+2z
lDAkqWFKG/uqUgjEukqXyrwXGNUPUeVMaQgsWGU98rfFycB89gIfb0HyfPpcOdMc6Oj1Q2xLRFIr
b//uNVrNVppcoqKL/DeHBOAS8R3vbkRODtKhxbj1URtarmSWOLgk9Flg8UVToIxu5dUKzYf4uW//
uvLVY6JGe0WsKYKVxxIkMxPO0mdtjDrKA646/a7MpThtl31GKGRQMNJFFm+zeohM3/Ve3cm+Hg2d
Ms6liFXJKNrjtcSOzIFLU5WrIj2OTZabNPbZs/0KrPIFuPRpi540tR+ZqwUKatCvdMyf/gFOeyd4
ip+/3lMsIETix6D9ibaNTvG9+JM8RsVFKMY6RmQLTAXNRbyT8wdcB1JbjtR58hVVPFvLSUan0ptM
03bE0Ijp9SG1u0QVQ3xVBDVt1DVYcSkYlFB6Pw6Ed18lOtaMIhIPdsiNnog2bLxbiC5jxE3uXe9s
P4rPZMKe13tWUu1n8aaKtdVzTGvvlc1SG4PZe1O4tCgf5NQ0nURYD1Rg9L9yjF9VyvaZx8uRlk+3
XoR9MxKFlSytXutBafcoKJgW3WUyJRzlfsbBmftodsByFUYZv7J3C9QFk+Itk4oI6rtq5rUskaLf
43US6W0V4O7zii0QiTkkqtUnyWeJ1T8VVGkPFPv5vF1WwGRwsJVi6hIXiHV0RYg9kLA1NSJTlDC6
/l9+rv6qSF2P6NGrqkMEhGIec4TcRu/4rkZTIZLHXsrlRGQoVozNaLOwciAJYmfoWcZ59poLCPEl
80L30uEVt+5aHbDI33IdESdbUT78V2OP7jF2DglP3x/92vM+5M3LiG2PMD2Sa7sUBKHq5hpn+SJ9
Ir/VGRKxPBOIY4/nnreNfJZLTfhyGt+Eoe5k6/+/GkwLlTE606DhosSW6qZmqDeaNWZZWzQzj+iZ
1/gcBhdgwridZV4+YnlzoLYlyq1d1s5mgjz55c3nnzb/phHXF3uiYfj+xl3YDlb+htasuXfXTssf
SjnL7MgPCamdBS1G+WIZJ0n3IavSpF/egzrUQc7zolZLIx24GHgVhYMCrd4E+hHDSYuR9bW+uEEq
aRhFUziMtQPxF6XOPeQk7XMoHLFpPzuJaUgWi1jsJULoRnXGvjp39tVNPFEeen5Sef2eAEKt4X7N
3Dy3yW+et1++wZ12j24uFxoj5zf8XeUnahKWhTRXxEYFvumG4Lu+iRJ69Enz3oGrdocwiCntDL9I
uh7yqK6WIqDXzHe2UNV2d+HGg67IXR5jFow7q9JsJbvdmCA6eBkDD0IzDK0kNnjrd97qBFYhkZ/5
WU9JKPEN977pZWCXyAy8lku11paf4prWCGovgVQfr75R2y9d/9CFvbxV2KXRniYQ3yQwhow/tpSQ
4LJ6NYFMv3YMSGOrVD//rMO6esJAxtl2+htBhpph3dcjynv1SLZsha5dYuChc4oiMPNn9BZjiEIw
0tcAzqZdwfX4gQU2H/iwJUjcteBB2rzCnlHmWj5/uOhPzDGD9dj2m1Z3DPiJk8wihQh2ByOI6gaJ
B+NVhHgO9J6r4yp22EogeFh03BOvWEpQnljC7ta5ZqeU85M5Eio5hH4DxD2TbMNElQcvTWUtFfZ7
j4VYWcBTDzCnvtholJRz/1XIL4h+1cWDsZ6p1kQw+tXot35SIbi4Gps2DqvGU7ZAdp3zcOte+FgL
9SZeeYmFjKVzlbl5Ol2NeDhYmIFVE23VOZghqHhpVsib9blHGRIM4imsV4fQjnEo5gJMdVqohAvk
xpBSaUG4tkKt1K9YRCMnZrt+md6K+wj6midevA4J0ol3bNhfhZJ5gIjMpN/esJmZ0zQ6YMJwQrcC
eAR+DVPKE68suv4m2VQkZru2wjCdnTAxuoCyXjFZE/WQjmRRo2GMsFTsSfWG7hLAmfXkS+wXDIw1
ZyrH5PuXAkR91YnYYi3D0O6zdAPXQE6tuTGStDMmDCD/iJgsCbgGGkRAJc/JtwlNnBipyciRHWk3
2q9yQ04pUpcy7AxmzwA6K71XFue+kZum1cV+YrI0tzMB/zXM4q3gz482RjmJFoIyzYS0nlktynrk
eiShSzGMlcRW6NgguBZ3pJJHJSC1TT/i6u1X2qmj/JpkixWfn0RCskks0tIrU67DeWBJP2hwUrYv
pnN5dmf6M7Gk4UZnjkcW11+P9UpXsbzKucDzw9+RCJDRRpD5jbdBxx69t3baGvqDm9zd/1D4e52J
bkyS/1dAzbSsa199gQav3IxSSLDfByzs0Fbft2WrRxwdrdFHpAUqlccMkOOkBj0UaBzmQk3kGgcW
CCsI1oolstsYfUzB0Ii9AvMMMSvnxnqkygsX9NI7mRLJaczIsOeE5bkSim92l3Fu3A4OmiZ3MnEW
4S2+24e1ufCzzqmGG/SWTQX4TiQpCVGpqbza9rUcc5LPT7WJyOqgZ94m1GkIupa6yWfbFqMip+oK
qNovah0EU3db5Yf5DhdqLqoP+eE/+aGw9R6GL/o7eDibj08uaA+/ZFXlNNFB10/4g58s01gG53Lb
N/ECpMjYJae5UJ476rakVrmh+YdsU5mutQKbaBrJ/IJscmp02aEu1IllA4+f+pntZYDp7kNdxUwE
I6YrZcGIEyDMXeZHl+b/RYndqE9Azu3m1GrslykeDsc1SlH/YZiHGU4Z4pFXjncM0q4+q7hC91NC
WDNjffKFnNad7djXw+VjGNkb2q7agMBU38xDwk5EpbszIfXxqOxvMza8gFBd7XbpYF6vPSSDiKYq
fxaacwYVSe2E8bLyd9pH7a+6Dj20FtA3Vi19kn7Qyu6EWSgEBBiKqlqbZSwa7vLtHayMUsVHR4DZ
WvycntDRZBfVeA7UwYxDyzePWsitZ3gb/JgSzWkcvQlQ3z/tjz/MuFdehSe6+4YKmmJ4UB8ThF99
JZlgBGcz3+KrZOooIIx/pmDke+Gkk8vpeY/XaHXWbWem0F7XTM2+oo3hcwxgdjlpX/kii2g6fl0d
ruVwzb73xm1bdIMebXAL6+PTDdzPDE8gHUIkAyVyWi9P7hetfipje6+ZbKr+9+FEjMYhZ+Vt4XO1
PDweHg6jKez+/fnq6hbHT5AkaR0PRYFndn7qLzC5jsLWlr6DUPhiqHN9rrw9m4/oaV2OaEul4+9x
KWagNN04Lz2aMsyYCK51Roi6sg8JmITo638Y+NSTrJTN9a2Ti6N0wJ/l6c1vNy3oOuPl/Q1Ki+oK
XgWkHkrnSFk6vobir4cZTMrLyIcM4PNUPDoSZHmr3dPgVe9H10/ODZzNnIw7KjWpypoRiyCpf80I
2nd8d75MSRpfhTQrMqy0vLXWLhODZEPkNUzp+7hH5yUoe5H3sHBhmtn0GHCfQKkjRm3atw4X8swH
HuGXuShiGuu09lbjma2fy2qbkHTW2qVt06rh5+ishYy4br87Asnf22Dr2Zwl/KIW0uU1gvIDnmrT
lyrJt+ljvonyta8l/sPD4A2WHGZk9E4PwC8BWh6bpNhnBbgTr68B8W6TmlVgQIxRKYaHqTAqejHp
uEliiW/jjXIogEKWexqPhAPn1alq5rgm5w+axP8Ei6oPvc+djeI4Phy+dIG5EbMMBUWVVJcM/ZuT
Pe9SU6yU2q5IKym+7NPqMGcpEyUZb1EaizQKwyWSy4+FC7OsG0S8PtFOiR9ozpMKVfs8pBLMNZqG
cRnC8owTKX8yrdkaThY0ZH01CvhWSX2JpEYQujPZZYDXq/ROo1dDBwqOsR6Fo8O6PMrH5wWb00rL
vek1l7FOdWLXoZ6t7qo2Wf+aJi+aqJcZA95gD/EySG7ywqTMxvGOtUph3ig5HVt1OyauMIpyzs1l
SjbRwtv4+swL2f03zbi57a/9BZyXG6KE/qTwyATD6zeR1F19KHCMR3B7o2qLnu6Byv/u9YqLI+H4
UwITuLCB/Gs4BkSnHiwE2//tkYPSEf6r92JOIrWD6v9MRlhSR3cIxQpiZm+CSJ/R5EaG8JyexX7v
XuotWHi9RqittsL1+WFM6yKWVEsUmcBGW6MW3DuQx6KPjrrc2aUrfFmd0Glvv2Y4T3eyr4z3SQww
sK+SuBgfXSy7+bsCfOtPj0U/sYe6WFhie+oV15c4o+fumITURT8inmLJmEzrwGAL/t7aSXhnJ1kp
i8j+eid2CwLTjugZi5sUIa7a5IVwfkLdgL4KabToEd5fVis4CIBMo7Aptz/nS/5xJ92puuct/Aoe
UdW/q8K4LEm1ETxKnOPfDBEKdddv2U+VCns7t7l4cC8wJ8tRQ4EyXsjy8xSSXx0T7ZWWonbZzJ6B
oxUHu6w+wGK4DFoOQjw2Svt8uH2hw2jeCoWBFOoMU2brexKVGQJO/J70Q8POhqwT81SrjJIqR1er
0N4mMvyc538NXsQ/+S1ltb3cCfiRRSFRd5X5J1DZEfJW3mrhLu2+nz6mLHCwgh1hIBLNV1wDdsfl
FGGIIkDEUivx3yKIAi+Jb/c0SBnFz28tH3I+iHCvsijzg8hX4Xw6J/XVrgMy9Djcr9x9CSNun7dm
Vdike0ox5iHt/1jURUWbkTdwnT1MsQ/RbEtGsOQ+ncxObu6xGN59091ZCyKEbHojRrWARYeDh8xe
UGsnLRVjz1gR16Tzl/WOS7VvWRDukN/c0bIAXIou4f0dC9SE/ESkgV8ZUgTXMJ88w+XJ6HNTWPQn
SMp9uXekqPeSeA4dBitOQh6cA+vrU3lURzDTbLV++ucpDmqJ00bykZcb1ANTDn0pNn02CZlp/IYp
NbzSDefjs+n/pBVAnIHT9IhgPUP8g69pspmX/PgYUpeWPXOxDyFPi5KmDEq/X2ZVvcvSRULq/Pqx
NH9XdQbzcGO2LDQZib5+4yrq7ZkhQWbrNvNe3ssvMKI2CC/JNI7kOz8Dv1GfAljWEBqvt0n02R4i
8B1+mb7MUURivdLZC5LsuYO1NF+aTlqGJtBpxh9G7JmwrtqRDsUNWK1F2vYyfSW4P4/EgiHGHrBq
hzeVeEBJVryFVpql7cgPeufpX+pe2bkYWeNQ2BL/upgX6y7l1gZdLde1k7os547kQUaz9Tu0GEnu
kl+U56B0+YUsrFByDLVO0yY3sy5R/4YwwcSQ5GqAW9L4SWQ6uKKuQyQrd1Z0S2+vkWEEg2qjYqdM
eJ/Jhl7TPglDqfypJyPp0ewDoZd7giK4Ufa1e0e8S4ljAC83ZjVnm024HY1MPDnuldciFobHsdUz
JaJw/aERHWYdnMl7QLRYigy/3iIHNSEt500yiT4kIzSgpC6+4o8AMTybR2MphS4Pz2u9bdLqfgob
p7924qUWRgy5RuDJKo8PJ4gP/OE=
`protect end_protected
