`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T547rc5zDOerCe1OavV9oe127A64Qyjl9cRjKnbG0Fw1JTeAGcnU5J6hzlKQqmpecO8++i4VsnfS
gVbA/wQbbw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JU5iuc/kQwse9wugEIXtUYpy46gpWfwrW6Xc/SIzL+T4zp/mm3kFQzWAA8NgXVOIuH74dz38rRxH
rk0+sLcL3R2mN14y0TgKRJVcKLglkvO3ThkTEnkNb1+lJlvBv8dsQNa0SoPxswbR/Mc6tfTVgiCd
xmvW8RxkilgDEPPOaOA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UIGc/ouGHCFtVN6eZwi48jJ2YkKhZTWOAP3Df618jKPRyZo2MPV/+QSFUIMXIR0iQFoLIK/XtSOj
UN69rhY9879vhc8I9YSJlB7T+HQR/YpZf0fNBHVzQsuGEIWhkZjd63WVcZ+lNYFNrICoryYazb52
SsGFHuHQs2SoDWOcDfx1trW2YuOIySx2GfKv/UwKLExkxQqaqdXKhgM9N/2/EZKpIw0DhXa/EQox
i5e/kU7CJjguPTyRG/+JSqfmsGGLhUiHBfCNDVX3fkdEEgl+ZWeLps6M8Y56f+EJVPSmk4ZrkbTs
yhSMiA2m9C4/EDr1CXt9wIph7ay21ULCy3Qw8w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CERDAQKkX/PSjjx/erdQvrtLdQF1eIUaq0lCSbAV+ptOcv61bykhlz0NfCudbjFkmgBtk5XHyGai
hWxAMNLePyN73NyZSlfnYwY6S4q6d0uuZAf82NdpLJOSH4+IX67nwCnv7CbINNpeN6O+yNtKJBaQ
nsTaa5FlupaEiYpmisU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MekCaZ0UiQ+IrfzAZLwnEO2MPam01qIdbcdKmh7CBvtG9P8qT4KPEKiSZUNtXTnvP+q8o5f90fOi
eyYiZn1ha/vbUMHQdi8xbnnAdGsahW5iRKceBlK8r+1pnwkZsllKoBOd0ixcXCOzwltVM2KC73DO
jC4iIiCbUECE1IW0xa6CTyS9YHNE/LavsSDdKZ/vvROB5iH2CjsqRIwQgSMNmduNX+ldUmtvb8Q5
CJIbhWOzMLa/lIrz4p2B3h0h5MytfqGyya/q/PxUU/WuJbM155ACQlzvqkzkf7JjEK6/1GFE1Sq7
X0X4DGjfDznb515Pv9rLpDjky2mbrGonETlQeg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19584)
`protect data_block
c5SdzVPqMoAcucjj7/J7Ketlx6GKob80Ekt3p6JX0Y+QZBCZhzhEP67xKQxCdt96R849vIrJ9I4j
Zvf3IcdEUpNsV+r28FOWg2dxUBo85BO+xdC/3QEsLuPTC8c4mv1LJPttr/6MJXgDVLNMai+1jr7l
/VKf3/46hXu6kScBHen2KphEEYY36ORjreT4kvSYGKj4SsIfqQvw8TIzyEZ3MhLsOa+4UtiJ6U7I
dmLG3/q9IC2orwIB54jqF01496J3iLOgCZjebHBLyLyIeCrhgNxslWSY93z8hM6Ki5RpIsSiGjNR
H6BSe7X9HuF3JTbp2O9NLtm6KPeNEuoqn9s/mYU6JsjF9dRtGV9MRUvgjyYSwnFg7g6egfXPpfKz
mwtDs+BYIZgiZ1MmSK+O7NaxvqLXbNPK218zX6Fimkw15QxhCc8Y+/yePz2x7lYvEwQjCdfekZ38
O6lzhzM01IQnO/HnPA9Ug1bZrL0/qNFQWtcoL8WaNj0aZ6J+U+ixBhRX34TwnHmZbWKQgK2VpRyE
/Jn+sbBw/jznll8LQRcFAgYYqYfZfmn++Vz9kUMRTTcoirTzMTu4RZ8UPf3at6P+lv3poB7vdZ+w
lTfFQeXl5vyaZlkNdWHEZyDUgiB/03rhtPEVY7jEF8PLb4ndxkywlPWe0DS74v4t+CJDF0eINfqI
TcSYevtyMIkDTKB6vwPfgUYQEv1DOJRqKftiBSb0xlz/7WFFN7G0cIR6NOGwuNyjCwlLD83io4O0
HHFQ2JZDux2XYuZADliBCnzVS83+AQJLqW9XAYXbpMB6oajiIan8bG2lddWvJkPOR5FxhxqHmA6d
QEupVSzfC68n1v619kqWJyHW9R7vwAHct7XrHPOzJ20PSXtxqjtLI3zTi/69hx/k9CxTSj//qym0
JHGZUi1u0gaIFYp+yKAFWPJCOkoJCg/CVUY4B341DHvnMpIklxpFlYO39tBgGEEfFbsdQruQOK0Y
FCW36T1oHOqHqieYHSiIg9TVy1J3U4GLDTt9MDanG8AbDaow4FJbvXAAVT46SU/5h7XGvL63m4Gp
T/Vj8Sc2Sh/do5gMLFxI50k53huiVGuGi1y5/g2Wqav2dT4wpamHYr+8nJUlOL24wdezueDWpNT+
L83fMuR5NXfiq0ItG0oCH8ERBFH6dMWs7FJjEMS+HO56OzF57n/+A5oV/+5a4f7yNjynnVjAyaFJ
giCBsd7Oh22U0VE09po4Z/tBjhtQjWa5ks2vdBZYF/cGyO2vS92c3k69brej1x2aVRqy7jX+hBOr
R2bHL+S7sQzvxi5QCQAcLJByaKqNP+ot07aeS3s6a3HvOJREA7ejzxcVoarsslHkVrGDwZeRtURX
vyxBDjlcsmBkELYRwcYsh1caKVo1XCm6IkfMnt174IlSSsNHfQlVeqYlcvOjKhluiZDM4XOaezOF
S+ORzhdWzVYyCkIL3xd4t/EIgVu8KtF58r9FTqTUSIJK80FoB58HcL5GYl6GG+oCXEIrCygFbUia
Jhs6oMdfSufsInKFhuwJ4N2zo9ZLkRIVYFfYdQGRNtmPOFB1LT1vRtTajZh/RaaoX/plhWZrtean
UGLn2pBzRWAYI7A/IBjLkMRmfwdxY2Benisv7XHIL2xx5OQKq6vgi+JEcEQtwLtRtMZLIu+SBFnq
aGCOzf+4VgcaoRHuwUN3KbdjSPy7NmXNcDtKggIZdS5xTrzSfrWidvQ8IjnkOHftHqiEV0DV6oc4
cPtDm9guOi/KpSzEXTnkERPMZdXRrgBZPrkK++08BTIsYihQW54hhHwjfF91OKn6yYPRPtSnRgi0
C2t12uBTDsurG8fvXYVWvSB7/m/Jp7otE4wKI21FCLIEIBNsTSnYeGaJG+OZPX6pGa0HD/zdohU2
eV4HCrveFXTPP+uWTyOpqCvmUQ5Sbth+RIHrddRpS8vrWG+s1gk0ppO/t3FMGbz/nM9x6V4xQu12
KAAMmmKT5MZYUwaDgyxjRQUebdlo5dYygHK1kYk0UZi21RYcDOZxdsN2NUkfiOGrtralmCuwFdys
BWbEw2fFWXBLRYB4Ip2VMP3dBRm/a/zUZHMKiVOA8hk26YDGXXuJppYDb70tvAfAT3AdaP6nc1Ws
HreIebePnIrOdAr84neX/I+l439NRrqrU54VPltVdwFpWQFD3UjS1TMHskI8E16faybVtOruUhJ9
TzdFjCHVNtZ5c9ssFv7bfB/gEuV17xbe1OJk9MEFkl8rDSWN2LlklQ6ITSbsB2t9mQqGhKgrixw4
kfygj3eq0JcuRr7Sg2TKjWkxU06G+utz8OLb0Wkn8+tITwOIgc579tRwYFQqmdxm9/N6gRtLvZ1a
KNJhpPit5OyHYCkfwHHvNeNosW9sF19om/hutMtSO0oJFyLeKPlxeCS5S7uL76nhlsixza9R7VZO
v6qLCtfgut5JNiQUnIpLLNqldn8vKZONhQm9TUNAhKjVKAvsfvmmUR3mY0J/ccVPaKhmlMwpLAI1
6o2oSFj/MKKhCJ+BGDmonvIGc1tDMNVHi/lBMJrGfNlB27V6rnkS3m2IdJmcwjVZjenVMLzy/pFz
tspiIOR9uLpBd0B3C0CmH7GrPgTBpHFZkkzob82j01mc7+Q67bED1mwYgQSzPEPCZ/mEKeT/zYZH
C3je/nNQ4WXqPEpkBCgR0of/J5MOb8cTY3jH03i9I8uzy2oLdacpmGtfXqAyn71W4cTTwSZuf/DX
mrhyvrfYajc9tEaK42U7ZpgAVQhLLAXAOXTHVtMdALB7xsK1GJmdCDkAk9MNpfzssk93UkshlzOA
XE2+basHlrSFINyGhvB3e369t5HEaUgDHrS+A5h9J7k5hnySsq8Q5KtKoffs67H/sKb5NayUdgD+
5pafLfXAdQeJpHz7LATS9LmZE3CwpTEoCLTCsiI/cp4E/RWGP5QnOa0q9lbV7V+c9+IA7DOLt55j
eqLdr2O72r9dEI+c01ea38nf5TNNIlOD5c5QOo5UY9Aq8BaGdtELxEoxpbWS2Tq2Rcon/aNO3oxO
w497lulkj7DAMn0Z//XGqaaJnc5BNE1nNy2b+CuhQJzyng2FlqU36iqdC+4j4aKXDkEcNO9dGpJl
M6szIOJpQF8JPFZaDb9U+9+EyyJMJGw/HEzuQ412Rs4slUAMWOHLPuU6JBsQwRfT+/HYbykb4Jjo
ylnkLQgqRxdQY9yh8nH1qwAf8DZ+UaSms26yeXw5bjjgPA6jiVW43rKJH0/8JlVt0c4AzFF69JAZ
lGNE9R62DSaS6KAqoOuou5mbJvhPomlk0340nSsVhgAMn8TtFVHGI9DavpVK/Nv2/J4kTA1El2gK
Xc7pJlxNQRCx5MsEgfebd1YBYplkfYlOGuy0hEzw9GQS0C3bSDmqEwWgv/xgnI/RTyJosX5zVtUt
NXFg2WyIpDcQREbevv/WLrk0iqmGclEb5uYhfNq5uBJNq5QEwd91IjoiTGp9wJlCcwgRcpEig60K
2srXtXpMWonJgP7yK67LPemXyQF86kCYEdp/Jw+x4i6QwwtfJ+iLEiWOlnp0R9t9lBvOLaNHFwqW
jieO0BJhBZYkN0H7I7rcR3J+qwQKFwPbUmm0DGZ9jJR66vP7E/dVpscLBc1ci7RAaBdHkVKtLtGY
TKaLDwJ3V9H0BBtJxh/N+Xktx4DC8MehUnhzaWDcCkD3avq0gOhjZbv6YFmBxVQSavujAV6CvEPQ
vzZOSBTYq1WO85DTI0/i2mZ0GPDdHH/G4O92n4T2jfn+bfy0RTA5g7EHY7berqv0PXNZrFNmM2nF
v2Vl9E53hIfvLzmHwB/LZ63AzOWHZ8Ngi0lYLBs12JIsOnAABV5llHxD1coZt67EcfHE8iysAM/5
RyzGhr+BKwvEjIkt/d2XeYqy7Ylp1UBuYeTkuvFpkfnwwRhHZ2DnP5JjC/RVpkGA6fpdqBoQDSjW
6RVRf4JxrZBmVvkTtR7rkGvsAEJAyu0Se3rX2UDrnY048tuT8XtCdRQsaBw8y8ArOjqbhd4/Xxma
AccFpWXVZUijTDLIQA8HYYx9DHBjjYOQ4422Wk+syBKRYqEj4yF7TMyyuZC3LVsPp+YXA/4LXSY/
FoIjjT+AGhHPP1uliLbGAiqO0pahCYXEIqX67AAlbmzpIoB4e19nXJ5ApFDs7KHQbfVZAt6NhaDE
z+4/OfiAi3RCzxf98ExDwoMTMZOEbPp6WAH2tZtyJNdBuyolmp9WnLdymKaI5ytgBaYfNHMWJ253
9bqa2TOWgIwv2rakGvTCr2VYpU5qWzlLxLdtFlunrSq2vxWz4zl7FN7LNVgvYfx718xr6uJhaFbi
FmxyleGsLlsZpCZ5/6PzRD6BKzUFdWShmBQQmZB43R/0OLdcdXihp8zD/B4Cn/Nuqfx+PDUBPCP2
lALuUgeEK7dF5Byn5QQNPXJZ3wkYHI8YQMzmzojwra5O8EZnLvyH9F9HTD3lPkaTDERlPmBO9BDX
T8UNBHPFE6DbYM9Ulh2e1bGuoSYMNdx+ytZ8IDGWs0yNdzMdq5dJSLvLzd32LL5AZLVJW/4/JWs9
DBFNWqv/oFmciGO93+vz0Y2RS2IMs7dLlD+xnWWOuz0iZfHt4FWRZMDjz1OTPf6HfZechC8bhYKo
xUuI+usGwrstk+QOYqW+FJP8bnBEoZZYx5Ru91H7Smldoi3nel+Ef5YhgCY/PAWwKgrF6b1OQInI
wcQg5Te4OU1UAc9K7Y9WeOXVIKDqjZrXxb5xMswyTqRprg3nzlycflBAxTeOrJtH5wGLSaHBDSNY
m82qGRlB6BHhOpY/m4CQtfWq3dOSeYfqBniiaCgoJYrPnwgqk20cz9V3xvkEx+7alsYMS7GNQf0t
Q/GdAyfC/0vespCUSoBZkd1iafhQMH7d3MvscBCOueodqXBFWYU/I40F71jL5KsxnsUqOCpOjCtu
PSjMkMNssIuhjrzm3SLsO3amXeyVes83iCQRf6DqPPWma+Zq50TNRdKWJCDL0v2Pfx2KLJnO8G6J
BmF7Cvf0BbDHuBHWEiuyWUj1OFfMUvNc1YEJitiO1UOtqBT+9STQNsbI+kYG5mz6OT30C38F9biZ
l+pI1qqsrFXcFESC0QGCmgeR1O5aBhTq9ZAoOEG9U1AnWq4Kxa4v6dCmBv7ViZLgmZ9VJxioqGDS
G8lc2P9QZbtSBqgaLtfkHpMNUQLZZQvLE8W/VdiOVECYKPEOH0GMaUxpm37bbDokRgGkKnUST+if
k0veKwsb4f7zt46dYLdQ5qJ+Hn8LJJDBhNFxiEK9Q4DqaB7Q+A63fbsoV8ozSNTikv1D4HSyhANx
acvRdNhmJ4yzj+U3q3ebVzyctUl8qaX3cBGgSgQ9LXmIHR5HTYx4Rrk+/WWWPLi4JlCSs0DzT1sI
vm04UnXqTbsK7HvuHe8LVGsp9Wfof16cWaEUTE5Uk9z3uFz6LsDBTS93VyqSfXBoGuSRKVdGejou
YTJJOE3xJuCAWAzTMZwHf0zDVsqwY3Y52HceU4CHZgpD4mhbGL3RNtIg9XKXd6mo2nqe+aU+hF3W
cb8cNohcKI2Fy+GpxplfRjRa36WpKOMs8j/SS7SIUMhhu1x5uxXof1O499X0gGjatUYDaevjKqvF
zv+zPIBgn8m5x9MiyMb8/fuvxnYEgMe0Pw+GOTzCLEbN602Xh+8kY1pL6SeMBVzhdXYJX6Avdlzr
5L8uSmZuG+cnopGoz3+tT6W6zqQznjPjhKltfP9zonWpFcrPqjrL+TllEK/tAjFcYRR8qIIUg2h0
3QTE9ITiYOVyyDmtZLe6tdBK32umqyQmg2fUHIyKW/c7iOZ1ckvm9xtUu8kIZyQsvHmEfKR1MGy6
EwEKJ+6tzykvRVpPYOX5ZbLBfaC07ojrQkpUIhs5NN3wJJKRrUWlr7YVpsE36KFmlJLIJAH6qJOZ
6NLbdHwXZ4eFiHa4k0Uc2tZG1H/m0ffRdZ9JZKW5XCSOV9QRjBoe+iI+oKYRzlV/OhCtkNzQqlZr
QyerAdXVymyCG75o9tBUXizVMCab642IptH6BRx1JJ0uw5x1PLPtSmRyhuvKR7SDfuvqlG6Rzi+Q
n741SmzWBeBEHZvvZRxKe908OKM4ZmIUYbfI7TIJE2wAfq3Ej6Uuqc+FF4IPIco/mZ7i/+8eGVXq
/PcZKWifWTEpx7AZwE+CTcz/y9SX36prHeqW+gRTtKQcoy456N8QhELaPfMYmaCGQ2MEakcaGfP1
TW+l0WjXBAxQ6SsM+nW9Uvs8PJ+jFoBHKjlvYS8ucHV16uIjl8AeK3Uo9ewriaINxg4yUKtFTJ/5
2mX5ex2SF6PQ9OAmaMebLluYqjpCUCjRbo2K2kVZALFT+LB5ExKXcqgw8pVa0mkZFMyMqnlgW8HP
MPA4VJH00vW7PTQkKNWsYptfTV6ImGBnMCWbBsq14Yod9bh/8e+iYBg+D1PjrmSHG0VgsdDtMkbj
onRLnjDkCpHH2yEVwTzWQALKAsk93qlnlFqD7ROKdAVrLz4fFNSdrDNeEaOgLCcUXLbsWCcOAm/W
HsGB3DsEGe8kBEE0yeNYg0f1I5oa9f0Ou6J3Rw/E0F4pJVS0TnACMoexkLufUgEIp72jCs22A/aN
LiYYHQoe6LZOEjEA3PTK5t+IS1MKg264yotQ/Ge2mjfcFgJndNooslu3ElL1+jJh8yDffGCmSvaY
YFTbTAXlQQmAR1HnsIRLDvkpHC8U9TEP/NzLZJLnY2qZ9GVAuEQ1UTogTXULjouAwD+R4bgC/QUY
aI+kich8rmdMCfV1E8YMo5tlAztz3phZdy/TY2bvAdAbhU5p3Onpo/qbG6p/LZVxrKYYRSTqUnRQ
lALrRbz9lPY+p14/TZ4siPwhqar/V23nBsGjK7yufsiNPpPG/0D+/2HAMijNFX35IZx/EZxnCA/Q
tabeIpY4zeXMD+V1AGNqCt7EKcJMqvt748FapbQrcJkuVNnJb25KMNWYgdPziTVrsyKJzTX1XwAz
WkGK4mKufvWZX2A3QhiB3TyVqMNUN4gtkfSDWQ6IWsxcuRqktScBfWH2VY3VmiVahajt9Ub7+BNu
FQVvii8DH1XR7XtIh8AIzb1EoL+YD7+IP/4gJ7D0isZ4cALhGRSqQfxjLTc+7yOGHCqfBR2f1iQV
OIkXKCJCJ8c8+p9fgsCuWI/iMVYdlbcROx74islzxSHP5VfjNY/DBDPeL7OMtX0AvNcScC+vqnVN
+2NY+j+UnSk+dF/vyy+aHdzCRXvZjrj4bMbsL9+dRW8YtpDRoF3ma3+DMG2h/phtX/ztYXp4iAnq
kpU+9WyVHcyF+HjTFbgA3gL9XbrgxlCwAQAIZEL9T1cLKyp/s44LUfmDNAVIDA/YmWkHm+pAwO5/
2X02MBK9pcLdPU9BE69d44f65COjbAcVUiEGHJB+dDAsTfa5MHMhpGENUg6bnGhBfP/9oZH2EjYH
HjsgX35nbjFRNjHkAfwhS2jDi2cm+v0aSrdzFUdGmNympzPil1mx/gRXV0cyww9k5d79hRKzO31R
jGv0bFNMn7Hgj92ZEhXzEdgye5bAhhLzHtU/UARcG9n3gGTF0b2IFcC6pt7fGWo0AwvR3+ChoGsz
5k/tl3iE+XEPAnQgKA0ZOX5GiA4ShVVxD9mGWdmdRN9UosHmqVu+nEmpSp1lmfYUEyROWzb1L2QL
qvdt1c+BfkKj/CR25vP42AVMQltAGiA7Y9JuFGvRX7/nt/FW8qcmEbWdSPiNfduut1RxIGmE1N0D
xSr45dkI6Yk6+1LmUpFSr3DgqwrKtzQJGIfGTDclcKSQenQskSBoz5L+LZU4lqHVVDUhf4OdQXLu
bzeR+diBVXqU5aH0hQrYnmQS5er/ofGB7Mv1FSU8plEf9TkJbIceKbw4jAc6MTCAkGxtQOW2i1ZD
Hy2n2OxwodPCRZuLTjzDz1ppufVJ9QBaMq3wt/iKE9N1dxxI6TPr+/MiNuXDJdaNR2RIq0g7AVQe
/z533zWS/a7/KpWnFKArxa196M2RnOJQEPxacakBWYFKwtft1e2PPGTOu5g3ZfJlODgvHpsvsUK8
cVXkJ9mD9Tx2HFaH3xsUPct+ltpqEedVK40711T/guPXCHB7B/z3+p955Dj2ibWUwhvs2qjd54Sk
TEOnIOB9maz1FcVk4+lA309mwsJHgTQFeAKZzCbRUqxw5hkr6j9ESP73oNsk0F+D/X9zZlnS+QaS
JjOM4wLHcCMq9A/IIKBmVwII7gxQglwezb+nDpxuKw6OEGoVgBdZyut2xK4ieuC2Ihn5JlI0H66j
g5E5RbgPYZG6M9A8LCmemKFUEwRaMTQSSPIzzoZkfvBM5U6GO0uWdRH16epOgYSn0zdQlRBFkP8q
juo6dKd1+KCeEw8JCJFaVKI1LurU53ELbgQONJxjwzrrGeCAiBzx5zLkWX1b70tdR/XGglKnlm6F
EK/XrIIKWvmyUxbFHqg+P5TuKC8wY2eLkIVMOhWpZbZRdYyEZ8kubrOMZBDoj6LOyPKUsgyl0OVR
rDpLWwUiTpjYXSRBhGEXReImY+mzRQnIDZamXD9HDCsHPAb+udov4XEkWGAwqOel2dq3H09ZInc4
85+RpDqrblFLC6Rt0WQqZwdVoeu4y20PyGf2lSY5cHdJWxZHR/xqyr59eh+dZB/OEPy+DMNiucp+
0KQ90LVKcwHSzSinVwWX8yJQeskOa9o+6BaGYU4vDNkwcX/6sm3i7FuwpVT3MxOlUJZ6NED6mx0I
iFPSkuK6Shvbx71Iz6sr+Qp58IDjlqmZCjgl48rVwPG/xgfCp2mL8ZtNV1cG6k4K44ADC+Okuq3L
TiZOhEEHrmMX6q9mGi8p3vfle9U5YDoFJK+bBIMw9COZHkRkUrS2I0wOAVMB+El6DyThvuUC69Ez
/7GHgjkHdcemV1xnIzWLdF0OX4EYFn7QBl4Yq+ySG8K80PoXNuhdGDb2kHwrkVrjXq0pkypUerlZ
5eaSNeMUSeoWswo78eMLwPIcB/a3F0jX0Zc1q6znHuqhvK8EGSpAuEVTKof64E4mBCcT4eWUq0dS
gvJLnHY7F4cZVQLgwfFr6o6G096pJuk8Oi1yAXJIq3y6XNLzFa/XdYTXqX3530ENtFlUSnRA4691
DzD0by/NQfUFUYnIOLvV6Szy6X21BDksSfVCMXNYnmgUAc/6K12vLzkkSe7m3Uh32YdVS/QbgPvb
TktXtv/2DWN34PIv3XrPOvoDelPaDr5d1JYQL3HUYT38k6o3oe2hzTgZs5Ac5JqdCmldoJFxwW8l
0B2IqwGYQaVhNBO23Rf6P6rNJbB1DyksLbe408QgK2iORTa5VB/bbYYuS0cyNyfiUXYkv5eZAPyz
XczAmk+cjwHPKTfzYETLa41vpckr4oKl1/E86wEIVg1UwaDV+zUqHj6jglR7mkD7OSl761hcCRcS
pn4sBIwg+lsofrp8pWHCTmTLTyqaDsdo2t6BawMSUb32CkK8aTb7hsonM24+8aUa86KFum3Z+CzB
vUCoH+2KUq3WONpz1k2WDY6pWODEFfHOrx0EmeUy7LqbEcE956BdlNQiFRJscP5UukMC7Aa3G2iy
RWTCfQR6Gr2CZKVvQ7764u7sllIZVcbnZcv6xjYvC4W+4N2qPcIgtJigodmDXXMP1+2/wiJAGOxt
UONOtxby+Yz0Imu4wKiJHfIKayaaCjrIJsAe4jVwRqMWcaeYnEHYzp5LFwZQY3bWll3/aQnxvifH
kuv9T8vJd18K2XwrYEv94Zd00ZamEz3mj7DFSn1y38S7cNb30+VHTeASAFzYLqMW3NBj+Y+KlMcd
GANZEQT48OF8KV0hJG3+EwEbcfI3JKmkJqjJkLNnWOJJPcRlTBnSKxhXaZCEX6hv/qLCjnUkM3UZ
BBqGRe03RdjYMOF77NdFNQyws6q7bVaxcXBSyH3jiMIOvFfrxOt5gmvF0YnuZCAWWAygwNJYWtF/
5faBDJXgj4N2Z1Ejh1bJAXEgs/Uem6ABv9/lMxsW8mfhlu96t+IKi69YXxL2sibIY+uZS2Xm7gr7
p9MOgpcswofFWZmAHRUoKO2hBaGBQprQxeqkKv+ykl/c6WPGPal0WP69gwmksG1opivrIiMvSdOr
b8yGWqnXc1RGQaLLy4OlIsPKfvVjSK8Ovwhh+7YRcVgCVBA7/4xlaHc0L40bN0yIA31Kjv6Qw592
UuAQRtcLVW1frfrntWdmKhJa/mNn+L+anGQ2YNfKqSrv02vVpFK2GWsGu+8E0kRTCY1Vq8cztp8s
fq0xTvmSedjplCip6bMD2Jhz2nXo3sY/bWPz8IhQCokmES0gIMZvmXcJ+d0iSlxxeTYCTnPuqHqU
Yn2Q1IRK2FjT4lIzWeHNcfqIER+JFMKnKjsyA94m/GE5NG7scMZ56fCp21RGuyp5JEatT5TqjTOA
z4tzVIT/HwayqrLz+GZqfURpn44s8fVTRQayUxtufigwMk9NPhXypPUbbpJAsoO26oERuvpjCemo
JZtZMJXHJnNngD+gBls8pdEEcyB6JqvUW3US6jJrPhs5iEuOfVPs1DQlRuZ/XmbNzbJH/OvtnMKZ
nsIm+WwLyDSerjxsgGa5KgQVhbWkf3n6h9vRNxWGZ8JumfUXdCGkDHVDaVXtBKfVv/hV4xdQQtx8
Uvqc7KZsI5qRYbEu+lSLeGEzf1h8c1dSUkZn3pAHoOUinZrtqXiwQA5TPkymU9QWhYnb6+fyKPg8
iAUYyYLyxtnLvB5/FnG5xYZSyFInCvWskOaC2OEaJwjkaGMb2zVoYIE1qP+2pQlm1i3SpcSK7Evb
Y0ZL/WZtP4iTdmsWmZYKkADh1xKTLJN1eVKXwhzB97NcTfX67cMyT7tHEcDCPHUxAMAGS3YWnW1a
6WfAz0QZZb+MWCcursOM8mDEwjkgjYqqDPnbXIKIvPTqBPANNIEkcuX64l2FqJXMpT807S3xvZRR
EvI7NglzpwKoaUMr9lLHNs4jGaBIqXT/u+ZVvNehKDB1dCN/YnFe3Y66gRoxCLf0IyV2HI1FgX3O
HORedu/e9FuE8gxwCGN9c/817TV4uzxSJoKnAGLSe3L39EkCpedgRDDahQfC5l3zzDNIHKWiHJhY
S9zvZuDvPwWuDY7e8HIxeW1QJVAY3HFCUWAAof2eOq+RdF/Y6XtqgVf4EaaCWzjWZn4Cv96/Jmzv
AVyOPbSxBxaLW/WJZI8u//fYDy2LDWcxEa8pbpCyWUF38t0k4FMVWQu4GevUmmQssQxYnWUIajxz
v55p8eMHJt52UNW+0Xic4ShB5jemAON84nAA31zPJRhR4G507ifULYzIWi+9tHTRzn000nWPMWGH
F5ui9Au1+f3PGZ+4rU6IiLsH3iFA0MVOtwWt5SahCdoSopmEWIslwr0Fj4y3BcXhX3OmcwV57h7U
jDIvj1Lx06rSd3GPZn/8+G7iBfMTC4t8v6Iu3qsxAS1byp/YX6AHh1BgTBxbb6YC2wAss13mtDji
x7E3PvQcZQewUJWVhiycHj2Hn6fMvSlGu1UwXKvx0OmozAUESJ93NWbxxC5vPEI7xfwikWvAGhQS
IvlA2m5HqUDfxzsFUGgcxob+U18qoe6tWRuK9UhXTDUmdLvoloRHIe7aWpbeyFR8/8iyAAuNBAEw
vKofR7PYU2/wZBOZ8vd5YdsIoPnP8Zw4x2A5y3tRiFmWYfpMDo1bhShF6kfyVFkcrHPZDzPG2rvj
5PhqSUk+/KbkbeOuFr0Z/ewXOPQml5AaJwWZzgbdKbVkvuHvlf8YY1U6+SsZGnDI+g8mtGzdM+uA
GouGssia0c7hGTBNllw0V9WTdG+5iyfQGhlQ0PtIcSjuhP+y0PSRFFg/MR2ySh6hWqoyINVMpUl6
7Q4KvS4rDtBLg1uaJFMR+Cp//OVqK0fBKehwlMj+5+6k88/o85i3Mn24o+NxNceNvSdGQ9lE65nj
N7/Md22SNORu7WsCX7ONpydmbzZPfJJvXudL9z9SltMKiCrOyiwK4Z7IuqyPkUAJHvTGECQYzARv
CxUdjSjydrGd3fl31p5nL9DS8HzFpUzcT6Ql0iJJJVDLdqbblZ6eCuqvqe43QT7jMyCL74cDyOyx
jjsdCwCDJa6z3JryXJy6EVzUF3iZc4FML1bqHpNmWT7s2iOoCBY2hGZ4MDE+2FVB1GcWGKvpLDxt
34dLvUg81PK51QitffNWs8MkQumBeRT7JB72jkkUrbnQYsu65lYZv8PUVyuVfDmNJc/EQ3k1oqgE
g53GBCg97O8Pf4Pkt8pmFNxkbz8TnigNuif//1YLIcwQgam2TF1LleX6TL0hNaeNLzNoGA0QkiF3
V7Q/x6hyxUXUIMUGZTbIwbBmYwMF9N3jhq5o0Syqi7GLn9PYrHwqiAY4zMJa/gnqvU/1gv6ijn/f
JrF1EPv+U40AukAufRFFMyy+YbjoFTbHL13clB9cKF0mI0+P2r6vFcOhmd+2JygztgJn8w++kL+n
wL1Fu9JByu02jSqT985kRXsIjfzc2voc7rv2595i+dtHKbsu3Y9DbXhva9pQUBCxpMJEh5cr96kI
W5rNnIip6O/1FIbpODfn+mjkTXFBMpjFy42ywHrLeMFkuDrGBy+nCPA6YJN8f5HvZZqP9Gl9Qtq/
3IRdKd2nH8phBd9SfQLAU5On8/IWry/ZuwAwCl253/7TAxsjkTJoRRJOu0w9dA8j2a8EQ619sGX6
eCL73okpUZ747jsyfL7y3ulPs+G1xhuPGi6+F4rEcX94bWYhhuKhJTvEe61KT+7vMK6V1DK25jtx
nzhzogCbXHarslW8JtwwlXtMgHTc9dMlb5is965ILoRVWAWcnS00CQcp1SqJIrBbnoRay9vwoQ5C
Lu3GVFggbmLJMwbr+qPTDT1dtlMcm1KOiGgo8JUOQzTnpoTkwLFxt1RSh81vNO7PDAqt4PaFDz1R
Ha+ABlLXqilPaKqTfH/MC0OkEtKGHU0QdM1I3RaaKkrj5eXzVuFJinZ0Ec/Avb5H1jYrkuU+Apal
vAtKkcD5p/n4FVYRUSM0AkPHCkuXHjTdyYQ+dKNAU4NfRHgDif9b5aCYlViOkPijoZ53GWMu43+s
q+JxUfpwZ21TddXc45jm8cBniJGIywMa40IprLme2kD8rr3y2eglrKkaqlfaQu2M6EbW7oaJLlmD
TcE+cweIFcp+nnc3FhBU5Ka7AtvBwFtD/PpMvFXuPXKECKuvrNS64WnUve9h9H1Hw6yJCF0K6aAx
JAvO3XSBujvlqu71ucTfaYoMoLW9tbEeW7LTNRo+nFZGWtulapOnOi0yvRDsn81alQrJpw68btLe
P/kr45eU86UyVd1dMz3+bfNj2PbT9K4NeEbW49CS+70G2pImzVlFzOSk2Y1P9MZcSmRsb5LEW5P7
JTfcGczMhBSGIbWBb8MY+UOF9F/HiV0tTr+jI5fV14NwWfEKYsmmJVMjo8vPDDP7RZgDoMbjkI0+
qeAkfnVGVGk/6ecI4igJxg6Zx0smsDwtZhQ9orQAltwYVeIix80q+elURCG9OPtRv2/0gxllbCV0
2Ak6tCzBpGiRIy+BiRtbPY02Z6PjrOfA1AL0it8hT0z8NW51Wwbmqt9I3VcRu6aYDAdgjzom7tj5
shaMgncKI84+JdgAFmvPQD6w3xUEC/TmqsV3+fEpg1QVfKvlxDKp8ld7zXix4x0q7oZn+vEgaIbh
/ZZpviOVZyiOol+hJLiGc0SK/n9ALpHUjCnrGyssaZqzA/ca/I/ere84fIz068si1FqQlqpBNFaI
+g/B/6gL6JDRt2IdYuCTLV9LqTWRQxJyldySC6gM2ZXnZl3sXgrEtfIJRFtSHuW5xCKxDv8JbRVA
ePngTjwoGG2DlJarRkg+br1qKILE/RGk+ccuV2TA61WQnIWI79h59JsgxIMIesgfY+M7LXRORBXl
RXhffnW8aL2fSvmO+wtReQXu65Ayx9lf+JuRGur7M45kvylqNhXZSdmaiJQGzMuRqGkVuz7/Nhac
WbGnxhuNLrEpKekJaAo4cvf142okzc6+jDdMh6O620J+CQJDzvxG98W5nq+uayAvGDrHTIeL2qQe
kHW6fwHtBQkxlbQx9GbwQYgREm67SeenV3mE+EvF57FCOdbQb6l29ToktCu663M+Inj1JWK6BdzY
JZgy/TVPJBVtmjjMpfJd04z+YyfrXK9J/mI69ht/AuhGufBfwL5l1zSTyXffpRTDUIq8E2QBo8dY
soqjfhTObwK8wm8nR8VbxLVz+MLsD3w9Q53axTTLPC/tduuQX0Up1VZVxWPwpHx65qZ5ca7m4d3m
VUX1w9DLiPgGm/e6iFlVnyLv9c8PTcGIu0Vez9xvE9boSC7VUv1hAnYsg7fRkFxRWx6BvI5YpVTa
WFmYlFB3+Xweb/8fC5w6bKTCq7gX1xXiNqxbG86WNdpeY3DoMxydB/jGqMi5efaW7TalCY/0bvtA
ytOzMDyEplISbhGsNTwphWL7xUNtaNzShza9D3Ky/MGZ3swX0QZw6MV0LFpS3A7WqClK2Sdt4aY8
Ay3IHygSHDtFswww348zhcvwriEjb8G+p+cmGy6EnAGO8PTm73vcUW0AqJmir57+Buolu0yo9l6Z
4Q+DcE7pXfiVflXmhzg/uMUGqfe96x9zrAPP9NnsZsnF8mvNZF4wcwvbeFqGjF+tjn0sQ/XjCQhA
Gr+r/xVhZhkZlRoEFwwNP5eGKCwTN6HrDyHqlDOmYnePia+/4jAR/UEBGFHDfvW3f0rSgGf+T/NU
6jGCxqThFNJQqbOwrBqaBruWVLnYrHIIRSX3clTn8Tmbfu9DTM+54/VXA8vi9O8Tcit7wR/VEOsF
WVIxgVsIfB+n9fcqfnOO7nlHHIR+DKcqfV6ueLChTqq+xIk1Lf7WedAkM9Az3GDFpyHlL4cEhgiB
oOvB04moBMxHLIgKh59e1mHIzObQqc4ekYOBIOzps3TwXna3BFUIWZlyC0bra0fI/cbnZ05JmHLu
flCC/c893tOkwoFfN64GHsa+Co4HgTJmQTsSW43h5TKfJnBaxzEvo0dwSrbSZKf4z/iYjMUvycvE
ncibK5NbjHJHCyw38h7/Ba/GUz/IQOKFyb5l7EbGu022pHREu1zdeCC2xkw17UWZXqMwgX5fpq09
5jNZ7h+R+U7bFYOW0TzyzKs8Ca3gQx05MY2atxMPGotZsAD4gXSNmnrW33ykN+tC7VEdpFFP516B
aYlHt4jrgqCLSTSQOoTqwTuXFYcN2TiLBsgeFAarDwGzout4gW+vgc8vEswy+N3aNLVj9rM2tQLl
tjSXNMBTDnR0RygM2AIPywnEschGG3+yW3Mh+WLecuLuUtG8SRiqPVdbjSAfYkRqGzZCkTTx91ZM
qmG3lKMjb1U758frVWT/hW7w4YjMYYtbGfGuRowbdEbt2kY6NVO94XVO5H1MdVf/FprCUMjPPqO/
jLB8eKWV1tIlOql7GHG4YSMrWfDHvSPIpxa9NvHmSVvqaGmDJPIJQRMfXMfkeqIdYLMhGCdyWj4L
8OiWr9pG8uwfDCyyiYkdKh+w4arLx9kn7jXq53gxah+hRe6xhPuXIOacH/4B6SUQQgrlAHrpfXfQ
j6joZFtwNSmOpXswn0cQinMLm89g2R/xTvCkvDoCFq9gMqXT5Kxu2NTJeujGBL/DRijPTBdNOz62
ruTtzDdECC5iV7NKeUH1KE8s3kgy323p43nivhDtTCTaN+uiP9qXneAORVKnh4oXEqNx8xkfita+
aUGn6wl0TWRwbMCFfBwZxF+tdymEkLuaPxwN+5SZGY38Zo2e68tvpzh0R1n8O8gi8qIrwlhg0HQS
2dHk+e8x2uMIKe/KAqzPlHdRS2X3ykmY4pGe19Wg45gj168kaei7H9MvXLKU1HADbVHj24972dPg
weVGgTAUivvSnh2bEYJj5ewa+QwBijR+ZoNdRl7SQ5hy6LlFJz0x3BmXUXgmxp1cFkU4YvB5gnZZ
l/Rgij+NmCrcNmd7jqrxk3Y9mt65NwKC8NZvzCsZq+Gllg1Y9ptMx0bLZzPPpVeJM/lQCx99Nc1B
aIObVODnepLwmDBezK1ZoO0nVUKxSBZqCe+IfCMfegywu5b2YJWHUcq21r6Pl7wCPHWClJTHmPZE
qisb1mB98VBPoJQuQRyYomY//YaIACFeWtZxp6FpE2REJ++fkvo/TbqJ0D8Lhhd7DlZA6VkAmwlI
8HSybrbgphGitJ1w5Va9/WC6dNvKT1ca/VbFBr5JUAuCA20gW9SCuxUZ9DZJt+LqfmCEmKPsq+Zs
ZUUAzfL8DvD/ZIisN0eFYL+J533nmU2E2tjB9kJMQuVWED6ujDPt1lNl3i6zOrN5Sio0g6J4/pFV
NoMrx7YcBPT2/7SHLANMXxLptc/lld7zha/2DJoxTwWxhmhWNLRBDLk1jEABq3xEoBM4Ix+pjtdC
jqL6CwCRQpWMaM+MCJeBax1WzTO7Dy4DGPVeFowkWvnLuTtj8RKKokVyiUf2vaWH4Hx58GIHSk4R
ZKS4DwDqxg3HuzrPKg1GWIaoBQIz9IPQp+/yVsAk2aQeNYyjFzhibHivsGRGQgjy2gU2KHVm3dJx
lqPxbg8dLX3jcVAYdoYTv9OD7WhmDDKd6sf2oM4+7DWkOeP+Md3V6WRxA2oxBQ18jej1y/5iWyQP
sOrWI5jFeGvE0n4pN0wJJ/7d1hLjb7IGD/2tq5w1qvGqwP0TNAhkjEdZmSyIfDEnsOxqlYvIadTD
nDmADglVznJ7BZVoXtLui5C6833jgCZNq7LlixMm5zYBopm/BkNsazObgwaKh/CveWbN/hJy7k0X
25KBUICaEg8bJ/Z5o3M7Nu/mUWTPq6Z9qWNVRcO0ee4/5gQDHZCg4AgBIV2XsaOl5uFCaQeYtnhV
ye2sk2OOcnMDvBUL67Yu3fEOi4wcL7SdpjBExEdEfnI4qIm44y/NQjQNJAgZT5dnoI97Z+Dg72/p
9MrSQmon4C6aCenM7fxP33LIkOjBS/3ywVEkWC1NOXzRM2ppCmGXegtsVa4BHrNNZjjyg67G96Z1
3oSHZbpOWZGbOiVdRd2Lgsjk7tpkLWBPcKohFPRI2n18Fbj2B7JW/SUJF3roZzsPD3m5YPG4QCeg
xzcTA95ygJKzch4IgSfWbcSi+NTIvKfK0n71bkClIaZVsW3XdgNVy9v1jSv/9MjEYCTJDG9RFw6s
nRC/u89PrWO7wavH3My/freUvo9fLjzr85rreFfKPBTH/zPVIwPpHyHNajQ52YHrnZaOcz7pXcF4
AkG6L8BGAvSgVWxMTPI7eLM+UiKMmPCm1lg5dbPnNSvcUlchNe66zbAOPVAoCbhJZLmabLqI5VkC
DgoJZSpZgGiLtynk6dpNBom20uNnCLVAjrroTTA5mNUP8IBDLZI4yxxdj2rvYR06A1gEcmY3fxGz
dEiGvm3ze5RjbfrxDSwHP02MP1Yg9lB5C+y7bjLWyAQPoytimgz4g0tZRJiK5KvuIHT6nYOo3Ytt
XTlRrYHunojZ0zkcGh/3DvGuJz8fa8xIJfTDCTfiF94g9ZNozJREFE+9CGBTLF9KuaLjOY30F3tk
s4Nlupoq6Ote1xDvvR+s927ioupEG4aVZJhzK0TbWQirp+RJXBI4j4tpnAJvvowZOtCkEyVRo5d4
DX/UcexWSpzIy1oxlDOmvzPOdmam+JWBUqNER5nL92te/JeuiauBIyiuL17h/dF5JXbBkp0aKfAo
MTkOtAfIOVbKvyQYrJqwqCPeBcFtRMvuhniZDFme5CLCWpE1UrTdhqMx89iZGlc5vQxA1QKft53K
05cwpzvD+6OWPR07hInCawVSQ+l7YL96bwznuzgQeOgENJqNFjii3B6cSna/ad07uL40rPZZBPZA
LNlOhfIIozDgfjS13uMWlLAu3m39MpYgjAFRu1WT0VvPJ2KrUG6LIORJGazG3ZfaCbJQiGg9+AUL
yFu4l3PO2krWjux7tO4iBJH3aU7RYFBYfbvfbsmblY7YInysWUERf/uJBJhYnoOwNoMtxpDNbTQ7
Z48d8O0rKGvTpF6Xw9IqocPAbExxDSyq+5081oP4NAWnPhwbj1VNO0LxulYFVepkjTUahBVEVEyS
QjpCTC6KzIshs65W1gHrx0+vHcX6kHduwZF52AYfEgVlAS3PjbGfuI70T6kTs2x7GWT+Yi43/TBp
YejuOIVP4XxXs4UnupwpD0PLDmkbsOipRmMpMS+Kr5J7vPs+dt5ChkthKVHuLuSFnS84+6m+nTWW
VxJhFPOatdNsQFD/JN5RGyS+hyIhXabu+aVyPz3wC2WNvWFQ28Pb2pWOtyO/STV8gZSOX7NLOilQ
HcKYAlTBXhjg9oMal7bgwGYX29TdwLtWsAVXtzgEez3bxXTAUl6gVAMqraVO8XyOIbGCs5l4wQGn
VSd3Gx3GPKMSJhKKGr8DSXAmHczO3RH7xoChwrCoa+fRn4Pb29H2ATkSpM5tFYNH3WcT5u+Pox2z
yjoO7PsJsMUgKvs8XGnaCTsIt6TCX9o01N60gTqRwYOVEMUJRnodRsfrjVKd//8emUzxzDF8kAmf
BkKrm4TX1dFET5WphJTcpxMKdMiM7luxRA2B344yKMdzfJ6JJd7PZQTsmhor3mtFNG+0nGvlWful
Y2yvjM1IyDVvTjoI/coE95iF3wav2cmP3EYPj93V7DipfSgVWW4XuOJg4/m1fBZo6WYp2QvrRsZF
LzoWuK8RphCwf98vLzutOIjUQnp7/xZt/XRs2EB1qcdKde//lzDlO0ygV5XXS+M7vDojZudB5nmW
OEt/N+YvVhYot277EuYmS626EShJPb35MJe6iGq2QqwRSX4ENRY/6Lq8G5aG8JwdgG+zxxW8WIEg
j+RhYh0O1BY1mdPqseJceSpFQPJgNsdkE6Q6RNNv9tdfcSOXzIkM/Urafg3UZ66yAxjDE0VXJGyq
aEA1M4Xg6jKB/nyxLj8z9ucL7cHOUTgNPHhlfGP90US4pM7YB7iCOEvaMXGS6wGVJ2p+8wd0rCks
7psCzopb79QLVf2CArIHrxyOwp5TS8Ill3k28ePutqUc1xtwb9X0g6el79fQTrjz8Fes0WIMmbSp
dlGabsG5djD/AjFwh1WldIgzjnm0FtlQpD9DoYbvktL/XR17Dpk130mcx/nDmBhIDvF12igR89mP
1IOu9qu2aQA5ihS2zmzeSALH+kIc7zYgZNyGMLJL+yLWxQrLsAdecw+3GZDAnCK7hQym2VIBXWrs
Wg6qmgGE3TFGC4OeUHJ6+nfdD4MRP/i2S9bvezX+/fDXPbwCm7UricHax5xD2QnEBhfq35+TRmAl
hrnA+h5pqOQAfGFx+SVsh33XMjyyQx1CE92b/bQb3pLyUs1b0zG8tuVryeFCQykYDoK8cvZ6YHWo
ozD9tO7N7XLN7HcfFkTc/b3Tr5+n/v6KaztocgLhxdSgktt5AZ5UlRSpEbepL1tnyUiNTxPLQHrD
uzY89H3FXHn1A8mPZc0LHFlqI7s7s/IDvAwVmfriBlJTJnZjsN2x7biMDJPgLswUgl1FROCEVftM
QP1p5OWhyXQ9Jc9uDYnl9MMcvB2cbHo9KIjCbp6b6SuS5dWetexbVwcmQzePbbhunb5d7y7UkjJH
/T75B7pg3qHAsLAhGDiKvS/wW3DzuK0Y+cc/rW+q2FuouMGyezHpPbAT9ABozEixun7w0KMTf7n1
hIe9fDWaT5kiUOOECsdulWDVq9OGDbGC10vzNWkJG4LG/hY4mbbvOAc4s/GsEjgS5WusKklzWNlq
7MGLDKPvy8FDc5WUNE3BgPwJStfYfDR2nLin4imyhGkHI5ACDzzNAJf4M3cRhRQTODAn4TQC7JRM
g8IpNUZXPduYOnJ/eloAIc5NvgA/jWLc/RdyaTho68hECzHioNH4KxIRUg2aw98HHGuQWz+jPhm1
Sz1oayGLUG0vkHkk2GLbMdaKKxix/yGo9VEyK29xcQEm59/A7EIwh4PGL2wWBA6ZVq1LRqnvbndO
4DSs+2W8Ui2Y9gM/ks6H8y7AT7He/ebuneXOIibi1LwiQjZz4WNfBfY/gXSY2ilypulSdNoI29hx
nQ4kh1FTC63jLAId7mZIiUw8I3qsyIJHfoj5mA+PZUg/lMGLbXGfWS2mh6ZLnyHgSXcSXRlN3P45
cUyK/CM1Lf6Gu7eYAMKKJVTZGsOOnbaWZfWWKjsTJg5IH6EAOTzBmyt3R4vnilHjZzS2pQdf8DGQ
TfXrAuLBP6JePifDEiRmleLJAUs9muDQ3p1tAn4NTjq1RYkGkJ46c7BIehjWNUZNSZ09hFtdFJcm
lC9khTqu+UBVPWhzFdoTqiodX/Tth+oW+UuEwyd8rV9R/nwx56UruJlKRcjR1ctE1iSCakRJBf7o
h3cDCBbSFAQzJaTOI6NB/cN3DsgHHqhydY5QqyFd69dU2cyn8ldRAGFK54CKaq4DTAbJ07c7T0Sh
anQiYuf2kAHBl6VqZYC1gH5LebrdqpESBZwNCbROGM7f0bBW8UoJH2NrjS8w1Slb0wLYjvNevaMK
rS8TLiaqgb7iCg+q7GLwLuEdAVn7s++oNmTeAMvB4YKVX+LdshLXf4Wf+pluMP7Ad7kAKFHz6JVd
DoiDhaOt5tpLg3oDEFMLxuKWZeGD4MzZ9yKXc/Tio2iHlgZxZn0I6oqMsybttUtfTbR2PITwC5HR
Z+hM7juT2F67NR7HGZxWJx1HTqzL+DkqWwvOCJkeXJGRtToDnq3QHifP+UUbM+3e5dL0UR6GHQOq
3g3mpPKCFrAQSE4Mc9UUwD6X2DIJpSrmqmtH9Ir35gQR2RKajKfUOmE6mgtemkwKox70XOCZVeWI
fg3H1Np5pPH0hrGuNV0LEYU2WDfRSevCcsYx6saHR/yAVNZdufwa0CKLyKkql4kB9UoeiKnW+e6g
gNV08mfvDIGrcVzJ58lGagToD2LkHE3Tcdy3/1WqXmxiOMrjthuJG5Mifow1P371LkqPvSQqoCfM
UmFkcmNwJYamY6dp/cXmQnlfVW+FZdUFyKpyYxyMU9uvUsbga2lrLvic+Xz3/+R/K+azuZM4aCWc
WxYOva5evchuvwZQqF5rqTlT7cKE2gMH4TvUkU7mj0O97jnsCGvfYOqVmoTHwut6xkohkokURZW9
AwVGP6hLRT4fNm/JKiGy1lW6/JdZQoqfbJKujVBMoCD4HSaRPkU2tyStXMliTgTl+ztuy3HpVGMW
8ndprFiungIzpBDwD7+f6e8kDdpUvlCUAp7uUT+oa+/o8KNo6QviTw/kLPjiM4pf4VHnhgoKxY+h
YVOthxsAZi+g2ZerOkhNDvh6xem5niLyXSA1LtcG1poyNsBEhLW4uhJ+DglmOMukVluYKZh0iq75
YUc7m4kcI+zHBQs3MZkjuSLb2d+o34BjAQT9XOGUTWq/ZfY5HT4MWV6vGcBDFNlMzXbxQI43nbLu
1PmYRDqTEQtsuClmzhVLlI8T/D4tzYkB0PYgwrH5jSHXDYAjPsGH1TPTaDnCsR5gSy81ZEnkM6qn
69SCe0bNRl+sgVwQoJ/rslB4FRNlsmPHZYsJBs4bLqrJL1dZoCMXzjnAwFEKOGSz6pd28bEJRHYl
itNqU3+fhbxtncmea9Rlt4pGG8nFJwdnN2vV4zfMmw0pw3BeqoPMI2yWbwzCORGtTKaJYoSy0Cb9
jxyCT5zZ02PzI6p4j0xg6YsSIdMLiiS4d2HS4q4gCkvXMiCgHR1tjBTXNNPS9BVM9X0PUBsBHJSE
hm2iiR06ju8lhdazuVy3kaG/Aaom106BD0gW6tXxa0pycX9cRAMiesGqwg/6O0fqGeXuZvJ3x5vb
g1wcMChfJjWVe44/+1Wvo8pI8vW+9WmkSPSmu/S/GRuPqqYET0FVwTahRJin87TlQ+EZXQ19+HEo
HmbzuRlX2rzLg3pN5w50pWVhKWK4vTU4nwRt939wksVxGs3dFk7EivOOsTqtixXTe9G39wegTlmv
aLNOhCmXCIPfQazsQGBF2SahCz59lRAgIyPUZ9G1youl8qp64WkRCFsp204/40nrjGxnd0tyQ/DP
xYt/swguoCwI+QbnyyA6ZU0JgDHcM4xtLipoVjuAPD72SMKbedumNeWHjbi+76jEeU8c9O/OhYdY
YT7Jx197D7w59egpDf5YJi7D1J/m8EPHh/ftsou7lWBoFCx0m6hW2jDfFpYzEvJ/GfbpoO7MkJsC
JKJtiX05K4C9hqmFXDW5ltDfVkLQh6+y/u7IafyMyY3TZ97vmnkq/Jg4SnPEW+WpxgAlejZgYH4Z
1ST/OKhSBhaPfqvecN7JiiTrH6c+fATYpqLbjowwhk44HiBa3VK3hxI4Bo42NCH6YOroPQlzAGaK
F4EBTTakRk7hA23keh4fjgnd6DsbbfaggbxxbXD26Ae1mrGshI7uwIlEnEyd74euP/IVqWsPt4LE
B8Na33j3754W7ZLwdSZKxo7PTOb8xFvstkLLI2UaBZ9JPT671OnklhmsVQnMmsJ8cH8Jw4ypAj0i
cyvG7kZNCQVrNSAltKrq9Dc6gpzw5tLo93+oFzhBOcghDbf+cAeTeiDHZQoKk4KpSXZCQGi9kjfG
bm2JfJ7NSsoQHIyBf0zG9tp5Hdb6Nd9rpBzqofCvm4sSprg5d/udoWoBbZ+Eoc0loQRA/UQarFhR
BmbZpx81QKlrup1zuJXXZffiLpo87vliAvg1RfLX88mrayUrm8sUPQcFEw2VSDz/K6aivfnySpi9
o5DftFZLv12KT0g/c3N9kBG4R3vIn1h51uXU9jxXkS2DFnwtdsSvd6cJrtRbrHppFQUj0R77UIzn
CVTy6elfFZWOdgsqdbQ8Z9dai0SMXZo2hCqyEtrhd/OSVre6qpQMpqdVGqi6gXpRjICU4r4VfeCI
nmCBUz1VGbicusoxy5/p+3dtv3iDYAHQGzdWco5qhbhd7KhyufmpIlpoBZvZYj1U5+iPwpqhEoDa
NQaioWJyvKXVLiYo/2/TJsd8pdOkQqoIx5iqYZRfGnxUVXrGFxUvL9RUj94rpUsUOCBgQ7/Y9nuk
YndCLInhxmJm+1ERory2/qPnGlBbYKTR4OqXMCpZffXO+90xxlOz5fb5UxZC87nczFHhueFrU8mM
i+1dxbiwmKcGYj/2VhbVr+oQ8UZFHNBdiuZFL6va0e4Awl1b2za9FOvKHPS4wPL+PnDoe23Oq5Wf
MbLJaMCS10iGXYmDd9D2oKDdf0moZCx6KQyGfI/Dc02MObSZlveZ9qXn6Fz4DzN1VPuXqrQBTgLJ
A2xoav7FycpkQ0hlosHzJaEwDrYTFqyL/6HwIeUHBfZVHb4PYTNeMRDFuYdijPqwkPf+iDmUXCxa
mc6mTKtPTTXS1oJ1VJT7NoIO/jCI8q+mPJq6eZAG3n5SeIhzlShSJb898i2Niki/VhxYNonQOC2K
sq7nDag6LH5CxXQD57UpNvtKu6s3sq8X1IbQ9aAMCvlngMYGbyhKlbItFUDGwlyK0IIZEOFTSCoQ
Czliz07FlWOfI+wToY6lVpknq5PuvEZRx2H7W6LW+yMYCCnMNG41t26ZdhjbqMO1VRZxo4zWV/fG
8bodZ7Odpu40g6Mdx/Y0AC97FbZDg0iJVO85EmMp88ptiBsy2aMsjFMksuw6Ug2Crx42u/qehSPs
5yjX2gtDuQBnnt0HtisAZBbAeh3nqAUHpskszkTAEjhdYrZYEp/DqVa/nscl2mu0VYMmV/35PyHj
gwmuZabCgEF2T/2KNgeowyvtjuHgHS5BBi951MVS3vzp3Y9Fs6+rJRsEGMX2D/yJ3y7Z0JJhpshN
gUXrYXL4vsVpk+lNnH6r0bO6VHaHnM6evqmzahf0h3ZSxB/rUygCHRIBdAg+7Zwl0awbV84rUyqX
HcGvE/w+PTnSRz5kFOp9aiddTY0zvtQRI16ciZ8AQB0rJQzfWEPO+V7POHLth96dVZqxTnHk+iAF
7Nt0/nHDv48rpdyz8KR4cV3D6yhn5UHBas3Y/u922i3hpuVFm7v1CPabGhYE2AlENL0ZC63SJNx7
hh/2O4XB3ztLbKY5rVbf1OENsNH85kodVnkfvinwley8CWhuTIA2OPGB42kP69KtvAO2mjysfM/A
Ah1zPjRnVHTiOHURqZSxJhwzg+4palwP7Q2gM0Y0JIVjXfAU7B5CcUHOV/54p9Nc7vx/uKvyR/ki
2X8pJAJhdePVFQDHKfFjo8mKqBsde28g3PWNZDx5gCAoMg+CS2Sfa9kEjHXHCRYFJmKSrnuwN2xn
fuHTQ2L03+S/DIk+iKn7ShLgu56ZYbI9OpxzLNG73oz3BL3lKVt9t97w7ru21ElyJIFZ/s4GsOMb
1AhASepbqeaET11s7ooe9UYLfx18jKzDkQ82GpFqCPxpkJyesVbevfJHcNXWfq/gKIqOqbUDQqjK
i2A8wfznSSLeUF/2G2Aln/0Ww63XpB7KN9yg41Yg0CpNP3xPgMohRPk/oEWt2V2s7F0R+9nkqg48
Pl6geXxBaisUYK//xjA2bviKUef1uP4LuSi94CHkNOr0Ato961Ck9rphooNbgAQHMsytP5PqQ9Px
72cWH2S8mU9Ea34Nfh/TUdud/PZMFpXQ4IF9TogDAV/mjuJF9tp+GSlDRXjwmeMgY9s86S7Hpzs1
IiAHWcK/BjxAXJPedyDZ5mw9RM2i5Sbb+BZD7PcL7xI68lQEGnZzMbvk6piyTOD9cyPRpgCxAvQA
1aUE4auFL+AZLCVGcVRmZVmw6AWZCxptTpZYOQVPGdPBq2bi84CvO1YLkN21kK502izW2BqJj7Zd
GWUHkzrN9VU8ufJIHF4pNg64b+WQlGMbPQZL6+Ns1Zm5Gne5xN8N8V7GUKDhGSw3x9FShCzRoQiJ
NNd6TbqWJzqCVuuQRDK46vcxXCY6OX/flb+W0QyeVan5JvN724Tg0yiOz/A66uTlKlUCumHQ5PMu
CvklpRLdb4bSDjLlR5+KBc7SXuJptBNUxTeX+Wx0WhY7m9BYf51bcmJpWgiiAUIwHpSXNl1oebNe
lge2/Fs/0Ggd/m4n0GyMIqWi21OIuQnYy/DRBMTr42Ds4o1AOe6t/HqPyVzo7tK9FoVAhCtjBOpu
Tx1+ctMQn1JsePZiT0IDG5/SlkD86wa27u4b6CKksYKNZpmVAgWM2PbLa7iTLrLAuq4U6Z/iF8ON
EFi5nms9X8S0h5uxEOVlM9Vb7So5e3SHxnouCX89fp+9ZGyARZHjbNgYJ0IBWXqY8BlPl6vw+Q4a
daI49y/qC+QTEfPc8BWEFyB0TOIS+F6DvnTJsSu7czLvwEmyzIy0OEHANkz5H1/a+gvXrym5kHBU
dldoZxIKrmNkI8EMJDoBmdqJFaSSMcJ258jFedm6QdUWThy3yNqA5/sZwtjtkCKCppQ/00sKLtDw
uOrbSVFcxdmqj+3JzxTv+t5RntxJ6QZlYg10U+sJZPPRGh/5l8+lkOQrofnQ84w/5M+USzvCm7aY
rSQfkguO4btfWxejquRqWqqHPYJ/6XkGtpc3SV+q48nNbe4P902qWQfP+yOZBr8WQQR1UMFnafNT
evIUJ57EO59o2ne/IR3DAzLrm0gUHEbeeCwNBrJ7sWbx3YF8QpEc+DJeqJMcFnfxTcGrKmnGyZsE
fglq0cpwPGEGo8FZWCqjB8pI+kPbRpkRwGXoQrzcuOyiQnD6N+rzccYeD1H/DJ9WmeaAZDYyoQ4S
R9KnauaewLPfIyfkSGPKHgxrLYWistgF8pT+QkZqnPx/umtywMsFlFjyQu5WXTiKQcF11ZPQJyM/
n+727crttx2XKUiuJYMzYaCWbLsmbDDnHVqSnBQl8w50YoNkl6Vj8O3+OsyoYJhCdXh0pery/D43
MaxIw9izIDJAMmtX2nLLhCzN7ngLDz2C2/UkZ0Udv4OnM0ArVx+JyZlAgLvXFR5s9JR03nxC75XI
RQNL4C8LI2TxrR5yE0RM8Rz0R90b7+LBkU9f6xxO7/8GZTZGYZ/f+igkyZOC/6CMJg1WSKeOIToR
a4zt5pjI96vSV3sbEODUh+Ea/XtDvDuzWPRUOoCgCLXK9f8RyJhR0i57K6sI9XoTxZHjvFAsOeJ8
dwu+/i7zNaTdGyATccZTvAjQLzFaSsUFyUaE8a8uHZ4M
`protect end_protected
