`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Uqfmhhe32U+grK02JBnFtloD9R75vrZwSRuZPqR1VnqBr7XmHZ9tkHJS1sJOLfG8Zd+796XYlEPr
esn8WdZgAg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SQ2JFvkiP/6Sc73sJ0iKdnS6VCowgR1u3Z45BvJSh4oM6G9yLO60+MTHZ6334rXMreWy0IuTJVfx
YsKGLRIp1v29jn1JqL5X4+K/1XG0/oDdQD8qut3QXA/Sr4fQEfjJUYYMqnTvQt0dKUWt9V0hhst/
25yj0qy5VOBC8jSzi6s=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WJ/I+yHH8FvqqFy1co+ttqZkj2uaQDeZQb5hC+1bA3SuWwRCgvFumZLJdKX2yfrxkBeND8BSdhek
yG43nJnIKHgmtCpSTXIqDmD/8cG7eahI2BTK48q7plbNzSW3CZdXSn4RL3CL2JQCZKc+m/is7KXO
DSgsBSMWyLrYMnpfcolh2Lm4vV9btRLcaBz+68qYXExE1DCa6DpgDDy4qv0YETqlkq93dQ0ha/Rt
H8A3DG32kmMl7yK6s9PMAc3GlAp7xwDBU0GPyJOd19glVdCAAIBSPFIBIQ2HHLdJSYL1Xp7anroL
tgXNTs8HJ8Zv9Uh6cWotDFfPYSYyjwyUnbn+hA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p63c4l9Cue9D6FDOAkQMAJUj+Hg/3ruXtR6nWx6J6ktFuaeu2QHd/dww6hkLZbBhIyG0LXCXtPD8
y15+0t2dgRkquT+Kn7umI+RIxYI0YGMDxmxNW2oeJQyHBYUIcGC3Imia84h8pjT/V7z56Kr5XfgL
xs5UhHtArBz0OhWEXuc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KUDZm+F3LxExF2Qe9dGMQ9l+lzR7Z9eJz2jl5fXRWxdXkwrIZi+J51Qb9ZqMTVb0RUwoV1+zCLYs
XMnqhBhAPnrzL0y+uggoz92NQ2tDaAWGNPBYI+Zh6/HWnieo7Pi5qDrVLLqFq2b3vNyr5775+Kop
x/zQq7CngRYoihhAXk5plZioD3eP/bJQRN37016KTYtXod+OZUGLS99HPEEyQITYf0pvagARKeEs
kVnvueeuq2ktx6eWYJFRI/hTLJV8QXZZoPUMdS/Zxc8Fi/9yTVI86xCXA+ESM4U3OBGxLhJQLoWl
vjV+YjEDbxzMzWDuHdg7cXYygWrc6k76gB+Slg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
v0jjqkX5YBHW1GSd4SbkWQ75fs1avkUdjZMYzmET2csXr7wGkNxlY/CAvt0ToFua6xyeTlywtDI0
F8p5j3umE2mwUDDCONVj3Aeuv6FWn8r/IOnMMeRWfmadS9Rm/Sh3R4OEHAE7U57WwgiHIKPK4cvX
BpZdESmiW05dh1IBrBYs3/Qsm3n4sVT7ie8qFDk5cxNK8o/DUzsuiyqJehFyt38RW8389MHQ/XCz
uq/8uEm0jA1tq4czQ18sWdjsNpEqf2SqsuKqHYKcBKFhTMGKUYnefg5U1+CK3wYpyrhg5wUsaD96
iUFx1wQXEl84ik3qRzq6hv/TSgziiiyWZ19vA4vAB+YQgQkUDcny0txE2c8106EOeyJ+Z0h7mHoa
9XKL2mqYVUs5iJ6V3GGOL8PCaCpa1DIeuTH0JnXrn4XuefgI14jhqn4NZfSrV4YlqymfPvAXpuw3
QuAwWd+a7XUGTUzlLsIz4Tvj3T1WfGe6VJYYROPN3WCwYfwjniEU1gEcU5MpesQGLXE0fBue8ylE
t7JkUHJedskRxH/St8X1oI/ZBC+DT7ADw0GwZHaHCe442kKbaJNZpLtziwqAFz5Fefqu3hBHI7Wz
87Xrd2cvgbHCNKx0PASmNO9mAIqYnDP7QVqB5DO5hH2JjYaxUHclkqPXRXoEygnN7oxzvNa2/ng7
GBpquLb267I2ixn4JWa1i8Vih2MTHL+Wk+8H5/1OhAnNS2+fb/ysVQg0mEDdoKTMEkUD6xq5K7Ji
NZZ3H7bd6wzXUXduzMZNlnx6B9AIOGXl8ph32Gzjbs6nhhjxBU0b+JlSvYKj1WzieOjxr0iufPTp
40E3qWeaLpKdS7rA83IRg/qZM8b27zbCVmLZXNNk32uI4Ptq7xyxaLCkZFUxOhz/EmPJFRwXUQRT
LRpZ9XyebGE9jB0CFVEwDsrlSW8D2FMrUxLUUmdMhDZzrnpQBTU9xXPQFy+h38cZqAC61GupCKaa
MjUh+JlYuVSOgdPieHuparWbVLbGgeQK722szQUTZ8rg5wKABwn0UTX4HilsVf+ySvw8wTIhfRwG
+0XFUhAtJky5m+HGevma9DBipvAQ/mlGsrTctkUC1OpMZX5/4Ws1nWyYiwsRUeLHnOtemZT3Fdbw
DOzRJIio2wWDQd96ELO82p/t8mjzBMYTT2nE8ZCqqCDm/6yl1G55DYclUZsafGRUqFkqiIOWYD7r
zWolrEhAUVcPrpe5I+ZUD8ullGpoI1mhOqxRPECrOasCCl81dhLu7KJbEEpMIPJ6kGaH2MFg4SZ/
V95+XdEKvCzKLvpuoqwM2Xd8LDTl8yAwHZBodRB7wHl2ivSntGDG7IrdbU07K0faFKEuHUq/UOMt
mb3ws2ps/bnMH4EWSOloUqiGtzl4cP89/5DsOLnT859LBERkywyVBjIIBmxIpV8MBKCTJKpQCbuo
th3K7zMZ7NEcM3iatxsx0yrYGsCjiDRzFtscWqw/V+6VEy+YMjXO+eeFuCEug/kaPRlvzmSp3G7K
EQ/MZiU6nrmP8POzhF5icPhUeSn/z9GtEj/Jaqw4s0yx5KHHJZnAg4lC4LoTpvu+L+P4nYlD23oy
Ylb46sgwdOFO5jsXKmFP+zaSKmMSNg2ztz0z12+R056qryP0LLeMubDj29+Kaqy/wAhfuPr1mUGu
QapJ62DMxS6ofMYIEEBOl5oUh2rp2cih3XLY3yXoQ+84Y6e9mjPZVwO/ChIgHDOdsWIwy9h6FwX1
se7zLsIRvi0wZKs1u4CnMwXj/fBTk2dM55NlHmZJ0uit434cOTHmC4o0i5aJ3HzzNUcnZX184i6R
Bx9PThOxzsURZMwrD44WWD2teEJIJ6XK73ny3lRM6RxU5/vjOa4AXaVp+a69VDjcry3NGGRTofO/
VXnw4F4L8fcvBHJ0Wnu5f2kEbmM3N7B0oH2+CTl9OoqEzs0ahfu6xGFkpsDMg8m91LTN9LS1gFPh
pUr/Lqq5rR0nOPXCzZkGWdAZEPM1ltM183BaorMMYhsa6vB+/DMUxjTFcB1ExsvP6YrP5DmqqF9L
VKES2ui5SzOWa4pfaLDHgBkuEW6mwTYDNqaev/+SzN107jKE2AZCNezq+Ol4jbVCWtN47t1fCEXs
+riHZ6I0uqAPOR0GYQ+WSBhfu+BP64lWHDByjaLyeHTt+2q2wHm2dxInOUtmR6cGyzEZR/IjGPox
forFsj7Z86ePnMziDfFDLvCLPooYUOapI9W9O9r4gltX/JXWU+f4cqIOBsCQDjqHx/NdksPIocMd
iunQy2mKZzb4nCEXAcP7fZvAIIuE34IOWty9xYyxvzmUJ52BUWo0JTrdwYXFfcA7ik3w9GTn91vo
QB1WXVmZEge2sklcFm4Ncym0O6j9jQWufjujJUGCeEcVzpi2aeq/BzXuySgc8b+vcyXli0mEm/x/
WtERMzY1S38TMn1j6E2IbR2bIguKIQu9xc3APp8AKpQtt7hoyqCw2cpFS+DdR+g0MRdiaFjbIur3
3YqwTHvtoAkz0ftwvtFqjX3ydO4hsgW8TmhjazxYbYB2jj2ehRbL9ZwWGWfSFZ/iMGL2lpysZGdm
5CSXVOgwXsCqZKS6VK5m4O85XZI0zx4NW0F2Tg53XIX/xF0O4uSzha/U8V9oJhq4jEv4qxs/KZcO
MxafCE8A9NaPzX8MKnT12iQIopjMX805JKCk/0ZyYqUih0B6fVSikLGnt7AkDAdsUMhL5+HjJDyg
09wcj0wnM/zBTMlbXMx0UFa4Zq06c2nMkpedL2GEbMGmRb1/G+EZIZTgc12nVr3cHBXYA9NUanLy
3oyOHvhO8ckKTrmH9RblZIZkrc5G98droz6EgI1W7Hy3kZKETTGPwfqAibNpEZyTkMdxl4fTpXaa
r50s0aIOO8evLlJ5IgXvct8RHe6qHfHEJzB0CxKwUWd0wIQM+ZyWwrT9zz7Zb+1PDCj61msnRsZl
iXW0mTaCo3S7jhmL+7DYLpIir4ZtUiWvgIqcLfCf2mpppeyakKwpFpaKGHX9DCiBtlVBvkmfXMVG
YcQcRPt5/6lfN7qzPlgW1bH6DaEUwADR6CY4CoDAZRjHaze4fLI4vmTYIfjsBbp7+7WWHhGFGeHh
QplV3e/hmRdUUyNyMSLCEc2+hP00aBgxGOD/tY7YJ8L+MVBxDSbbxhmKhQm9dEwWC+xy3Mudp00U
QCMJiQzgtN8b94wV3RVWzYY9RBmMaFTLp4evr92JRq6sTUFQOjyTfjJi/InGqrDJQTfF198I2YNe
SXgYczkgebsAzjTnKO+tJinUYt++nS+D+2i9KONrKv00/S/qeKuLjqbISB2RyxmgK501mO8rggqT
15aX+wuC1aOoUYN0kmh4N7oInbLI3iZTBezFR2ojy4A/Y6PJi0YrZtGWtvwoG+B3Yg1roT5Pbleo
bgrpFT3/vycTemdsG/SDkc6Ojr/YMkoN8Psgx9SLlvG+WWzSwrBfYkFwltFHRdKGngidP55QAtnW
K7p+tlwc6Vmvmosmf0ngme27CMTozu7ue1AEO+woGCo7YUfhuonVL3AMgc2OnyvuOIlZf4/QfWqr
9PX81MLrWGJA1YMpjT2PsOorbXLPPo7PLtnwYOt4jn7RwJjbWPfyY7+Ln0Xuh2vSpOiUrd15t/WS
M9NW2ziKyFrECRLa6Qie3IfQXj9QpvRzbJ064AAuFNyrQCl04k0zQcunVeQaXGar71s/Zxw5RVnL
FM+1VMnrdSRDyqRV7K3rZakudbkpMIzL/rS9yQkcK8ISIDO7fFuID0J9fgvqliORZ7jq8kM23Qph
wEfg+pyA5qqkf7DSR7wqx+b+Gnq84uywN4YG1iB3jN/Who7HYZqRW4K7+5k6thmMThUVR0blOyhs
zPSZY7/o2UC5s312JfUt6TW3Pn04NNQTIpQCpoWq3+kuOjuS5ct2UMvrvI3Ze6fIroUo7RZNGJrc
pKhZykA2XCv6A6qlfvkKCwN+I1p+tQdm1toOV6ksfVe29UBrWUshVsSpl3du0c8j1onB/XDYgNgh
ovYnrSZRBatNljj2pQHjMxqEOz8EsS4a2xKSe3bQfqvGOKxqnssk+vcWcZLkuSWel1bphs82MwpH
uRYiJ4Y/64XPHwDp2UpR0VIIGlRdEljuTdg5IU5CjAMJ4kCFbEQ83Kl6xxyxpmK0vMQuGEz6LFaP
GfJFd8fRJHyG7j1wzT4b6oMeffKOUGCfwh7PehyTaasPL9KM9RoCDERr5pfKr4+GNW5vcfMXKC4H
qqBVDU48iMJ/XbdNJAHVaDVrFlUv/bk50Ec0wJ1sf/2ITb5Vqm+Rej0+SMkTDJsooh0AlNCY9e+6
8DSuQxUyQ81DbtvqREp6AnFJxBW651zShsDphaHQhWu24I1iKoDYVJ501uz+vbWNxo9CIl24kPk/
KbrAsKkir1AJvuGegZ6rkTS9Ey/CXM6C5o7x5RkrQfKOoMdWQl6tSfIk94sFacE3GGE2V5MinzAf
xQLwzAnD7CJEWlNC+THQF1jJYkMdzl4hpZWSnFf+rqCtJhMsghTvgCBDxIFYQO8OzWtt9G7/kBQ7
QpCkbRsEkz/+oKRZjLf+I79PFckws4XOSARtv8ZxWc3ssis2uI3Wyucg6epjVeCGU46eJcBrVMKa
oSO0m/TQyTyK11vvA6L0CPS6H9vcJCrwCQOIPExG1Cp3GbgHGppE8LZPk2hANCZmjCJLrU59/4lO
66MASBfoa+bqHT8KZC/Rr+S0CGU6w75e5KWbEjHRXjOVYU3ZIu9NM+6q5gb7zHt3sP+XmBJYVgBt
Aqc+8sVX+0KQheLVSQyB+uHrUYlGMGwXWtr7Ukr3Hc92Xalrg3DJPfsCat/KM+09+VYxnzwuDlZJ
ga10moUiJZCxgfMY0RhR9Wwinget2feUWk1MSODMFbY59mTL2xBb4b0WQFWIByHd/HlBIRKhg9Zl
2CaOEt+Kr1wsk4c/YhkgKZQwzvndvqNQixBhnSb/o3De+f6MxOH5ZnZqcyRd3NcrNa1Zsdd7rhpB
x/nuTL+aPpzcxVIke9WMoqFhMgTnNbrSip+tRAjMK5j01XtQdEQtBBW7xLJ0Qb0qTPpUKZSae2yZ
kIaLZIzx6KRV+CQlgyqbBZFvtglgFgBx4uoS983zdApYN/3y3eV4IuLo/ASrSl3bVfpuX8fNAN0c
D+/IttJhXT5cGoObuzH/lme+1U0AUbC8vu5fhkih6H0xrFrG3DXPa9Rw+xvzt00zDde5dAabRHOF
c7/iBgeTNhQ9aj4dsSzAvqqyZZC5/W+mUYCgpaAishpUzRtkfLXO8Zj8zad4oNUNU4ALGbzZpUaL
5LMoXCcknvRYFQOuxs5X/2+tzNe9RopDClURf5c441dy/elVyapyj0n5TpGJ++Pyl+WQN8jHoDZI
tceXcBXAyRIabjnpqnAbSgOxs/pmLVxkTgf9EmlINEAJUHzXIS1s7FpPc/LP3mFgqn17RYCE2aZ4
mdUM4iBPgh85vjEKhUfWxEm6LJ55SlgmnW7RXPdX3eWUObVbzkR4g80OU2Sg3DF+xYrXTFvOvN0P
HDUbJICtN3U5k6raJNVhM8s0588W0MjlbAW/KyDWnC1L+OgigrTOEMKA8K20ZugpfBX7bB3F8Zkl
hqr/BWLoeuy6PiZbi5l2IGiYWfEs3R1QrGakB6+/nOzGzIMhBDuIzoRaq6S10B1bzziRi+ApFdo6
wflOGFoGRhalvRTAYUDThiZWnWwbAb0H9KKVsF9aU2yQzuCbQuyrNgQnFFHpLgHSh01KPTvx3tr0
XJrX8X1dNHfpMFv8blY08FOj+AKsWrMkBywmyCGgKpKsDK/66gpxgfvOvzkxu7+kMkO0MouRRYlE
lJw+i20UvjGqTk/tUIcTuI8cNgAy5nsWAztbGV46vRwx82L/tb3jG0jCyGXAAwxl9XJq1vtPzlMg
kaT+y7foB+kHcj+l644ex+jIEOfJtXtzrml4Mmd7B+l5lEHn4W/ILuS1+2nsk9O4zxeItXBPeJGn
7cXwby0T/ZFbZl7oAugeam3LRzP8N9KwmmEMkVsux2vSAj6glRRMfuL7tefUoryHfRC4ph34IFm/
yvdmMUt6kBoSdt8JvziIbc8AktqhnhuSaIyowL2bp3Ebnur9EDbpdTlnCV28uLPFyVTkS8MTiaJk
N/Q6bT2Nsx4PdrIULKaDOimoLiccpdBmrLbioWhYhyB0A0prIGd24k6L02ItmezTMIu/OkSpiSiQ
28Dkkr5kxHFQ7WEOLLi3GK2J2oh18hJ7LGwE5HpljVTFvPHI+APqxla/YhHSsyLwO+FvYlxWyjWU
IaWeatFGN1+v59DsXlCAp49xV68cDmSkWNmYbvmrokB8dxCZKONiIV0Ia2oq8oWca6cCNKJpGTK6
rQgDY1LxF9GvQihJ96dBjIBI9V7Iv8XABJCvrpPU4h1a5PRyJYWpfrNRPm14eJGfZ2mPEbYEl1kr
ozi0TCd1Ko6XPh7z2McPykTARK5/Zr0PV/UcuNoGcjw4TOBxnBKKlk3XHCStHtCjBHVjAWuAHaR4
qngI3LucbdAvn3x/nDWAvE9/iClYg9s9m9FXlHnD6HIFPmTbXQnrCRpFJTvHDJHok26ChfKde/8P
MPupIE2BNq6IWXn10VTK2wS5TNhbhVwZ+jUbfHMxUc7lk1589ij8pcvjZTBxFqA+63dXcZs78Hpj
7yhJxYTCSbizZ8pdox/TRhp3o/yfhnCHizmq8f/qT8HXikg+vkSy8Mj6qAzcMAKRQOgvYgp0EsZl
HbDoD6T/qYTEXVVKTJrRxfViGNteVLAKYD8l6QKu+m1r8DaHKrTKH1zJRF1+br+cLE2Kgp4uPBXD
RbVpjCkyUHymdjuQsmxFVzgUAZdeYCBYWTHl8s9c0zvSI14GUbuZQd1vip2E5FNVh2hDxt1oBr00
qJiRCMIa3JBuGvTpDmaX9J1LRKriyXabFBY/rjLuap4igYv6FVGBA2qkTeaWHAqly7810G78HKAF
BHNGgqa3xHaW6ZMxKqjNm3UBIwnOOjMJxF9YYIWdbjvU8ZKhB4BIU7BYOkcjdT8UokOSVO1jG2IA
y8zT+TN7yToZ5J034wYB3DLQZX4FVfFlNszAT73l1iC2y0rd+XXJrlgiWgnrCz059XZsiKgBrJyv
RHzYvCn9COKFBaupsO4y4iXU2x4+yDJRyb/5TqlMNHfqYLcsqba4TckGihwZs+VeQnXFvyjLBJsu
Nj+WUjYKFkXa5pmIF5iwaSpoIM8ipfAEBws0LyWk2lzNK/QR/vVXkGlI2IA1khxK/HG+Qon+buBZ
nFyvTNYwArz17HpjrYeVHzjBMLauT7OrkqtrbJ3LPQLSZCbTe9niUiH2ylsF0AR4lzGcqbaYkQfu
ewTd8KEsC8TEnnTRj/An61TPfFLHMidAnkN++C5VVmBjNZH7+gd5cQC9vlzQhgQ4sSWwiioGsLrK
b8KSmIGINJLBn850qFzEDKvD8e7Ngqxd1MsLLXZi+mHNCf8SPbsMD8w7EjMcjj0F3Lh2tj3oxAPC
CLJoVdsmyUTTjpvTIHUPpxLU9BDsaU7kXV7pCyqyMDvNg5Pcj5MwsCmyf81A1TGU6Mc9pMymdoVj
Bu/zqgDE+R/fcdg7NDFg72xKMIWEPjWsEHg14lZJlpVdamsRsLfcTNG3qmnb4T5xsjoIYNSC811i
I9/4298hGxaV6HI8e9Re1k+cjmFCLoHQk0EmWss8ijyorDGCVoAWVmF73ojq9GST7pMlz8P5K8T6
QX5gT2xL4ySiGkeK55IdE36lTmocT5TDu39w0jr5hPWe4EBo+tQ+OjSKInCMv8gXxUi/hk4zrbip
ayS0+Fj3nmv/CIKDjDwYLzia5msXAHrtg6UksG4vyJrnurh/GoqHSHd9/fzZIZCi72n3U14nL4EE
LB7jOge048gslmsP7KWqXvPpR1kqKKC0y7xwn5fiGYNWa7fVtLypzpb1BqjvO5zC6IherFatQ6Jr
gPMs8MTeLeTObkvSqg22DlCNSJOJfmwmL417v11hbbdn16MQUMozjJgBpks0J8EpB1IUVhOi1MFg
frZhxx/xmiMyfGe1L6CoPF+3Ka3XJHoUv5dGVWk/cMun60Ip+mPukF3gW9FfK84phu4azRWo5EDY
SfJWvgZ7v9W3HzZjZ1RX4O88bItGuvRGETKL1rT6Y3rjtqePKgedpbezSFdftIBl0OCZ2o/gm6wE
dcNvAWoGASL0c3Vq2UvrWDeMnVXa+XXQ21e13nXuf7MPvZ9kGhBb52IMY2JbpE1/IEbXC02O4ijJ
zlQIdxO46w6LO1Hi8a8CRVow6xE8hUOwkerJXc5eZfWs9NqAdluMr/dUu0PO7Mhsc23+8h7IQCWw
lQ1GXsauQXSJgbJVSlRy9uWCZpzsH0yb7r+vMZelgkIZ1jEkOkRkNj967rhMFD8yrgGjP1NmcvbM
6kAH9wG5rYHPkIWWy47Q7UmxWTNXubMU8kntTpl6a/juZYO6PLoTztgLLa+R5K490GqeI/EpBszH
saY1+3qYnn/j7vapOwdMZKgk4X78NRaCIqAZoZWS/Ruq9JdkItaUCZTO6oMGrWreKfy+gugKNn91
CS6qeO0soXim6nKgtUHECsjsjjOjtBpn30CW9rLBsJfz4YtW5BKpuT5OZZ1sMBOccDQcag1Er6XR
UjShiTZRKponwgVO46yoldd0ZumB1aO9YwvQ6t3piEPSwX7M4dWGMrVlnt+38bBI2XadbUuDNXQX
YsAYg1o1jJwNJdcZidw2J4DgWdYugQcFmmQ/AzP3q75yVuwO0uEC4oyRIvBHYHtKa5zDobZpVggb
IeDSfea+LYAKYw0u8k9fGUX7P3YUwe7fpZnpzz9xc8DKWT6gnnMFY61G7Aus0/jMz5VlgUDNtG4y
KHjbaFBMwg1ybUmdBJUm9eDKuoW4vslRsx3Ofr2po10RyP93rLXPZMnm6+UJs9kGTNk5TnjPrkJw
mXRsGj8tKMIjVolbRege/W6Vu//zgSD58rsw23W9cA3WlY18CIomY1RZTLgiGXWWrOl2PB3Csm7v
ie5PGph533jgUR34PEmmsiJQjtnJ61VfYt8VN/kQ3IzOUn40YOxD/tbVu4C1QS+bjuk1L3i78kJy
659I7MsA2QM6AY+Vd0B4UB9gdWxdtS614PMQN8qwC1+l1by3kcDYFtbZoPGtOmLVjQH7sjEOD3MI
9R5cUovdH9eVJnQEspljsT273GIjGFAWG2BLBl3N8YGxP0S2b8Gcsz1UZHU2klbW12Dc4qkSHESu
GnhasQ2UVoUbdwsHBd0I31Br23exRiNc9GnBoE2G8FHoeiXjqCxRJtWg/tFK2VZbLGVMvK5H8p1+
HqI02+vkUatZW3K2QsE2GOtAy6cbrIWRiyFuaNlMk++H0xxKQ1i21n+jvoZZc2Uk+ZSCV+ppH1j/
+GzZ+39A7Wtcj5H3TTTeX86uNhCLgJK5FtaAkEkwNP983oJQuH09enJZqldp1G5dOl5ygxLtjLV5
FRTRPZNpfErJbXptNlBHbSM9rJvLuhHNRtIk8zAGfzm4r/pA/+twKmwUOmTrtVFjZjtDYqexwIpC
TMJM9s9k/Rap5m+cNKE4TjzWTcJawS7a6RFd8yfsbyWTeQXU43cxwASOz3+W7Q221ltQrotQFXOs
pjrma3h25xZRGK/NnIGvC9JhhzVleGvhwPQSJ9Ic5Oy91QiYkKgolaBBF7nUClRAD+/b1Ak5prg2
78rsN+uOKRXxyjDG7c9FbXpLFbWxPL11BVmkZHbnk5ZxwfrgH+Lq8K9aqtbQ//o6RtKJ5Xoe7xGr
+IxEJHSLy/QwnRYf9o89z+oXjIAxSb8khWqTvmjaARl28u1YtvaDFaQcQM0Szf76QOavILGunWFP
cG5zhUCYzCJxnlJI/flLPl3Yh6WCmRTIAKLK5JOA7CfQ2HIBIn2a4iZ4veyU/nexGaI36fqtKVt/
YA1szf34JyuuTo0MBhd6iuXzipzs44AaZfV+9GZDS/+S64Zau8PXaKjKN8BJq09/fB8rqU/y2Mz9
jDkrnT1LlcvFFFT3cWfT+zzurCceVapqqzoPVnfvN9/CKZvYM4xNrTTSBq4C2Cbsu6eet1VNI1LV
Ou+b1ZAFXiGUPMuzl+hqFkCvuWsIoRRtbUUO6wRvP3H3DxFW+zRX0L3fuHdGvbIJofeKhKQuYvCH
QpWCAJIoulk1TA91A9tI2ZmM+f5xpqw40CC/sdbVKh6apR/5fLmTVZn1OflATz6UtELJF9NN6+jh
H76klqLStwTGyZRckvpEup+8Mm+hCofQPfzE8JjxdLoNY9FsZC1Nt9McJRPUweu4ODpIWn/w1wVj
vkrVKkJLbQsAI6qXpEZDdh/FScwl84XEu2RFm+WCHm2MjumUEwctCYAbdOqogITlJbGX/HJRrQJ5
SaZQ5pbkKVHmw8lxJrNy9+1ytUGXb/k1wAqHF/ZfrSbSXh2hmDjrY+BJ5W02Vehh/0otHuIv2jD1
bTJ+VCRu7+lDnmf6LKcPnpY/hvd2Wny520nCAvgKdwQ8smtM7yfTSbQ3UFiqlaD/zILAXAQYBxZl
Ll1dnlrA7lvTCz4bvNSvi/7CMeEWUHf90ZS8JBS6Sn2oMKakjDijosfOI30G8OpP9F5KKA1wAM0O
2UX2g29TaP+vcrsMUbgEBFWawsVP+d+rAXLEqMJIqlZLB+uwOWNHD0j3ZggdMiL9wTltRhcHzaIB
qEJ072sg8yjYeQAaebRJ9PPj6XDJW3mkucpA633JaV557ucMihEZHnSbF+LnxuwZrlo5WllbfGgr
WS16u4Mb52vJwzxXvqVRgLJ58qt7hmBzW0xc9kxTFOrT+TDiiNYTNXJEzmLI0nPgvAnVbLs68I95
s71didG61G2iNHvtmTthzXY3ej+mXM6U3631c06pfpPAoORKuu3Nqx9ddQvO/6Gczo/WburBNGP5
zgMPtQFaqvnov8LYbfLzjyh8JJ0g/ZelgYxM+S5B8NhxSk0eJc+RZ1jI6n5ihW3nf+fQ9/hgQ94y
9456Wbh1/qnCCj2drvjvNz/mN5fBvzuB4M1f/3b4+8SFEzgBiGLd6LP+rrezO7Wl/TfV37gCdwTY
7JNNuzfZKU/aZ7Nfjp7exUcuIAgautOpWxy6qgtJzVtdYIQ3lLWPe0YQnEvbAPEtGW/Rkc8eWmbX
s/R/mt7BFNb/PGUjq2c6C9jDuhrvFeKa6Amd/Xf4clYp6a7NT/W8HSBGBCtRmdAmi6IPdWm8cIjz
SNAFi1V5klt/AdkeTmjet7C2VUJb/Y+eP0rclLVgdBPLduiP6Egcu7PN5+yu6NNr+/0HgPE19TCm
6NW1HnLad3cR9w98djdN7/4nEzewssFlQ15iBGMQDKD83+I4Cntb0gMvmstA/Ov3/iXf4cOI/FtN
n4D+lfyZXUp0kd+kHAR53eM82yXKZ4Y3K7UOTvepHO+54YzAaFJJ56u3+yE8cD1cVMHpnHogdkiX
Z2ZrS1ttmlrZTEi1AWN+Exa3R4S1ti9nxllG0dEWB733dZnCcAp6r6ldDJwv41e0NE2WKjOKWBiY
zWT7ntZNnJZPpOCqyfs06hDgRqCUDjwZvd+R4c0sXPDqSsqDBjV+22rKit/pmiEYaiC2adZQjdOr
qBv1FYABwmA5L3hbXLyHpoqnVIR6LqJpvepzlzoSjgdLM+wWBU+RcK2lBVPKwVYISyIwPmlvpwe7
2YywefzEjybe5HI37S/slQj/acuMWz7nHoeRx15WemmX7t3wWj9bcIR9WLCSnNA0zhM2DCJHLKIM
ZXedJyynaDz2E+w0uwqVmgTiyqwrBzPz33csqbBv+0CconbR7mszPh1sHFPaoKPxLtyaIux+pznB
PRg7OMuX/bBlhlplPIXabGUnWNFs4QQ1IuiGSRR3ULHtpEl3Wu0S9gpQDuDEU0cZ5bf0E6zuU6Ud
uStHDz4IIQiepaIV/kPfqlFJ1j00pc+/kEVOMxXazRKCMp8kOwbcMGlFig4opoYtdqD3t206dxb6
+BAJkunK4n99HQvWFr6OjXn1QfJnpb6yAfS3wVfW0DvrRDtnOsEQy9TZhQ11bulEWabl87u0KlsP
h0n6p87Fzi1HGhSTQ73J1dXDhWyyD1nKSarXecPKRzUfSWHq5pUz/nqJxfgZHudXo8mgb8jlarZo
cV2BNT5uFreguCMpSaMjdaxdld/UZ7tSCi1PyIAG1Cvh4Tv7c//+azi69BIb2gl/AjTht1lC5hXQ
QjQh4r+C0Hy3k544tbA+IOAXagXOxhYzwyw0Hduq28beWwK5z+w/PPJ0ATNjjsVoafHZhWMjghmO
F94kBDWdpJ4j+RtPQfMJPlLiNVqPjzi6VQ2l6iN8QwLY6MAIhk9wi4su2V4C5hqwBvO2SpggvqQ6
efjol97NLW+25UKeOfV65vFFNWVak1CoUGe6Bxl6kDiVEHh3bDCeawmSXUBfErERwq7cic3CK2jQ
yV2YQG3SMXaZJodOmT6ShCMJLSHAW0zVxoArBlayjmSQlSptBQcVJOlcJfFudNu7z/pPE4QG5vz/
AsdFK9nSDfXX5kTPxvkUF2pGH1xngIWqqb2pKfZyg3d8y1Pg/i3c4O2vUbKRMxk5j220b2QMilKk
EtWmQFs16PLli56G63E+ktc+8XJYDAdA9heuAsTSHWvNcqDZyv+Lc/kSx2UoQh9d4WvEIsywM/RS
ginPfcC23sNPjLxMSzTZWtLVSSDPMgXx0W7SV8ZqFR4YqL8jcDUcy2uiNFUkkds+/67rDcjlzsSb
tBzE/MllYBukRNEEuRwPWPl7ZsLZ9fOMlbCDInsUjBcp7eWVXBYdn0F1/1Yo51OdZej2KpGhYjTL
dt9WIZ8GfOed4dtgaevdP++vVKj/aTlyBiZjhFMZqcRsEO3uT+5oOqXR3uzuIT3aednRzTvQAy3h
CJPNdCKyeccln2yvLBD31KwTU4DOqPNYbrBQ3gbiNPczn1yKVJ45Z2/9+q4UEel5oOr3W9cNuB5U
O+t5Ki9CajzEW5YneHoQAXu8RRl2dJQ3L7/zjuDyQaPnJ9Lg5Wa55bkDu9SWvAwpqEfehFjSHBql
nfqq4oOxDFvHhf9rK733p486cTgBRxwk3u0Bncj/eD5hfnHm8LKIkUcr6eoRiOoy90JB48fcrZ8M
BdkW54qdM8Xm7zfiPfNic7905uWGagYBiL/wEq2MCnAC1AwI9YV52RFa7SULAcaQ/T+f9X9cnwAA
qGRNkFetGpQosY1ikhYi4SFo2fp+MhWx6eycZYStgr0s/Dw8JtpRnU28xQMNUSuMQs8c+ijNgpFh
OgBKLR+FZR1NFRdz0WtdtJm9icgLZZG0IZdaWrNeki6kGesJ7x6CJ/WgNQG3viI7K1Lq1Sy9GZ8G
rcNL8MfDfRAI4gCfPz0LZuu9zmA8XVYGEjDaSv1VVrkRKGJhxunp8DiIOXDhkekpYyThqdU/Uh7S
OElkFi5G4alTP0oTWKXIIfEH0itCaqL5dYj7OEZIwQYvkUp9QiiBQw19oe0wVyfI09Z6jIP6ZzDs
vRxoxIBM4g1WE/rmW+MslrrGHa5JZ8oJCQfSGKtlCpaBnX95Ii+eUoHKxqDbBA4S79F17PXt2zkH
RJ0yci9n7MwLn0iG51tx8IdGOxMzmEdSYkbLpBK6Zr2frdM8eKlBxe5kbhCBSOHEisT0tl5znVLP
mpAKQahoYXDglW6pTBo+9Gpab3MoBVepi6Q3KWmHFmVVzNyItwuWF1WhL3UPp3pgEiz6aH6kPhxv
+a+JsreKyWziewL5Yic/9uLlqugwYhLaTPv+IQP7ysfmGEuS5D4Mvwb8fuwumsXYqvC3gkjeAqBz
YhLYJyXN+5YHXK7XgHmS8NSDrjpCFsyN0xb6sH2h/8fY5gzpknInMQTQnuTTYBb946mEPVamycAH
WtZ9oUXuI5XqqB/y2GU7kazOhFchEosNzL/c4hVqfzsTRNphoWi594TZ42LYI2ey+ret+FndjNsR
Ogcp48dBYKU3vncV8CwApqE9xXcsRGKKJMHLsmkjnxc+lAiL4zEdR0x6PPsv3tujmgclUtBU+gHJ
t9erAl8YN6Zp6GcXCYcDBrpPOV9rn1TpenkPo2qfm2/0LwMS8k52Flp6GAELCEv6px8uzD7CAYK1
NdgMgeJjRKsxG4kbFPOoXp1en6OIJuY03kNsCIE7Jp45B0n5XuT8UeXCQpjY1nrhMWb5yANjJ9f3
tXGeh29oRWPinytkNAc6URm2X6fzEADu7NsKu9ZWjN2T6p31oW8EeAicLnXSf841qENZkjorQAWT
umq00NKSC3wgYSdNIaKzV4OqfE4k3fiuNLCNt5LVuO9xAt+3zVueRYrvatFhsx2BLURDp/l9JcEW
3MVPbptD2YSaqk054pSyTj8HeB2kaT8seUBEVtx3aM3eOQKutikEYvvunoWQ7AmZW+PAPheasXIf
svmjZvqrOzY8OtMjzTjdetgOmr95v575uW5YneH81QaBV36J008xpnFICZK0Hv5WiCxHkjpy6dL9
7PsZzmE/fLnFMvzQ9EpZ7F5/+u15dkHSvIxv/D3XXqzV2uqKyPD25sVcvf4fSroyjlO2YNz//x37
l1sZFj1QnYZGDUVTVR4g/m8cb08isXK3bgclkTmul5V5sDV/BO5qBfau9yZRFWh0TS0BGv5um4mR
67+yf2qAVnLYdQ3Xtam60JBYgi9T+eSUsW8VX7RegkzdnEC4rZ/eh/NCm0JhagqRoVBOflUBpy1m
MsOZTviL0eaWTGytxJv6JdlyVUPKcqmnRqe7J9FyfGm9Jh9qodyH9puRY0px0YrouKZVWyJkNFLh
k/6fvsf2DAso+c89xEZT9207KfkSzzQ1QmnJrXYGtIZ7iD+qRoJNd/YmtMnOhufEaBbzvJCk/0re
o1+Rx5LuRvtgCIFVrWqv8IboAjgGolKPTw160JMaSaxoKK21CPLuN6XEf8KaYv7t+uzI754JaA75
IDSyNF2NpidIsQjhHVa1gRQn/buJoISKuPHbTxS3HYQ4SGn2+Uu2bEWvn2Jg9V9x0fkh3XCmHU7H
Ve2eRxuILE5bU29WbK7vFOxx+zSB131izl5Ar6H6b/D+xSj7/DhjthaJh2+5lstt21gM0kHa94LW
9HaOT8fJBAVH/nhQ20pn1ZUGZ1Z8GOIeVmhA7VgQYBqWzzpu1GmGuqJAVROnspt2h/eJHygerbel
l7XjCfZFZUBbowOx2DA3ADzqAQ/ToMgfp72KVxCcJicS+z0KKOfwmQkNnrBA2AaohfFmw3lY/Xwt
7vETA5pqxrlFvZdk2zcjnT0cPNf1JKKenHc7G4oS65e2ZouJt75pHDbjR6SN0HC5R4FlZjlIcTqX
xZcac1iwBlEOP4e0IF4ZM5OT2FpAP8btlnpmd6WO3Q3Q7Ggywlh8p6YFcE7S2NM3mHLkAccWBxgQ
Q/uRGSJ2SuecOiNBq6UWx92662C/Ao/Mm88HkPhexbzqwUXWzxBBZ4nvAman+UF1JbqgnqCfvCNC
zPmC3SacgQ6OeyAxGrv6ltAxyZ+MYYjulqWYcs7l0NDwFZ+KMnndBwOpReXQpA66cxFGZLeF8laK
fRCJNcYkkZsIEJA3hyovPfRVY2FO5nhZvIhy87yDu4ECpcE9dt6L/AKPxDi3eiXnXzjcXNnofmjD
mEIC03oHuz4uQyKE4JOkJz/lq6nhbj6N0l4vz/5W3DKAXSkEPI9qVLlCAzoap/AFHEnNj/M+FKsW
OPtyCaimpu1mu+PM8plVv5MQh+fgxZYyHAqFzUh6Vx3RmDR5vmySsyixrpT48/bqrtbSBMsFBeG9
gb4xm9yB2tfByAU7MMEwfTrTXrsPRg8trXSabG1Mx7qzgLYeEksrovW1eF8QOopk5tGLa89aVZpP
BexwLVRMhY7xdE7NpIQtwtHmE8nJaYku/g5z/Mz8SaHbbGpuQf+Yahvbf99bAjXL5EyckX4sCDgv
Xi0EhmE0wrnJ3z5GAdSA/4j2ti4sIoufSxLDNEiwiFl6UJIdXu5U/GMrmJdAGbTBJqze7eUA/Cem
55bHuFwTnLzdydJqWO/oXeSPQZLpNGeKflGj9w38R8gdOnqhsY0syQIsXSovLfOjzR0Qonw33Z9u
mL0GxuWYQXbceVyedX6EuGxmq2GJYWRvIDB86IPd6ePE9l43AeY8SiMSmncxt6F0qLsTcxV8N6i/
nBvl9Q5VAqSUMaaK5FkGRd9Ew+4ePyrEaNkwIa4BkvgGslFPan+g5IZGFQcF4fQMBS3TL0JH6H2L
3Ga54jeGfgHAllIJsMx/hsV5AUsQdus0k4kurwEU/kc266ZaUt+35kgNbol2NqRiI/NDhUeUMC0r
yi8SqtCrSNpEzFIFlW/9FFbdF8sZuiDte4Q0hlqlKsWoi9zdwDX6KxGBOCuOha5Kks/5NwZnB3s1
3dKEoGZEbW9Jq9z4CXW3fwchOeIIWyzWBo/3TtzezDvNflMhaFR+dfN6Nu/a5p3CJEhFdhtcEcUd
CIt0ZnwNormgoekfhZzmNWwHe4srrzXKallaqoUedOWC9u3tBCeCx8loP5PW7so1cGQh0biidAD4
/Nuw7SXkriLOrD1wwJ838QUnBDQMotqGUbJvdXKknK1V2+rmBMGEBGw4HVKU+vTAtul/SkC0gug1
8VssROFlmZOZnCQ7xUBf8zQNxHAMqJP7p4X9o1BlnTPQXCvHNUxKpfP+tf4559UvWL0npdGJFIcy
lAnowB01rlbwXW8PjA5qDFCLwKY/kwOgxtzTLQcuxx0RTn+zcHlBUllw/J84EDvR7tkqLDBE4jhr
oLnjMzZwkF68WaLCSy8GkT7wkw6YJSSBn75Xf4QjXHE5RJOQ1hjdWcF1rkeqgXXGavV+vDCzbsBy
D9j5CtFWcFPCMHV9nQVeRYBssqQOc5igxWQw6ykDavbkdxmwDvP23/y0+LWicrOowcLh4y681XIn
gTb6s7Ekg2yA4Y3X51zbRCq1vcmsq4sJDARsX1Mtj+Xzli2hMofuq5/ZDcehyKvYRTO1fw1w2FKe
zCYH0DG6ZGSW9geiBUnluVahqDVEmuc6m+EDfbKUqrNqlK26OG8DgZqRMfFQX28rmF0GvdiNh1dD
1b0zcPkkRWccmF58sAUqaNnF2JwI8ZtPGVdkcFBlKamp51E/Kb1b4vxJkqg8tQCxYYj8+mT4/Sd5
dZ7C2zNUuQUj9NC3EerL6RwGY10+nhZmLDaL8KBwMobNAEKuqjl4TCZUIAuUdrhvcZa5V0r/lJAa
NwojAiJafUZWVaIVEzShA8gL5QDNxrD5MV4XgUe2y7WlKx6UxJdXXTI3mvDXvpU2ZPU2NX3JGRdE
CFOvHGQ5yxbkmbDD4/hIuEFITt5v3AGnC3/ZtIb+gBObg5b7JWXKMV/HJNS8ivKrnFrzNxFZhxkf
aLpx3sbPNnZpiFpXwhdEH+6qseovG13LyfUmMzRtnx04ZtBaCZYIQwzgTJDDuJhICA4Zix97ljNc
85mRAFwcojrqG6p4xvaT+8tavFna6HF80T7Xi9z0Zug4O2+QjLz9cxF/eSwV8uXTERKqgZgqC4VN
hJCvW+4FCFrh3NqRC9g2wdA4M0e5EUjRoDgvFse+bh4KH15bloVwzebQPShH61HaTxwLpSFbaS/g
LDKmtZoE/RRzNUiX6/esaBrSbeoZGt4YSROQ9SW+pVssTU/Kl07hVR8W9m4FV3g7n46W5My+0z7t
w56nTHknb4kMg6TNZqTCDfkw9xxO406k/R7hfBgUbFrBnLWS//Sw1q5D3ZBq7o0rHYMnzWzgmRgo
fOfyCGhZBHrS48KG12sMDUPL6/nYY8kRohLd3+A/PjnMv8UU4iYMWjuQazp9en+i0JwnyE+1lzKP
QH7w2pxtwxbdwmZ41eqkxAPPH98oBMC1sftdcaYQjyHuuYy5vIpmjnLwE+607x+Ggxyhn30OrvQG
c2ClyRja/K5xi5bwfjcPbYg2EY/G4z7jb8PdBgIhAMLIang/7srjyOeagLY4O/OD5uKrSHiQuHfb
VCa3vmGuHMJHA/+hHZeEYcYbacQnlaxGx3vRl6QUOrNLtJCxa2ODUefQVgTxAdhUVBQ/vrkkBot6
DpZ6WtNjdeNEPfjLpf2KHehRoe+fYIw3KJzrfJSRQpA2zp332wI4sy+X50X3c+luE55AAF0jx3gA
6C1xDYXh28Lk/AHzcj+WLKHNz1vmonr2pfKkWLv2D5txXtRDTEO8sB+xuMRnCr8K4Fd91zWpJBz3
Ytrs0UylEK/ZEH+Xcx6RyMulpUNnjfoPBOzkcbuzqb7AEr1NPmnlZ9lsq2OazHLvPBPa1hjdOpbW
WbAzNVpITYE0zn7gbj92IQmaSZ9t574j1o0IVFfoD8w3nYXLrA2qvUQob3EV2NGGIru8xGTe272Y
UcodFRTEQDHu4Q2CcZcE2WjcqFEmVswwAXDoiG2cBaNBND45BXz89rI0a8Tv3+SGQt5JzdlmVcQi
vCrserlABtDFxmpVsUzcCcH5k6euijtODvfDb5BhrFqb/lkJ5MevTrnxnUydPWr2tKo7phs94ovI
grzG7anaTSu0I8unjixuIxEaIFLHfOj3xLkJKov5TNzWRtdCT/5rFQiCbQuVUh2Rqfx4gVevSqv6
aoEPjpS8JxV4jUksdCb1AoQAvtFdlubS6bSORgMX9D7tkGjI/7nosnu6a3rEx/lqgtcTc6/AwKza
y8ciNIsebxe+Qgu7Ywf6hQ9FIsZ6hF2JrqROfukov6GBgxgXLrRU8IH0YQ1enLjy+wdWIDHwWPl8
x2fmV7vUzQyBnfrI01m2u5pIA8CpTliscRxdqs9oZyonzOZuwGVqhXL6Q3Ke1rKvOwZtx+8vbVFG
7oTrpVuRneX1iy0acjrGpomlBb2bIOIPAh1kOBEEfpHZ/7wBIPhxwgDnDDRIlRjR67pU12DS/CSj
ST7YKccZ2g3ezba8x3fEq+wHJ+Trg5WdRBbg6RNJmVybtTnrY1WhvRCK3n+hTiH+BUxiNkFd71dH
vdFau5DNkT0Q/kfRIIWBDCE//xuDJijulUR2zp+/nHCfGSxyXYHxxRMVX85bJ7lHQs+bpOflXU9Q
E22Mog1KYhW7ph7puwZxEo/DmgR5Mt/PQU9meIaX0YN+QByQnEl+QZZ6Ad/lPaYHEORkgJQXfK+X
RAUTxoWZB2jfUy1ywV+dmw/3U2s25Mn7v9b1aoZZIVWJM+Gv+JOmF8N+K5T83PeCPgVszLI3UNYb
2/ihPvyONXEQZs7YA3asXPdMdG/o23n8z82oT2IFrJBCvObuI4H6EmVKNMOmxBk6IVyJkxAlt+bI
U9bOgubhJEzEXHkZojAZBv1W9A7L0LVqWdQo1QQ02CyDeaBrFKiFq+y1GwGPT+3OuCx9nn7Tpuqu
BzF99Y6Bd+xsekaFc8wPG6/JT3iyNNkCaEoMMTHmI12JCh5T/U3/2Kn4rqSs8vGIXcJkg7jDWu2h
yEFaAFxm2iEvFDG1RO9/B1eOnfCo3MyjffaO59iptiOPVOmLXJwTuGi0xFd2bl4C3NmuTkZNgASY
JxJ3B0bGTOw7WhCtDlY8Iw6TMcfPpCm8s69vFcq9DEbACmDYQf1DvNiwXRIXTOfWzckaDcK7tdLp
RUqRfoPwP/nFYJwu2LJi+XLg2akcHfIqtjE1pu32l9dfPsZfRKnEKhDmJS9NSlVaaIXJTTlE+RJa
nwi7wgtGEshdgwHUYpzu1gReTs5VDdtiQhPsTmi1MReJ0KJrhv7CQEpSuKrFYKkzfFwQZugIyTM4
OXyxyYYu0ToYK4WJKRUXsmvuaKBSMOLJqxHIC26fZL3+LiptCrtMOupAiqRRF3kUtmKFCxj0WiE3
PdF4LshMhtI1K/uK1tLkA+zciPWJQNwWHltELNrCUaelz8pvv/irfszKi5lnYFb+0JhdAoGKtdNH
vqIgP7PjnxUHr42/D/GoxJESmStesvT9wxD6gjBVdELJSVIxhW6iUssQohrRgZkBnO7ciVddl+QX
jrCiWW3NLWithM+OqHCm2YivAmKHXIQFtEmPRO2ci7mXGM6swQlCO1rxKq8DSbe7Mg09Suu8bGtd
npVij9d4/N2myhgt7eLX7tzcvsFXgHj0qJz1fBZe5XnTMRqlyRCnH4fK/cWYsDjYwXsj8v2n1JWo
9gOz+eVlYzJdlkYdEoB7n8yWbhmemYg6pgv0B/9uIpibMSEQjpsEDXtNyHITn6gmyb6PsBRcNuhl
sGfnR7p4TJfKl9HvN7u+3RKa9JKyXrSxX8EV2uf4gQeWukoC1w6n+W89bTBnZa40O9oknweW5SKW
5WRa4G8ohdYIdHVS9fmG1xOAdYrBnP75G8HppYY1p+M7EZolePNgMB55TS78XXt5uJ+umM8tVLuE
uRVkYfQTHQirckIf0ONkRCHdnhqIJVXkdz1b5fMivJbhI4Iy5Inx24X0YDvXdPvizbrcs317t3vA
67NmvRY9S//q1VQLSrAUGIidlm24PA4csLE/IaOg/+KxUCQZPUB9VrRKe8f6BJityo2HU8w9KS0q
DbKQilvZGVf0xI9LSB8XMdK4rubTqt2LghDfhhZZ83gaiY7wlKddpcATCxjGn/EJyqnUiQ9+CVJ0
HpmcFniAjaQVPlSu89yZSpjVJY7V8UqABr8FTnqmcirlU3yxBUxm+781gz/0JScRZcJm3AytHMcL
CFBe0If3Imopyc/AnlZqaJ/veZEuIJk0rhmGV/iH25iedXRqXWO+LIFNWRBzlcTQkpLMYJMPK9qw
Jn7mmcd410KcSx2c+7WyuqNrf4SGbCt3svwnosqwvIKhiBvZqWJHSQKEA9VMiBEovIgeA9bbgJp/
4hH/K8pHc56KO1/+W89ERTrdLi5jUTF+KRK0En8+kR3e8wcZcokGPCFLno7J/Z53a23u0riQTiXV
hOkfOxiV8+XMaiFqTtv17x+qk75sOrG/LK/TSv9ME3tabggE1N+9tiDDhfmEe8V6ZntA9zPNyiX5
nbg/AZ7K0U8Su1EegYhNB0kI0JlFC6qzu/xeKwVFph5LHMQEn+FhS9iaSWs6yFWzjnkZhc09TAva
1Mk2OH3Usa77Wml81LocaiVvBS4I67EWKARTlYvqC7dzq1+1IqAJTvAwoH7yuIP7VHy8vdlKwlHv
R6jSnUGfDWQY82Fx4wZyFSM67JE19TuwoYJqyqqL4TkDIdPyby7lm0tdJCHmRVNQncadYoEfIVpm
/EUlz7Hex2fOeCfQWh8Uj39BOAAwFDc68+jaKPnj/zR47o8F012gDcs8CDPVKjdhwWFd3Ah+VkxJ
ffaPKEq7OkGuV+xBsrbtdgwsuiof8K2tUWhXn45GuRZaYaJmtEiesEE4Lyki0uSGsWHYn/6Pvg7E
ORkcwOSS+K8EBXySvEdfu1DJ8bX6xHYUGb+UFl/WNT8wm1Tag8lfl0MDiztULU1UROqSaUFLYg7P
C3CmaFoPwwaEGs2q/FzzEVK0R6OwqqURd3L0+aSETGhtO+UqDpSM5its7wQgP9msmSPSIPjRhfEK
qkBJjXh5j8raoUjZnT0cmVgf8HNt3gT17v12CXLLI3SVeqv7JRNQePDjpdMWczXI7CkDanl5k9LM
w/+5PGYlNESMqItU6KqMDZJ1DYt7w1kcqpj1AyF1PmNix49FQL0IIBts+HJxeiH+8k7QZOejFQZG
NQ+2CtePqMgY3Gq0m3e45EMJIJZHNLYQc6JxWMYhXj5g8HiNePqz5kMg05iavGQchauLLPcYswcq
1zjqShd/tTeO3IqBMBcwpC45FpBbL4Ck2CAZDPTIjqN13871zize1gluXuhZBIBJmX2hkv88Q6na
DrQjnq1uu2CDJEE3LKCL6GLeBZGF3B3wWcFI37LeqAPsT6iNnNcBx6QQLAUDMWfsuHyZoHIENl60
0PYEnqgimd9lxbIyjXXLDsxXqvbp0G9cQYuoxkZfPUi6X+QZjZSktP3xofXqKD4Kcvxc2rIQLRdG
90lpFfe0yl2sS8jArDSEn+dLIf2koMdTxhzPTq5vyXJVUwOc9Bv/BfHr/W2MQCCBEuTQaFSkxuOc
/gq9ZMmkM6PXgTsm705ZnSX9qO0uetCJoa9mXVN4+UccW7lghr/QGMIKcG5z8veHLuAyo5w16bcM
BQnZFE32Di5aOi1QktNBTJ3j+1ZPCAsLWb8Ebd3vkd1pcKQuroO+aXqJ4qkKdcOITeFpQT55K7nV
/19EQObkr36mrMfLtkQMVVsLZHZEWqF1Oddt2pBh/lClmC+MQVnGvjpRTPcH51ZOMaXGmA84OAKX
i0N0E1COpwk37UB95qcCfiEUA5ycf+pDTIQEnHfZGchIqPafW8iZqadl5+++8uyUHX4e7XQfSGwm
soYVJt0ggmqVbz0TmBWRW3RVoeMKC/6sN71aRaotw2yjroNWbLx3SCqin1gILMz3VDdRtnInfnyF
xlfOeOHcVQ2914Qx4/qVUSwVLCyLVFwaD8d1Me3lYaD8LnHsZxoFRs3dixFjOHC0IcQ29A3s6mJ4
PlJDE4RrCkniNeN4wtvlfl3KaqwvWpBS6YkPkqtt/qZZAFnpUnOd8xoVtCsiZsgOK7NoN5AI70+q
9CrhDiGG+4rwjobdtlJx+fxmSwxbkUgNW2enKeSf4z23wb7i2BjRHu8VRHad0lx4R+IfH3Pn5Gt3
o66vT6dW/486JyW2n0D9oal9s+RIYeI7axP91QLg2GMTQBSgx0Q4zlaWF8DBvjW+061Cg8w+1ZwT
JgtPDYAeEMasQHRaxReVHkg0PtBMoc9mm7Jl5RYQLD5SBuk3qR0dq1cfcVZEuu5s5AeY9rIv1n1b
Ti0W5eks6H515gLKy2t5hVJcj3xqB39ad3995D3pMl/OUJcOHkq6wHQvI3yKFsWMr/8IDi69vTZU
7IUIoZsilz6qXJEdRpJ+Wd0xHPgnkvi8Na0tRBIWUSCfP8cr7mAUwpkDRKwSL9SS0s4HS5H5Xrrr
hKKs138nPohovbhCwRiCJBZ3+5LSiVmi6Lan4hEZy2zvYACwNCnDgi6QlwsdkdAXHqQI2mzXx9HI
TxMVb6FVoGAeCIWpzcss6g/QDrkvtaZfIlNC4M1jJaI023UVRR71GkEgSOQtKHgV+JWGQakmPM9F
oHTeaJFE6vjo0LNe5507FPT+7khzhDpwm7RjEmvt3YMjrsISJHuyL1Mdhjt9ssGYZIDy+lC8rCs8
FTfOKGAjFfqW5zTl900e6WsPq4cETnHhJ8a1btTb1+/ziFNlz8tlGFRM6y+kl1wVvDmyDASjhR4E
3lxCf5CEuTq2Jo9FptwpLM8Kns6QbgIqrtzY7yE5IGX0xV/Ewa/DZSHp8M7zXIRdNiCS30zYbFEX
RvBVbb6chV/3LHq12zfnzxoPsLWxT3hKihRFU42qBDl3NKAnuV+OaylhmkyIEOH8EKUuL3R/5IGE
jKmB3p7yoMXR/8wzazIXvK+zOP55djh7b8UK15yYHZfTe7qMgss2f7Kljueym4qxkNuoTyAQciUJ
ZB6OfyzAhtTW0LeQ+0Jaohxw1R/XXo4salPkiqjl2bF/zFqM2FpzKkeoh4Bhn6GOkXKAaa7LBkch
avTikfIvne1l7R7BdZLzKnOXVChP8oFqFHE22C86rQmY1m9v+b0mGZpUhh+VSz1UoiRUZih++zje
eriQjEv3wmBQYcEyNH+et1erXbt0D4FRF+taXKUPQ0L1Pm7kn22VOC7QgztuTtjBjtljmBEeQo8A
RVQQxiy79Wb5DbSwgWRIVEBivYz2ZC35DXd0OOUFUt9OjYoRZExRFkuH6p6P0LvndaJAuhJAPGra
t36c/t08hgQCQ/fja1T4SpzhPUDYFKlCX25HYEPUkcilNZ8j+iu2ntN91h9V6525cYBl0T9pd9XG
Vb/hWf+m1r4lrHj8pI7WiJdvQNktX8xDpBQ5WovEo1CF5H3IJ4HBGfn0TOo6ibSbxrIddsWyGRCn
vNABznV38TQbjWSsfhFhRrw2pS2ZLYgyw+0fZLB8XXNwk5YCXmQ8fS26GCi+RGIVEXcLD06Dkb0K
Gwt/ynV0p3eV6uBWLM0I5dOXyxGF0XFsRjGE6uRU4RAldoZiBrvzSimE9BSW6zvf3KdzwHtSLwAX
SJp90SMbA+IwhLzYWljI97FifsuK+cyOwKbEJtXak/PHv2lWzjqtL9eHQRxBLgJGqhhgLqCo6QHQ
m//ky4TXBOFrxnP8LSQQKGk7qg8fvGU0SCqvCOs0LTAoCBT+2Ftcb5LaIxZD3O5dTsq/Ey1D7O9b
mKhTDLX/bL2hIHd+47PGtXOb02pNqy6LN+HR/4grhBMJ55d6CTJwovSWgzT/dpDVwFpR7UGyxP/q
umj4ek6Gg/AYIxa8LxSo+dHTkPPTzcT0ApbUJi0p42GYWnwhoLq7qDUAM+Pzh/w6xTn2Vz2W5eXe
fzmQWczZuOGuk/ehhpaKr+xc1jAPW4HhCa0iIQARidsTE5q42WZDAvOxDYToy+kFt/KbtNp0H7wI
4XhEEKp39ynO7l0vAXxc1Y96fSqjfyDsALX/0d5GG5BVb51arPFTkvhl+K6e4WSSryMauB3xxNQm
+2h2mV5pZicCaTssRW7FjISICrelc+Yd/KDUOXRSeDPIy8qOSZeAl6j0edV2cjejUfYZv1eks6cu
2V6zlZR6TkwR3jRGDQ9///d2P+OfW/364Y0OuUBdx0u3/2sEg2tqYkOQ2tb7j8s4w26soHMRWIaK
q/Pej6u4wlcg6JliM//URD8X4xwBRu5ZJER8mq1Cc6ExK46iI75HPvh4lyRBrmyUA4fJHqNA/kcq
MJD9txMoYFCc6qTpLPyOFWdIssW4zesaY1TQn14aoJtxsVM6qC6ogE3SNBK/NEbu9R89EONvQoFI
9Rc4nnLLYF1gUEEDxz2p3brLlEEJNhIr4b2lt/ZCaprAOXCKlno4MQfcnZuSzZ5JdWu7x+G7Dkbo
dlFuK35OdC8aC4fvnXzjdc4uEVboPfGoQhB3s6HBc0xWbrWBykgzOGOUqsB4vpZwNNvP/91WW34B
NhTEOgPj4nqag9HPYHhqQOFq6FDXJVDEhxsij6+7SwB3Ea9u9dPrpCYHktJsCp6NSYNBsFHBWROQ
MxmlbAwx95cI+IvafGsfJatL4YskkIE76wbY6xqN3szpQeXVoeNLmfzy47cPG+ssIZUD1z8dQaUt
for6xbV7QzhoVI4BRi62nI0JYpmBmDBgRixN+4PePvrX+t75JCJUW2JAXT1zqWHeVvxqdX/yw2qW
csokaNLFoOpUsxGSRlZrgNBSpG5lYQAWMGlWas+NJ+7mMwY/gcWplD2w6cF8AEP5iFgi6GJxcDpQ
8PQEc57WgKirzKustXFWmfrrLhf94oS6aYv0MK5uKX7kN3gyhyyl5mvJGccuvQ/jd9HmlwyU2jAV
9hXMYQ7wnnV7bhBXL0W3SJajoYSH+kDNRvII9ZiHVfNV1rjehK03moJeAEBwm9+ebYUQcvq/Qebz
puMDcpm1XHbTt19fMSWhqMdZPBICVgHoN9LzGEOUX0rVRFS61XBeApihpuOJGLiwmZI3SxwRlvRs
APE45a2iyMKI0/c00eJzTM1E9qodMdI5+EmkhsxMoh7PEq/o/9TjRNCP1j0UhgMn7T8A+aGIBtfA
MdNRYNvXGbQO/178acZkSVtFzrT1SCHihdk63s/ChKQ0rsYDPVyNQzHnjuH3sv0blNPNyAc2O5+J
6kN1L+jYJ+Rp/WKYKcsn3O8HzKR1wKT80MRILHVhayhW2hCeJ3AI2IPytLrLXE7snbtD4WJkSgCF
+McEDPubFMcncQHuPGlAvFSBerhGZwNJ9CaLnUpExS3Ib2hOODVtNF6c52PkAEPfw4xyT5PIFNrY
SF9cghDrKdQwq9rERvYU0lWfacXAoeGJqZrCRk+5wd0KTdBmDzUtInc6pdLGbUMy7vGQ21E6s1fd
VzYED2IgmvwHrBfT+3KnUualq4eTsJQBE9PNU8nKARcBfs6Mfj/5RLRiqZiIybpEj9x6VLsBVOOT
GkRXQ9fP55INrpVHt7UENmqODClKt3dxcrGDOEOwT8KuYVJwSPqYVwnnA63PX7gAgJejMc5+52RM
CWHrAgicHIlouOfMjfnvhoRgzIvpJ47k1YXcTUAdJN0qYn20liW6N6SUJVyzqegdL36ei3TWZAaC
EzqI9B1JZ9vFsukS0h9eigwcMvfxlUvzuSxq/zomDbbEgE8m8siVtLLQdHgm10xGq05H7zcdzbX1
L3CM3bitdLVTD9djZcdHNvy7hF20OCSmx3xXP34H/XR3WxtkNm0d0peF6MKJng+oTGFjo04vvnrK
kg6YBsJ5SWrD1Qra6AWojKISSd+TMHEMMbZRg6oNM4O1jrgYZb2jYDHo8i4VoCPgRWQXWXPHnQMj
TM0p4SMjM0Igg/zapZq7wjGZ/gxx80F5B0k4UR6AfeoGfE0rMbnqyabLzNYj6DdKhXeogjhQlnMP
JB5HE0oAxdDMLLme72FYI63XuwYs9LTqrKndr3hxw93Dkk+3Llb/MVuyXdGbIyeU+prCc5/iIf5i
aVFjLC8tGPpAdTo55Bqnxixbumv5OKxElpATcjNlFk6VdBwbk80hKKqjqDGKjMy+PT6WwhZtcQ3o
hsIkOln/jdLcgzSurENoZAb+k8k/sPPpwmFf/RPDD4njCePh6yiHFKvY9sgtWacI1j3XiP7N0RlW
egp7dYeuCRUTVZ3mSnU3c+lgN6jKtP7ZMaH+E+DD0kMakC1LfJZ54QY7T/22eymjWKSnxM1+uY4N
dEZfzlKgDGcdAhnrZK1m0YYhLLe0YIpgqztOaWYoEkysEhjbh4q5ueAje5r9VdpCnFGJtUHjP+6G
vQCkdpv7xHtpM0j2rQrl89zcLzJ8w/dkKij+2URx/F1XvkaZnoeiVo31BZt5IdXusYiKRyG7pMCd
YWUHpROTgQrxYzAamzv85HwBf/8HUOvw8e0LWTt6ssd5LGuXP2Wy06/22qOFU6YNc67AX8IXcB4b
wc+AOhPElYki50i9fefvFoQb2gyIFopFRP6VbC6WaVdMyKHXz7waLiMNnyKUuAz1VQEZs/IyRAxE
372zk2y8JaojorloRGCVA9RcmhywMMzwWRck907CD1r2RSWUgxhasWvUnVgvr8Zg7HKj/miVMzRM
aWQy1EMPGz8k+VzhArLP2E4aQ94GK9hS89vqHm+PtSoR8eoPezp4Edzz12ewToRuBYAP+NrXGP7g
XOpPGs+pZbwSFvm94tRCRuqlGe2y+rq1uuWz3HNysNGU4H+Z+tyN3TMgQAxJ+19/+uVEyn9zF+yy
HtyOus7M72t1IlMrR80O6fcx/BP3T2sMbPUhD2oGbKAQ65Vf2r4ZDYKwRwgJ2trbsJZMwO/ppY70
enqU5rbhOmTO4XNyTopXN0nfKWsovxs+hJ+TV52p70c7CD6zzlRDn6KdY7Cj4vtjQHmbGgwdLtAt
wZR+unzPWnyyJ6J7s9k0wicgJLF47VWuAfLZa7RODdyTR1TSEu3cqEF5CwtNnxXQtUUXNrEh8fDP
fALwnVIbCmmWAYzjhEYO2RlFCLvb0fiohfc2ZmQc7Pfo8BbJ2Xu152O2v0sxhfAac2IbRVlIGJF8
TANXG/Zmsfp2WgSJcWffsharzmMIgWlVbfZGWO3+bHHsfkvYIjWVOIwM4JEjY2nsTnp3FqssBgEy
EFZkQw8GgZhV8hrrQPtDzdqDH7UyHeX4tOo1yH1Yad3PBiTjhHrKBnDbV69AWjTuoBnXUyt1KInA
oBfyDdGbjdRcCgftG/JPM2eLplDmO6akUfmDPUj/9wucFPQZ89OdfuP/L5YR/F3o2x3/c5mBvwAX
UDl/AND9uWnCHVzTau+wEEEIFpbkvXnu+PZ5s0GmhCUFhUU1ymH6f/sBVdR12CwdxZIXoENsEKG7
Dvuz9mGrSfqLfKwk4c/82Yv6YJP6ZnLpUbY0l3iurWKcjDpKmxa/t5BadX5xSzWuzr3lkNW6ftBf
uzp/8QGDzSeTkDaFI9TSlYy/vabP7gYKL4GqP2kZDhMD8Z25lHdVHej+CNfFPInDZZPEZx2XQbdR
nAAjv7rxB/i9N8/r27+Lk1u8Zt8PUSfE25Xlj66R7+qfpqMaGYXvjj18/WPCezRiO9JTlq5ggOai
XvYHSa9N4CoYT0TLsIxvng4OsKRfbx3AZFo8R8031MySbGYI73qTRPjz0aliV8wS+vc4iyeM7PyV
KrEsSkKZfXEbdd9Rp5iot4VAuYdUznfWHQbSys5+8Oi897n4DMr0gCA1PhgaiRVe5D+m10ktCulM
mQYXirn+bt/hkuJDKKVnPGxqKdbF+O4DyJlMw7/didVfMW5Kq1CHoYxNq8T60QS48VvjLkaK13aF
pD0pabM6hXTA3VOaaNFIAkDGsmHRMvpfr+ncnWmMtwjC4Cf1QZwJAFc1olWxa4byAX2z4XQdh96d
V8jmG0P3XqbDcHqmVoC83+TkVcrHXAXBoM+GcElOmh3Q5P3OfbyAsmDnv9UyZ2zXiuBqWmwWAo+F
FcpzmkO9QOG0VtZdYi5AImvQqoMDmryHtmvajqu5aGJiFJhxqD2f6zyGNZf0IaTZMJiadDMcLiBE
5+RNye8Rvk/jMTogAyB/m1D+t9gemrlFvZrqEZo0HUtzWiXrYRYki645OzTM9fE07pd7KxExF/IL
cLawTuIPi4F6ANExuRnkoOkc/vStCU4LUX7R46l8Z8A2RdcjIu3fbLRFO60TJaZclRHWG3ruwMI0
PAOB9gv13hVaH91qpb/mZEpEGM0odwtelswzGiploBfXIkCnryw6Hs01iGZONYKtonWZkTLj6G+l
4eEuEL7Ar58USz90BRmLzdbrAYj7jVKGdhY235HueXU/kpOdAMXmvS1SvLBGLdvDB0SygYoJI8nN
3yOupiacvnVPMfGs/L3fmTuzs4Sa3/aPMXq9sizkZfMPHEYsapSSMIWaA4rBsRFlZKytzl6YRQv7
sx61XKH0cyZuAeSSR/F7TSNljf1ljXJDPMueVXV7qwILKeUkx1932LtP3gWMvKxiiCv1PhXPkrld
GJasI/rVSgzAFf5nCEj1aL00YrZSkqpwdI/eM24fneXdoav2QTjxOxW8zbaW2LCcx1kkRfIWOpP3
M7yl4KmLWiUtIIIZWSG3nKuNwCKtjMyFxe2hSAZcAeeCXPv4m2FI4Phki70CcIJ0QAfHW+Wq07S/
V0mtiiIv26tEnK878sJ+w8V5jpSd54TKtMDmPp5kjXOD1g4JgzIQwb02zYprDXqUflmksE5wGqNz
vxih5Huly44ho5deVw+9pAbB/bhSOYLKq+A3/aT0DKUynEXUKXm2RRuNqXADRKmIuQ36kPkujrWD
z/pCO+LczedEFBeKDf5pzZCSzdXH3aawb4jfbLOfash811qqz/xa7x7FpGFRXVQdNjKucmVysTUm
mhE1R548OliyNhhHwW6h4C0FxGqiamgnHzSoetWfHG4/Qg0F5hIcDxg2CnVyURryzweV66ebW76y
70afQ57N95z2n4tdJNDJzXnh/7jPv2B8LDV1oAn17fiQPzeN2976/Fz831KAPpq/17lb2WJrBOfd
KLkgTr/KFhsySGWZQW9XDK12lXZGAW8Z6vv3OH+CcwQlWf7u2+I+6zvHGDDxSkoSFsDdXmNMjosO
LKyPi/H7jR8aKmUk66zuiqdAD09HZUa8188/RO59OZIKq6scai3W8mxmL0F9wS9SfPcSQegFLuBi
k3EuMPvxY6fNqUU0l6STv6hJPtkUVM27+0vFESWkDq8gSm5wLsvxcTN5jNZlEyO5fBNWE+vWCBFz
IqVVsdTDiU0jJOp0/powgE01Bacn6CRa5gJvBxe2cBB27L2OmlKjdjE8L5od+W2iyShi33LW0CAr
wnjuWaJODNJfAomb2nIl1d9SolVJr6k/ezC3ldbHyjgYX1q6zfUFXJLwMrqYT5eUZzhCuNJDm1+d
aR6ZcZ+r9Kwzgt/R+0/lmJPOx3vKiF4j0neBWBj265QslY8J+EPmD3nFbvhKkK+2ldjV+M21Xpwg
qvjRsMUjV5iJH+ayuQi72OhPU/h+zFSRNvQ8pDjLl3OxjoD/dC0LnI+0L0RCWbNctjJkqXxBkbVL
CKs9jXd3Lt2ccPUj0CWvSwN2BWyriJNi5TZ8bX2VG1pPfYk0KwBgKWAWGSdlUKrdnmBABgPEpcSF
d82PYDDwP9CT34GxKNIxmbMwrMxHN0Ahrp7o8DkswYMk0fxfXiTH+SirKisfIcqZB3YAEWRQrqZD
bwfXiXKQdlFhnh6bVwct3BxnSJr0LQlNUvkFuGX8LQ6u+aWpX5hPFLal/Gxuth4FVxu/pqXJTAYn
oOdvzUnUxdgy+X+ikciKgNZ3wR4xQ+AU15H+xqTXs5g5T1NwNoW/Qh1hwfMj4lHWyRvVSv2wrXsL
BIHLVXekYlg1UfSVGkG9Gns82zcIWZXnjE7uMzAthkhnkVVbB86vbpFLzXfZ+PHEIXtSUb52C8NM
KC0AWeD/xSdkedk+39kyAh3cMMYqm4YbP7ljs+npG3MSMS8jjA0Xbo6JZFQDpTPaJhqB1+y36LJx
2Mc/936L9CeT1Np4OGfuEZGwSSTEsmNSrsBFtnBHEIRsLNTPA3trOIIISSKcJq2P+YBL/+s1Bvp8
1G1WgyYMjJpVF8zZaO5iXMU7lfPsUAvoxn468uHkfKWNNcEJJJpI49xtlLUD5zJ+vDwcVPWUzOg0
Mq5tpLruvKwyi0vHqgtEBYB8joxsuE34JFriu5Wp+qfYCnil0XW9FqWdN2SYvrXUud6pQiOrpt1k
HJZ1Hn6n3GfxPBO5PAgeaapJAogbY8oBHIGft71JbRwIYo2JE956tuAGjFuTfjg+6hhyfHZE8tEr
7OcS/hEwbdKvBXzez832DZtcArIM8Zgq4AlX5IdGrb38ogoeZkVP5pNjHNgmyXScG0MBmKNtNlei
YXVO+kI+/5U13eArVvvU1ngAP/M5NQadqLG1e8nAI0Gcrg2c56XfADTHPKDPCQ8unStJpQVLHfGL
0ga/cEek4XEDTYVwE3a9AESKR365XqBgUjOz+KFsinLrB6kpkaOi8rOHy2UnbDGENIiws3UEW+R6
GkhbrNw73l/avELPjirc/SEUuvyDoW1GZZZQiNMGXISFH/7wJR/cZteZPZ31bBXoeqdVG7GOkVUe
FUdOPkfmtxyAmOnUepQGlW/ip1p11wBkTgRS08bWrh3hgUxBCvD+TyasUu8ufv37DgXg/g3HyA1H
NID1sieoC2oOndMvNUMk60Rycuhc1B5e4l3NC4ITYbLYaN6PL64LtcDgQY0fetHc14F82T+ctQrZ
U802YcMS9xWnSIwPkq6Be1VQ3q71YOEsYJw0walIgIZTQ3ijf7RqkTmmf04uJUVNq7a2Ij0glhcw
9R4iF5kG4Pczp999VJaWLfzbHIqxSZcf7sLrcSU3rw4ligAsChi/+rSqYKWOBfCRQd0AynVt5Ncu
NTDeW34m5ReH6nlVXrBYQo/VOY6gAUTdD5e4jUmLdnY48iVFSIuGPdQIcMRREpwpqR/5hlqrv/Wr
1HxYRrFhEszKn3lwehpHo9IaTFUnSDPcH/HG4WjmCbl2srVrpYiXpRGd1jFiTs1sAMkdbKlayOY/
lVlHBUax0D55yYfzegnDSf92qM4e2enCon+N+oXe3TKYFyyTEwIX/65F7KhxIqJg39XY2ykEEsWB
hoeFeps7LxU0vl/1Hgzi1bqGG+vkYKb75ULzo4HVLVEJn2dhI1NLp4YG+lpQzfkJr1pBhi6LLgnr
+JLITod9MSH0HYSZGBcLXOTZNu9nA11DCKXdqNhR64ryi0K9Z8GRzb/0CMxxXj1RopvjzZVO7gXe
RKKRZ42lLslvK8C7PY1P1itGexYjL/rsAjUlz2Yn0o8r+h9/hzm0SiMNsEpU3DlCOJhs0wXzlfxu
7nP90QmjTGZkmlYZM9qlB/OnFxLOoYsWU5fDsiUQDJ9pIw67Fp8O5yQmU/KJPZrGIW9Jjf1bDd/T
qqBcfJY1nmjlGqB/gFzaqIDqrrwVoJcJp7qkFR4FnvIzB4E79CrFpFf6UllMOxhzdi+iUhq7lQiQ
xZSzjYHpm6UjvNBFqN1WTURdTdWZuyOku67YYNT8oCQP7WMypTmr0z1l3fnP38ATJLEpmkT5msSe
uAZw7tNfclig5C//k72gRI17s0LwHXgZTqCKdolLc2yywMRTkrf0VD3npDQVx3MRhadU4yi0uNGk
YQBcTdJ1yyvACydDH8UEKwdqMoJml5Qkdo0rWedDb1kk3iaziHnB+0nB2thXS3gpCQphDOlkiNJJ
iGwfAvbjYxKogMKdqKJxio8zeEbhDtga280xKwWdLa88JCLPkEk/TRHj/IhA/jRS+/qd7CsXQMsm
cS/im4Iwer5my9HEtNYIztnoYpfu1ZA5ZgXrBKmDY7C0dUBLQJ9jl5x7DbleoFwKqD4ohlfxMpEm
TOSjjTDtctUeoy62eYAiGWI3byMGyJHgOVG75juQBfJUdNsga5Znom2EgIIYYefIQsTzKtRqY9KA
AfeMZGkW/rSNsH+9eXWaJ9fTX1l9D5cld+AMUEq4lyC6QdO0L82NoIHaqW+VKGeeBbud21+eUBXb
DaMU0D9iq63pyex8d3Y03PgDPSxaRptTas60YvXSeAb16maayu+ex2AqPDzGBBaHivVTXZZ0wwmC
JKyotZQP9qMUSJXJUgOQ1wZ/9XyrICnZm43ZICLKDJNIhctA+Uz0ofFK9E3KcDtfaxegpIO4ObXc
+srDEZYhZft3F+cK3cm5iMMuVhdCXO3Fs2gSg+OUxwdh/evJehInb4rIrMUX7JHos0GKNNLvC5tM
ywo86e6nN11kbuRIlXMkLRw4rbvQg+suh1/ntdmqjx+iLLwTsUL1N1vJMwtqqERVmsuPaT0Ndmjr
zu4bBNXOoMJxG6PMIYreqO/kttak0D74eapWDUDnNrLEKn1z25q80ixaWbHC1n5lRqM27AgRSSE/
Yx7vEzdwXBg0ASnrY7opLknLNeZz00tEgLJ5P4K5byJX7mN9J+MVCSEwBhinVUjrcifItP0JHknW
11SZLYddfzy4sdU94S3IzGgIdKOKGUS/pK/Ifq3rswFncZGLHdLNhtuBmLzU4bytgTVht5L6SLjN
C4WdTcbPXyKvs+xAPau9e4T0UnUSlTZjY+3WXnSDDhZ9hbljiZlyc45TnWeHt+z9ct5QU3EH5RjB
CS1Sz6MwtPz+ozaXwpNDb442TgDOB+yOBH8IuBLoK3PtZ7fSHZwBALmH1O1WCW1yrFB35nfcoc8x
MCDq1CSDFGd66Lq/DUVEFtuw3KWuRU7njZlP0rF95sZ7nZBc2UlO6ZfRXsUyUQs1CJrpEZnIV5S/
ePGmX7vDsnPMFtFULF0Iom+oNmH7uHWZy7IAEMEs9SjfsIC1mCK/hy0lSe1rmk/cbAhguAnoyC/N
NFRJ3CjJaa0x8vz472BWUKRwG4XRy5etyUkQ5fcFD5cJjyrveSS61psLOJo3Ad8voM6oXLAJnMMQ
bTqFndprsIFXpSVC7P3HzD6dTFHtm/1vKuXxuaE3JT7yRw20dX6x4PuCivGiDgzM72+IuTwuFEMm
urNTXYYX50BHJqVORPUjpHNcyJb+XD5b0qxTg46xUajipz1NwSMxN3A/dJNrrLfNj/1sUjfpfV9J
AdYcUEwPsYNRJzcI72hSDs7edhLK/GnRwxdyikd6e8FpWe6I9+RMx07jd8nyTnnAvLB/pNeV4lSP
SWTEi8hjrD9p9jWRD3xi1hEQnaby63QcRIoACBmb0l/dR5dGYmSYdV2xjNvVjW9JRb9X5uDev7K3
wMzYKOnnNxynYWPE80dbMwUXAjRAbebIZrLnYzTCWbn5K//dXvi+J/FS/J+OMKhJVrCrPoc5fVOZ
LeYD0LA2ji8I6uJgCvVu5VXCZ+UFxZZQ0XXmOXgmEvGV8/BAjW83ld9pagEoeekRNp7XTEyrNjKD
4J1E5y8GybjZ582r5yk6MdPf1mazGl5M/lEjPhkuHvVZOG+ROeT+HmDQwi/mKin/GBcr1cJ+FBhD
d9Y/1QXa0+FlVhGf0f3lNMQ/AFTNgraaHCssxESnlezTy8elMwkdSafeOB80sOLGC/o/S+CyLljG
ix3BjkOAG2vB4BBz8XEjW9fVS9udDtYnf2j33tvqtpEWgsCaR7u0sJSBix639eqKppAeWee6XIsr
IfoDymPpWPqrnMjLVJQj9HMb6TF82OPWudABxRB6fOzVCHjqKD5Zkdza5CQD6xuzqrVy/seRPGmB
SbmRkaq7+cB+d3TKgSeONwbuSjzbQBIrhyAuD8e/PbTPvSskJkMkMJO+XT/FZlDPqte03m5i39Nx
EVV77uIftvXrw7CXTSBlcWM8Ktk0qj9lrbW10TpGK/R7uni+Nkm9tgku3PcyIrxEqmPdbnBFy2+4
9wi37EMcazRrM7Xh46f2GQs+PkFW0avboCwWRBNTM2bgCzfTZgcqwP6YNQUmOwVd9kx/H6lPX4wV
TODGAf8UUuM7lKFyM2z9QojbY0gQCf5E96DIpZKAkrTdT5+zADkIN+Px8zXhmrGDjUglEd4lEKz7
oZq9MmD/75Vd0CjOpbpJlf+J7eF8HzFEYS3vQpYGmdERtX0T4ZGM9uHMf8fpEHrtpu1RA1iSlKNJ
fwwtuF5Yqa62fiohmcw3fFsrOkiYeiKSae847b7x6Wg1AwsMNjh4CTy+9dZ9EodQi3D8nvQKduE/
TR0a/z1D+xK5fmDWch6GPAJwHs6pmmtwXRQF8kJaVOpdJTxHOsNFMkpgXPFaufhtnwOrCnUJOJo/
JrlUhJysfhuhrSl3nuebAErq63Q5JExSUPXdY/aWA1UJGqm3fXSk3dq/zaQ9Od2zHDVE2EEMzjWe
CUeiTrl/dghzi64I/40H9kpLMDAnUIlejHETFUY38y++NwyMn0qloe1VkOL8ll0sCSDNq+h6GEJS
H7/NHnZEVxUhjomFjZIn12t4KLuzuNEt3vTYkX4mPv1kyzUvqhKo8kaFsP8M0jX2f5OJdW9uoGkH
F3gJ5v7pr5BiKOIoeM3fSkCZO+9iQMFaEsJKgpbQSsTzrURTQtzY0kUuF31RSGS0MZLy1dqYomq3
vpv9ahZJ0md3qRrlVm9JFUn/C2wmSwETDqT9thAQnk2jcP6uf2fpUp9q3lTE9tdPG/AtIA5SZVYD
eBkwJ4fNjOkQCGo1EvJsYCHebe3ByJgqW5dQF41VpVH1ZDZd1plgkZz70jfaQ5tdmR7TXhfe9+z+
PdyL9iT9PEz+isReqhP17xeCOwCKrcChP4fMhEPeT28NGfCHpSfCjeMQnGBnaYlZ2VKx/lAn4RoY
LAA26LLTb/23p3dNuPBM4jrl3Wq0xpTac8kpWQQ+Oy2YiA3PkQm4pNtGG9DpCAhqAIT1kxTHsaA+
xr9aeWMpIuxPcfZkb1dsYa4a+Hc+y9QRBb7aUNyxB94wwJsNOzXtd1Hbz/Dj599N0rvdXzpro4/r
Lar683pF3c3d3pjQN3CsjInT9ilm+czc+MhPcb2DlPuOuhlOAjg8pbbQU74uHMyX2e9FqC6njmDP
/CdwdHKi3tklzFeO3v0kCVJN0lgnwaM8fTIfJRaBTtH6gLJDW2hkZgfXqPPPqP0u5rFeQkYxLAta
4Vw2lCs9rL7qxgyg2p2RpIAP5WLcXRg54VEM9zhi+mUMB7EpNjy+WV6CFMu4NOtYSeftp8yKXfnQ
mbN/VM1pGfqMTwAJiBTseocXP3+otCqeDAfbzWsZNOxe35VOTToFp/imq6+gc6D4WE3OClwIy0XN
xYTl0JmVhPWrgPxwxfkzf56qQgXy+pUrGzhf8RsSJQDWtdQ18t35trIZSCt6M9YkAMQJ+J25l6OT
N90xsSY5f4A5B/uZqEZzx8NcCKmM4OMWuqW4DScDTkP5NUl7zR/wxjceFSSg3wJdH5v1j+ZP32fx
GgbSmYr5rcJy43FRC9Wp4yVvXnjD7TfX8xz/lxHNErJRW6QsOmGhlVtST77DmxJ5ZTBzHpIpvYAl
Lu7yxAD5MedyNmYWmxU/CK03EJkxdSug/V5hsA4/fxoxukR1OvvRmvWYwr1in0vOKAtoR3tpDs35
EKHyxyncxh0YY7NwWSUKbuhCV/ippzZ1HFVkjyp7VgSo9o3KdLC46yXw3Yalc6IXkYr+b8O68EQf
5iG3SZTMNU/AX1Hf8jvjHKtOYqIlHqhl3WyxAJFp9c87NvNKR/ZoxHcS3zmLqO3TEhu536uxmGub
18SXA043axJLnQUlZcxXFYvD4i605Fc0LHfLUNjapAGwfgu6e9nbm6G8HJCBMyRHNr7hNmVqD2A1
1vTxW34c1IXlffc0ZVDlnuhsJt1iItyBggzME9HrMcwXz3EvZkLuj2KNrG9klGLBBo9Dyjwduxs+
Tr029Zosro/tkE9siFgvm14eNLCXY/DHQqVzgKShgr8Gkbmw+iYCduFrEdOBGk6Ay5Fi6fleJC+8
VhJJVwvQk7ji4wC+VEN2gLUgPgc49eoXYUr5QqTNzym0VxTKb12HKCZh4+vORWXojQnHgtS2aoMS
hdbCyYy23ppmLW43QKfPo+v9bjPYwwCrYf4hTvSnSQLoBv1pyDebQinROTEz6vy1YrMIzY69MYIk
yfhFJZJa3jfne/5Z6kyZxHBwiAZPidP1ci1gFxDlypNIYWAeVSfWfeceIolze2f/i24raDftCdtk
gvQZ5vCp7dh5daWlRByNS0KCWVL6cpHhQ7n9E+Yulfv0P7dws5bnn+cbznRuHZr4WZ+Zos4Ir+Jo
nobV4o3MmAvMn6Yi5JShK2/LALT9K0ZiX4kRh3NlI84dII/YETUkMjtn2YrQ9lT0XT9C7WunUwEx
fh40PvYsxEK/2NpV8r6ksO5cYjPXPYj/NhnNzvQWsCMs+HjQDib8YJ1rmd6TO/lueeSkrARvSZeb
+20RVCKH1Bz7d7umY74XMngV3T1xBfOpC+CA/HHecA3GEoQkmROLt8tM6cQWMfq8ceyWKxlsutnS
H1glSTK1eM+1D3QFZshDuyH+yA4vdxd1XZMztqYt634m356FO/Fv7YMm3lerK9+nzZzkuOERQOcK
qIkJraKqr0dbghaWzaRnE9Ym37atrZXZrWHb10hqYfA+FSTVYD7BOF7gWtq698CWDczBK/Zqxhyi
eaZMyKq/Qu6VB8atgL2+/BQMveamnaB+IcpciD3QGfmGrM0cJ6lK4JNtSlC7JTXPFYcVNmIfsaJW
7a0lHZlqZI3dUyT1lVWKs2Yr0xE7BiVZw4yfLn9ciSDAes8L0w1zr0D6ddWdTUv+SSVcnxTQ7bxI
3/MFSvwfRsxtlL8DhEFSqmiN0pvwY1UwqaZ3TCkUiagWrt8axTT/1HcXwYTYzZAueeaqGyKptbyk
CWvB2ILR5j1hRBkolap25wpUjsjbNiXJUZAb6wYRynkdDZAMosH5rY9jJ3oZ9bRGwLc3Gt4sdbrS
vRZCZNZRlWH6EpU1V3u4dcpdGzmdZINgc4dSdW/AGi9IKjwWZngXBn66tdRs/pc5caK1Y9PSAqv5
jb8hy2Rv8Tb2zn2p6c+OLmUqtw+iUZ3L6voUvRCNknP7bJ79mnu+FdVvigeereAkE12iTXjHCK6i
MZV7nVR51Q0gFkPNNt0kU0dhEtfB1lZa0FKnWayfvWFPvbHDPnUjMScd3O/KrVKDlj3V3eDaLRGw
kJ520QeUuhG0OqgR5pXJpiAtmSgReMvy155LfEctVPc3WHSnCvbPyYTZXutyjlyiBLYWPRD+k1M8
IMy+a0dxIRolTlQHo9M8acxc0w33tFwgw+eojQ3el6EYl+tym6cRLLEosWzRtlkpULN1WNOSB6QH
bU+18CMPcRd8hceiPxdXowVheOYQx5Oy2oe6pPasNFns/IyyiWlylWg7x7d9CWlvkDA9TTFPO6xX
wU21iMMitZsXmLP3r4yxUgBp2gUIuNPlhvQGVg8KK/Lr+Zd0YLcsOLhHlfahR1P9FobZs5UoFdGw
OaqG2WfeF7w9rrIpmTe/pGF3LsydKpJUpc0kGEv5DadtuQk4UIFW3XvjFgUX16cwjzB2P//8L32j
kvnogm2UFxIkF3SjjmBrtAPtFq5B4CYi5/6Vqqa9kMU+TdbF64elkOaimqXHUJhMcvtZI3rZIQ11
dZ4ej2b7Owu2AmvBRs5dRkqB+VtnRiUwdVhaoNkOuocH1Quy6EkviQf0ykkhunjWAxG45tOwroHK
Uq/pf4xaQfDu0zjJlpu3L9vAc5CtyoLzoglHRTugtLLiOh3NCAGTvasNMAJlX5kI58fqpQNt52KH
LjSVfKYSkPPJ8YqlFF0l9Mj/wiSDpPFi3ovhnnXGGZS/7/jeFE12bcnampHCbKJdBkJrhb8fCCkk
OdjOEualTsiG6kZp24IzAZNgNlKWFglGkZbWOV6JHLKf7EI8yMgNVlOTB1iyJjwsADXsrxy7erti
6aAq/3mhqkbCTAKW1YU4qjFXj5Be1hlXh70KLVdVD3Bm7U29VPxv+tU6SJntg0/XwfxOxC6XgUCs
nM7s6Ddvv6HfyqkXmbOGxjc5edhTuWjQHgo6sH/PUHZqtl2aVliSNaLRMvNf1mM/QBXkJ9tI2fmA
68+waHazpqqizSEqhxS4KUpHnq1elcbNC3URwApv5nSUzsp8K7gFIsrIJQqZ1M2Jtt3Sgl2zQ33A
puDhd7Lv4YU2noX+VfuJfXhSNjG52ohJvvNLYNQVYaXYBoMICo94+zeKmlzpIuKD/P88mH142ScM
ZvxLI6sHt80O2ZKraYL0zJC5AG9Ej8LjAwCx9rDjkE0cdwNG6+WkFREc2HPCXa5UtrQdKHZEvNl4
MR1agMTKLBN+Ok2OctOjYrihL3EwN8vvzBk/5Z4Pda+yXd2puELSd1j8Uho7hIe9BcSlyYu8KiXe
vSCD6ilvK33751vHxbvXwhm6PlnQnQXpXYXZ3d6q2rYDsN3sYDUUSQWD05cbHX3qcPob9QKe9mVz
vvttQo5TuY63V9pK6KAZs63pwfXGB/wBGdbILzSqJOAkFcS2yZpl9AdEeAA7zU4oHxFN2CkSkOg/
qFbfWWmBJeEX/KJc4CUaFz1oPGO6FVV7LP9O/rG1qCgNdE7dRsrcDCNwcHYjhi7S1pwC5h7aYsMd
639fzC/MoWTMRhtsswXEs2EBRbuWlH0PtqLedybB3l9bPtU9XrDHunZYzW43vufp0zKft1y9pUar
xF+OU+161kDAmGFmdvC1QBNvbtlCSffhKWUsurDjoJyGU604G04bPN50aoQXNEdbm3Y5az8/hS6G
/86CasqF86zyKhIBw/JUGO0ZTgXqlWicsFCJG5/8UwceI3PGgFbXPA7YrAc55/6yK0wPispDp5Se
193D649MD7AykLEeIG0RFv5jB4jPtSaUYjfbUHcu/oH3BEmHofe6BucTz4QRjfKSIXeBv9QGSxuP
eJI4bd1Q4zE/ETGpPv+l7izKKg+4PENX4WZ3rB9fWm6/C1ocLGls7Arx+lF8bVNk1nOfeSPW/bnE
UfdrMH6G7DL6C3t1uTl8iImXhCfscqMWl10FEsjSmUt7qwklZCviUQWANpZcMvH6ZrboFYV9JxzF
+T7wVSnxcGQHHJrtgaAWC2ciYoq6ablbBMljpKqyEVGCi/yuBONAyn+Ap1avVtQ3sTQv24O48UqY
RqJ3+ZCkyt/Xv6peR5FuGg/0KoTRyerkN1R+K4mjgNsuVEUMa1aHUBkpAaZVMyX0/+kjeMdkJV0d
mon0a6P9SwRlcPKOzNfV8G2XW9gVhbLLhItaOP6DXAYW7Z6Vvomkchxq3CKCdogTHBnMYbf3B59y
GA6ejchgzY6Mu4tLJSGApfuA58HYhNRXs0InArCAO5VSsqXvzFjGa/1P6d/tBpe+uUX8g59dY/Tn
bRA1hnmdPfsKxkHldxZ+VYWj9eoABmXZngSPwbE6IPu7dBR2Xrfu4VoLDlpfgrH8uCdsq1BB6aec
/bHOBpnrM1anNHBqoTXgaStZEqo1eM6HjajJPCC9iH6+ew3svPODmpovxEnjwTd+2EfYw1j/d+i8
VMZigxg2O3UGwjCFvwyoBif+elItZmHRs6oLg09NxfC+hZiY99pjmRzBZl+kYRsfKrZRaASToWkj
6QUQFm8Hmr2NymzN5U8CuE4LR25lQAbaY8FRie1pskwGOl+Jx4KkaQcitsloCshDkGHXBrXGAagT
C0jNTH/R3J5jWYNYP80OXKdhLn1xFC50/xlqd+jZuKqVxY3Ip+leD8o9NQ+QKDZSxdcXnWJ1qpX3
zNrMj5XtpCzCPnqgnq4+ENdDdjeZvhn4ILGl6I99gqaPVLbHdJGUYf+z+hOwA3Ci/DD/SXMpjfdx
p3UbP6eGrwqIVOWda24bTD/2QthOGHR631YLLdlCFCrYtIw8ApdsRUmQMCFypCmCIC6XXtCh6rM9
zm2MJlISJybghWM0X5e/mxt2CkAZeFqukug3Qr+9rdsbi4OfWMshXIA/jZB9nP7n+8ORIxo70TSg
QFSMdtJRTvw8L4A6oZgEmcyBrn30Y+t4UbmHl7Oe6Ubez3hj4uaq1uf615at6ZqOIPkUfB4rw1Qg
lzIkYSTyq5OGCcVDshf31tLnMU2dzbtHwEboyrYohcPRD6KsPqVoR4Rx+kTwKsrcfeLvQFZYVujd
gpI8Janh2uVOyDA+/TMVHQ+xirV3NmSzGvmSYj3P/jozFV7eRasE6Z3MKoaC99M1PREl/CMYlhsG
dGP5aKhPmCkV57WScW3/SXAvCxbeXbjUWKstzH3ifEl96epXWfZcw+xB5qD7ztPkcpVpxcKWK135
OpfiCAIGKVdft0WTP74qHRFdCRaiZrWbcTWJfo1e5ElMczZ/209BvyiY5GmpP0oczSgmgZg4Xr+z
wa2K/eTJ3edK00HmRw/EQC8XNruXMPc3R8f+oBIu5MMCW293QVnNGsKoH4Pb+H8Dx0rlRP9elwwi
Z25FsbuN86AvezU1iWGYdcqIVsWnv4+Mf8ts4+iuxij9O0Bw1pfOVEIsV9bmvFlPMmZXqJGbkpbT
UbC/4smEoSum1jq2bxvXtawPKo27m0lvq4aGlj0HtJW8EImaiw6FkcYS9mAIyVX3nY+rhBPYM/Rl
b+gnuqbML8iUHya8vMci4UuTslP/Yqpi/Lpop6YcF6lRu1yFeZY2s1z0pcQhM7H0S7UYOFcE7CD7
L36kRHS8tVGQMeMKbXHIN3JEtHjsABKBtRYVfmVzC3TG1HqHp/fqbQE2oS6ot0BLZod9VP9CpI1F
3j4IhckT3uMAGX20dPSZF7iZs3CFgiX3RaVEvsVpYVOubMkIouIOw8OTSGtoqNaZhPHrOg+HXH9M
CVN7brCehHXaXwXGiNcLc15dVFPlS+UC1UN9CWMTW4vxgfyhv5uNnjwKaYfL26KMndnt6SiqirrB
XSFiVbb0G7IgfRI67ZtLv090JKgzkV6PaWyMyRjb9jmdmOurxSPJaarZ27wNyrnotgEB1bFHL2ft
3ZtIQxC/OCskE0H1jUDIkGa/aTmpjSuIbc2nY5EP472raYjDEjJhdM6dUUFx8JxNiqu2PF83+is1
ICfNdZCGXWB6raNFvwm1Sy6qoBb4wPTo0Ytx8olrmYt/etyJXCTLN+8++yO4miHoIVHDEU6zXXUV
CHXnkEOcAJLtEeJODxOZsoambKnK/tC6D/DRk+uLdIs46nbIMKj9iRN0U7kEpZqnzQX2iLXnKeJu
8udyw89ADaouSsG8xsu21gnYdDIfsw5xc7UPgKiY6nswhmU6h9z0pPh+Q1V0WkTEX9Z9QKTzYyNd
fG3gaOhVtsz8uiJ39RGOIxWCngCyVuVDGy/Mvnqda4K08xGdDgrapAuIbxFQ4ZViohkaWOnUCSej
PnuxN00a2p9ievCnDs2b3tYyTMUdh6MfE0u3fQSCT5oxA7o3yFDa+Ze4Oi4ygsY0pP7NV8ezEZ/M
ox4Z0mt5OKNKstJ4YytWvSIWZYYEldvgdndd5I64NJ4B7Of1uLqAc4x3pXesteqRog5lImg+5RwE
NhbLWr3CYs/yl91gDqwvh+N4c2SEXdmb1Zv+BlnuP8UDQ7dHCyO++bjxCCaenyNe05o3MSy/ZXzJ
fS3vowJFA1yFBV83auiRQ4s0gmYkOQ/Pz5Zk/BanTdxPEN3d/A3CtITPmfIuKFZurSaTF6YxA+6X
tqG62qOSy+6aQ8A1yKTRCEc9Gm1OmsKx/GLMJzAv8OU2xAglYHIQDC46dIpIAq++vuSTwZbW+pU3
+Blk1KF/BXKkv6al4wUx3iR0J2Tx9vgNYftIDTIo/8sEdj7uMiWt+MapVcTmqxQj+oXWRRNnO7uw
DrVA6b8g+TNkG1fEEOIaRL1fEEL1i0lvrldKaPXTabx/ew7jzeVLLSXvLbLJVKLqq3RFl26/pRKw
VpglQz8PyfgWQfBV9Xwbd/j7jZn5tvFioqpJjNF+dL1WNh+fzLQF5NJV9YTQTvIsT0ExuWogf69k
hRrfYHyiVya7aFH4FYBZJiG50KB7flZXbA3N9red1JeXjCw1BiS6vRG4IVSNeGLkhwyMrQuLpqkj
D2qbNWdnI0bFC6Vv2dNu6lOpG6Y/kt7ZnA+g0rMrLR+GRDp3l1MmfddhTMmTEstIvRRon5/MUkqT
vSjrq00ThLCu/u7dUBQN0pt8dAueIQZrzLzrqu7HFZWrniiKK7Pk9mHECoA+F1Qr0XSlmbMtfvqn
Km84Ro+11YZE+6r8epZTmvNDlErQCgi/2aNEA5JimsqsLRoedKXane1edKnafLgeIsneeCZKq3ck
xD/0OkP3LlgfaEtTxcq18ToAlv99QlV20XwYutUR2qU4xniX1KewjuCLH4BNrevratOSZtOwrIKp
kriVR7ODE0X19qfhmoDU4Smbt8kWQk1K8SUObU48PT9ffNLeB2l/VUWVXH22llYuOr96NmgNLM6q
FtoTZXaLQmgI71mV67qd3LlFtQCrAmMvtNK5XfI92tSjPePbvtJmpuvc6Qr8VuLZ/eCWqOGUhMWe
bhNbx3GyY7DqGbtntWjPTs1GOB4LvF+KQZmn67wZoNQ5AvCqe7r+KTopAcg4kv3q9l1YmfkNVq7L
dlV7OZVdcQichVG/vzD6WxuInXwrWEpgm9KMBS85/ZooMg735uCSUB5cIeAQdmhKFFMKvYbHPAm/
Oc5OQzEVToqYq+aiiHoz0nwRy9sijoOGOKEW2SG+FqxTR88O+5M9ohBfMDj2SSe1QfUIqOCG+SL1
NyLn5/RIRToUhZLOGuK88cycJxUpxUBEy++I1SL27fICAPIkn/lRiptrvy3DQc1lPKS9dxsIWy8i
auwG6yDFcRNpwL3RDmLCXsSDeuKv1tmDmX3TZQRCAWyto/uHYAFi+43uxKwZoCIVIFcSzktuWZW5
1tjIfo4yxb0akGh1isY6XiwXnAOznjg17dgMvR1mBzE7/mEALAtgeMJxqMndAnKC5SkNKr91poDf
GjiPphqn+Zp/2uB+lAjp7HV3uxLU2WtsN93/sLBDgvaF+llTy/8iY5cZtm8ByIVxGHXPv3WNr+s6
KdT4hU3goS0b3QG1l7PAn/M2oXcZniWCMeJm50LyuwAPGyd1Uknvt8AIJE67vJdc5O2u7exHHMuM
HVxnwhy3KTHxcs1DQVuj8fgyf81drZavUzPy+9ByOXg57vVM3l2oAy82TV78k/qrhUJv6i3EyN5o
Zu8oxRaTLFUPAvLrD6YBETI8SA1JmBzgO1LLB9WxXucxxyp6TwuUpiC3BT4t8Vtuyp9hSsuQ75pS
hJPFWMAUNTp8P2xY1U6gaCdlJUDDz3lX3WnFAv4OE5sLECx3qnzocXSnSSgmr7wxfO7bfZum2XK8
9pRFWVe2CRJRK930II+x5EidHFbFGRhx8UMdrz1XsDMbHzciaTaGJSUEnVX+XDezhYRwxChD5sXZ
dBLiV1cKDCBkbvCyHFmI/lQ30qqbe3v5WJn6Rfn8MrqO71hfyfxx1WjYfZEdRPU6ELHt9iZ0fFXs
/TAwugFn58e7L2OLPTXAVTzonTIY2A43dSuRcz3MRACJAvdxk4duDxTrA8dqaXCeVPvsqpjX2xlg
d3xktoMPhkKrni6IFjEisEYhEawZESYa8KcaEU4V8GLGQ73L8cEYO+IVKL/deIyZCxKBmGlvExN8
E/Hef1y5wDzFgfv4OzOary6YATPRvgJRy6/kxmqHtxQ0SnnbeQgfuYjenvohkIvatmpubGWfLcU2
GedaYxRLLij6Lsa3v9QCM/SaLQlx4O9tvGfkOnZHL8ahQjbfXIJLY9FWF0tdQAzPSf3OU0K+4T14
Kr7r38YfC3k8bAXtnvBwbUBDgkY7QYQS37fMsDo4jV9l+/n49J9tjnCIOvr5SV+5+g5xLd/rHWxF
pm7FCEC1KoQID0FoLMBf/F2bJyC4Qq2DUkgvGC4IVSWLp+WAODYvmFVjLQ1l3swvaeU2201OLe/s
MUXlr2BuI4fJLYarGbHzN41Uh1tfl5KC2OVVHE90hPFi9dXv4VRwmmEebYZuzAiwCS9htVYU3Tp2
Fy4v3VUY+2RHGS+i5GCN+AZEUlSButBChx+VZYIqiKYqGkBvnNqrN1T4HU9CoCq0luUZatA81Db9
mSWbJE1o63OXGpUxE0HZPKyRfAOZowPUwwrYotEYmeYPHWlrqWyp5TtOEdFd4LwBTqCmoE4oebb3
NFUgDD7Daom6QOZBheSsKYmk3nuxkmsC+wPBgUhMrfccroYhStSGSP9Cn3cXXDcp/0witnhojW2G
SeCnxX2aa+1PjRRGcswSPea9CFNTEdAZWT2RZFHpa83U+CjkuvIk1UQmxqngSEAWqC9tlgzSGaqB
MkRXv1aNECXAv1n8MxpqQ1EJ4FJ7xNwM2Bg23ooVr2oQYiimJE5OBOyx9V5x65zUEYTxNNVCrjbf
+iwjHcP19sFfDkYlF+YoeYmKwTn1YqXTrZfu3AI8A0FH3n1PNASKqWnFouLZ+427o1NknZHrRbOg
n89/CX0kSICrCa9hfrg+zMI+j7ka4lRKpkBeAmVp2h7D3swfwoABwJkTtoLq8XltmAE2Ac2Xs1+w
xhYvOEYBs0wSs3DBWn7OqATr3EQXL+fQD9j2SqX9TE5dKgY2ml018wcvvBa6cRwEmsyHUSzoAlDB
hBzTjgXiEiyk75JK/P9MAk18lEA2+gG31miwWEjjCsGKbGJAl+z8343lXa4SyNQTr9Ote9w5tzyu
oi+d4v+UN8L6e0+I/YjuKaQadRwUtJfWrRCWVjlEdevOjyOD+cJlORFzQpYn8vTUv2J18rgkX16f
RYaoYE5dKeE5TB3wgoid+JOPMlkryyOoJycNUXSm8bvop+cAjefsCZVEolL+i93UQV5ADsKjT1mu
NRVEp8vNn9i6Uu14ll5ENY89m3/FS2IaKkdjXJ3PONhJCbQ06MxkH6pCJ2VhINp4p4Qum+lJ+Uzq
nMnu188WACeQxD8/eSH7h4b3UzPpvFYXXoxCdGGL9RcegE0dA9QQOLydeJffEEVuHmZucXdSkQ31
2u+zLXVhRhDV8wdxkdAqRwuiQxAowarQn/MzCt4lbvr0xEeEtKHJ650tSCFQI7C8m1MEjkc4/U3a
6OwshKPQl6coPl+6HngxJe+WD5Wvvs8oFunu7daYf/ziTaDs6bG1yDJJ7ra5GRyDYcFDUOGdqAvk
pGXWmdVcTaHbzCiqitDx0PXhMpnoyd4gqSNj+oyQ2aqbjCDkNBq+PN/CIxrsbPES488cicwJoGP0
YV0SKWY6XT1IofFyjkOOFWydPOXCuJ8XgUmfDlbq9lpNPY+QQt8zDRQuDWEsaQMRDrunmNohK74y
ATVQ08Vg0kfumCOz5v7C7PybDHIhD3JX5OIiipy79juP0++MwRNsCl712ZSCvgZ+tgRdPNEEsUWe
Uc0s/8Yrw5hP75mK9ITOmxhrrnviC6hjgmQptQxHVgl8PWAMFZPTdB6N9lrWVgsqWmOw2Hs6b8YX
M1lMvTM6ryPgP9l2V1Mn+zHv0Vo1YPkig2yie8r1FiN/5lhG826Jb7ttCqXcbotU8RX7XUD0M40N
8RVD+/sl0756wTD3PcVbOyW2ypwyxvQOWYcmOPLiuoBZxPGbvd/KHMvPEH20wXYCbC4Hg9Gi6Tha
U1RsxP61grL6w4jH9qSsldiQhSCELN3DPYsoZ+DQVKqTpQD+Ne53O9a1FzGA4pBvgpG1cZ030JDn
/n0yW4GOVJPfHEtiIT1qDpU2NsODzxS5Jz5u7BHAJN4o898r5ErC8saaD3IPddAvigETbICazFMw
PJdnLGDosVtA6/vQgQu4HOiR0tBQRz+2bdNwLlzLo4Ouet0ZDQSAOOmIeRc7Vui+pyooka/0Y0+n
hpuxsj+Ec1SYmTXPtLSqagBfAE2D6sFma/2hUCU5MAgq6hcmutrnn7Gu8KBUCbDsrJoLE6UAq4nm
yfyyYh0BA0g9WdLzYa2pgEpoQd9ebcJF5BAH+U9guxy4RoYAz90VuefkIK8IkWe9Z3RU7+FqmQZ0
Vv15F9cSQO5wu0fKiIRTQuekzy+VNjYHkpoHZ31X80geSNMkiYSsxe6ODBJxQ456ZVcz+S2j9Zbs
UfIVGMqMYYAUIUigqWJU8+lv9ASfEjjEldOnTEsmn2aPRNilQY5O6afu0I7G9Aqm9FCRA5YqEBfO
Hr/PoSS0XtBfVJTNgNDEEmoQcijOEkYy5kcwCAeOLAul9gsUpHsRkIePBLPWNxNFOJ0H237vhego
WaIf+xWH82FvC1Z0LomPSgt2wcfpEu3AXNBh92ctp/I0Ul81GSU72tyuWOPqll1nTxk9thTU4R7H
JiZxSEFdxrwhu2EMRj9mkvIKZ9CKebfAj5utlSQttUUf5acuB7dqDtF0K3twZDGlYVX18b0oJ6zc
YbEogANekMYKJyAxxQqTrePNgRzkvDUMPs6LU4MaiuFC2mKbFr48kj+BXQ3NpDkk8ZRVafITrWwg
iZ4WnwF/63HfUsthryDIKbcdphWBFEuIHTjl04svq/16bZ1H0GlQGM/17rIy7ijxy95Tl0T+u7ub
zlL7ivKUW2weX1yfH0HUtuucrRPfrtrQCWang5Ah62J69i8viJ5u9g6FdDU+DzXjCLobD3V9YEWf
nbgxaHg0PYcSp7/JwquW8ur/m8jUYBkiPLDmW8zXq36ddSat+yMZHcp+V328+gcsk53dzdKnE0mR
LoJl/XoXmIltvusLRfWgP5mH7H3Tlt1rwY05VBfWp1EHfu4Qt/K1fi+EWday3dVnR4sQKUg9rQ1g
fR43lWCIA2qeRZy+18Ozvjs+qIVQElQzeP+8fZ7r8lbla4z8AJkRZcR6XqH8hZ9GmXema0LB6fro
9X7PC4KWxC9LDEob4ZvmPIrLrYhawbZLI0f6f6fGKU4mS0+DJUhnKCqde4kO8+iH7Tyh9ges9LFW
L+2o2z/OMdOYnmum7CyCuWFs3oo/FM6Z5EewzADXl3CAsXZETfWQzOh64v2HZxkvHclJx/SCA8ap
E4yJj0TO18g7YAFDfDGjCRQofHuSVX0Ae9raSC3PEz0Mh6hT720icQt8qldOZtfLYIu1KzKB4zM2
1tfxFW2sbYh7jF8g32pag21cZNfyBeKs/V35llXaoeVdt4tqlVnDU2p4SHHokrhWZhSUvSBs0ep1
i6TEHwF56CjDYK9i6yVPG+KdIylRSSJMAwFg+KwPrV66OjfYNC+TmhYr5qIWZ/LqByQ3ypQY0GLn
arS4lShKpe1mZ7KGLLboU3Ev2WKkQRg3G2XCdxvCqFYd0RAJ6x4u8O5jNUFOatg7kx2l0bngdtXm
dwB6zcT1GdVwrYS26gzIVrSadCWYMTbQTMXsobnmRtV5/fyz5QP4VkgjsmqMp0StTK68ruLVtgMv
XL0xbKKSlfpBfqFbLhRZkTN6BwEcEzdiCa4tuL1AF7+q6rDHfj9DmeQun1yePrdkCPGY/okp2q9x
7B9io/ImrnE/+A8mrT1eFSfSSYPXm/Jzsw9f4ZLHnuslzchsTrg/xV7h2XvCvPMYgB+usGxnlPVy
HBK/Ety5S5J6hPKykYC6i6bRBKK+JN2D2Awmv3vAW/AYi0L7ZWWfTdliAJ+zFZ1mcldl91wVp50G
CRSQrgf+ry3ej2S7siJVUrCkQMeg3FC4J0UqNWGgwW+Nh7afFnO7RCnrR8qTtpA1yn2ZyT9AGKGJ
OuAeJLwqGkiK5AsLkSzOMGx/wsjTmfFLxHOacCQDta5gLQS4FTEie5vf0Ul8KvK7v8N1UrEKGEip
xDqLUtwvTlitQO+1kKWDplpc5VulUTGoDHYsrXbbZbBxDWFFVjT1u0uUEZBzQRLx97u2a+wo4HsL
XGqX3bOfmGBeK0IROpfogWqE1PwB5qU5tMEaEkdGp7LqxbmF/kKfB0cvlNyEzH1L0L9qLkolyfh6
mHEv65jpQMh6h1gEslLSApyxboxIQn5gwfutuZYhQAViMHjQxmWxecEU0gpRjR3lmF1s+Zs1ncQE
kdg0bnJv9xzg2wRxbbnv4Gdn2gfR6N/Le0ja/It7b2TB9ofoHVjxdz/wvY+EiQtv8B5ezuF5FM2r
oR8ShDBtwptuCjuXh4ChaEi/VpaHGGDKGc6f3ckFAZb/XXVmni+y529WVXlzs66bZv2crzAms0ZH
q5KTMtwWR3NuSemCCHt91SCBgrQhxdtTGuEB8Sd8j7hYXf5X/XH4frF5GW1lHNDJY3lBUpxqmkiv
E80t1xhP9oIa5BqCwx8TladzaW0aY7iiWHmuwx2ADgH0/jxV9ka7ZSkJYnQ6nn569BOcKIve8DLu
31+tFsW6dCLvaOXAw9O7WAWQObZSbgBRnKPkZwiUlKEw0jvbZDZCFHYo7ejET84IGb4jMTCSS4Tl
BQ0KFiabIIcdjSVr9CMQlEInu4H1wPEu4YOECHplr98A35pwrqUEtdDuWmp8cdbBqB1Ov26nQOGM
kkXmc7hVIpdZMMUSsZAYVuNbWoeytcSHMQYzyrrjWD0RDyhkzcmgqLQgBnUzMQehlR5m+ZvvjTr2
cl5K22/3WdxltP42yIAvNN6/gctMxniBC+Ui8TnVf9Eg+kEOaoG7891TDAPYcy6Dcwas2vk/TgBk
486CzhrbmsFmZqHNein15gXhebn4NjnDLCoO7I1Re19hKtr8KfNXYQ5hSUHliDQ8P3ZYOY9k+9mD
4PcdthNKgQtyYhy0nXB0NsbpZLFY3FbtOlTNOBnF7utZIS58dUrFrF6Wy2RqnG65UVUw9ti/TaZF
ouqMusisByqoaWMl0BC6YLRz40YNi3t/D8CMhCBuWB9NuGp5RKyHZIRHjWeOOupP2ETP9j4eHGgm
Ohr3L0rtqoc0dqPuFwi3vEaz/fy/S/6KVZgR71C7cPZmOrTfdh9VtV2ptQdDDuYsWmyZQ3XOCyJb
ARCuTwA5tdI+CZ7zTrE9PmmSd7Eigx53gWdUK8xhbOoASE5xAWtEJ1T+60eFkUpeh0rX1FV1orVN
iW4D8SYhMnUN6RUkz7alEPmQIlqNuURg799BKMtzzs3C454YIjOl0kBDidXCbtoMsj/XfI9FZi5/
oj7GElEmtUTG3enACmr+cChK71OI3xS3XjJ5TzF1EYmWKMSuxLfeH9fdya5n5ABKSHj7bILhdN/Y
L9Ge74zi1QH6YwgPM6Y+OkDd58Q6lV8iz1SJ3DvGbdMR8h1RR7DasafyblXuDhURNUEJV4H3M+vT
SSwT7TBTuaqecwtd91l5E5p8DAzXI2r2E62JCc0g+dveuXZ2XIbv95pPF5BRBBsUdh1eJAb8QRyg
mqZTrc78dboMfwz0L4Q2ZkEDq4FOcC1jORRuu3Ca3cb2pn6rk1W9EHgfc/QuPhXsdkzbRNV9AgzL
za9gtU4Q6iGcxDg3rCidHimQYhR5YF90iszf3Ygyd2ffLcatMmvdEnOSomNHYdIKNw7zZt6Epjol
uCEWKNVM3duG1ILODQcHP+sjQFNwyzD8imON5M8qKLBOk+6BCs/rr2p4p2iWvzgZIYrnO1G+VHr6
dAo+hVlSdXIVh1Es55RZ8ZlvSJl+oqREYzFRynnWXz2P0/vyjoPP/WJT4ninN72/stmCCROB7xnZ
oPg66r2lCNsudXXjAVNAvtfd94fe0b6lDyEOUWuoLbMfGcnnBaLro2MU3E6eItYzzTydDTo47YR8
VLAVV78inxYHhdBaZ73F/zSs3v8gGDWKD8C5ANclq+42dfnoBKG7izowP730kkQthRcUpcpXkhnL
Uuj2fZfa55WBGCgfF/Xy3eCich0maAt/qXZDpMX96r4EYJSpzXzjGJF7zrys9lTuIl45yAekA/ur
l7HJ28Cp3vlKpdawaQDGLu5IPRKmLL/i1iTf+XfMin9jcIpu//Xg5KRavedBfxhxeOHqPP7k2C9Q
Uu48qkvTFk0wheLsGvXpHCxuE/Ub1vYeKGo53Shnpq8Y0nIiWVns96jFUJHGrmnnJm6RmFP57t4Q
oNGUtZYNoUOOlfZE51yncCQqkf07jXWu9pvy/hzSmec7/biVUxD6yvw7gLV3EGY2t+0Otpq6NObz
QZE88bR6F0omzjxJV5xnQVYowB5JpA60cA4X0rUpgUPeh1RF8rAvmdlD5mbjKRO4IGLNJ3sOgxcF
fSS61vlmi8kPLxAZVgEGFm5TUkC8O0iN3nD6GDhuKTLPdG0aATJi/Pq2nFVTwZrTgH4yk6F4ymOC
NrFU+WiWz9nnM8MxUiD5OruAuvnn9sLStGiN+wEUifnEb3dtK5t5CAvsjyktcsZthIgafeNCPtdy
NAWjL6l7ZjjkdD9EnRLjX4VdUPvHWlqRPjwMNmaK49AR3Jdoax4MFvKS8LElPQ4e/lONCIPkOSJb
3xEHkXmzkgp2GaOVhyjLSpLoVpSXolWhH4Z1diWV7KlPtgre2fczD9CxbKDyE6O+Ligs6XTktPcn
T3VJT1i9CSdllnuRYny+NO7gNxYQPllo2uRMVlWB/5EMGEyKvR7vkaRKsJlKpEu+vuQr82KX/h8f
CRA2091skx9ZNyAGUBDoaGcPVXx21IxyGb5bx7EqldsqtehZd2sHqnQuqQbpCutqPfJ4jL/J+r/R
dgKq12nB4M/ZCLShroOWP66NNui8+sZNJrjO9vW3SF+BOeHAyoFMSBpRAWWqoWvtP6EKEsx+7Cun
SCxrmgIOQGmC1buWIdyQGVxRLQCopCr3V3YDmwXhQuy/0/rmXxFVOfAMHIXZ0vLA7XS21ScV16j3
pqRGWhUM/hjEmkSsdAiI6nOSVVoh9BXPoXVf22QQWuF1Jf3qpmYDwAF4sSCEylJEEClVoeS3tH60
m2IHYk+s1+VaZlBiXyOelv4o8cHdPnTE+odmKvfchxvvG9LAcVJMgwG6s9BcOLta/i0X3X3cuNlB
q9w/72sOF3CcC711GFlpKHRx3o1Nl8ac4CAeI1gYOmRy/3kdxiZeS7gbo01ifU3GvjmmqxiuCaer
+iMK4dxdOAbUS60RDOG/L4uzrFiRmqGnckLGJZmaahmgh0J4shz0EMGhWXAwGpmn0fHPUoG/ACP9
+kkqC0N8UmUXIRWMM0zPIpF5EDGhLhxLLIK8elYaT7BFXS3YTFy9s8sZ6myulELfJEmuEA/CYUoq
sXfWw2c76V9bYSQnBCcAV4cWeMIMY9/Nn8rwXv0SwFLtzh17VTXYsdx3warLYfJ03vcSHvijzTVe
Gi5AYBcFpqBQXhwJrMIe1cQSA2JsMVrL4VfCguEciSEvP0PVDTmfb580Cu8ZERM+JTC0L5feEtTB
kCrg5MdivoY78uaSpMigNi/DoMqbd663toT6ywwCquAfzfd9OnUHqKWTlOdtZfJJqz2gWcL6kNds
IBr7unnbZ5lZNDwE9I4vnJKrSh9/R+vx4xC4DOCj/TYUJYDQ26I4yRh1iKP2oUNSnq7I+E0LFb0d
RWOnOCWLEWM76PFTQqj4bjOsk8mDP9VWjIGEdSH6I2v3g5hPPws9gXGXRVI4u0bJfIm2CNJk7a0G
iqCpKxVhLMwh4p395d+WFmfEv+ev7bbWOeCgCqO57C/2HThJctRB9RvgvACqVpX7oVfGk6yz7waz
uPQueoXKPhQ5auAPLBxrr40KA3skX347z4cwfNDNAm/uH+HD2fneOI8iHPUQpXk4q28i+XKNot7s
TLxkWID0HqcUUYwtjJm13dPl1Po66LEwhJgJQfMiIxdsIjCGtXb/Svyz8XGBglSpVyja7OOjDOws
GTYScfAyqRQZ+ff9GNw4RqodkUQzReV3mxBY6HIg6Z4ME51E5GRfdYHaWJBT21xJ4Ce2kVTGWQFf
8x/aeePG65KS5EPDhtxppfkQkk4yCvUEhfDRd+3T8Qx1i/DugI8KCNS+0ohMKUeLjHnZiQYhpb2B
wZCfaDag7JY7/D6qy5qjRtLPRdj/LyrVg/LAZ7oktPZ+W3nyuZKcLIdTvmiWYXdWgB4hgL6UrkXa
WNekl8fwIhIEcJe7hQNvUXxL+adaA9rovNJSXEjauptioAdw9nSz+j2V2CRCdO+K0Bl1Koav6F2D
mXJFjzc5NN3F5fMlhBHJx5SxaliUxIkZZP0x1gKdu2xZLKsiP5K5Unx48SBIN0DddnXEM6de2p0K
CtpjL4Xv6likhGprXGmKplZiGChogMRSJhSu60ol6mcaSps8y45dv+vZuU/rRsuT94Hv2uzgCgP7
rMqNtjhi9+lFSDWx3yuA4kaKTbgfqxxrQBIvrUYyuOIs399Fvq9qquNMx3V784oE+bB9wkgxmg/t
tgJql7ReYDEjoGecFb8Fn/0NGoVZ+mDgmCFNzFJ0UKhkrtg2gX3MlhinlKP9P3o8CbtpGqpVq00H
sLvgMsMrkLkxqAh1ocPGK2HTYjb5+/fiwbyG95Nkae+WIZEaxl/+IlxHg5bJ9vBVe92GCL83cM1r
3iuyo0YnRBITfCSmoBzc6Y4n8PC1k9W2aLYkkiIzLDvMWpmDd0XTE1AGx9ZqTIwzBa1Jdop+zPay
gaTs+y505yKGukIrachwiy6MGC+zMCbqIXsCERm5jxRxyUOOlqqcWisfmKgU3pc2noCYHeSAfjW7
gUyd3esJlXHY52IV8Ow3VOOW2xDNNVSfE4TGcGpyJpvMloB//w5h/GdB/taoBlvwEZZ7sOXMkEYZ
piMdN44+3mVnF8BYIEeKnXMPdioGP4fzHPkqDjWsLQQl1+EMYoTFWI4HYESrdX/uSruF+qApMthb
LZLuBne0ScxsEm4pa/dI+Qvm/1g8lLergHzHLOCdLMYBJSg82fIkHfzl/I2KUvpojFG2d+KVP7SY
XD7bvUz0JiIJbv4SS49Mk9+rqLEVlwDqKapeFeBupje5lpKPqc0VC+pneuFzaG/XnwqhXwTNFzub
m7U/ceCP3uXlAVikoqadG1tmejijA/JLDf2mbXzdapxl4ctbRHJQdnpYK2TwUzsSeO1MpCiA6DPL
beaji96CdT+kVMETQ0AuXo9NB4Q0WeiBVYbzyIEnYKSyz++cAuUiKlBJdUFgC0riZoVnw0RGmT+J
bvoMHPzwzE6e6ASatZNqhvl/GzYHt1xNTIPrTo3CVjz2uWX+B2lFf8fyfWQF5vyUivUGYnQZgZAJ
aVNNnUBLd+eXLWGpx/NisCAHJRVk3TUQ3KF7iSZB0yok2oy2kMfnh8kvjt/aOJxnpF6eeWkn00TE
42OPLQA5rd99AtjlY5K/oL62NJTF6xw2/MlOuOBw1CmIniLfK5zsuCJdSKKi394k5kZ6PWKbCNaE
cedXhb2f6jxt7oXJJD25+GBTqkFesZUlOADor2Bd8QrdVl8bgHYbKfB+/C6wpA/N3ThFGpUvZd/v
I4q4WEqJLlaIUjTuY0vjqy0Ui1Qa3Ji5kVwNtFN+1QL59K/DedL8qCkkPym5znlpt4JQaJYTpfV1
tPbzGBuDh42ZVSFUbu8aIyhuHSV2BiLN79Ei7rdbC3iFtal5MxASWEIW/tIGoeZjBZSjSzIkMTl2
04rmmQ5hRLEaK8YSHFg04btxJa/yU323rkGrhJ3vWQ0vKUdjQmf/3nE4bVm2TVxEklFlQYOGFJoW
OmW2vF5yW36Jrlt7p4/dG6pWSvnLxkPsKDNzb7vgK9WxpT+1xQJF7GS6dSe/sftSluF6Xn+IXzKV
oeBW894sAXG3YI1eLSfecww2Ft44CQASECK1ZP52D/EIXSq8IyAmT5j3gw6dXh9IHc6br8de/iT9
um3b6HmJ60YTngTquWKunrPz5/qUX+AaET8I8E/lTH+lrGqfzSreWSyyX/biaCNdB7y9h+i3qCj6
sRqTUFRImyvf4u6r3q8+A5yULh40nMI0p7xLv75fjmwtbDPsltgfW9lc2vU7CnECQGxONO9KbMgI
DR2FYzh4MzI+whk82IujURUTW/6RAUsq+jtAuDbiG3IfkxmUfXbSXs6E2s52clOHZV8RDyrfws7x
oJn1RmSS7eGUM39e06UzETinFuZ8nJr5q0bzhvIEN2SZWgZhCnPh8gxR6wwfiLkOrLATGlA9U+1G
pSV8/TZkHHTp9fxE48r6hyYm+PwZwqo1ewsL//HBniv0entYQKpNcgJ6Erd0QKNaIi9vb6yzOoHq
S9EcMKwyDZTn7fP/Om5LlZbuAUCH5w4b0OBeEVULcKBNH9RMH7cPDREPJQmllSaPO0GKkSYD0f/e
+ZknokK6hvAm+2tj07RjAUQQX5pn1i9SAwMyZT0CpCL0eELG6Nex5fcpcLSOUGqTkWHqp8aAOgxq
QNFT80js9jmc08BcmM6ht0BWLBaGacoHGA1yFNxwbo7roh7j//jB90lOJXkJFIz2ejXntovLx6pm
R+RlNEzjOPCdCR0w7Uux3yBCsfZwlwsnr/hzqwE0NF00xybZ8yiau9XbC8IJud5FZUxyhEHfaeBL
q2i7hpyRUSzrbQGUuV9/7S1mLUa7NQ2/a2JJKmOr4F7NVgSjqDY+NBUfd80HLmsNKuuUmnf39SSv
Yz1gCpFrPfOSV/6Q4GQOxDxK/nnbsKSkt+ouXkfumOJVZgh1iW/pDwNZCbikEuKPduVOh2F8s11P
dk1ktVitl7YPFtcbRUyjyKJFZLy1Gl/EqqKiJl5GodHiu9sN8zYvpI+ft4K/AlDW0uzuKU1hs0Zt
S30pv6UTlJgUU8dklFD1ksG8BKIpm8kPUfmY7EGK+WshrBdHlsSS1A7edKe3/Yt7cwOca85ye/B9
gddA/QREb6qtkzMBnQCRbDZ2AcTpMz7Gui1gEOigHkpJ6VxAKAl0/7ES2HWtMqDLUCF8G0CQxPLd
BCXKXU34swJNiOfSV3v8g7HOKa4+3TIEBtssvJ1WCLQwNGPmyDG/37ebJM8+p9MXnanzfE3ikBYx
vPvCllCCHcfKQoUgPHIKGNmyUc1duE0CCGRAk22wDpRBW5/rAH8m080UOSgfEyThFGYaVfD1ZMg3
nzpZAnvnLSIK6zRuVh7zZEG+lp31VDZdiwMrsqbFAdKLhqaeEgtZN0mfZtyo4JQDLHzv9rV6m4T5
Td7i1VPRaKoTGZ2vGgavFa8kqeHRNgz6VplY/isuMdHN2T12WrSwqX2gN5VmX4Lqo1MX7J/wA2ti
inkUnlghuzdZ1C1PnIJO+Z1JePuQq7Tizmmo3rA9cPpoXRz506EjnAPZ6lthL6TDOmf21BY1zZIH
jpduXe4P8o8dg853EwJ/nXfLx9wWbfFb1vdxTG9arlh9I41WOkimJq8bHKxsboX+0+kWWrUnNvjs
rbdtiy/SWhYLvGehU+zP8rkeAtsARz9k2VpXJU4b/oUnSFzHvDevnEj23I1Qp743hUcwb8N2V21z
C/l8Ukd+1tU4X6Z8p7HX9KovXKvHSPf3HvTjW08bBQfvvYoDM4XqYxDBau/aEn0vnA8QAz5BGj+4
FBW2AqytDuLCFT4m1GK5yQ/D73CTLkfMeEmxvuSAcuirNi/7ge0nWZ8DEFSZyRgwc3/ZB7TyMcdl
VjZq8dCTdpx5WbIeogclhAW7VAOdy6PQRMi1lL29dgQFpDd6zzi9P38ph3kvsOferT5bGx91SeKE
iOsqzLtZume3nzyffPtNDxX+jgdwgSK5lhhQKJNnfdWFHFVVl2ZIiDDOPYgV3BsPWASCA1QGOMak
ka2M0+JA/NwqxD8wd+M5fvEUHTKsI3ggVO8NWrW9QsQPihhpiAPTAkdOgc6nhSDg5wWsMQSONJuP
3o057eXFr1PlGCtBPdqrSzoNQlQzSGzlcB5+Wjbbt5XPS6eXCuNT7pK8hQiLnLr66jf9hqvW7s2O
8awdKiIk3xG+9sfDt1SQNZ4Jk2vygmm1wFGRREim9mLWhSBuqYiQtSMa79CoRGGaAOXtCCmMClQ7
CkQfNNSbkwNCyRuC6z3Tr4Y/zOuAQsdmrN8N/wz2rrVMQDzHIuYuLRrUkTOj9zbjV/MhxeDXCHFr
0fqAREHy0Z7csBobf8FBLEQ4vV7oCsU5/z5Vy9PlVX1pu0mu09rpj5TwF45p4gLydgmOmsYisQq+
6FE2yuisMnRIM2x9Di5R24UQghW8f0ZSUc3/XaT06JKhVeivZ5UdX/zfDXkvALNlGR/Go0gyFwcM
UXM23vLm2YhwVj6Fj7uqNpScA9N596AFhP2PbjN5YGgHZGLU7RjwQ3gzdgKqulBu2mri+8tKvP68
zmu1Yq2iNeApwQOJHg8NMmYZkYqS8bXc0RFGG8Y1Y+EPO3YhR/QLnftLFCWOTdBs8ZRUIqlrncej
MmmBiAeKf7Oe9eCqPDY6EN0LCw+LBBOTQXVKgFHU9fnOKYz+0rO54bGyQZmDURX+10OVDUotR8nN
5gftwHAaBKP0ceHWDbmVveE/29/JcvZNFGKDh9nCGTu4u6sV8f5Iu0rY4RK59mLXOOdgv65lqdUr
W6mF9KmMMxA6hhmDMhlBNINBiZL8//VPqggfc0dfsOlUG9fKELvKH9aoskXTPUlVSPC0zell8wBw
cc9KVQb3ZKfDFpSRxQuvaH/psgkGSmLIOPcQIWbmXM07Kq/XSJGBixRzwjaOgg6WIWiwg5lxzWIK
Y3mXFr9viabOOuU2TneMy/AqOEEnTAI8VruyC6B6k6HgoEfm5ZJBGQkxDUn60ulBP+m/hY98AD/B
ZfXzQXNEeqL+1CP1CSX41yCoJ6g4YVIK6QWuIfGQeDOCcbzdtvuVdp7NQEbuofjAzyjqNLwHQjHg
M8zf0JyPKAk8tjkqKdMhPSAZepYfsVfx9Aqaq6uloVx1hWADTDxrCspzBF2sWPAzzKVxcr0vPDPD
J6htJxNFa4/AEFW4jhxf7KvTGdFU5B8m28ienYxUp9AvEUQMq3fqSwwRlCSSazX7wsCHgJ0e412l
Xh5AwNepZ32msSXBkKhyy1SAJT7G3Japlzdkh+1ZTkIx0OV/7e79wVqeHAUFTWXgYhPqFgAN9EKp
Cl94EQ76+6hSphV5izYhPHZXV6aKUoEdcpk7j0j24yy2S3/63F/HF9+xohSgSqwjeJOJJjYRCW21
oVCmEJtwc2DBQH/AbD6cgXUf29UYZH/y1c66Hws5XXMKHMbvgbGgF+WOFU0BjsrsakyXpBI3bKwC
J71vJlL0Quu4p9xhzQFiMm6GVeZnQycKsXSeISHBIE2lZc8D0SNR/drKM119yLikAVh8BtB+NMbQ
KglT7snqOJ2gitCsx7YAxPtSDb7dOog710LB0KuXimJ9M84CQDGGIOjoBMO5TZfFmshNwaUCIklw
pG3+/ePUFxlq20k3iFlZd5CHmH/LBQVDSW4zKSG2JUqNMvzvgnIED2v0vEbOCCjHjT0QD7cFQ8mo
ymE1Grh3s4b06yPV1hTZV7cF0dzpfE5rFugJih0M9Hyzz+J3ppLCBEENT8A+HnV7ewWa3Z90FLQ6
c7vkP/+Ly8aBk0QmTjmJYU4AdnWSEmNUzDdeK2Tl451O9hJzy5GsFtcr0ZGbBYSWyOEOCqN1WsBk
TnOMNRJVU9HXkmlDiSVaH064qUPU/HgShI6vbhVH5dPEBxoEy/uKxyscsXNjfC7FqhK2yKQLFW3/
e/xmWANl266Y8x8frqNfxdECkgX8c1SPHjMvkBAJZNxfGEEDE3g9NIHkPNPba/2QynCEo/CJgaB/
g7LcrPUf52PSRecgnkQm12T6d33zL24zD3bOlInL/0U/lVcYKjl5vF39cChKvUabrz8pMaKnx3ot
e1AbhPnMvgL6XcNjNNmVLWwGoT8BjdNGOW+9Jx+dXWai/BeoNe7OPc9ul8mxSR+nIardR/eIekXx
TZHL5xs8LdDmCS7kzDMaG3M9kvAe/JW3J7uO+yMQQg07lopRtL2AEU7t1tpeJvu3pWIv1wXp7iiy
xFius2gF+FTcjsH2PJMTWYu9YgLb4sSUWIx/pEveiWHk7Zmk63KhmvUJgxsXcyvR9oox7NI03+3J
xoQxlNJ2g4+NA8dTm30vOI2a/SLi7/FwqTm0UPzOKAP/qHKxlL//s2UES07s9awWE+UBu15evUDl
FqHbge+SExKbCInbdbqlKKGZ9TCRPsKO9wPqn2+47Sib7k6Omr2UuVK6S8BgdgzHFJ7BNeO1oUmd
En8tr6ff8smmcZMmAVPZV0/iDQMn+vPVUjz3RKFhAqMqKIbylmzHAGBX3caujjzU0xyszryWIHi2
jZF3LXdGaLF/ZetBhkd+RwkXTEQYQzN2Z7YkzQOrrVMY33Tf5j6h9Tjy/VLxLxvInStcGmOMuMGU
eYVKap1DVHqDf7dQIK2twjuRgTnjzcGQa3LE8UD/zpI5k7StMS+RQdHPpJhCYH0mTfex+RAsaLFn
U8lLnzOlfLY1RAGfF1SYzr2JQ0s8J6bamkLEqY4D0zbPmXRt1YPpy/S5YU//9xWt9Lj8pGPAYL0u
3r8zlc/SgBuEQ1J8e/zc/Quy0lvV84KLHgB77lHnt8Z+W16080vmcw2RKnmgLMw7TsykNAkzq0U3
DeMpPZOqxLGzy8vVUsElI2sLpujoWDB9SmWhBjFZ8iFJ+7jsFfzSNeyEKj31QemXU8unUUKkw0E/
U5dRmSbTXQscxGBEFQpwOSsjilV9XntVzf6S/1lPF5hY5I/xat0RpxjckWm4Bi/IZnlDVwNl8dSf
4p9ho7benUrtdsJztH3udo8fJY+J8cEW4lStkHcxyr5i7vpslwliJT0W7GUHaFww07yO8wDx51F8
Kno6k6xCmS8WYiNx8v9mSMHsPkzfZ4+NDAe+tnXuNhz1UT+xDkSJa3fGZGDV2A8QNW3d1F9qY20x
Fy4NatFNZYFbYlfCzY5HDqZ+zZgABmbhQS5sraOx9Tf2ixzF7ZJNb5BsZuMF8h6/5eaGfz0fUfxj
cec+MKUVee950uWfcIWdf12kxFOnyjGULMyOqfykSMDa8E1NLUBfVRL17j4FJerO8sMxYiDMb9pa
Wit1JnVt5B+8WSH7Bab1kZ3fsPtTJTYMHixtTspLb18VcMjuBNvr7W/wNJM5GWOo/CO3C+hzzppr
3lOHiaAz98oyS1s4JBSl3veWssU5dM0Do6LKUvEPEGJcLmJKVNhlKUwzxt2DRNdW6Hqj4xQbAqkf
B3LgJ/tXbFT5VZNP0AWGP+52a9ZlUasbwFcqNNLYyfsjWHarv0m0aa7j1mXyOJkot1m1WXrZnFA/
dCSw3/QBh8/D2O0WPWxc494oMm8FY42nHQ/OOgDwU0Wt6EzUmemFEtIPNhSIZ2op7Ipl/L9C0knJ
+LOxLCNXwRnvb0ClktnN6Ycnsy5Pgc3JuaUTpSuBk8uEgC7YI5owU3uWBwLxbua1S0f5auKCcKZO
o5RHTzrHqGkYqk0XqC/VFx53RX2OPK1aA3XivKb4nPHGFZKmQjIVlEWrM8ccWgrFllSfRdipItg1
VQiPOvbU4pLfT9rH1v+1ukz6AxGHnFZr23ErRaULr3v8AownpNFKJKEPPNkefwovHVundiZgvOn0
CcLas020jJeGK6AF1dUL419ZLRuEcxddwsVxw8jPwSW5bh3WRVdy8OW9yfHdM59QR7olKYuOLYm1
pWKtmVjynCCGO0JkvoFvLhXcgO/XroQhbi93LZv5NV+t2GMG1iDFvvNLgM6CPtmADW2kgCkg6iif
JoC2phaS5tC6h/I8xmQJn5TK20QKReemCJjgZIfpVo67ba8UW/SzC6vEqib9vA7GWOrwZiqX3czO
bK5R0v0ZgT61c4NL7Rlu8zGG5gzuCCQJFLFEu1KheSNLs4WeeJFRK5ITgPq9icaooVIRuEZ47zuX
KtJM6egEVl/RS47CqQrWmKVfZx/JszL6aIYqtLsydq/MuawZ5uikfUqrPQ8Zlw+CmiGTLdb1y7dg
a8SrOhdlTYTJgJ14Jpe53ZyOX1oXWXHLQFDGsq/mAwnAbvUqRQhAcb14BziEiBw5PYIiOPR0xEwz
L1LPcsshWZBt7e0U/pPwDkt+ao2tdI2h7D2wAInwrhq37R6HXcCTycmikfTN9PNS9pxLMe5tIgN+
0pZiu9Zgu4K+xzxfWhlphhZNtaP9XJ99+k5paHX6x3dxlQ6t2cuhL0QHdq1wXnKeWVo8pBNA9Q8u
F955XJtJAARnnsCnIqEr+mOABZmxa3YJ5wdRHYyn8M4I3JymeF5WfuY1O11vCpRWEx1QY3nxlNHF
Tvz2gVy303MTt64nBOod2BnBc3OpricS3m1Oc03sFSwIJH0Wo9wFb7p5L2yhjQwUDWhrLk25QY8M
SDZTTVMRnJ5zbGlSQ77zp5Abyl6cyYfpO0JW/Dv1d8x2nAyB8etyuTNm1/x3PoPCSkZMJWG0gqbQ
566PSYLtDJbVV49UVbis/2aGsTaYsOsp0ysOmkoCtGtKqBdTGdFwUr4YACNcgjZ4a7ddjPf3jUb1
O8RF09Lfl/5b//YUx6JlQ9nPKo0HsTsKhvGF4qFMdqDQjJV6I/YgNviKnkNyPCJnJ7l5jP0t3VMm
/apn48U0WJrUJ2d5AypRwdZYiORMiXEfT6wEyJey2eb5hQ42DgpHp9fzQb8k+4MaVlCOkWDE4FHz
VPrLkSiify1xDD1Kheml3v16M7+XAbC/leEdJ1O7CiCdtn7t9ajKEBUweuZv1ge+fVy+FwuUj/l5
sl+LWljLppDO1cAtK1ZS4Ok2oWkRnwg4dusk86zeJrHSPXRbCwJCO3f9gGBSg4Xiop1WV1QV3f88
YnfWN7mmJxOlHaYoGgtivO5bQW/pWwKdXbNPLqU/ID5EKYqG1UBU9mmcpFGwn7YM1oueirXyes/p
q2DIPgLa2aiujOgTl/MfQMhB1u5K7UT1aluR9GsAZUnfS/V144a6rvUMJ/e2+gOQDbkwyFNbrkGY
+ZGhEpe0+4IU9JW54UM7y5VblEhLezAcgvuyE2BJVRh4QrUBqumjRe7EUx5X9qDsayE2OMX7JY7P
+ez7KudVeCknn+ajBFKUs0ENeMjOfKfiZ5CXTNPDs9QjYbdGny1qBtSeol0pKMX0xafS8pFzTw78
ZgDuQKn1wNmx3WME1jCNHm5knkALmcE4GoJxQj41exkdzDbT1Fsjxps27XQ77sNQlnKJGUsnT/4i
iW+481tYC3/fonb0EBs7dLgnZyQra4Zin4vRQkgplY4Pia+OU0YU8MdgILl/+ya7HERbXGwV8iQj
lnS9hlo52I/UKHx59ppveq1LlTlpYKllmrPBkVXYU0vRbOFZJN01YDFc/MXYPd4jZDeX1cbYMchG
wpWweNqLy17uS/csK3gjhVPPNxXjax80I/h+hkevLesAVTxoNGV6qHW8Xjl9IPq8I4doOEhBxEG5
e+D8RPv9zopxs3aUd8goDn8pRsM68cuv3qmSh4UcauL7F9NoqD6mfkmYqB4cvqnpqNuQ3eeNf8Nr
yhOTo0z4pYiYNkUnVZ22XxqyjkK7eyvMjL3flc4lHrlYeh4RcH46AlTgG6ibJgYF/kE58ys8i39f
igHS0u7CZAUlA/kGqDkZWyLUw2iJIi+VGAqeC0iQB5a3kWiHIHu42vSKRuQSTtqKB8Qzv/h2c55R
fe8UFIKK9erJ+pZKMIkjkobwmkAfsg3nv3GfCahorzXZdSSFcBen8Gv3wHLy+AAXMnFXxX/mWQdy
v+ncsVekwfvhMScw9shAYdA48Ep+AhAq3fDZ4FfS5C1a/Tv041C8WGvS4MTrIQwape0uFKKz+QrO
p0pI6DuYglYYobgg+gPPIvNeMPoU7BsVDH0xlLy8VMS+gea+pAPFHZudiXrqRHHjLigftKc0Edd+
WBFdkZSCuAVUaW80Q0j6EeGc36tGZ0D7o0SPKQd0QuZIBbth4iq1e0dv7cn9fJzuBIUIsG9lZ6qG
0e54fymz1+MhAHcxj9d4nes0CObWI9sz+AOQkUcXQH/TOT7aa+hEgWJn9nDRWZIWDH35CxRuzCd/
hC1B1jpvHM6lvZeYJSP3GHr/XkUwXoZrbM2ROyXEhOk7sYYmruCOKdDl/eg6mWxffelB+ftJzFSh
hVlji6rDMdVFx+Hp6HuO4p+7GEroASSGpIGGm7MTRN4ISKAPBVfNgwqdE7Yptga/m6+1gd+X8ntq
O23GhXvx7f2Rn7rE62GuA2oA3qyiQfot2uKYkbDq+qmZSy9Ey7si4vMTQkHhbDJxXFy9VJp+6b9f
vgBo2V79yM0pe8soEdIq4qMbL8uMN6wOUkKOry0bf7UxFtCGoAhi4ZrDapMhzMFOToDXC3TNmx0o
zFyXkVE6F4acU1l10cV+oPVBnrHOZ1itX6XoPL0+r7YgI8guW8gQE5RGxx2KOl3gfipI20VnEjZe
sQzYSWLZqcLk0yHEn3f7Rv8IGvMX1VwTMy8f6TJntiLmKpdcrs8q5aWANBZlEXbUbazi5nwtZwXt
6/HFy039/26Qz0dnx1UjAuEQmfn10dMFZMcYMTsqHbVYBPl+GtxwwFm8l/tf4IpEZ2DHkUi5Boee
WWh7jC38KYkW2FROa1uPpXfyeKK0dHwLeTQByPda4GU64ylj883VvyMYny3hC/hT+Ue5zMm80Zlh
sgufeXcekUJD1mFaTXUiLjbKJc5cky6axjbzpMF4F3V7aJ7RQESYAJCLLviEn7x4WL7dHyNul9Bq
tz22LFk8kzdC8CIWgUkfZZjmDMl9tHTCXqZrowloyjA50XBNZT9RajkYCpRSor6CbxSEnZ8D2hjJ
rp6nWCg+eQUHmo97/iNN+HXv6mCS0XuJSh1BdnRXM81mQT2XxXMS6VHAwVVzZxmi+XPzfti0dJRg
Edk2eNU0Xnk4wl8QnegWhf+biH5svy66fpLCdjjV4/j9sqzqDO66+uW9zq6nx98P0vkRwB9KNWA0
3MagK7caPy0n82VYVcmIQv2Mx50qLwg1ryNsaLTuAAgQcuDMngOCIERJW33fMox3ZPklSxP91h8v
GyC2h/2p+CgHyNH9Nur2dmEwDzZmqMcQDF1RxzkiG9V7/NV1+24kXAV68gS/VT/53EhOHmTPDemD
aIMas6we08slK4OQey8YpqciyxIiLn0kRokKmqxOQulqgjCm9OdYAJ+h/IqM1H7rF7posIuRD5Eq
2ivMZSTghzCdirhoMh3ZvWcub6fgEnl0GzYDr+KzKajHWiJK6zpJ0QiPXLMyIMYt5qKfr4OoqJeH
ZWTCDA+X+IDUy5Zg4Opz7e1rn1lXVyM7mPI29LddTz/OAKYldakML0HM3Ry31pQSdBu7aPvOmUNk
6KmFVieB0YtBc731NQoQDvZWx4S+HMx4ywZG4oAUUz0rxh6u+OC19LHYjPVXz2TkDis/DGKY1ChD
fgA3AYBC7BDtyugyEWOIigBCF5iL7bQk+D4y9f24iW3QMwNhntuKB312dt0/aAK79lR9kJ7B+mcV
x/3OcJ5vxtdwSD6ZFTix6ZYOcSfNMJoaTdYchOJmjHGxmP3gXryKorhaqZsI7q8KRu4CvXJe7Dvm
WG70uEjdHETJ8Ah3asFedriKgrxoA+L0RiRXEZpMiw/pbeq8pacYBP6dTWkpMlKrWVfxoZ1cscJt
uoC5cR0XixWuBVhM2OVYdS88Akg/VfHSVX+b0O2UFIRhg91QOIc77/IEPuGk5LmV8UjMZ+hOOkbE
0H8RcxKiN8S1UKAx7j8takHH5oxb7QpUlgUBNQTh19/mk9mYZwLdOVVjSzNU3fD7YQo4096inxYO
RqxVzDTWFO3Zvb4+0qQPxYwRwllTFJG5RKfZDqQh79Lqcas76LL0xvLYMPaL+zym71Jx3B17xvbZ
YbZdcqKtO8+VOPcrVosDQ+t7OdHJ3cKkRNfDFdNDWQ/WsEn21Ff/xaTOlL61/EAvasN0gCNzBQPE
ZIyOxsFJD6jA4Akb1V+DDlmN8zSUrLHnzQiwhpO7fhv0wJ6q1m7zkOiAPdgj8OfwKzlZ0GAQdN4Q
/+Vr+dq2+DMhTQX/bp77JX0WRzqDlp83jV/T8Y3BlfKbdRjIrYzpMcgqmDtggmwMcaQ/fi+8oHuF
qyrVPx0WMtB9ZDJzKBjla++HgEaBtMuevG2wqpYPLnsMGcT4L9zJlpuWOk6SW6ifLflcc/ump/tZ
tJIVnkYAP2eOAgAtThkh7wV0NdZYMYtSOPtwlAhBeR7dlTMwlHo8UUvHnJbumoHWOlKAGypJ98Vu
E1GQpaUWEqI1ZM0hiQRcUFb0k+W2eUf5W9GQw8PxaLAHGPTIpndYAsAH6ojnQQx5G5os546RVFGP
uUCXVp+dr2BB20CTUypc9XdBWo9wpX4jD/3Pz2/IgQbmO2gx75ccm1Y+QqmzbG86YF27Ki7YjpJM
NygzSLQl3xQnAFJ2Xq2SQj3lPHkKduT0H4AGpqKUAWNTzIKd154a4zQGD6+I5sW/WPy2L31Rpotg
/szZ64+9S6x+BIM22Y1Vg4/MLymQ5q9F7C0HNFz9EvHPx4FZ4SrkZ+wMK9vDt+/yu2BFKz+w99g1
fadPrVElrNcsO+s0NsLVMFOTBft58Hva5NxwG+DudTFYF3dv8YAXIySar8xNqUIn1nuh7vPNIi+s
uFib8hSWnLZZHA0bHvxsSrGl3x+rYf7ZexWqgLBOVxtXPvTmoXctjyS95iOYlEIDrzPZi5gDq5Tk
VwV7eB1aERmkvSFolE3ee54Sq8ATMZVYvkoSEqFgaGJw10SXt4nFZMkaerKnK9yqqHiU5q/vqbYk
BIem4sZrHQrm31D4rSnH053gUZyDhZmU2ZgLz07BJ6B1ostL3UmWvsbEeTJ0BKaEQWliz3pAu4sR
HmsxQvJrURIw7GSc+GDmTlS3qP4+CSbc2B/yUXhpgRDu417Ip9FiKkMj6/YgcRWv/ZsuJekn95sC
YW/B1R9lZNKSfyocL8rRtVWRI3awnRhBzNpNCSttDm6E1GXwqfVKW4G+Sbgzq5DBLHwZ2+0k3ZKb
vINH/9QIKLGDnfGFs5zusS7HcfMPFDuscKvoS8aY7rhUL5qe+6K1+bB4AYEJsNXyUOV/WdvcrZst
vGylD7c1iXk4FCSeM3vpEcifU2RWzVANBkkMr4b4MM6xFEpe0PXembZGm+Li0gM02cB32om8yFkb
fqJMThpqpfmv5hDLi7NfxykTZhdbsUbl2Vt5aXeUoR9ehDNKSNBLgjy5E8bsadoP+kgfFGlltFPT
TuyQrWeJ+pOHBhvo0c4hkS6AvejwWuykW1x205h9mFYUIOoqLrLF/AVjUhoJtAGdsoepYKKp1QqG
Z82lgzZ//npumv3PpcBWYMzuYIlJq2RxLpl3/aP+TXAPAwMqrTyGZt4waYcYuFPBVr9ikimhbKjQ
Urq8bNL7tEQcLDB/Wtx0CDQt+JJDEQQ8Ia1fNOno+Qev7aclqb7TN4HQ0t79tkQ/Jg8fcV1CLtNr
GoquxbI+hnDxT9A+la8bdB+k++nV42yg6OUn+R6/mjBw+Wf5d0i7dnOVeKmxvn28ammjtajVA7pb
uaUc2F10cbfwPJ8Sc+nW4M3ai/hnkDy8z61P0HTC+bgcDkVfV3geAQ+hyw2qdVHMnXF7PHPvWc43
8fXs9z8Sag048boVRXVrwPskcR3/out2jpSAVAUT2DUtTXLFbcuqb2pPOZH1AG4+QRNMTJDR66G5
ChFkIhaa6EoTX9SqDibGHwTi0NNQpbk/KF4O2ZZ2vinreBnPizmtl1APID2StRftJQL0VGRQP+Ce
KoXHyNYX8yz3W9mBDVBx3ibvrn+ZO0Ve5KZ6k6pOwywujHRNzcwpQfMLU/b0VxMI6McHVctb3WIt
x0WF2ikNvwCeBvExgEgs195wPzfHjVj7gFzbJD6bWuMieMX1LJaBErwyUgdCo8RQa+qh/Ek07B82
tuZZKaMzlD8lZ+S/JjOKW6dn/u/ZUXSTJRIk7XoBB7i7vcatOFIpU+rnRsx3FxcsLVd9qtezjceA
kEW7jjAV8nm3hkkn6LZ/H35lck36NLdW2cnxibNCFZnzIsMaL0cA3YrKQCb/HKn5Y1/nvqnSjvUS
PnHuL4D9rkZaHerpLZvfSY4x4kqfX4no+a7+ZTl9QO+z9IwqIXEeyjimrBeeMI7djrRo6k2EKmqv
1GkTZ+NVPX2tAwr7q5n4ruN4aPdBcEw3Qi4JBifmvGyQ3+wxkJSSYP0ohTq3fkRATdYtNbj7gChy
D1RIt3WiBk2YsULItHNYjWUP/UVwmsWNZ3LezpapQcz6AsjtbIqz6zpwjIrCmDKFNKpns/xSAJ1X
E1pCm89h49mS/Kj4tRNthQjbd+ImevVJ9b0fsbK9N7cNE0Kh/YnjhfYMV9hAlYH7z9lDbioP1KW4
Ps4VZW/9lKnSNczO2yUj2Z1naiQ5uhXDUUvbtlCfEuEkxkgXkuv1U5F2iRjQb3MSdJgWYKNXhN/8
9WEXYTQgZY3vAr0eGilJIezNPjmCwT7J9rg7DjHVUpyR8Vy2n4uc5v2N48++hp9XBqvIGl05BNXF
H3c7xBBDbkia5e4jLRUvctLOh122BxzrS6rgP2hPcquTPtgP4eymaK28EwkBektuvoB8RTW/Est0
scCFTP5k40nKiQXq3ZsFegLIsEcRIFFovQ6Q/TqGUC97GC5Ez+xxfOuEPYWFdhZS9hKKLbYOsUDu
1FPDApedupli6M/A5gQIw3HTJlluW121hzkWauegxszRRRI6w2CLzManW+8A5ytXIQsD4THYUAsF
+Lz0Dr4VamdPPz8lSLzno1z6IYCD4r2KWKBUDJ+OQCm/uX8AW1i+V3ECngnAGdhpUwiL06zsM7FN
flRul6/zRuUWho0fpIT6qeU2dbBfLBPTD+oSN2Xu+WRCWDdfrfY34v/bY7/dqvHHRitrnqlnaloo
tavap/JIGlfLLe60jskng+PSERtO9gRfxcjy4wSTFAgiOjFdEM6rkzOtQMV+ZGy/J4BX/OE/iTBZ
ZfeLw8xrzQMjfX6Ga+zRKgNutzZ1j4oOJrrQXxA6EsUx3Exa/KtcEKCEw/TsKi5CQ2WPupgRSgkU
MXJ5E3METU9UYbHJ0ysyc6yO/nNdl/1eTVwPFYXbPVHeNloE1tLY3y64tPL558rbpFxt3pX6XQ7j
VBdK/cTTpmxcdSUq6EaSdq4aXAPlYe5ZLU1jEGjViOWj9hLV2HG6zUVOTl0u/MbOpvSTmyJcWpkZ
2lWSp9zGm1wtc0YOWHVzTBoZWr80rlDDLoKdfPbGW3llyzw3r7ax+GqQMkVeOIijKPyOY8w2E8xK
+J4b0IDwB37LH+Jv5puNMl1C+rLwA8hlHrBPCdXloAsjGle23xOx/lGC9YvSMXxjNUNm6jLLRxFg
NOoUiEGq3ES4zc/sMbZw7nFZf3c+yrxoegWWwS+ypxNro1QCryA37UneKfsrDQ/LF8+EAvWFoDgm
IXu1p4m998jIJ8jPGaVV7IkpobTg3vOF2Noyv3cH/4UogXLgx+ZPbBhwz9K2PJPNi3AY1EOeYt3w
/CkONvoAnsp0dM6TJV4/osTf+ij4Wo9ictoUi/CVHUHJfN/aKsDj1wqny+p4/mI6CHRl8RVUlYDu
UMDvIe5WklPJkgUI8jhhdJWCZhUpCJBTjXgflf2IylrpnL4oo41gWV1wmXr9nWT7h2gmi5QfNZwM
KlLBW6o3X9V7dvaX21U0wKLVHqEA4vo0CtDaUM4evR+PpEFXnFyHRN5iRMyi2WBDRuDV9cXxDP9e
fh0U3j5eUZ13UseL1roiDM7ky4yGbKsB6YobxuYggSSALMBYZH9n0qglAh/j2Ej9t1lS7Gbuo3mx
DlMVbpWK/31S8dSekap14B12paJO5gHaUV5W5O/zHQcWl6jvv4ZB27fCJwMs5pI4TyMwXRTpm76c
kOAmhIVriJPMtPkt+wNtpKOx1W9D/hWWq3HKamE0GwHf9QBBiPFKhp9fLDv185lTPRk7XW7JrLL1
iBo93QTrJzAv7LNp3DQIG/zDRlpryXTHVyJC2c2dgEhw8P4bJP1ah/hZnJNJvzRQR0sLaxwX/I1Q
cpFUpbrPc74zhZnzENxfKDNs+b19z6P/A3+wn6xx0V721X+thEjL5CnS8bPVHAuxwHR18DKOdSb6
Kx80DDDFK9lahUbMsQpEP8trJb5Xyeqgugv/PJvZxROFYiJuTmB0W5pbZ+Ro/bSn9d7sTw0oagd9
XdNFE0ipwVFaYxh3XONw8xkVkSWBPBeUnCxdD1AMBVMmh77sLPjnWoH3KV04hiTkfTtWQqEhLNfm
PIO1S4l4VwOK7dNfF8b8nwyP1DQJQGchQ8SVuPRfixSQFBG7VmvRbdtfeD/Ka4WCkSmI9QEaKFRh
ZFkdeOfiIoMyKWypJG0viQNSWtKflRaSMEb3+Sti/DtpSoKIY5mw0PCohR5VgrfoA1smvGB5siRR
QnKrG0XdVC9Jpof5SWYTS6qAtzNigKH5/wjfkVVyHgdiRyVMIbNqfZDpKxUnKvM4XLtNd3w4Hq8V
5gg2xCRQp9IUMpeXDqAfnWjFnY0gtU3t4y7A/Ner2dty1k01GPTjxRdpCmXg4RkvxJI0Dya2xNxh
HMFeIlc7VWwZIJFDukb07Fgc+ZdBD3Jj0AC/Kc5FTPlfSDU7hjMO+qbDoAQIn7VABcpUI4dyXlr1
K+gQ2knkGuKP+PrK78dyFNH0aAGHfpTkd1IdPxpcKpo8Velx9XoBsmFWoS51quLh+ehNr+b0RXjB
v82lBMuv0FUHWXIs5UoPEL/+LFHGq1Z2dISg1XmMSb0onkb9ma+GZVJQ5tmTCej/TNKvuNKfuqro
gwnKZe0O8yXkWEGGnCVdXW4F/+UyKPxTStxT85UW81/8CqSOnErnW5+oN0WR3oswRNBPYQBg4MFw
vPs4ZzFNJl7od4uDAF51XUpQYKkH9jtNkb7a1SxIN0giCN1OT752k1U0aTijwCc5vpPWI8u1GPcx
72KnDVv++Khho1Lozit7oJQ4Rc5dk8kp9tizdGFrL0kCAh1tDroFd83psi7jtlF8+g5JGpOkXqBq
5KmPB0OFGqM0++ZXcwAAGN2Buj+4dNp9IZpTIZaMHCwTciflvCdPyXnkMdt9NRW7YYUbYhba41q3
u3qoko6B3bUCpk75pueLn9mu37GhdDFMgNzuus+0PgmJu6GIXQro5XMTT5rl3F8GgRQsb31dOD2K
KKfj4QVZbmD9kQC0jDhHg/VJiO8WPwdAPLoOpXHV1Ow6THKGN+0ksy/EDYYf6BVmVXzYWLOGm3IT
risnL1h7bbRXmHjaG5Ys33LLY2n/fPcEljYdcyzuSKoSTK9eMYRutB6hfQWTCqq4Qf6QnGcbn7Wi
L+NRML1s/7vcQQrk+y9m10DzFRr2CJrv80+fR9pxFu3Vv53oTc6AdgDA55uLYz0qBCQO1i4H9mQl
k7sl4KwnpGHWeT9/TbcgvzMqKy+6tNX5DZVNXI6F1uQQ2FUZAv6vTsNjHFp5npHAjWt1wzXyMQrG
91PEKlUWrX8HO3jewqzY9o7kVXl50TKZYEkJKBxKvz3wDM4u20LJiMjRkMFXcZh+8QdT8Ii/hQre
AzsAIEiPVFkU4Nee4kVBBXUY1bNLXR3gGXAajUmgr6+Z4SoeWXarEFRc3fXDtLxT18/N9lij/U+q
Lr/beXmud8xFjbY6O1K8vG/QC02eHuR7bpKqeLz/6k94mdViJF89PEqJ0i6b31M3KziJwyhFmKfG
r06FDoC3k1RL9AqbFk/E5Ymp4u4XmC8xkJzbrih4jYETnstXMmcPMkxU20LSNUVGNZwygRbFX63l
5l23BNz3icvX2BJjDxuBzA+9U84FD6/mxhY9rdxE4G+SSZW6m54bNFCPs01ispBLLlsvCzTEOhWe
IFTfF/8T7SwIssiuevAShC1WYvJ8e71OsOPdjYGlq+shYWxIBsX9aT015eP9yW+8F3URC7WwKc6S
f+NOZWhjxBemepMBURuhIjfiEvE/lsEOD/iArmIEI96WTaUy8RqhrmEX9mf48yaf+xe4Owa8mVDl
nrxLTA4eozlckhlCjmIvRgOIhWQxHNthEjTWdv8wwWs5IKEIqVPhPSojAe4YosbhcreNiRH6/2cz
oXs8uwCcXalq2H+RFBePo58DjU/KKmckHiUXKGPzVul9UnsXS9Iq5FpgEqaqOW2sFgpETU+aNqjd
ezEmzCGmbijYlGmgwQhz7mr9ZU1NhyEgUi1Gw8UAvDC5Vnuk/cO05yErbHVwlBlRNA8/vS4TIcEl
xHI8bjMCoyI8AEQ+AQ6xdhxBSq82D+PILeX+vG1hyS8PqEBf+1mDa2/fPRmtUvlh9eWU/3F77iir
V2vjm4PPLiYjeqffyPcF9ogqgP9RGgpANw1Wmb2m8W2ZmW4ocqK/+kQmino+QgrDhmuFawclFJPW
F8qmfs9nbIetXkYGvFRG/UVzfSGM1+y9dsmZOqR/L8YmlFmRGoNxOyJooB617buJkW/rUMR8bnMR
OrEuM3BgFW5IVtqwKqOvt17AcpTcMUFiPkOynJuAKNiGtP4hqkz5NqCLwUxbXi5sB1D4kHLkk7gg
UmTGA7ZSvg2mNG955ELmgXYFc9w4PUL4fduBuBTiS2tYNKVqJBAhQrnw7HICr+uiAV/u9o5O7TGP
N19ToLv8wN53khHYWTxH2joLaeWkIo1K6MGLAJ5CzGQPd3wb5Qz78kND2Kxk6NYf6SnvLX1An35e
bCxAr87SmaLffe+bpdG8H6mizQCa2dNwzaQ1Mt/kedJwpGKdszSlgQjyiNpq4nIjTeaODq+tYN4S
SyR0NHFdZ5/PNmYS5zfD+BIQYmWffF7TELgdLv8/skzvFizIDx3CAqDx1rONUJK0PEHVeso+xETc
5BAdkwM/d9wTRFwlH4jfq/mNomrbPdbMzigWAc5qjgz19VsgShDqbDjdOeLIYYZCj3bqFtq6uLve
adQQxXp6kXC/JG7bXGqG+OSQoW67Y3ew5JRQD8HCA1KmFrp+oqleNsoRr0stc0Vo9YOHMYqeiGJ2
MlrlUEPvgnw31K56S4ynMMI9Dd8QF+Qy1KtRdPK+ZHZR3ZKkAYLtsebwbHlo8A6rA2EQSttpngxd
dZhB5cG5nslTzrP0LPng1LQdNfHRW+bTb+KbWXAjzjdMYMfz0dJmjnHkC+72qcPhtmYVNyO5XAE7
NQcPudEdSdu1ynlEwM4ua2vLK4fmlI0MdhPcEyP33JVaXcEsn+JyKKrYZ9y1OVUI0jfPCMnLiuGX
nWSPS8+OTaSS5PWbMryiQYhtrMP618PU/gS23KZwRdCya7zqRuvvEhcIaZ1y1uSGKFVMUjzbXdlE
57gFbEvruUh282y7c7//0LKgbAEX4qjPJvWsH+sOGmho+TiuhPDvFvAkt4zSfv3JxjIghP6ypFSD
2y70njn+qgrobRy57JXv2bmnaJyD4GGAWZsku3qYQWuXFwejN84kiNKydpO2/+e3cduzoLxvRiNb
wJ6z/sDCZ7rZ20rTD5f/rm4qj06xybQrFyuQgjnxzosgpEY/RSPeU86v4aLlz+lmVuDY8g0ZPLgd
FOGWxWwm2j502ugMDmT27+6RjZeUH+5pWY53mNg5YVbE5dACzPk8u8OFZBttEf+s3EE/KsaYjIdd
aEI3AJ8PqA/7p4KvQfkR5zfuCGTq/B6eLiIQ6nD93XFYy5uZclwimATSFm+0k6YBp5i41PS+J6Y5
R75TGbw+JrP1zPm7bt45C9Z8H3oxwZgCF/QAHYO8FD0AT2e8vYSe59KY0pqqD2l9/qkC2aXzdum5
ywo4N0iY5b0oSVyvjVWJYqEYB2qYiWhrzu5tIaaY3Edgo8UoXdJjnNBr744DkKC3CtC5SAVqwWxP
OsE5BqWyhoBDgqB+9CpBuU1weeuTitmG7NwfrDZS6+zVuf3LcHZNRflzMlYSj0ffur13maxXRmpC
BFQV6ZdFCui3R2IvPA6ZSpQol2zPTsXeAfTvb1oNR0s0vt9rmRtw/0GRPUpmvNnCe4FH1uSI0Myj
bE5IeRgQKwNmRRE4Apk9Yjub6wgx1Sy/QkhP5RnBCeQbQaR1P6o9DRaye9veWGXrjPH5Y7GHURdv
Y0pzONN8fvrfVcNBG1FD9AHdyMimVOYAdSSIRIovOjgLiWiBkzG5uJ9OMfdpTylQytjea6MTcDPF
PUGYdjYnZrQ1aoKjScwM51P39NGmQdPvt0hsGXkdRnzE6zkwkqPVdlBpsdIXVG8sONXVivZyc5hq
3PHX8sbfHsFr6UHCAb34l+sBqoB6zoL345CcNf5zZHljFf30KN2bPQXLK7yUIaNXoNR5wvNTVpok
oRElM+0lqTxtbE8kV3nqWydCU4x0rWDDFLNkJighYepscS2X6sU/mPKjGrv0gz7LXfu072HYF/U2
CVfnOdk+8XKlbjAAu3nB8IUHUdJ5LnO+av/vqmM2m4QFYbm0t8eze9zy6PtPcm9JxAC/+qC1lDWa
cqKUl4/DqIyummBTCNS1wEXYbeIPqTzUVP/9K9wDp+A2JDEg2os90qTXwswgOBeNTHx1DqdWKtX5
Hze9stjI5gGKdKfKSW8L3yB5vtstJy/T1dWMI9anZgJPuDpRXlLBXXJ2SW793TpRpCetOugOq+qW
hk1SK1vi6ZzScifpFYcUfqBfWXQLGakDEcxYnXzgsggeKI7rPwnIuBLrTBIdKtufb2+WtBjyJlH5
QmfkpDHwfXhxr0qFjHIAT4Dy/DwT6hrmsEwnUCNf48YystfZW+LK3h4GDlU7nipItxgnczMDOl1s
ymzL6hBLwfr9GhqWyylrwtOwh0zq6haBi3mNbKHIJW6hMb5/H0GUHGz8LDqCSV/BLJh/2Fz612Cb
WSQSWEF4mHtNhylJEZ4dDWhKgfOOodNSrmV+Y8EnVDKddKTZP44o5abT1XCtA/lHS3FBuNIlX72M
D6YAol5pEuqjRtO9C3+oTl8Q1USm5ro19Q7brqUuuTmAv0YDBH+mSj+We5Rq/W2kUsstFea7mYOA
qPmvx/qLAWKyQqm67nE4TWlrg/6+5E1KK2sEqsyQunRRQs+UJhJYhaGgqvSTgYgYE7xWo776GQp7
5IXmfQcTDK0KZdQpQF0KaQtTTxr6AQNuzPPUuSjTnRPweuCc/ztgpEq0xYuCf6qAKU50osYsUAV1
YK7eZbPeNDYl4InwSQ0Zr2wJveBVJ34K/JtGO+ru3z+XRTkG8cYFLipRkMys+GgUsGP9/0hrletL
KIo5+z/838fqQNv1PZtRVVchZctk7hsiQ1nnlbBJ7v0W9c55ktrguNz7y7/mS8moq1XZbv+pD/qO
dPWyiKP5dkXLXKBSlC0Cxh0iLRXCXJEF5D6Ek7wl2tZZzzHqwwVRnEDH3KXW7+VzoEWLXfbEtk2F
hvSqCbtV9K80TNbYTAiS5Nz+TLaiB4J8YB7ZaxuxSNWBVzkEyGC1qn4EpLG0ZeYshupt/OSyZQkR
gvCIlQHaa9HOTpe/vA2jK9CPlIhpyaYMbKnUsa5RXNDYSYZ3toxNYeSLVudwKkV9gziasFUHjOss
SeoQu+BDeDMCW+fl33do/ybW50nn2yg7H6Nu16G5UyRWlPoUig5KOpUxTQ5ZkbkfjDZ2SSwMfRgU
eOAGR7UplqGqeSen80M0RJvSfRs1Syg+iFI9FquMT95fwmpv3wk18VB2XxC1VlD+A4BjT3I8g1rP
l39NCUMtYFbs9GRoC65QaCtqRgvWtF2SzL5SDjhwmgikdCFn2FRWv+jJ9JCZXs1ENwqa09ikWZsI
aiX2sM+jFSWB4o668+9cWdn4CEfk1DB1TnULEjLYPfkT8SvA3k8NcB7oJZFGehmlc6CrHEDxq38Q
SbQBH5hGmZOfSPBVkTGCgfRfTEWg0F5iOy4trg8s8spWP8mUs5hm3bzkwpBbhNUdnDvQSNhbpkw5
DoAvRKfcp8OXfAh8I9tp2SnFzg9JzynguhnjkbNh+HvRRtQsnbuiIR4LEQqv0PQxqXgLUMJDeXue
vb+ovihPCgXQKw4r1CLKUfPWf60m1EC6lOKAV3Ae1RYi7Awu01Cv3CHFUPVJwo+gPGAc2rhDA6Am
bKtKGNOQLntjrCa4ICAdG8iuDUtj9dPa4zin5pa7CGmZQr6mPG+LbzQMiqCxCRJfB/U8IXMXqxTg
JxRt76GKKJ2bdpLLhddj1m1Il07fT78oLHGMQi0BpKrxUr3s7w8IJXKjnVj4/VKEnksNdKEgTJoV
GhiX3jbLxiwsdLoDmmhV77RvAndw68xNnW25L1lG2LiCPbxUiZyzrADkBarLtmK5IZ4/YR2rjAeG
4gum0GpcmCTjVIASasvDO/wjavkFbHr2boKSxLJcd7DBy8FH1czZESV/glS924VuGxVjMZ0VrVrK
e/yEub94fulUQH9fYfvlRW/C2MmLRDjQ1C3qXI9doWUMN1IgefcsAGH6AUEIf276bkgtKHYwjTGl
knqp6NPnyZC6xzwMx6TmG1Jb3MkivFC+YfLHYafOE60FaGnXdetvnXq8L/I6X62YobTgLZ4UA68a
i6GyJ5ty+t2FdnxGTufRM7bva4tLq4njDdE8bNwRQKN6AQuTuZW8979zL+V2yDhFqYdJgiYSqBB2
fGWoIeHgXLShcyBrZxyndBBgSLs751IIh02S4S8jfTCKIk71NDhzxcAcXXKgBDAZJFH1586k0Q6q
PKrjPdfX+hGUlICzf8IapGoEZ3m3DM+0AOiNU3Kmoe6wT7laGOuOdbdBDUmlOXLh/67LYIZWWqtR
kD3ugisnF/jBvrVJNOFoufKEAXeQAUG0omUx8v+0f3274nEbepbTQjT5stgDyP5BMym5knojGM4U
X8E5PlvJAiMFMoZHTIO7j9ffNRXQd78mHb6LA9ECyx9Uz9zF6+g4wGe8KAYhf9BPdC9R+Vvu4A1r
OGvyGZc64mpnypi0/NxSiqzW+yDO5E5uD9xVnbUZZ0AUYOehILN0UMZ6M5J5uowyJ89gJdg2c5iV
51UtDPjkxk4qO1vkM5Qh7fmcMdJHMrosx5T4tq3AAuV8La/PEg0p5nNxkvhuLDPUzHMPt/toNouE
WIG+XSE4q0ggNS2TuwnJIAZx6NCcczH38rJTs+jSA1fx1x4fHEQOQ8RZJmI71FKNmqgfwoahGGNI
YSPdSS+nFXgNx1Fek9AVc3GqML4wma8IM7gk+wPuv6IIseqdRkOibkAJ0SJPVRrW7rEZwysk8fpv
JMs3njcox5N2NY/PAGCpLElMSobiUWd4XCDRbIn6q1h1iNjdXLElyWj9mNj0xMZBVT6abJTO/Gqo
m8vPymbU1SnrTAAv7sPyWsrPKI69idcXtrhZw8eIqiNicVodTlc9s2kwSExJungQlDGj3YgXLPCl
OWGSMM1wUZMpMaU+htNTN9r3IVUqyZ1ri3es8icGPiNE0EsR/xireDN9XSKgcmC6paHQsVFFtuRt
gY6rQJrbQaMlqSOoPbJH8s3A28VKudZMISu3AUEs9E/5Out7biUem7pHEoJdccENpMgVJ/GJhISG
CRYBM4Z47TUuGNh1C9Fxj7iHDNTEu6DgAlcvZ+wmSDrBDFK4C4eSeqMLFJ74pP3rVT5FV+WvHvN0
Gz/4HnXbM5IkOuFHaWeu307W20AtozXghsnpPGKN7eRUlEm1eOdRp43y3+F52KT63TSimL9t5p3D
/P4fa92C/4Aq575+sHah3MPSBZlelX4CrsMngf7xQapKaS/Yq6vyu7uPBnfDK4KTFu0u5r4JeVJt
ncqWWxG4iZ/sCD4UiNOfNwR+8lMcnTQ1UMlIMjhBT+/RXjb1wfHBDsnvrhkTpUxiJjKOO3mzniZZ
xdYMU0PW6FqJ+EMlh1LkgfIFv+lQd1xRgAzH9xYMQyMX1NX69XRJqcIk9GJIMMngkwwAts4iEDeE
xzMXKFcGilBXm04eRnZafIAzR7Sa8sGvilXYJnkxk4BlQF72gUM91OJBwkxt4XHCnVRtSQr8ZW8M
OEXP2bHJdmcwupvFZXm0FfAvWCjRjhpYHgIDXtMG1D8eM8g/5/nNO6amAdwqXpvc+HFIVvtCFylF
L2bZ8gIbVyzrKKifaRZQdCkWPOIovoAB33iRtrY1szRDGldAIi/py4j/exs1mWS6khwqmtKlWmz8
0ZG8L+VJVZM0Nq8jev7TiSYuqCBMFWKRS/hS/K9u8KVuz2FBGyfySiho8+2PgiOuCpY928ZiHqjY
Szi3zUtmxPWrTnV8xnO93Cr0DxhewH+OTSAwKI9GFYqtmNodYLfxAgNPBnzyLhtnIhX6in2TuZk1
MOBOLDIIQ8bc3Ojmery35wFVX82GTy1pYYPCyhU3lctprTh9LzD4iCWyfhghNuhuWzPhChajqPTb
+pEu4hWivjoEHaJWSUPVNbySXiuVukpfHZJPqy5oRpaTLQfKUZOjh3KwiAHTolJLa5vtXXJH3HTi
0SdOAInUMXKiAufoqDhbgam49OXk5iLc8HR/sexGTp2BIgrodQ6dMAO8PRWyb6Yw+HdOtecYOq7t
Q91eO6C0mfOR9QA55A+tAhnu9ik/CoCtF+w+eOqdDqWOGZxmKDPbx5qZOtXJZOzrPOHryCLwCiEH
XRld64QQoyDMKg5k3i9tnFwbiqIX4sMkabErujjwnJssf1rWf/2pwHzHIEAfOQ6pLrGOXTWR6i7e
Ed+feRLsCM/NZ7d5wcBqsiyA8UDfdFdIKoZ2u+kowjB1e2mDzG9aKgs2QrjTwPlxPub7Ggyd2Dmw
QKX1EaxAW7K+/Q1wC5VdiChtRszYWQ0b4M+oUPxISIH9N3XF/5+vMrYkYymDZG4xLEcONqM3RYmw
IcVZlNyOu0ba3SeKizx++lt0m25MnvtSRa0Dp1tRSN44Uk8AZV16HCZ2Ncx86i6AzTUjkpFuiUgH
80XtGkZM211MYoT/fyojraxFU6mVu/k7szCFkDKIyEzBydqasE4TsiCdpgWfLZ/6MNs+eR+LkYLd
WfTaVQF7t0a2hOJCJ9xA2HmSHfRlNj5MCZ7cZ6vp4eyHOvURFMB7rrIPi7GS9aKVjHNqypdy5vo4
gFVCNEzkVOftuj6tPI4C38DVzWwOJ3h7V8wKqj61Tx2NtCXPCdlS39tRC/ZDHxXHQWA7ifp5HIVE
rKXDFn7AmQGNpCmciRadutmAenibB+6Z8ynlk/X51gp+Wi9b4F85OZDcF421d28RlLOv9x5WatI+
zPgmrB3R8PF3TeTSiUVltvXoqnVgR2oOVP7J3vVJF4tGnpY3NsLlO/CHdyYlLpRKcXskceD62NMj
eBiHOCgF4EGMG+9nmZF4xzFBR9cP24GarbdRYDmJWaJd3QqTXg0AlFcBczTt1+X2atsrUQQe608p
Zbsn9Uq5urOfuh2bD44b2WA7REue+Yq665GIZCjcC/ybwBHQ9qzJCYOi9EjyBu7hIrlZn/lZ+sED
QGV+0gClA6gULOKr5OdBAkipLwgUPpZfiUUhAGcpfE5rQOPK6IqG2p1VAn7RuZSy7Jk5Fe92DsED
DIjYuaywGtejkeCW+DFm/3nOTkyU1RSZe4+94+u3t6e4FxmKTvwUkfiRb0svOgsD+cfSN88eLpZc
nL7BWAGkNNr96uX948SFcFxsN6faCbtibV+sfCw1ddQ6svafh/++3Z9TU/FxWmsS7FbUmXPJhb5t
bctvGC/KEAgpcLvnK++jowVMpV2zA5O3h89ozxdhIokw/AV2LUQMq8EshpbV13S20U9moBxfDPxZ
oOqvh9xJlQjDVk0K1ht/Em6KIMlpVtjmURvfcaTpH9x0VysmXK2fhlQ+7nv9lYPos/QUXMzdO4oW
LPqwDTjvQERg46i5NY2/SBLA7gsX3PUr9bwLz1iCGmmBSGXkWCtQqOSNdJbY+jU+GRlkUk93E01K
kc0aDea+41PhumIjb8CfOArHTY5yADJjY8UdvG6uZCvCVhKNfOxJ/e7CzTIlvqf24ArxWwOlCJ8r
HPg6sf36cqA/SsCM6Re+LbPc+oDuJjWRvYYk3ztswapX1AvBne2ghRyOfkuh9H8vdF+h4Iq+LcJK
+aYnv/zvqPL3Lh9fWtm6o+kKSFBXHGH3bl5wcWOzzGSkCQqOPE/R0ApmBRoJO6iUL1+Mqp2Vtc71
8yvEyGcTXz3Mf2acQsRgQFriG11LBtFAJy7xb+XALW0JZfJyza6i/z7kYuUrz+jCYM9XsP2kO6z+
vh611HmUHxHCktXuv72ZpiZaeoTWdN4BB96RHk/4dB9aSr9gPIxLGFpossL5Xo/yj76yuYHrq6rg
U8IFJeOF9Tji35nJFEoQ+4mYXdmLG0hCbAtg7ksGP10H7ePtBJWgBkqCHsHoFfgVasIZlCQB5+03
H75Md6WVqo+oYEt/Rqb6dgV+pWwM6obM5l7lPpr+8RCidVOXJq+p/BUGSh635cgWAKhG8V2LCzN+
eYwb8QSLyEwrPXLjKZjCsbqK3nYE+a15LovAAWZdjKxyP1AGb6NQ0n/ZZp7WyIFLwlqpHMZ8jkgf
TcN4ybvMJv/CgHML2MTBdEAzCd7L4495GF/3Be7j3pp1ex68f03CT45c4s7Lt4WlY/J4MAAHz69h
LhocJp6D4i48RsUeGCtfL8NlV8Lve7si1C+tJtZpOv9e1j1o6dbIGPhJR3ujoj3Tw+eHaA//GKv3
Gbeio5BuAa5LUs7cUGqrLVK8oq+nv0QmZMz+kpVWj534+N/JOSXJ9zGhCO990QNqtB18Ht6falLm
NiKPgSeOFysJq6U4Ott+oI3QciFViNUj9igVSZoc9nQHB7ApebuQOcJYJs8E82YwepZ1TB0GEAGf
qv8HldLXLT8I99CJ9qprY6NUfl5t1TUyoLi9gzR2gNi+Ou4RoCeoWF01lVH623T8iS5NmEBjXrmN
3q7QAJWIN+5aa73L7gtnYqzu9uaTAw19UPK4gzO7MKTf7Q6fOzDTKud+807XK98dxCaFkp9ufzCC
NRlatEeg1IwQk+GDSQw/ajdJtOjMe3qBVWcXhkslGILUVHr2C+9SwJn5/mBJ3nBL9hBEnUGNf05Q
qREu9RZlX8H6zRx43GU50ZoEOpaibXygwxkYfy7tDMAa4x3NNrGAqGuZQCk6gEAWvQlkc0TqgU3F
5KA0JUdPpny7CCte8u/Ch1U8rstE1YmldE244tpkTrFYHbxQlV7LvtgZqZRsBzIr3BvnDXsZHtOc
kBEZdYik1J9gnv7HGRigpdDln2Y5H05gAtDuljJMJJLy3sz0fWrQZWNZRBIfSVtVZbtqoLFnS1+P
H3DsnoZnsebFjtwrFJKu5sqGnQ7bJIOqchMCOyskG7oHCXGLVs7Q6Y8U9PznrObgVHN8pfWUoBec
0YwidoE0dmCg+2o+3Ck8+dS485muEIQpeMtsJje7he+NGG8GO/7Cm7BgIXpVCmuS3IdGIVG8FcCA
k6INDv6Cs5k6HLSphwF4Rt1bpXRQptnL9UxkmCqnjVqqb8Xf3+5nptLwphqinUnQ86IGKjN7XRoF
ucSK+n+tPJxGX7gIQEYQrEy6toLm2XzRK9SkFuZVZx9wCXA1qkFUh4keeSpOvmkEY9G3VKsV+huu
Ot73GP8pkhmJ/qBQxBbyRUqmueTmRreXF3YROfp2QUEY5AXw0wydU43lC26hyJ67e/4GC784+tNJ
1vFPVNbGHH9+B8uYSoyrYP+5M72EP655olUrVNLErJSEBiDdWQPjAT+XBSR3ZGMAPg5pStu779PV
agffptqueTHuE5bX22ZVuKRbTAm8grN/5taV5QBD22k+oYoM0Yh4eW8+yJd1JxBJc4JudRJxcRV0
AaMcH0Zt7BjmkGh5aRzgIhhmu1SEWqT9Z7b6PCq3/mY2HBjwZE3dIt2xySUyyiplUYw0z84wSh+7
2Yp0KfG2nhomy5S9tz8k+1iMa0muNvwPnH6+p4mksGRpwY3Xrdip7FQ1PwfTwdnykEEwr7oxsuQ2
cRshcPML7JNlqtSmMa8R4b8dYGOlIT/b47tP8+7X8J8V31xU3eZgAMAQPazmUdGmXIqKNHJqKsom
u8MJ1jrNxCMjdfMIfAoF2uVDBUwgRPE+HtVSdM7preMcf3Pply/OLcd1Rb8OOjsXHYJ6V+Bpzc8Z
PrgX+ctJzzXgRhsneYHlZS1kvcNcTddz1hy0SI3TReVecsc47iN4YHy4/NeXHmsUNzcBaBpEKJng
R21aLJ0Jyys34iVA5zZQ8Bds8EFFEBqA8eBXVDeCsEpSl/FO4NOChCr4fDhQBI29AftuyGCoXB9c
wIQUZvyPXEp8f321o8toUaO7wLl8lLngiUFrtsAxXEW3Jcdzt2LXtNPWsLr9izX5iRbsgO1Nwl5W
BJ7cwnSkjItDfgliNdYZMUWrKJPJsMA6TB0SDaXbkSciMAB3ofzppsg5oegI729N6y5B9z2yyrG6
chv+R8At5jjoGvvN/7cXyaweJkz1CNNM1KJ4RrWSmsKBWejUduKJFmOlZqOw05bNs6BBw6gyLwrA
zc2gVYp2sGyi01YZWHbYCemTqZ3qlC+qQmNglV3UYUpewNQeErukvZcdWBOQVGTPjCOdentMkeWu
f9FlFjelwnFk3rb4Y++aq5xbUtJNNufedDspGIoVdpcGCK9FOYZu1O184I0A+f8nOmFv4qjAh246
R7WqQwivPUF1gtVxq+CdVa1C67ZywPcXftjLDgd+UeoIaMLTVDDL07tgI4BcF3bH5Gr61bASL5dj
ibRO0A4zYdRIM1gbPL1AaZxJT7I9BOIrlFolgEhKaL1j/icKy3RQAlymXQKwv2zHV6Pkm+5sQJSG
jqUwGLES1lXSf0p0G4oQXe4je4fME1f3+egaXHmPB0zd2Y/+jxxynqvbwIsbpmCWFynxN1g4XBtm
94FoHG6Xv4jWIecokOuYdnzVZt4zG328UnsJU5aJEEMzGI/gIQkJkDlieZX00X3pUr1rznoJwRfL
fDNWKj4//rHIWUQnTJBkrRsHOMh1wHDOquyNArlpaVaRqT38zSCtzGvi5r5lZ0nLXpeqaJxDbqkO
yDSoWnjR//RUF+fLa6q/e76ujCdsPYIo6wHIdLmexG44iRmOI1WwM0IF54ggWu5NXv/6p0cxpuCh
+ZIa98Ggc8uj/LCvftRZy+nLeY4OPUGCmjVoWgBwlxRLtGgnVpG/JK6/8lErKCoa7mifkF89QrrI
aJMFu0dJ4IGCqYJPnz2mCeExtlD9VcPkw6yQCDUIV3YOY80muAeihbFU2Pb9uyKbULnkm71OEKul
NHDZuw3QhkObb2a5xgFYSbtVFhLKDDrOmuUIK4cp/yhMtfYVl7vHKbG2adCtTD/lcB5jJ4j7d2mH
WOUWFMsnBOMz8QEQzQHcLJ2wFEKkotKfP4cIvT3RJJ/aZ066emTLJjmRh/QaI7FpmzW2yhWFejqM
GJ61OdL/3Mgyg1cDPJuGL8GFP5XFH9S0mPx4QkJypw7LkuWJCfCwK0QodC4NmgsrR9NoR6eMRaQp
79bLmg9f/Pvi21Fp+RSaC0HrCLYnOKoITpCYahb8YvfeMkLnd44W1MvRqA9Mucy/ZFRa5lBprNQc
r44wWKqbn6/qch/kDzrw//1NZ6eYUFlUj0zPRYWkQS7U0vGl17pgAQzdosL5dbDtjvU7NxIP9Qxd
A/34evLiOr3MH3d0PlqEnipsmL8pOvCmvNuc2uynugYPNEhyxmDIjBbnO3AWGwFdrZY++23nEwGb
0mR8Ub8qHIjfJan898XB1LNImxsn6rSin/W5tS9R2cApaUlDUqHq1acwPuqYnlz38a84X1W6zztt
q726WkYm2voMYsPFyGwZcFbJT5FSyX3qRII8m8seXKqmBQTuxEiY8iSjdbF1DG/7nwj+33nOM37G
5+iJqZBrvr85kWlXpPiWXWAmQMvaFuhr420rLFdlaBM51agiH8PDStOB5aJWJbfdQ5PkCDEOj2uO
S79IQ84+LJxs9c9L2AG+b5FUUEI+nOq2jH3yrGq/arBMW+e7wuZFM4NUF9CGMKVj2Iovu0iW4/eQ
M3VZogTToMi7KkHyrvyWn6O2Q9wF9o655u1hy5iI+gphWi6P5z8iHsszZjxrnOg5lNzty9+KeXZZ
fwPafw6keGwrD+7057M2rcVBFzwJ2Eh5BFE7z7LI8tRWUwIAbf1qm6sAL7T0uLRQ9pcRCKNDY6pP
dWZj7zjRZi8xdAlMd7OYpBQXGOv6yAZgCtxnxaBCDlGroK4KWTx0GFjTtVExOLaM/ZYYjrD09x1p
9t6vfadF5SVgUFdC+r9eu6Mrh71umHUXSsYrgJTWdoEk+0miOrdrAosX9oHx3jomIjHyvNjPYOkL
VzfG7I4ia0QzViaOH8f+dMotu6y+6PTHC5du+Q5hEoveiyN/A+Y0UNuYNvYxFF5R+eFvjQcsLv4D
NxCHs2W1g9o1Pj0ErvWdbZhEuKpR4tl1wMSedYpGbOWDBgbUBfFd9r91FBXvENiJ8Chvj5usiCQT
CkkvKUcHQOEm5MxPSvQxE2eaZhciL6Qwk4HRJNFHff7xwA8Exm3RcatoXc6pX4WkLlOuScHSLF8z
ttIOioUvD+Xg5kOOX681m71oApof20u/EXYP+htc8xiXhVDu2NNU3Xbg/nqi5mPXM51j8pHzAOsK
JiJd6l0RN4h2i4V21wJe8B18qiCXlFxHTcYqt+nDpgVMgXSFI8zGsuzP/+N2NDHNdsxFr1X5OtVy
6qZJfmHROuvTFLnz/L2imuH0j/gJ51CDSa3R7CxjwwWyR0d8BQYn8WWSbpWw7ziG88yDKP0EImQ+
eufh3t2FZQTUcTVwxQYFHH20knepacD/tWmzUwSn7O6OJdOE/VR6JzCB3CtSvgGsDoKC8lD697wT
UHehaUxJhojl6dop0cqhdbIyw1+MJK3dEIycNuiYt4LJ8+pZrDipSe1UX9chFV1NvuqPBf2diVhX
sL20s0Ks0KkMoIAGQWu5W3Gokgzq9mqe0QpJdDVDhAgJLvrGNAT8fpBTZpv7ZHrkc3CvPPDrff8t
m7kPGZ5rCkm3vNYd2nYfnUO26PRkxPMdbcBsO3QkgGS+iyhRlsElVArLaiRnDC6qf/2Sexa5IczB
o9RecyUJdiOQxKIguBIKntnfNcPJKwiKLfP7YxXW3Vj1AIeqz/OoU7Yx/ul7ffuNnDCG5jMslLRZ
4RAXrgPB7L8j9h2ucH0gF0PGCjiIGf7XmYN4W39SFWFHRkJ6zogGNg0jVgJcOa5r+lpV0RVwqQ2z
GiKn/KsXES8vG7EjSSubd+PnHB/N8GrfrsIJ7VqeK9HoPfFW+sADjrr28pYLjGeiv2+EBRZTDqXD
fL0pLsSkmocjuHikaqhPcvThaSMkVPMPJVoiDpIMWOiiMnotpIIEBFeD4Rjj09gDahU0XvaV3epo
9IbUhdSA8NAoFjwXQXsvBcDHW814lAS8rWuK8TEu7TloITAXUFMnzkI57eBxX75iuOWvShvPiuDO
6SIRBb4VEUA7I9OvIlv38C+++KO588W5KbLF5Ly3b0ETq3oAAbnl1WCYAJ3ZME4Jirhu5bIiqfot
CBOu1tTxECQz5EtFhaP0Xgy8+npqNJI9MX3J4cEaMxx9EPsLIcRcMkFRmRX7uph23ANjPBDd2Xm5
ztktz9HYxZZ2w0jm7RfXfqjIfWs8j+VNEGcPlnK5b0xPhXesEbDAkP5rNSSKdgjpovLOfIBX7V1Y
C4VKciO1bVcrXbRojnV82rc17kq78sejN9v9Vs2cT/LVWZPEcgB3UCfOUX1w96sRlvXYfvaVPnoI
vISycS37qQf0NTvgOgUWU1mdsnhSc75MhpWg95ri1fcOuzBr6i5LcaeD8zhDyOUxU8rmLBbUzSso
RidAXP3XHu4/xkz/4hc9RHfwhyFEipHPPIl0zb9QIJQOC+k9hgRXMN4tvnukDSb2h8R313YzH9an
i5hBX0rpBNxWhaNZtUJLfrlxwhoX7uhLJXJmcAt+0dvy7PShKgAPO9MhQ0jCnQCAuqQKQ3Cx+iQm
STPdfpwQvx+WJOkDQ6MnGaXW3FLuUsMXq7D1IyL1YikvPA09Clij0RhJCjqsdSJSBTUJIQgCZqBb
lB/j9E5Smw4Ju4fTVVyIK9B+mg805gLU0vBgPE/vY9Qlu9TKxVuO1VYAlOpm67/ja+AT0G+Or3LD
wP9bG3ScP4pboFnj/vAE7ZYNqwoytnbTYegJOq1ykZ7eMxBRrcsFMJcKZTaRtH5ih/aRglLtPpTV
lm8d5QpHZR4se7nvODlbqUDSN8cYD8FHn0wDWT0aNiKLqyCohiSLpF2DdwnCb2htg+vgUlCLbTvC
0tsw8sH0e1WCOVTCs4XNFVgazXxp/RJMrLs9CxicCTT0/QDNJQ2mGVY9dJ0XqoRqAPZMUMasyl36
LFIUmfpV6J07t95JvYPKZBgohUOd650YKjnmkxvSnEe0iGtlWMSsIN4/CtQulkDRHQlJqsiFUqF1
QgYe42RhQ0pGgwNEP3sLyYFgBKqc217G+TmTwacqNC7+xW7VyE85JibKpWvt6tzNrfh9Aqvl4eq3
70/9szp/bSERLgoHBwa4vExzE31NBV+abASOHgzmwdlfnnwb7NXmnTNjgxmLgrSZoYeu5HZF1hdI
ZyoraHiGBnnW0It921sbEkb1d1Zj5uB6VRpiBWslb7TZkClSaF5xnLhsE5KP3tOsm0zCAEPrbBaz
kZloNqD3aMd/6vuomRHeg8KAtWiq0JmqWyd+jX4WPviwhK8uIcmps/TQORVADIu5d4Zg6CXnmgAJ
/l/3odpRU2V6fDvkWyeW/V0giYnl1S71DyWfGZEkJ5lozo4CwrVvXJb9KCq3dWsXNusSzm6KHo4y
625pMxyE7015TYxX8/s7yyj7wcdzCAgzBZ6WdH8Wc0WAbL11eZTfH2KeqDSIyiHaVwpME0EkOPjx
mm4OSTGxrMcYiomrtArMrz6Sb8rDVLAfRbe529OfC7uXBz8JWdmuxFwETwlrCJww/ySGMi78JvIX
eLwGNESd1fF/Km/Sgtb6vaG80AalNH0A+dv0lbxO2WLBJz3P+oiklpwiUaIIwyPDzqM/ytJJqxHx
GnygdNYkLSZJo/OozV4GnoWaR9ISmIzRHW75oFqi7IEgwH06S0k7SFnPAQEtuy4yxV34tnsU4gFp
m/Ss8TC8K4mWt1CBN+RqTs+Bm5DRt7BueRlEPzpurXaicn1od9Fhfb6GlggCMd6PoeqJOQO7Nkbh
p3Ac52pWxscgdYoVAfIhu4z2Kn1Lyk9J0dyrSJtQlqtH6Wh2eenpVVRP5Z1fJNP5yfpu9XRqD8T0
UlduccAEc/y1lazSRROuDOt2E0mlvDkNOa39MsIXwxRhvG/dVHB8n7BLBvfOgdDGhGJXMb0x2Au4
Cth1mjK6LfYVh1eaXSxOWAPRVlqn4+gCAdabUw9H/iQULveqNAUcOrkgwTy9X2j/TFXX1RyAFOJ4
PastP+G6vO+paYYa2VfVgi0NVsJdumx1SC0lajhsqHPpVqkZo4f0GThUqdbAVLtnZoZrfy5Udrxf
iAHaUTvc5xzmi3T2ULmUacoh6Qu35rN/S+RmsuO+MAMsZo6OHt5y2/4+LvhoKMiRXxkCoVP2pb5C
Nis8NlSf92Hk7MjlA/Ghpz5MvqsamRWu2B+yQUnWnsi9zzjDMqza4ZZ24IlZv4jIZKML0MHr7khS
t+qh2DSDE8sPqceguqpN32fEI2TVAnErm7kZNNuW8XTd+mx3BsAYPrBkz8XkdSBQKg53LY4AXg+x
i2f7wGjSZteh/jQUVMPjPXOwgY/4T8PWlwye+ChLSZd38r0URwcUNvYyY8HyU9N/v9hl6hOzZwqg
WZuS58UHQN9yLPhm52HhoPJUJrlR1wGMWoJ3rmZC66cl8PncDSOQQjRf/Jame+lNA0F/sgiKx62z
zm37wEUl+3qYc8iM5Cxh093vsHqZfXNtkCXStZZSUzAR/VqnOYTkNmWltWx0P/D/iltoQIpvluc3
0R4TjtrSHaN5YXdikpgLWqn8wFRIVEufmZnSvqvGr+dMf1a9vg3BF9UUQuiKL/HJxj6JWKsWS7CL
s6I3O7SS29a9I64+oKZwdwedyNZaNMzn4b4d978547S9DzzUxLCvoSwVeGAMo73Ubvowd675W48T
eHNKcXbA4o5zWg8BqSqMKOcwuZzp3DVA0Fq6HipT8iewDJGnXwRTlEXhOCUgm5IcZ3+pqM0jA7u3
tFoO9FWyfdvfLaFsmmnoGablpUEpT8Jwwi3ag41J86nCJ0OSb7YTMC594AY/YH5cvRU01LHTZRYg
opaP7h983RaL3sSdoxl/VO/JFZkY21r9gc4IsvxZP1X0y+JUbrpcmAkvQvKPShqcgWzZP96wJvwM
u6n0MEjG3tzZ70bMIG8nFxH23xsc8iWDkxcYQma68wnyGiwX0QS//WPPXjZkRCIvpOS5lE+538ta
mX6/srWdI97t4gMAj6z+alWP/LCtp/wNAsCNt3DAYZpCjHJeqXdVG2P0WmiuAnyJ94MNnFBamK4W
Inz0dWNKOkYvVZdeZaDGiVgIu0/xIji2sBQGDULl2+5y4j38fE6tE9o80i+4Mi7EHRvO9IyAl6L9
4vX84fmofXIa8NDzNWsw7Awea/jrK6UKuOrPKbT8VSYdGnDJGcTMRiBaZg5ZZfZhwqPL7G+X1eE0
0SjCIsE7+pzOIeFl3n8PbppPo8NTqBmnZ+l5RJH0vZ0FviJOOe2wTqU/mWAGgoy5W3xe4lR6L8H7
uZBEaj+er6Oe8PrGe3zK4Ug3DS+3ODWwBU4V4RUxLT5sgfNZ+uZM+F2RoYd9VlRQEcqnVDukfSl/
ZmkmmKhvySVq5pBYg60TbWDbYkg9CO4th4P8gm+UDLj/yc6rnet/vfrgGgAPBbkiYBBX9hPK2dPG
7a8zqzRfjR2tHhiCW2wmz4dgnlUa8rFXrOP3CxU563U0LkF2iv3ULo+8SMyfNzu/PX6hUw+bRjQi
YbCFHF0M7UQT5x6azzgzmNcJE4r/BkLo7uztZ4xHEVjaF2R8ofx/PBHQY14Y1VkVMzplMnkWUeed
dj+iFQnTlyiD3LUFh1t6inrW3seQvFwsWivIWbnrlP5snQJg5EQ5bZ3NJzR6l7pxGZbBWOjQSWVH
Uyu3QqR37+gE1MUOhuYmiScUBqsGf5rAgqEOpsj0D3QePfAM1JHYiyM2F8qdpT+IPWImTPZtanYo
ZtPBgTkDxUT2zP4EeoJ0Rp3fk3Mz3ZPf8dzynNLYv43yTQD6nuoAcNiJ450QONPiIpS9bsBRNZxc
/TzQO5mjfVVt5Zo3chRrxSRAyOucZaocM2gP1Se3ZlrM9PRwdnUoT6d3+qkSarooUwTjgvhyAYfq
lJdXTow5mYLGCwceGVPYZ5Y5RTPhXZxmixUmrMjiTC+eQ/EToMRfq0qGSX2Qc8BqPyukhRIoFS7C
SOtsnHXFGU/nCvXNqcCLq9n7z5VKDcQKUh2FmAPood7XD7FNqmqOeisEeRHE7Br9l3XnLmnMa/Nl
QxpDbRZ7NlCZ7U6UsQyZIppzwgGr+HQSQSHRmrBMx286p/ZM/CmqUumkkqhPrHrn1l/X9OH5eTpd
bgF4x7+FyajI4mlvVJCCMJhCNPoOdLsF96M1QPXgYIit99OOzu7FvVpY57JJp7nfZ5i7gsbHC+BS
b3Lkh2vNKHvwjhxnMlr7M9ETrU64IZ8b8aMNZDXsz9sa+TKCQ99486qMxgBfv2/7YduGCYzVhA6q
ngrNz0k2nlzXJMb7hCJa5ImTyv6yIPcq4nc7YgK3ja7cvmqcsRHBp+uJRHavWZk5E2lRmv23Pfg7
LuiMGo5xhG9P/gf5LZZIZ6z81g6a1di72BsHZk7dOJ3Xgt8lpVTed6+6rn+WHFfl6DrlJg8uuEBh
gRNHwNLvLjvvXSq03LcwNVZmDllcErNqnbDeGXbDVmMfgMRO17pk2xDk5BJklO46fW2cv9fDrSOx
tjxv6RCIkTAF18d/Edw8S2mWfl9/Rmtnsk90HcJUlTp3EK1sGwTmyjITLPI0F5ezLQVglbhXXx2x
jxqv9hb2DcdWQQwESSN9U55iUJeW/5m8A6bH74UultrqJojxgwhTsSBI86faUb6dKBa9dvb3FTg5
28MEZ+BSdM1fRs5mINPvRzANsvWeCqFVche2u1DPHMKJPFRYNuUJve35RLx0EcRh8xWOLmxmsoEe
ZYJcKdT0ERwPDBLCgGQcIPlGf203AuH2cj8wlvVVKQnZS2FXvAzhpXszAi9/dUe0joaOx2XVYtOJ
IhVLArJLCo61CpfDWhFe6o4OJ9MuwtrEmOVfsNmeS+64JQsVgQsk70jrvwevVopZhXRK/CDAJUNE
BRb6ElBTqJZ0p0HYJP7a4WQSwZYFH3m72Z/owxDejZuo7OYCPjuFmuF48AsvT5qljPLkdZA+3WGq
56bsCGYg/oI/u6eoT9M2ez7NEbU2Pq859RbklZCoswFG/FLNZbAyX4rpXbUdzflmhNG8NYrQMOET
0WKhcQwO9VFIF2xMdYg9HVjbVTmvcL4mORvkFrNQHOIb6cY9VjeRCHngmis3kht+g/iHcDfszFSG
XrBmAWWfbwWcX02k3dQbhTDozTO49X6u1Hpz0yS/GcSHptvb0e6a72LSNmINycXF+1tTP170/aRx
uq/ucL8s9V6oGHeZ+EyGmr0P2eyJvLCACWsZ4XcUeI6IF/tWqwPK08bwHgecpypBkmV1y8wj4moE
RTmaMkQI//x6rgWKgaRL2wF2DvNYNKrXFebJJY28VuyNUE95A54HuuXhZQuoIaKlhiAS3pbDfTre
mV64Ztd7pPtdB3rymu2wACyBXxo77Dg+bEkFPNTZNZ6EC20O4vvAQAM9HUxYf9Je3andl1ODE1Kl
4Oet4MjevaHkLl1Nwy9yH3sDAB6lLZcvOPc6it1tv6dDQ6RiOpZgsrr1P9LYA12GiWQ8Lql2akD9
uwgb71SX+TVNe7+FbtnXhwtIVVfmogO2uWwBxB+fOPS15FoAgNoXq7+azrdFawEoyvsBTsduSPTR
PgvPNyjXG5m6Lo5iVz6mapag2QOn6UGVXBO6LwMyo9912kH4+NaLtxzuWzNtQXyw4nZaKgw7sJoB
eM4xoBt7GukFmZTgXHHA/ilBmbEi1nW6iIA5z2WML2k/I9ux0V3nOpPZdx0mwiVu0nTz4Vfvf4Hy
p/L08Kqk9VSFrYHpV0d6HmrP8TmwGPjtAaOKtJCYwZjUwzD0YakCyVHApHKCXdXMi7X0dmSpHTDj
kLB31ll4a+eWlUwZCDjtasxiywAA+4+t+iZSEGlDUeTVCSIL9s/6+9Ebbg7eyXCZ600I0eZnXgON
EE5vQDxhSrynCqA32suuD38idvrmq2YjAypkdcsFiW7DpzRtf//KDYbdA+tDSySgLOa6BfZXGPUu
p1OhYOHF9sln3KGD3e7pbuyj47fjqu8lwqREW/a2J1zoXB5QRYCoHu8R2IwkodJ4zlc97RlyiW7+
HKjxibOh9YMAllIE2p6CbR4GCVV2pYcoJQQpkzBm1ee5Tv1b2VA03b9UyAk5RlhXzksfGOQcWQP6
3xWsduQt5oTyyfDB+NsJGDW8/tm6tF5qFpzEDi+ke9tTjS5C1oVL+bCfU1kIdEAtv5sMGHxzg6da
MMIzqKhLg05HqcDHFMmsew+u3xu87//uky1zZbO/iHjJL5jJOs1sf6G2DKLen5oDall+4xWxs4Af
zupfZ4chHLtDv0ciy2nJ8c5cAUr+h3tDf4+ofoQO0yWd64nZSfuIvwkBtq0DL1Lua6/tUg1D9VEM
9uQUxhF16Z+5j2i4xYLDQE69RUUtZwsiwqZvkUskFYcOrotY3S782i1ST1ZFgC5/+6Vl4UbY+yLX
4pzgSJfsX2hF6/Gt4/hh5xsTu8CzVB4AqY05oD8TIgt759G9yXRFW5m6i4TFSEqv/2pfS3Gl1f+T
VNtkdymRnNTf4LhUfnAPp+xLrxBYC6qhV94iFi6i5IOsPB4YiwJuX/DujZecxzdsSo/ebIH5RMW9
xXX7O9o9UYFNBEELCHPeqpvTF4M1X9Kurs0wYgqArYhzIOr4ChZ2cgCwNvgLnL3Hl/1nJh80Sjt3
zeldaOthjDW+ZzAdcoYCrSXiT9/9NqtvBSCTQWfr3JZwW9u6lQRH3vsHjjBbRAeQyu05CQ8Bx4+g
eMVNT3P+CjvEWA4b+rSkFXetf4dv/5lp3LC6z+e1LnTPgOnaFHCbnbrHCozitjHz9et2NR1OV8UA
S5UbmNv3lqLLr4pR43wgAIh4srkSInglgJMXrplHdFN4TQ07Ep3FeIpPzt/6YIqNc4TAXqzSW4pE
mkTRxnmGKphyz2yJ3pxUED1INvAs91wxhps2pn4xeANGHl8Wc8jsuLeAahPJxaor03Dd7H6RdPR5
z/zWv11SwuLZdyHEjAC69+1N4lReSOXTqyTMKAx4tpzovYA/1C7PUlP9VL9VUmOudXaCrDP6MHUV
d6NvdIKkkvJxNEUHzeFDK8w0Hjapz4OCbmMEWvmQEVBa8jPzJJSjY3ebDxm1eHXPczUy2z21P9rG
kVzCHEPIaJt16RnIICaQSjNrtmHzQ4rnp+k16kq84ULZrn+yMC1fppEjm78noQ8AQXUozq2Wb9HT
n06ipq5Pjd62meHFenqlfkaERaHE1ZPdqX2CF34ShyELJ+gsUSd0n76BulrBMtqJf7DqcF0ya0S7
d5tLF66aesaRY9oxB285ukt9KkTXAF6LIoZvtA/qnhmkF7CRkuIYO5jEfSlj4DZN+n5mODs5BPLF
d0Xh1Ekrsk+CVIEniC9NB5WrFvDMVA4DJrcuG/6vFjp4bHzRo1wAfC/DILLj0BX03QoBPLDxsvr5
Syaj8Rff2eICDsqe6xKQzJOS5yTWTWuyJ8lukEbepqyOxGYd7lYadl54UMTPkAHAn8ge+y2zQKN2
U+wnwqUMZwSKkjjVuYpVZ09Hx0ASTY3Yuh9dPRsJCeNUzbux292CrAGxG5XQDkTgEB5wS35haIkb
s4B8hD1107ea8NUPhPpFCDMjAWSHZGH9rBFUZSDJoz9QhB/30aoT/AjueyWuV6a4rYd1N7MqzjSH
i0uhegWxFM/iLMoLiISY9ur/GlIP6CvXCwP8XDlaY6CzV+4KJch4eInnm+KN5Ygimqes9bT9y2L9
JV87kz4XjXQZ0uf81JantjeaSIB22qTFvGT4e37m6+uk9dRlmHonPpFhQu8ThuLxjSMqdBpPDYvg
yltRYMAZW8lhz+dAwy8Q61/I2j9BRgHUpux/MnlKHzQknfI7R9o1E+w5JU9oHHjq4M6BNwm4khYq
jlg5lSZ+b8njiFAk73RTw/9WPs++CbnhFqyNNEhuyVgImB1VW8JfqBrFDhSBEdl/fbSAE3qz406T
/pEet8yDXZJO1+7OzgxgETPjph/36ehbRFpSn03c5Bg2ea17TKZkV1kC3SZcLK+MeupbjSkqihA/
/WWSGLoISKjVZm2j/lxEG9RJH1PHWJPCCsCU7mN47kz5Nk461n//+hWo0KO8vt3rsI8pGubfgasQ
SJMj+eltRVY9OgJwZLAcHglK50Ej5GtUHK8HrmRWOxEPa0NzNORx/iUdebu0EAwdTSCH+GbMsqSi
AIBg0HqmTDwBdZQcMG19Vqj06RYpy+NgGXJLnEJ1fHmS6mzXuspPJce/ExJJEWMTG33DhhOz0GzQ
sjaLaSz1dtGmhDUbw0xJ8DxuoZKnd0ING5JjYbfBW3raIjf9ljsiQTX5lCU2ziVUwz63m1+UaAGi
ZorN8T4zBwknUU5qckiUdrFw9dbLkwhCNxgxnuREnvjpco4uF6tHbTaFAolzHY4NNSNI5tTnU9Oj
HKciQHSRrVlY0j4psD1BngLMd4g11zKfuPINRGm8zgPyFVNoka7hYBSD/fqEBQYg0uq3DBS+EqIa
hzhb3838wmHyqLaZedz4B/AHbCDoy56Nx/CkCqw0QwM6HMlpXYOTySyflcKG/zPSZVfTRLb1uvDf
XdVJArl/V/91ZuIp1zGkXCU81Cxxw6pt64p0X1TcQzd6BZgGh27dW/kBxlBgLUjMhDwYZ6MgTRgt
n5Mq81OxHgcJWD2kzmOIbjLK2U3lgNEQr4CxxvokYaCP/9QN+yU4IQOWU0VsiTpoGAUbpqx5fgw1
mmxJYjMTHNcrdB8YrHT4h2kBs2Aq2SGvM5MmzPh6t/OWNKI9mIvY6XGB//z/UbpJ3nNi6jNSDrws
NJOjtlvepcN2YR6D1VeRgTrbGAIUr3xS8L5CeuiYzebm5kYJEqu38tNEQg9RXUX6oDfFj85auWA1
WXu914jKlOHCJPyu3ppZBpGp6yvdVT8pnfx6zXNdZF/wkwi4lo1eyPTsAqvw9VGzGf6h8LyZ/5xZ
iDQyBmwORdAwYgxdMbgKqKXtSBowWsykmlGq9LaQx8wV9UiP6fOS4EpRJEp10IiCXYevt35296xu
8Phbw7gvxxmgGrWfx2EVWYj7l6W4epKdq1apoiBBZbdNJc85FEHSSdvD7xU9dkAvEjlCfJwFp9U7
QeGDyB1I7U5G0Xi+P1a13zxaUlQ7VU0bDvIFIznC+56aOzXfKXwDw1McjRMZkjOEWxoAmTR9MpWO
T9ChCSbU5TawjR77lOj9g0kQjCA3nHJXIR7iFv7FKI3FFdseQeDsuuVSnmruKXSmGrLljar6n/Hs
utavr6H54HwupvuFH6Ecn3J4Ec9Nn4iq1sMejj/7o3oY8Cc4Gg2BHbGcE9CYEhDc5h5kIMsL5K+f
WoqD1EWG5GtugeZ40k826soSRWpsBuNlkmWK6soXT6upngVdyQpbIaAUCKEC2L5W04zQZX51vULb
3bcL27GjSYQWaBijBb0dodrblBkfB149QKYMhnVYwDvnhv2f4IHZJlADsUUtfISrh8F//rjvyD92
d3CPveQ/w2Iz/7NGUugQ1PchbTOrhOfl0S0SDY1RV4eG/f+Z9glxoJ+MtCZGXpcY23sYbjVXop/z
huXYu31DdzeD17d+UWJmP8n0tCFQzGSd2vwhe5agwukQrz5yuyK4w0uQyTfJUYc+MlkUbxDXMXzR
PdMHUWwR8sNlRnfAuKuyN6cBXV0toWRC0OQY7RqF9NMi5xYM6cjRGraQ6Tv0reQUI+22IFjBy617
JqlMe33Z/Ww9lf2wVOM+m5kgQ8ecln9TqwpCA2VvQbWlWfOhL0PhVX/Z07un0SZxfYUiHq2/aJkZ
s+l7tJWkAUzYRWNWwlO+cD5l4AaoBiO5hsGhAsX7vSh6/DeqzSOR2moDEiqXjRp2wix14h9AzZv+
/wBpTfMee2l8oy8HlUA1avbJ6lZO6YP77+GEO/wYFKEAGfd/hL2l/TaLRFwMdsbZj51aMIryFCVu
fMc8z0FF1oCkhYTiQpN1c+FzRLDWBRCxbS02os4aaUAlFQZALfOshmFxuN+nvnpmJ+N7Ac2eBt8G
rpkkCnsCtdZOoG1k7vg9PJVdw+8Nt71xcaPAZx8QX2AyCdKpAlaB3AxgdX0LYffKq3lEjqyKPYYZ
yWIu5oXqmWa2O6hYX+Ab9voOsfwzOZiveIUPTV/50gXRonWZ0B4sJ8qEK1VZ4om4B5IHCwNTkmFc
orOGFbNp3dmZ2oHYDjS3oA/ZTylwUbwf6Zxcq/YNHtE8dUq8XNKR0CHJJ/4C/+2W1/jYaMq/lskg
egTeFeF1nwbCbea23zapxq08s81I0Bjp+fBzr4MaATYy/S4BCpQVTZ8zfMtGFAdD3aVXgKkY/azB
6+YLwzrWWyFFWhjfz6npe/0DRFbjdYlLSgvNUq9aimHD+47UWYpwS17xOg6GfCprRbywuC0u9m7/
Esqc5jtnaHi/a5Dj6j5Q7dIPq4x/9ctpHWfYvlfMinjppC4tDD3m9oNCUUVKHIjDCT3GNEQZuHGM
SPPt4y+o4cqlEH45lRLgaYLKXQ5/3KXUqoRyUoLxKzNJKfKj7H6KYpdRKeykah2gj9xbRi0UgNoF
nw8Jm0tI9cITyyJQ4UiUJN7CwX4V3DNHGWsF3M1QlszF2yJnxsl2JNyG/lrt2D56vXLZnbA1y2Mm
Q4linf5KvL2dXsjX7GPr84+Ma7DQBXDEj4gbElJzFBuA7lGPlndw2YJHe5RDXYfy373Tgkl57Vul
pivht5xoleKxFAvBIDmUcBEIQw4aKLjMdWgDUuKkMD0ea1yZoj7F7/R7VGBqP82EH4TIlKTJJ6Uf
ge9tVHssPZl3+FDIb+wkqs2GkC4CEG2ZQ//Eq+r/p35HhphJ+I7Dx8LwYgSYHwtcty77hnG55Zu3
zXubavlvbMkZd4YA+Tb0CIaQ2Kg8b4RXITqWGctr67ObqXTCKN+lNk8CNFdR5Y8M3I9z/OKqFrOu
WRiEtOH1fLFQNnxOdfyPwIlNmtKwjpkkcQnTC6DKVyG9Ykg0tk4VrBhNWRNThkTsl7bTVcwBvQo/
HdTUTtEarymcCJ2QxqBDMslOV/fMqo3ki1dpsbtklycfpuHhUHrMMihmhrs+wOPuQ4xY4KNW1oOm
nC29yYCrBhjUZrqRDv8Ay2PoCnFIn6e0UauopHxc6FKIk5DZG/gvcBRHy8uoHy0TUEy5zI4AEzXS
RrwhdNJo3jKThT+mantlsAnPNHPWD03586a8gDVtqcacocBSnUH+nPNjukMHtyD6D82ouJxQ/or4
rU5hIflennSz1VCwNBnIoyUTiRoKrD7CW2wGfCsCcGdJNkVO/LdtA0dYOZiu1OtLZR523+DpDqH/
5Q5gdNruCoKkmumOOnNidUquzNJ5xSuF6/6efFX9pD1WN+Sm0FTVDkGQD47gyQ44hqnN9ge1Dn/f
s+9TisBmG2gglCKpuSFfamL8wTTTF4f0Wfc9dr65lgwTT6MJQb7g6al6+iuN6JtcEONzOc+XsLel
8gMpBqFdchocp2sxBfiYa6huUiG55mtlEtlQDH1Cn4eB5QuVCTSAikGAKTlP6AUWU2czYfjxEuE7
2qRafpdgmwa0wb9+M7G2MI1BBs6vyGp8ahl4sRYsH4DiXnst/KevytbmIdldCLwgxORa3qlHu00A
th/fS/lXoKSYCpVM5ZBOsv7jguQt1OXfIjuVE3JYSOxRH/wc27qBqrvJdVf5f6kphjiVSuNk90n5
WCQwtV7ItJ0Avu0qEBl+ZzP9VVjQg0TOcxZkKvTwPMzMXcqEYSnN5K90SjYZLB5LZCaZNgk8wqy7
ZpWkQoh/Kl4vUkruoEnesWV1LR1hObETY/hn9AfyOU8L2MtBB8qQsgODxdMOA96bKUQVDtovOATo
UiT6+mN82Wocm8O06Qao9Dju6wCB+XhTgCOcn+R+/nZzVbeEUjKQupuQ6DhJbGxv84Pi1A2iRDhX
daLwax1EY6MoKQMWIT1OyXtwqHSMhsAQuZ1i+YXMYcgg24wDrJP+/kHwSVTXOCG0aUKCp4CDoSL0
Rk8ZptNw9k1xMTSG4wJLwTvww3fSMva59aLlSEGlFR0y7kFgUH1kusVU1SzwRbM14xslgYMs8Jgs
4Du2pfVjVEfBxlLGZBVG04BRxxC7uDsXIAbqTMK9fZ3PKgNyTXjaSND27GmcnzkU5COtCJP00uXL
mzie0N8jVR4u9PUbWb74FORv8+j139CDeao7DWbjDNzVB+FSd43r0+wvN3pWXgJfaFeERPtYhzmB
Jzs48gQ5eKQbjidGdY6qRotqG1ciLHT/gUaYWj2FlmGm2DK1nRe5NoDfP9ldOk4cRZ/nScJ/LVne
beB2HTJ6N//f9pPEr7UffE6fCAm3PeTikyT0Gx+QtPebDnihffP/cmNeA91Q2Ca0Y/ZMrweV2IPO
32h2CIVfhsPttYw8gk97qZzVYz2qX8jwNPZndlmwKNUMAY2XXAGObKXM6UQCLLKsLzsHj/p5SRVF
ltnD1bbP03sHC9qEP0ZI4baPm9JBQ0KIEaPqs7HAPtn1LN02W4fLN+iIcg+wUMogftC1XObnmSDg
QGTbVgkOaWawqwfkJA2k+X+xQwNf4EMZb5eICW9dgVkT8zFxA3tcVexhzgWeiAakzRzCsb8A0rRg
m9JLUQdjVJFgU7vL4gKdkGSHVESKtKzrR8AUzgrtj05hwJpKKf7xGbo+RfXD018asTepdU/U97M/
Vg3kr+5A55DR+5wN2drQDAvmxLMmKfriTArHmaWPK3iG47nc3qPSsyGh2h9bGt15nj3aVbi+WgRU
x1JWLY6InWl9JJa1I7AlrudFn8AJ1tz0jDG+2CwtvQCYJVkKvJjT+S3Gh8lYQleI4HJMhSOYsoTk
h1bXhUFxTyaWyiLs9q6+ikEpH3CXMl/D8388jVEEw4sN0GVc+EA2DtgCBjWtRMQ+M/iIWN8Gr5gA
bYeFlFI1tXOSRh6AKnWOA6V4gART1UGKT0KW/XNEB8+ledOp9jvBkAmxP/tkOzQWZ2qCyAr89vxg
o8/fTddGdgA1NoRgLpRUCPuMjNM01NRH+nS3t2DUjdQ8M1YKUeItEL0oW1yQpm9RaLYACWnR32No
SLSiP2V4sSwy3wbQ/Fj6i0Fq11D0GltGkKU0fSm968RIh3NZxhYkamLe3wb99ZcWLUvTUHC6aWbC
92Kh/BkqW0nMiMkw7Sw3m7633l++VHOp09RXRow9kAKZI1DwThFUcTHp/+gM2713HONIPm6yHnZW
i0V/YJvZA15hSzi3NUxEV5iI5jq4bzAiqansY0wI5+Z1AYZRB1u7aoSl/QGv8FmIul3pANnxyNvl
F72/u9BX7GMKVBO0YULEL4Bcyf2DqgkjcQCBiBrycogUa8nxBuk2SYUMHh6J6JRFZ+sG95i7UPzE
Y7kVd2gDASVrp0/zDkfOcF1x4dvg7ne8q0GiPhxAxW/77my6WODK3NN74RKnXuSZL0AMB+S6PESz
pBYfg5p78oMl+KZ0o6koIKzUQYa8sok3qjb5afO06lLe90R/JS7lMA+J76BLNWigo34g70MA3ydo
LfC5bme9IRhQMTSiLvzo6EeerkXGnmSP30KsUBNrLVvX4axWXWdp6jj2wLC4SY5VzpLMMgpRBfsY
JQlzW5yshKmSiCz1mvJWqf2X+rErgrxkAtV7RynKMQaFvVtA5uxlJEz9l0F+0Ti09bg4hy7b55vt
cMKFTLGQIFbdH3Lvdg4OOihfeEFXBWx3nAzEYstnCyN5DuiUryKi3NF1BMD5yUlCGHuFtf87UlsH
TbGjZeK3T7Q4JktTAp4Ji6vHagecf/OnM31EZyppbvrUBTAo5rGBEhmnUQWUVDe77Aif4B7l9zhV
qMz2fQ/i+H7Ek1UlQSiAdTqlnmQmw09p6nAUZyo4TTmGkh7tpQuTmKzlFPgYAsPpqz5FO7Y/x8it
Rhj9iPTqk12h2XQWLFWo1/BNWkMVa2UK9UPiG6D6A8eY8ipXs0HNtm3txuBRwoESkPujkneJmjsJ
rUdAXhyfvdD44z+MUpZV2IDoybz5rNlUZWDrKh4npXGOSAii7Lm3TGngacvabCBRVTNugNm9r5vB
5tUC97v5h411jjxI9ArWAtJZXnmM283/rlA0LWQtbUkttSw7z1Vgl4DbAAvb1H/O/Ctg9JMFkywk
Fe3V850ijGPBd+Z8D/hcWpDzqsS+A1ic1pL2k0/fPSsS+W1nYNagf4PEKwrl0G/acXtOpSFrEaUv
V72q2WNDqxZyt17DwKiwoBVTfsIK9xhZg7F5i+jtGBbc3QfyMhBZI8zCZ4ui34PBvxH81Q4z/hqr
Lyrpm++EhRHgAX1ZlsDPsi3djf93tAVdPkb6mbpGGAjsPT0rIRZ8LvD3LkbqicyYy6kIP/d6DOGA
IzyHFwTy6WoKJgxCo1B5pqKPCMCm5bggHrInWoSiZqs4qHe0qyF5BPA60XvS7iOn3+cNA0boG1H5
yM1PhCTidTMELq1iv+U8UuPSAvuzvtngm8BR7jD4NSOpj8ouE8stgem8G37Cb0GkzdayrY7nqSua
GeMXbtP9tZzxdWz6A4mZQDz4ZRdIgow1MRfEfegJUsumYP9fU5C11YnVujXUy9wujuuMWaea3G/W
JVwwLIgn/tpCK4ZeznG8gL+yI/O0+FRS+UtYo4CNZjiec3lhp+Ua4QU+rE6UbzqMO74pWmASUJHt
SN+YDgRA+gsdeLRQeeXu7GdZcDqM0ls92jiTHlcTtYdue14CwZIadSGyb/EHIYiqyozJrKeRNeNZ
0oKLE0X4meVfWkgmvtNJZCCis6JriauO9WgAJ8TSaE5qTViXrqNcufJ+Su4SSXDB9QNDqxv7UaW5
7KyhkeYx3PHn9+aVwrWUbyBMa6E/QrnQt0gJSYFMZL0WcBhxqtTFHKaP/1X57nt6uJKC3JO80PL3
beWFlgEqNORQKKT6NwKZrvkueVLilt1sLbfzS5g5k3PDaA7KQ6jQhFiFujhTrAv36fJrL2BPuxnU
Wec/7l8xxBbs1Y9BX9D6pPxB7/L3+79+yuKWrPIbYX34ReSqFEB0S9Ux+Rjld8AS5iw40S8W5crG
O+zXnX8iLHO69BW+SzkkIBTAkfd+n1+f2gReZWbpoGowS2aE+Q7EK+HAJOf2ao5KDuMU5qVDeDiE
R2XJNt4au6AUe9XHEO00V6/7XWedmqqMvKGp+IRCx+zkgeUKXaVpEN2M5LmqcQDpeRhVKSX4Z2Vz
oolXSS5BQ+r+kwzwLkxkFKYVXnf/QPBHA6eMLd0mr+DayZn0AT6FhIM9nCEer4KUVi4j6Wq01P11
4OquBrP/Gm280tIML4Wggdr6TqwOgGT5ivxy7edQgNDfuZlv255JpAyRXyCGK2dt4NhiizCOsMoJ
GUVuHjzVml7YywPjcpVD//dWi4rp+dNY4GkO+waLaM+K/50jUJR1UzxIhK+zf/4qCJcXtR5/5Q42
8QOEDcYfyVzH3ESGYk9LplGRkTQxs8CCu0InMnfuvhZCVqKXZYG2oNrTajaS7j/F8+MZCT90Nv+Q
2Iw2V8VDnhddst/oh+H/xTfD9rm3B44QZGi/7K76pD+McNsPkT8n4iKCX1eGYYlTEuR/tmKTFHLu
XFHPYXFjkowomsuOPInSEM7/SklFpu0VdYFp8DW/siuhoXBNyUn7VsbKMrTbUerNcTu2c6qnnW/8
jvydsBktQVM2xIc/HmZ/Nk9Kxvi9vCGLkA/70niBGAuNn7WZ3OHHn4PcYQV0be98IONp/zMZFmvW
gESJ5HsTBk8JOZXjAfb2Cb5/fBEOK3YnjHBz1exITwglbccltwKWyLOsrfxcxEz2OwYVfi8yBuIb
/0a/n49GpKDmQPPQE9Ljjg0t68orIKixeKzfNyg0a1TFlk7uluCtb5sltKBuIeOfgAeBLBbQMknK
3co5nb7oQwc+uyzOOISkgctyG64pdqxFKQDtYEYPaLDhsFDjjaPN4+qkvebbjELB8zkiCGHiJKf+
YbG/s9w0Gsc8YxoDnXrrUTpto2u90J71Mt9Msn6vIB8vLh/q8US1uI69tsqlRqyznV6RrAY/uApL
UJhTq/me4ssOmYywnF7IQhDIoEH4CnjmEpt1DaIxEUKT1wYwPSXvG91kfR0oa/xrQwU0QUK4dF4K
+mWZDruqo1zVm1kRFzq+hlq6bzR/b/rAlDIn6nHv1vpa3i7gOwQb0QDRhDdQ+NRk70czAyvyugQf
U8BpRHeu/pk6S9q7deKXbdD9+32VQl90gW8QEthPIomr7uzFM/w/cWbyvI/hsnYglGhdpzy8y7f6
B5A97fHtgMMzCktxVzAGI6ZBsVzzJtW2SiE+4plVipdrZ26IQ1d4nEWeBkVlCu4h7h9U7q8Cq6+S
lwnCk65oPVlVTU3A/+nqvQHJBCQo2VP6FjqT7AIymB5Dw6MUtrPeCObqhnLDOUFaVZYbuQbtdSIt
jyDTeju4jbDYmDTmwn9AvksXTyvM4knlNG1jXOgTjXv/VqLgXS5pdsUZp4pjcTcefM9/JcyjY81l
L7Iecb8nvb2rOYf7BG/k/Sr2RIVHzEUNzutmN9YJt84S6b/JU7BpoRyhaZHp47IKPBy3t5RAuMZe
lUKFDMGiyMxqckAh3/ZTHNqbrML6Uy2ULZepytvSPbPVUVGZPl5XJSC4p/OosDod4gI0B/LpfrXE
5Y9TYK67wsk5a2mSgbn4QbSSN5KXARL5yTGIBaJME3bptUVnYVciGIE4CW/1/JpU2mkA340swvLi
1fB/dLxVga6RpNhq8aYlWA8V3hloYrDX7dKbavo2uQMzcftuSAejw7FdOPsNkWIrHIoWCeVlEHxa
p0hZvR/HPGcYE5dJU5Hk+41dd74yzxSp5Xcr+HWSTiaEnhs7NrtAb5K0OEvFbEqNLJ7Wiz2ADVuD
BJHhW71DPDbXKnebPQoW7rs65LQYk+rVCNQKRxlLd1UqPdriua2JgsS87GQ96X7A/Y5Fz7G5ERMF
J//HmHy23hI18AjiONyRJqvTigZl2H3qc9S+pN2+fg0WBmPrbBHD4WejUDfI0905V+Vey0+FK5+f
gXYMAiNcVVliR/SwuG2rOig43s9RUzrq1W3q0nFf5q/r5o+JhGW9wmIy4EkzwIEvnsHLnojS5VR8
o9N6HalsTtGAyyDM2n8CdfvESV4r0YpWJ/s1e6zJiaPZ5demyV109UHXd9vmDYjRik9+aqwuNkkp
F6IiGuOwovg6W+eQb9A87mZFN5soLcrx91MTd7HVAjo85B6xsBQI2I0FccrZeTordQRJmlffiMWf
Fi6BaIy2w906rPmrU1VSCs7nPOFPi8IvbYQLZsQBCQP1XaH5ooC75/m6csf4wnN5PSqCsG7nXM7Q
lXTVf6yqi3oVqCjbrlol0tGOVkrBtlQkAH/2V8Bq9Not3eHd9YfFKGJCnwnj5eyEcp+8x3iLMoH8
pfl8zCCbNUOrcPuuee6Ah8L9y60Nk0JGsj60teplN2UBb3V733DA1quotfiUKyxQGKzLKZolYPRK
xxK70C5uAxSNVBeRcZOywQpowNAKRQ8Ry5budk1XTSW5m0XBTM8tmEWirSOyqOJJ8agqCI793wk2
ddymK9z71aJu1VI1FcvE2mobzDzheqoDRCoeAx/qKDpfzotfzXJAXWwh2S5XI/+YVuxo17WXSbiC
9oFTb7yM2cVf1MwL+5amJ0bkVwiiXF+5evOuzuis6QUJrEGXB7wT/lZTSGF3JC13MDOlqcO31xCS
d+MJep4yaqnggIcVLgQRbjJbeJ1F52UwkLa2lFQRKkx8It9CIupxv43l/ThEdIFCKEcsiw8pAHah
qO5GYnJzoUHwem4dwAsot5zJUr7Uy8v7jUEaGBUnJaJP9LPh9fgm11Aj0yU69qzxnhFh620TeLST
8y/DWRRj+ogH29VnTn0Wrk5CigXpF615qmIcoKIArumwts4UfhAUIXXWhHZfJO7Lzwo5Xkxu52g9
j13si8rHZegSL6XssrVGNizq71oyF0tUAMsNlyyMdy7Qx1ADIzXlHMZe/mEnh78QRw5r1W5Vuv+M
edvRzXJ+rCFk055kyCoeZw50nYNuN8VE4ZA1CXYefB8HCQLuTp7Af+GdfSPqjXF+6ylAmLxopzFG
XWMv58KXcJ3E2TQJhjbR3QNAOBx74ucuRTITrwNAqRwhGQt8/Nykq1fn5KiTHMlU4eDqcMH2hXT+
s2a/DIV5vMyxngWK+jWZs7H10sw71u3HAvkBzFyunYP/S5oD8VTHqXAtgir+/JdL0j+VTTnCad0o
Ns4mLm1vrhuVYODpwLHUcAnROtICRUG6nGe1ksYrgWmvlYbV6IbH4O+9a6VcURBbOggS1qKq7vhT
EIOzuynrsfxvcOITZOmFZ74xWpEOdIAd8k9dulosVlF0UrzVP2sLp0W/DHIlBgaju67a/f+a/OtT
Avs1mUfv+B7ZTistefmQ8mNkvlRHx1k+X8PtoHMWzBJf8pNBuVpEX388tI0Mr/uFqKz/tZPMkUAn
GtKulFd77cY1SCfji0DKbUV6sXCHYQVHsPugf26oVI+WvUHFIwoFqRWhASQoVDY0yGEEyjiP0LON
CVR3ieAPwYRWUbL1mAxqUt5OCS9RAUDaAfeKfQNhjehEWlHPDtWUdoDPGto6HjkISpZQ0lRzozjI
wkWU4kvb6Nfm2x0xJGpjYMETJyzm9rgAeA7e6m9/mxDC+5NwVqNIqOwqbcXc3+KDs5StuSzI08LQ
Pv8/KH1GFi2c5QfM9HODoMbUiZ07yl1X/dX8NcUsigzGN/eSc90C3s5D2rbGhaLKAGM3ojwhKCdY
IpH2waToZ7kOXxJrOhoxJHpOava+OnH3f+kB0aEVvOlUNSntLiqbrHr4LjsV5Aa4y/90jVLGr6zM
+YfvscUsNrSO7fPzNRcTFyByPtTwUtZ16crlLG5n2m2oK0kpwNTkhhp81rPsaGtMusTI8ydhV+j+
m+go8NLdrc7FKYm6vpIaq+u6Ci68KnYRjDzqOmkSJnDOk3Tt9J683QHl66BM98l88Thmo74S8pOC
3N/FsEF+XPNVd0tv4DiVMSgc1sHe+oMT2FDtOEaxfBA5xTDwx67dBunX5ETcxSZUeDYlx5HxeQ7F
tzA8QZINa97f5NMA+xwCy1+HPyJuK1mbsSzajXFMRpCPSDG15T5bQTYiixNwqQahutOjomD33u0S
rnt9pU7CM1jRSygzord6tEc2jaZA2c4MuZV+0hcXsaZGUgN0m/y31a+47P+gSu9Qw536AHsnJhUG
AEqHAgwpVFXfJwFHeOgVUfgwbcFTV6Pd2fYoVG5pwyoqGq13h7PvNZOYZF8r8syQHMewuH/Ns7oz
xPQW8c8Y5bwdNC4fmEZ6MhUdFJkd0JCjw+VLyHoD7jAXzTSWbpzDAXk6gT4UC1/ivsJ2Im5ogiC3
+aehvWGbsuIeNmU5LfmsOsqAHPAfDOxlDa/Yq9jw7Vx78886MX6BzfTJLzrznrG0vcNNxT1EhB7S
e5M/Qsd93KKbli5QGSnTXrAiPglEqn1d4tR2c9+A6qzulYNGvJFdJ7ZL2xEu1lW4kNl4M0GSHkf0
pBPixtyzGEI93GU9+vwQS7/+McxZgPYgUn3fWTd3brDxIIOfjEICCQ6qN/0g7L7SGjSq9QS2DQeH
3aRF6yIkgrQZWMeHajJocKgCKritSo5PCcTNl5yNkTjDdB99gNTfvewj3dBBSN5n7HgZ6RDVSfUj
gIX1PtPGa7sZoJEI2g6t9FtC23RXwGnM3Oo95jJ+g9s7SkB7EZUscAa7qkQSdQ/oNCO9GZgvgd5l
9lSvgxK1NCqK1xN4jn4fm+pu4ACHNH3jWJ4QUPqIfnlOx+rclpygLcUhtyH9OgTq4ChmFBJaOBsb
85i4wME1bhbZaxBcN5dAOmRfnJ88bsInBIpKJHotl9OXowL7EqSiSFtosWY2f9FvwJC/OgNI0McG
Zue8ViMVYYL+PUkp/pW6eoxnmqxp15J10z4CpO8VMoB8O0YelmKAU/kGtA0zXTEAq/vGRFRawAEz
ynydWt3l3CzdKp89L4YmLwUzlBksGFd0Kqt+1a+Aoro/KBZPPq+ChkU/FApPATjl+YL6FUkbJxbs
FG9oWe7+oJtR/O6fRX7U1zmUamw/CNedlReUamJibVfeoFRZtIetgDeb2zZn7OGPh2GwjDN2Xrnp
oN+aRzWIGTuc9B3Vys7uagfHx51zJQvBH9IacMgJ//cEINoWyZ/njdCSReAlA3tFyOLRDvjdOrou
7flFhkHZZLb2UxpkpuoIwuJUAaRZwK5dEB5Pmx8m7GG73Xv18hrRMeBFLocb+Hd5ixIAGCG+3MhX
QjjGBTnrvm/7B23gVDChi+utvzDmc3qiLiX+9ZvV47lrjPNuYUyz81hXfVfYzRy17KqzDvbr/Rbp
EtFdU0t5D+mSduhQAAOarC2KU6nH1JgNwrBeIdoHgks40Sto4S97QPUntjAvvtGKRV0BxEJKvv80
CmuwyYb1ZjDSFuRbvPRyJu3QPi2apup54SKAKG416zfHwzwXgwtBRR1yZBh2U4kktU+8N3Wf7vOm
COEn60KSTfmS6/Ue6SPVPmxf0dyURDdU4YCyLhXqsjvfuy1YlKLullS8uPIDBAppBZ85RY/nx4A8
F/Wok9tFqjEDyqbAB0hpV3nynb5M2qRKlMqSsTkTR29Bs7cF1Nmfy+MngLKUxkfS4hjFLKvbNc8E
Fv7n8YEdA5c4W2vWd8mJPFw84zQ69rmpfWlo4DfGRO+GhNyWBJ7MEN1GcJsBpEC73OOe+zMUfEVb
X+mnImIjIrfRzCxDr+Js2U13nafZZopoG7PxIidalCdvsQJ7B3V4sbbdYDIU8vlSUO3Mby3GRZFA
xLqXR0kcHehkOFsFCK60qXXanzWbE17BTwDy+e2IlGgHIEs8j+6uU2QrXMceUo8hxPkgGxHt8I5u
Qebl5ZbedI3oTTSc+Ue1i9hLc97DTQVo/lF0nz0WY5TVrDnQs8EDHFgmbvZvZyC6KwG2bnD6kG79
FRAUI0rBHnauvNuJkyDBsvGm4Jioag9Bz+XsnbBGnTq7/vAglu/l/R+O1kQcsiknMZLT0X4fnQmi
ptxP/1M4+ehltVOtH1Ki/A4OPcUa2P3eJmnfTNqjkgRqR0UR4MXd1TMC+ozCYUFlvGRyLlKFi1SJ
WASr54R/p/OpzP5UfHvV7xr0xcIFrI01C69WvkFk5Pz85hED9OJNY9MOK2XzNVCRxAOetf2hqKRu
15fQ50aFDsCLwamDEoMSbcrC4xytYSZB+PoIswf/ZZL32Q8x71MwVhmhiU3f7a9DYEkTl0Jo2MP/
PpNETene7coM7N3UYlVzNFoC3lFr7o5oUZZNTBTOx3s+kFTgWwGiSRs68xPeJemUngIeJMsZkuZA
5njAGZLwj5UVz9njxF/mzDGGOG5CInG+6hQtQ7yCz4yxcF13xxL9XGJ2JV5m3aeDpLWp63BzBIPp
Vm8IOKfzFu2fiQt97RIe3gZXYUuLo5JqpvFFE3jTpJN1WRgi6C4Es/oeWscXaMd8UA/G0GkX29bC
Kq67XOWCSv/bxQUmZSYDtr9gZm8iAo2p/jD6126J3LY+xP8ehw6f/OGP3fcuANDYfK8bfXzD8G+7
e4szF17zrPM+GIrZam62MruUNfrR0zHpc76BGrk1xbJTbObE+S14F9avReLe4ZTKHkHgmPkV+QIn
HWsddwWKRrGBNl0pqijIcydaRoRhm3G9jt9rYYTwW4PohEAUiWdbUMOQNkF6b3wnhZ/IvJpqFaSp
jcUuMp2gB5csLNZibJJlhCK/0u4lJNh22UhFHdfJeMwHpogM3PHFmiFEUiJo7DeqGU3eNKb0WLHL
FkLTJNPKUsHsspt/2KxzfnlTPKVvXRLRInGVHUlXBU4zMCPULx+FYNgml8i2srZwyOeSpwC7M8CD
buSlnsOpR/PfCnP5nMJ87Taia2shOPM0QZ8Fm7smsNSJIoGqLgyd3eMRxE4XIJx0O47sDOAQMj9P
hQWeLK7qXofhc0e79F3Hj6OYkA5TjBaeLEcYAYT2Oz4XQE7/xAzHKaYn7C0cf79doMxZwdtOJzhP
W0zjflG2D4Dkv4H+YymhS31hM2iJzO93+WMVsUI7beR6WW/ypjGkdK8f/aAgnz/p5qGISWtafYCb
4CUaXz7R1C9mUNh74GDJimpQe5FGN7nqUw6W/shuWtj4fXH6A+xt1qtbl88T8wsDKRqw9nhUu8DA
dWODovANIEnHvemSkeuHuk9ah8LTlJ3ZcbarWH755N8wlj9+Hvr5ShtPoGZ5d+hMrFPa83iCROjY
ET4Vj+dMt5lVZNqV4hi/Z3/ZTDJ0UdBh1Ce5BphMqdNql7DBenX57+cqWmIyMFCLmIUua87ATR71
5Mue8R9poPBYbfAb5ErnVYlsya1TPtx0O2tzsiu48D13OIgd/bzjMfBphmEb2+h24BNfwsmIS5L8
TDtlveIG57G0jc2KH29I+3DAvCtDr/fz2ry4vp1DeHOfeHGeFh8C6qQlVopuBFKRedl6LdGjtbdR
WeKHG/kk4yOWX/dzCkgmee5fksmkcH0/kvyY7aDYbJYnpj0iwecpYlnawTRjvkQ3ekCNPvEn3XOa
+Lfy320H7jxG0rhOfcPp0CKIIcu4W3QZ76FJa9QseRbusUNAoNJvM/Xcs/FVE2qCA0iraabL6rro
TjjsLxW/wj5w35CB3ceQ3IsXvkjlIxb6foFdkRkAbvdqAvuGfmKZc0GgJbCusUtmfGNxQHHBR27W
r8kgXuxn4qSmlWNul060nl2WuNKwVII09C9G2ekQa2B4c7yJaCq6tT7r5KrlScxZiTkkg002UTdH
FuIRftOyZFM4EjYWBxRlNgQWZS8PGAfpE6VC3jeWrrdJUnO7bXFDHi8n2G5pSzUkP5S5/I3WjKvO
c95FUa2q7oIcfN1H0YtIdyjBkJDOv6zxDwL8FiTrBNn3bIY+/TwDLO9u3TGFPhtuzCCnS5Cdy5ux
XWbdDqBpi64YVpFBnti63slOLhyj36Qku0dduii5lw6gg5kaPOEKdFVIew1HVY25I9zFEqWj7hXL
nkxnZG6Nab/8el5C2D6FyHDcvDWzzQOzdl0Em4FZOGMas3z0NI8eZcSf1XHEoXEMRUljrNyPcC+A
16U70Zf543ZzLqTSLALrySumNNOHLnnG8elIaaTvMlUy/wOfufDgu6M4yjRAI7U0VkymMVNSsozw
YrAOL2ECM5IgOosSNbNnkLDuGOFjcXpkMlIl5ce+gRu2slMqK9ToCWOt+DKJT0nWDLa2Jwmnr/rz
PlNVkF9N3/FefDKSe1bTN6Lb5AxByUU8pCjbbEXqdVs2sfsVlKCcN0CkjMzxOZ8lkOlUMfzNlTtq
elZK3kNxdPBor1R3Fehpt8lwCzsVLCP1arjGYIIjtnanwuiVbmVhhl329QAGS8RWDOGtyQTIJtY4
ITBRC8SiV04kCkaiSrhk8hIv97Gr/NgIEEfLtNgxEFE8ZWiyB7S8NM+nToUUvSfbb8+8kw4lUMox
4yTNkVU7dBYzTLt7CrpZOo1xOd+ZspS8+k9A748UDM0YCqCTcta6Jn4gVTyhqkCidnkjyDxo+EKD
x53HWIvf7LxOGNEeBPaYTozxT5sxrEPRx7Y9U/olgz0dLUASvu9NAnIIAGxgUXB6YordZMtLnwQJ
zcKM039g1oE6+Bs56His3jWgwyGao4loH+81vEK1x4KJvfjhs8OE/CZYzHLvyxE4tbLu1mwdSSGn
t6ZTw7dGPsHHmlTumUwk2oGx+ZYticlDHq6YSozYvDrNpqNGInvBZqAIQtxHGyeJ5N9NOkJBCGfs
R9AjzXDLtxn1w7zJwktQFMUYBrcp9AAI4k7809DNjCUb9cnGFW+inDL5hpzllIgrNkLkEq2CWTFl
ejsxBC/0RzWvKiLTdSlgkWg5teraA3fhIJiI9H9MZ0FdRbmgkfNN00Y5KAIvu9GY2TBarBbKBgSj
FnaYsK39e9tSm/fC5vFilP+Kp+BlERE0QJF++4Akj9Eq6pcUnI7stKm9k2SAsFkMVTKbdinqmJEg
TiDnUQCmQp3Nr9FLWGDXby/OwDLU2fwn2tc8AEjfctqb8vhr3o1BpIOf6/ySC3I7tvFLYCKXOG6H
UFEIai1XX/QI8wAsfbj4jIenyz5cx56wousrUW3ACFo+G6//WCPc+14TESURb7aHQnpW/jmwLUVQ
ZCKTyTOUV02sicfzQjgvDmC6CJBKdWnLerRnYQ6/Xk+oSSo9KdiJsfzZgM0v8fI7aatBnbPobw27
GGhQ8bqVBxopUQsDNIhGNNvS1HLAB5oR6WdeMWleHZT2LROsT6lNQks9uuMB3flwOfdxr7z/9rhJ
0ppxGZr4sqAOHb02eM+PuCLE3CtyOo8hWoKJLMHxIytdyWIpDepJprAiSaYeiX9dRA4tGViy6lFJ
+hxvFSpym8vasXlE2cAqoYGS6ZlE5ZzKI4AU1/PYxt+Ict+RyCcUqnZlw4aTAJDE8NNgkAUJIR8S
KkE/aqraa2FvCBtNfVV1oSK52xPDz0HEZrjJkK80dPMqW/LHVaiCYAXgUyRjNU4JU/39174R+mHM
Im8VAywW6jUqou+xgVBbZ/qeNSAkQ0g4vpdQlKtg6U3AlBUZjByEwMPj70L3VwxZCtNgyyoBI3YP
F2S5/e2EKnAJVU3DcUiRezJl82A2W8Hte7p/Qe2ajOxbPH+PnYGIlI7qta6EaxiUkJYOPjtLIve1
FVoJSYp8sI+ewYGSY7YjgDZjDzxsBn/XZjk0oxnDtLeAKTcgxe8wizzX0nL2RjJBMq0UHS/b2oO1
i/IyASQm+F11s0jKL/CNMDJqsV9dbhjGGaZKXH9tQjChv9EsSQf9tHq8zdBt8XSrZC3c0AeXPRu6
1rIinKK453xU4uRYHbwdgmSPGHnjlv/7pxDGaFm6V11DvCy13sajw6es6zenL1SuCNELlrK567H+
60anSL5i4ICKOY0ogmw48CG7oKxzHo41+sake8ZMlMSQwqhOkXuciBzOzdmvKlWHlOhFQstXXoB1
+sx8+w+AALjsk4X4OqxB8VYga3XSnBJ6QCs11GG5EmwroLzZxi1NrmqkRpF/BGVaMdqBYHPqgkss
tvmZnsOCuDYGF5jppJy7++DuOEX4UBCscNQ3GAH9b8B1UNYq3zGMYwnM6pQv1kFQyDBWMi+EfVL1
0DircXKlNSWQsDCYyGnZhrRzmFJe4/B0w4YJvVq/deTCBpGskz11lO+Et2Jz2HdNennzzbOoXnDS
f/cWXgyJ6DEQkk9IGMAbCbZxgJC3FC6ZNRqhDn/NmSycofyzxSdc/2Jbkh9J9j4Prcq6/San6p4f
blQfhxiKirpL+dzwIGLBlyY+0GrmgEDysotfKckOtxkvnM5O5gC+np+nIj2BKGK9DZQoKYs8AxMF
CvAFEk3g7CKa7YXwCw30i748UzHX3b9XGhAYakVmlshwi1rbfGkvq3JR7aV/ToLVCYXi7VpUpAAw
aQk33wwaueK+UEa2+pyvB+hhwG5l9gCWgnOliMaZp1hjnJ7FAMq5yu/beWeXKNGj3yooKWnpjZqZ
WyQFGPWEYqvX6s9PnqsxuC70g3xTXDengZCIk/n1EBYv2JphgB4oeKM/1U+G1yA6ycuLzouNumXy
jr2MErZbOioigbfQkEkpKapJvX35iANaku8f390Db1Y4+BuNNRkSWRSTAjbnuxqnT81yup6kn1bm
SIlDTKeKA2/K+a3UXNyux0IMIYxIqSRh47XglgDXRn9CQIMoBnitLsrytmOc8+/EUlR/3CS6D7fH
zSSlcGLGMIGHgQJeqxd/jAdAl7Z3zSPrvaWxeQUl8qdNxrFJKvMkja6/xapw576pPl02AJbRdLCR
Ru92Brsr5ME2zEnPnz4QdXiKBhQ3PzJb/Pgx/r0v91gsjE/eW06sSY5rueLASa8qvFMOeKf+iHhE
FOpXt8KQAnh+VYeE8it6L5s8yve/YWbuME1vyvwPGeauMi2NPb5xmelX+ca22mOZGZYq7pOZbZ9Z
pPU7ShZcC+50YeQ6U+puq8mAIr1xx7fq3tBmvNzn8SJHuS0KKTFr6LHxLmk1bQ2NCNFuoyD/UXel
i1FOTFbfwNEdHAOCnzEZZCMdX7L5OdNxrFnoPPbbKhV9uuIJkB+AFGlA6Th8AKtic5f3B6DjwD61
ZVGsTPoHxDYlluTlN7J5YlCqJSxK3boBs38bGEbVzwmFGZsX7ej76YWkOa7wCZWL5UU29m02X0P1
nhCZQ0MIhIz+LkV4Ebn9CknBME9O17NcKSBzfb2ptAIHWKsCfQFbGDix9Tuj0v0SJyCxQspjtUTX
HCDAgKpbjb89yLVgEJ0XtfbNTZP6w0o9S5SF3RAv50PwjFP5LZbZt2AB/AQr/RJ0tYv7ms0jNPgp
+FWASsxdBVtKwKuVfggkhbldz0FEAWpFDSiAqVFtIjMBRQZEvRhREensp4fSX89R1jBvjHlXQ8HM
DhfbmEYPZzRZwWpyC/zwe78gZCZue5oENvTqVFiHUMbDmWgScbyhANGTsFQxcqmsabLIRBbQPD1b
+4rbq+NTF+KrAr+iKyudqy3ZolB03c9woSoiRaYxW/sF2Ja6lEfPIafDxs9Idy9mn9Fch34HuWc/
rjsqUPW1opQ/aRGML0H9ASL/RpFTYyZa8C425AqOJiXfJPljds2McHb3bU0nwr0fs4QqsEPn6G0V
vdGLbpU4DLOuq/ixOo0vf+cWlgrYFzNDSIml0cOOdpoO0lMTJz1pVlFZia3EN6550vk5K/708nwl
8sFWpy7exzqtMkFt+W3zgT1LGVAlkvPt+hcXkT6gW+JHXKsgim/6z9rqip9aynIGl6qIeeqBTShD
KFvAuCUH9H0/XlVqn8TVHdPjUI2y2E87cg8T2EM+6Rewv+UaKSGx1n7GZHFLWN6C/AF3Z/k6Q7M6
q6/PJsWHjC15Te5mzvAoXRXlWn9bJdnYX3dRLkGprwnXi+ZBJV+SDFESR1K+GvSBrwHRf/UQQL8F
cTA90jmXBwuVxbML3nBOI5WqBy8n0mA6faXsw5R+AOLLp6+qOEO5zzCQefi/Ro2buhd3HMxhviOv
TIHTs6y+6hM3eNdcXbvdQigyFacU02kNpcz/4HDN2Sfyy9Pms4H0KDT2khxgDrYo2WSA3ROYjXaP
pG3me9TqBQshZj76rbjXzBm8zbrVgRMgIam6AsISw9wq+F+VhrEwDtKg3tV4TAL1OxZLYhLqwNN4
5suYCClbF2UpQaxnpukW7+NfIo+FIAVsff2EnfynO9lH9C4x5vkk5UonKlm5a/RbDAdJTitugsag
QUt7zlh6Pt9U6XIQC33tawtm+H2YrcIGC1BELsZlcW+NUseiiVJ3MhX3w/AbWXhVmhBkqxLiR3ud
gBael8SjPX2OyKJ0jPmRDsYIMJDcs/z3OQ5vtf3cjpcGQvWxQMEK94XpBOQUyfeP6gKRWc7Gwa61
qexmcp+eljHHQBcGIpPHui8TyhGJroz7vN080bIRk6nfq0ILb53GNdpBNYEdHWpAg+VJiCNocok8
BhFLZYqZWfDLCwGDlfpNE9PG8kApotRGBtBH+JCrYpj11QrUBIdWjwLpN2yc9aNEe6TCF6nlNGzE
UYQKS8q5OHSDW6726vDXS7kFv86DuKow95YPzgqOoyB0nqSUULI4K0SNXswYEstZG45SH6Oxn6qu
dLRuqG4Fidsr4lSKbz1Uh3Ak41/y7yg6T555nC4TQHTfiSeAsVAnkSIqbs9zQ3/TBpej13Slknum
5oY0RTmmO28/LNa3/yApKtmP0dYwvdjngomu6lWQK4qM9zYsfuftwMDfHasVWbQuBU3Z0Leh3EDc
2rsRVH9ivNOI8p0IOPIzQAnUuisWSqT1C7XnmNXLzKptZCzU/QS2qSYHfWuGJOEmUc9EstR15mgj
9INBxgWUQ7EFPudBp47TQJZTx29yQD1hlVGsZxgNyt5a8PcT82xnIJbJKcXPInt9doWhobxPz1wu
pcto0A1pIc8uEqk57VrzC/ff3zK5TLyt55iMxJgFJmE5WX/T1UsFsXKCeFqr2H2hFe4AeyCE56QW
8mVHdOnD0X4VUDB4UE4AKF3+QGpHFEBwBWtkAPmweqONBA3DADabspPJ8lEO2E9VSObRq1KtJe6+
3yw/1IuYjyfS7h/L6Tu70mMphYjqQGaM6h791AvCn3d7yc6IfkHzOrzbrOw+9ctMcJn++D/hwEu4
0UtR8zH6XsTDp30k843alrDjilHTXKey3KL8zoZGivzamF6eUrnEUeyz/mI/PWGJr+4qnEsfh/Ek
NBvmjk70KwrllkpFvkNOsZRm3/0HCJfJy5jHmQSrJ6IZHFS4lmQ+a52u4Pj9VIeu1ydMUsXK+G0f
i7PaKT3W9In/A9ilatd3Xh6P+mtu4c3MGZUuyOk0NzpzPx7V4FolDFTgxUT47is4sGoC9dPfTN/e
b4+du3Ey6ecRALnv8PoENUTqKOW/iNLt3Gpe2VK+PRKz2Mf3Mn0pCJRfg4H5EE8sBKhBZFuN8Cf0
AdaJ8k2sg3+kMBSW0kWUypia/i0ebH7xKOjbdMK7msv5M/cFh9sQRH7otxlLsr0f5B/x9PBn9niN
aZP8OP1taHbCuVHodEEi+MBUcH4rXLHSwRyOLvMxivdkNx8OBM6PaOMx9OzsB41ZQyg2izLIqwoF
fFWOjNzq/PnzeaxcvA1S8jaV0vOV1m3grlhvNz9N/PO5zbcM6cY1NMyv2mjYbm6XrIy8PCKDJzlj
8oKXt26vI3lj5yK8+iI4Bu77s1hbcm66MyP4oLtAUN+ZPI49NiBsNkDvIMIDy13pdW6o05zDR2iD
RFqW18z6XAky1y0BWvRU7NIjT4UoiViPbHl2j+t3IeS7pBfPRFWDQbofNN1jqcEazLWzgAprmcBz
CIwetuxwZlOTAUXJ97jixPuExuxqPh78d8vmXVCP3U19QXqEFvcU17ygBRC1ukxS1tKCmCI4kMAX
0P5oVltAugDF+sBrSGIJfIKgoiT3ILsi/R8ro7/uTP3sY+YpxtqUNvelDbKMqqmklo3B7DSajCP+
ZwwpBxvHVzxxvzaHphGMrGm+QwzNwyG5jxP0xBTTgoDCJ5joYMgj9if34KDWzczJr8N1NTgR7zYZ
r+Q0pwUfG+qucIL3yxBGsE+fVIpmOx6gOrk7O65LBlj6s40opsURglWpv4OXtIMoAX+KqHJ9nRQg
SN/h7+ipzE8d1SlllifgeD1YeczMmxiPTJqzv3DR3k1MtssNWnFUT7ZonHjNBfBjRBOK4o873f2y
mZVhFSZvYnDbcn/vQSfsu6fNIwJ1mTLN00VWT94a7gDi5twJlxwMln7rXkMgxR788YhPLFFtXLHX
/qAORBd34aH8fR2zNeBypeqTn6Xm9HTQEFfuMuLBM9KJSaWO0EakE84LdlLcJJm3n7ce+kuFKu5o
uteK8Qrzg5YDI0z0b9e6wbuL8bnrbcthiISaX/OOMam2kV40pNZX9rkszJus9XcoeVSgzHFjnCSi
GLWogyoxfyp7vLiN28Rw86zaDL4J4HZp1Y/6jyZ8M9b+hhwwUUW48kSdhbQhPZaABGGMgTtXZyBc
lykUCt3DUiIhJP+T8JBkoPjXpCduB4sLxBTiMb5C2IVeUZutkE4f5aAgEvqGnx1IdCdQ/+9Wv0vE
/isSgR3l4g3edFh4v4dTV9XdtRC/WS3I+sRdt1eGfxiwADjVtJrMJBX5A27AlARB8JGn3U6U/B1t
Ps0XjbwndAf18tkSh99VxvNZhplciGMlI/XmCybNggLDZpBzBqA81E4juRrp9TtYAe3uasTzwLC4
iElJx2mwCIx0MZAej/iF4O9+KmYNss/ScYGrkWWFHofhyMwFwdm78wY+msXGdjdZxz4qXWe/s1HT
Q7ixoOhtqRRwgGJC70C7yUha+bwcg70PeNrF5vCosf0+0l+yZePkMkj4ti2XPjKkBzWC/1uv8dNM
k8KJhrYifT5+JFQ+xCT3RDtqB7S+/6x4K8hGmcG61ERQcEpNDyBk1EIs7VrDYwwpC1Y3Wc6/eXug
pN1SjcvGD+kqkt8UytpEm3fXEkvodoIYhdyTPhznNN63j9frt547qv7Lqw2iOCjF20WeK2xzuY46
A5Sw2i2wlNlJlY+jST9Fg2fPYFsqdaIcstBmvaLSg/wpFzpGMYHjGlMo3qATvmndMujHb9fdnsKW
XqEHujtiwiBAV+4vbvVnEw2GaGFZyEXClByCLk6PA4H0XQzjt2KaYRAFBMVXZkoU+Lu2fV7dW634
PdcWqIkub5nTZXjXDIbuAvDrz0NpnMISD4ujmcsaIdm//FePJl+N0kSzYIk0704i5SZPbUF1ifCT
BM7DsE5KGALTuHs+obWbKkilUadBfvXeAasB4Anb0SdNbngS9N4wg8fisuWovFuozWIkHJxeB7zL
KHDkye2ntIl1QaadjIEhSSf7+okSI/0WHVYZJ6SvDZHaSft8a79eV9ljh264jZIdvRw8gtzGzMja
LHFbgLIt6XId3+kQzybNUmytfjnLq5yzj6n2CEYSpJj8qd0XZIIZQ6MzYa3uLXl8TvW94MjDW3VA
bmBCtVO3Z142CyuIv4LcDb29mqDFGmQNqXpUC7IuzmXkNyBuNdF+RHExyYRNrSHVB1Ahe2NmMgEU
LyPPrxd8yGTcSburDyPJFleHhK7+fwvL3EDXWsfkZp1/R9nZAmifcJCYRQMM2vlxfrQVZaxSc50L
T5uQpKugTvOBNU4LJtizoDUXhLrgxVn5K1+NpXGh6J2Mp7Fb5NG/rKHcHUUg3PSv0YRB+o5mpIli
7THRnQB7TfSBdaubPlM1ORXKkmNUGRpStssQ8+QMMEkWuQbFHc6DOmaDpQmWMIYBBn1dA9TT00bF
ou1i+UcqQoW2NUBqZ/VHBDllpXY9GU+VwzRPTWTRxkz4FpvZy/nLst11ErX5p3So8A4dPekgGohW
GCLUo5MjS6Y1B1NA795CLqhaUeiX72y2VHkYkfJTa9C8g793UFZPqVhxJRBh2Ogg6YlszRMcsRa2
s4DjrOW4/OoY2Npx89JNW0Y+DuXdLJIWNyWqC+kW4FN6HxhO1Q3LwxE8qYE2811FTf+G4CQYQl6L
1QxXJU7eyYLbKNxG7Y96Mi/hamfnSXnj//rpviUmtt+7mavB/puDJWF3NCz9cSeqY48MqWrDPOMf
s5nzXFEXk8JZDFl/WqYsg2wO832C0Hmx52iwm6/2oMvmP4k731eF4iKm72ERo04PoTmvJTjCREsj
5JD06SwCI7cTBjoYhxu+yMXNHanFgVw8e57moVwdy4daXKGxmup9RNwim6RfUrAlx+G6Um6Oqb0g
GYYMFnL5P/ZR4wmJhWUgVEd35qw4hsuPvFlm+f86LWMBVPPAzTvs1uOo8gso1yKj/9H6lYthbpHP
UKVi7PkCqzjI1gaacejoWKn+ELEINUlBLzmMMpFUfqeqEhHEE3UCVgB5BwOflTmZWaKjb8Q5y8sm
FbJ2HRqYCYNtqOkcrxW/7ZKTFSiqVM2TbPaoVtAkZZ6AejfM03+uRKW/OrWNyOC0RbYQTDjJzYQr
vb6a8n0ljG7ZATV2eMxEzeuk/EqC9UvDvvX8Thji/xkY6W7Umjsp2krVHIbFvg0YJ/R0XDwawXTo
F2oI1xchvgRCAQwzbsCwTsvI+QEi5osI1z5PK7j+0Oq//wWtgS+LAYl7dD4Q65UDclsWitDofcRP
wWLuxh+rBQKvEdVp6yg76jRr2kq+oJEzr4Ng76ex5kf4wJ0HCtQSWlwitvNZBR1nIf0tcu4vQl0C
vAo0AG9/Bf9/v6Lu2c9E9xiAChNVLo7M0KiP+5+1ttmXgemrYjMjbugGMK9hv6EN50lFgXQ225ye
eGRB9r+jtuNpZNmYDW1Om71e4telv209npqnX3LXM9Gb0fYcVsZfrdVW8Otf24ePjhthNA5METoZ
6+hUoNNrrnmuio5/hLFAYVi4bSTgYz8BmbLmz9htql3zXC7HKsN7QZOL3oF16oJUV1gZpyqsh4B9
y/2wOjtnYKcN2seRpqmMBtNGexL6kQkoC+9uAnGLAFRiR/yVF4+mK8z1Exf3++hRciWdL2Ia3JGr
XbImpT1MgaPDWYMPCSUbJtjK4d+J/ccPERUI+KklDjzbLXas8qH6ZzAC2UfOFat+w+rKY3gTfCWN
rB5kDGlMknan4IqlfrvtoJTwEmt8CR2818ANo12LYNANgHZ9c7MJRw0ecuEifCxD/rhGXA7JXK1/
pROeFgvgR6FDUQ86elBSNdvwk/xEM3aToKTXGEOqLugezg62iRGmWSg2dzFO1NMJTgwxqZ+WEquf
cEpfQyPHKlQMqWg77EAh7d+RyEEfCsiAmeov4w8Q8RJ5Kbh76J0pZIykESuHxTfjopDqOsme+v0c
wbz1C/AF+Gol6mIRPugUd11mW19HtRpB1rAsrkxvkGug5Xh4SHVPI5V9o3J082PqUhNh8AyUeLMY
wlWPzyz0A+MKhMrf/4GjYWltZt8rKo1YpveEKwPK3o+sviiwfvckE2gjrc1I7qRx1L2lNBIos1tr
brjCsh5FQzmX1a5UlJdl/IOW0oHm43+z/BkC2HDzbjT2sPbaZFx6Tk+iuwNMLHMIu4bkiVL+po12
1Sf4HijyYiSRkLcTlEqg9ArMVwpTt/Mwgnhgad7uYC334h2Wgn4/EaRkG3ORr/sQqC+GZVrNiW+Z
wN1MqKXf+XzB0qdQnZ/yx8nQbYdv5bwnwiGa+7oCHM5VXE09VLZ+5E/kveV5/pfXnGDv+bPrO97X
J82U2n0ZZIXlzKDXMeFytyMrT5RSVDWwfh+vEvl5LXHljk8b1RSJRjqrk21Wg8LkQWxSCVf0jHaK
0TGs0g4D/ICA8FnBve1hXMzJeUxXvxvCz0DttwNMZF3sWV7A2Jt7BdSylfjOZ5gATptuIEmrx4uy
2ZCZvHCiBoIOKztBZxmHleuPmhkwOijgqXQWbWgKcJy4F/k62VtxUu9JM2XkIXPF4nttibbVQ5OV
DMj3tPW9E3Ojx9GHsW/3ze6IP2OmqMc980c6TPco+7GS3CVZVazEYKgcMhMXXeguLU4hISpqX7py
VDTrfpXlsGz1jD+dfxXxRDH/IBvyfpbI7k3K0MxvlBKOZW949P3tP6mIi8CoMmn6LF/gtmGrEMAA
bTN9CaYCDn7CATWZ7+yZfLQVlakee/RquOIm5Zpq+SwsqPYZVkx0KIck7lUar+dqiu2u1Pqnwe58
S57/pE4Gdt3+vpu4GVN1QGvzsiJHB0h0cc73Quhvk32UUGUcIsB3ntB6fuwwt6UX7t2/G7DevwsF
Jzp3PknkkNShu0jFbh5MThmJPtz027rVqxApRy359lm8ZJDWKdhSUxD5qmPZbL1lsttKwZ+CnMzy
1WBCBVqjEwcyq9QrbQjo69gVtH+1/Ii8E+C/6Qfxv7QfJ2NgvfU4OhmI+HNxZgmFFfRAW/JCThq5
EHuPJ2SwnkaEDRaXDYnC6eTKnM1rXETpWrXXI1Qd4/uTfGAslrda+0izpfjCsfw/rBMlccTWlgwh
HAvSWqNWpzkTX8MrH9TOLe+zVKix6Fc5insnt61tOfBWlackwy17I7/XQMChM82XKhdOwQiy2+iX
PwA222TAH5wd2EJbMfjhUcMfZZg7vFTGBOEQ0pajD2xlJcaOFTYgwmjdDuw3F0tGaa2gb1XLymzy
6CIOL8W73GIAj/qS/S2HFpP/mTgjoSCh7VHa3TQS1vpHHEz4ICyNAR04gUdR9g6x1kfYRhURl+OL
aXwUOnUw6N1PIcq5AbAhSPMRXSPhze51xAzmuGRXdxyoi8TURXGKXcg3lYveENib4Lw9R4HtDCDV
I0T/VPbPoeN6B6Xo1+Qdmbs+vjOI6hUqOH5kxcCehN/pf+6Si1YmxiGvfYe2QXhk/ILZk8UkUW+E
ajON+SgQ8XLWuOWL06MbWUcbfceNiEXm3rRkqXWxA6ntbU8V/aCgniYD8w1/QdIdBAOVIHrhIVq9
ncJgb2dPfK9kJWAuRuOQIWz9t0xen6XG/p5ldEv/ZA/W454mfsG5Xk7eHi53HrDqC1ZefbEAp8Su
8o9Qe+EDEVVWAGG5iEpePaybZ9XEA1AnHA4lNAKLjQDK0xw68Ive2iVzfD9NnWAiZzfNjjiLC3/W
KdbHZ6KCsk+LULQ8LrvrMirS2miMRRrPicoJMRUBvDhyFE8R6yjMJDoAqkJ4YUz9OOIxJQAu8s0e
o8cygCakl1cHB6hFrZWejvo+licniCeJA2rF/LIReqSol8txHg4Q9NkrPZk+Y4tVC7OZGhR8x+G2
qRHAITZc0EAgnGqvRpsH0HqJWUDCb+UeU+Sxb8A5l4PqjtVAEyvQBypEkTS1HTgT04dQCx8yibMe
FW2WV850Pk4w6tcM24XlVNZivPTfV+hTG+/Q9xPy3MuQU748j7DCUtx6n7ABVN3pFvUQ1PHZgnM6
25NQfUEFaN0Nxjbzpz2sjEojhBFURtIURtBUY8HG5iUfhXerY0hQDb45B4bM8oboumXUvAE0g+O1
AVaZDV3aLL1Zcwr1RDSOtezz7H6NmMq0EydsIhO4QoGTI+uztU1tYEuDFQXeWN5CBnkL63j4cgsG
Ta9xLtEyJ37St7IYBfzHLU2AiMhLTZYhqll4j2ahluyViJvwpDlr1LMOAE9jPbqyqbLn5vVjW0Lb
ucIucmDZxY2bod5D9TXRKmxHIZyeZ7nqvrP6Z5Jhw0H/3v9N3L7c6neWXLV59XeJUP25gfcElfOu
5kzT4tjT/4jHFd5CTyYdA/OL+XQJiMUmS1L2KC80KqLhkiOH9ZesYwn2S5z9JXYuAhZmRQcP7eGV
e5XtfWh+Dr9JDYpSLijO+osEqf/IOCP/xVb/y9YVtOKRnLTltsP9U5uXtzytfoHSN/C4VUbWtrSd
HFdU8k6MohjY8L5zMHlexeGbEetR/va1wmNQ7WSjI2dh2xdrTXvWDTim2eRdhdUBkZ60mqBFIMqv
Myd4qx5YT7TMtgdw9gWc8luIViWFUbCIIbVkwLaV3fm7Dfx+1hXlOcbhphKeQgr1RbC/Xk/bzUC/
nGhC7zQh0+fLCO4P6ebAyzjSe4A3T67JsIp3HUZlIuFdC2gtlu0rfAYmrqyKEPBKmIiY5zrV58cJ
3Cpbpn0Bk2xEv6TDM/K+L9PnV/JKQwjIvO2c1O2oQ+R+vyU7CUPeTAJwj4HHIxM7AXNkmDSsLsY5
iE6V0XWMKpYzcdrmN2o5+jJ9fxHto7p25/7+4zcGJ7W2da9H4a4u5qb0nbF2kYaBax2OQbJm9PTc
ipYgMETPNHzjigbH/4oiUgH11wcB2tASmS3fiCv7m7MStBuRbiMFcisugAQlrwWa1Vsolewaetp6
f8GhlRg4I4rsHfrgFVsVdYV+h+05y7IxijK4X3WGVOV2Zi8MYlU+KShXM+kd6/mwj99zOjiUbeio
1EtlbGrCtYhLp6Cel6rh9FvWddWsAZF1TksXBFDgKawR5T7rJcbWPhBhRYiguhzPwlHd+gx4eN5m
rOsct3xAyvNcNKOVgiic6TVI2Vmd+gJonAOn2ORfQdFTUZd2alvKgj9+NyPbBKAGzkSPFaFJJ03M
Yv6KSUSVJf2BXUEY51oY6/19k7rUHURujQtGl/GrW7JUdOZ6Dp+lItrDhSwKQ+3eXH7p6JqxamKJ
HIk7furqbV6aUB8IP0EZ+PQZQiyUgUhOr66C5Y4RuYJAs/zPCWNS7AojYdjx047MKZge+FZHHxgE
wqDrDzVkM5Ox8hYxXmREahYuxIJn/W68uPl48VlZNbZAGy89bTU2aFAV3z8EtqfITVIFP0F2MFwi
hOz406nVtF6AL1f3vkpbu6/axmxDwPwStsM61WBDnRCBv+IIvvDi84yn7rZgZpjJKm4dDbMdCB/x
hFAS6K7CgjUhHDuXsftld2JsvuZKZKFAgXlOYm7kLFJC1iUA5Gk7+sjwjaebN3osZZl/qXdgQgj/
Ud7S71T6PRyQfI5V6BZbTT+nSt68cL0twdFlJWBJhH+22f0YSnUN9qf9Fm4vheGNMJfwjIezVrR9
Limihg0uE8RUMh38F2Og3932nczqrZ9HaDXD4GN5NenKhDslbBYQD3fen4aBNP46B+uQplK0xjZA
AzDIafzbsjPiKJTiUDFs5+5MnBDCMuCO7mBMJB38pilxP85Zah17efcpTADjCRlfzCbdv7ctY6c8
habCdmYvt4kASp76Aw/GiS4uSzb2UKQN+WCiQbuQrm42NBuP9wzwffzf6w44kUn6fvYDLFRoSK8i
W2eLl6+1vgthLcYz8um/vm50LDU+ZV2xZ1ipSrgy3zRD2QNeD4Ssok4myTlXQDw5ljB3czyuk0as
nb5Q/bSf27z6O+qLPRfj1QM7kwJCysGWOerha4+Vc0swufm9MOBNbRD12dH2RTDzLKu1nAWnMKpT
OtMSLKrucA7mOg0pPMYqpjbjFLO6Q04Aw8EjCNYncBPY5jXApPaxjbKLkoboqR3/syHhFAZ4Wsol
HYhAdPY2dizxfZuzP/PS2BBP02b0VYFwJCEJ5Bsnw2dUCcX0u+/i53kDf7pNGjTZfAmYo3dpG/HP
Lp2MzpHjBbx4Yo0XU3JauzOj6puVhQ3v6ppqM4/tmnKhQosLXPL3ZFwhdjqlBbSlONDliinmK7pM
fBTLncnaMhDdwxIhTBinPPckHj0WZ3G/hoFOoUmoKL7/twIeSt+71oatziLlcdvotTKSK+smlxDP
17c0bR6LoYaXu+k/TQd0L4rc+dmJDT7MDFzc2w0A/DotEjraWjmSo3QDGt1GxPqx1BL11MVpaPep
RMdRaTWkgegxac96HBhdBR2ssSCliMnGaeVq8dPmHqWVAyvB3nRwpaQxhbvRkepmV3oUo3kyoNw/
8ci6WxTJZBUnlJ2zxSYUtIiF8QOx+YXru3PTANUKl8YSp4RI+7sfdMmFgsamRGtmNdSpmTga3BGG
Ym3BHmASQNCPomm+LnSuEJgKGaMpMI8PfyLKDtdmMwJE+ng9rRZ0VdliFhmWxcr9AQBieCa2bap7
Izy2QXR+00G58rPotRxgpvtM0HIWVOB/ZzC2gxFm4pwvOEveDUEKk7/T+DBLkQpHYMdMfHG2il/4
TM1y/jSzVKWBbJ+bNMOJ2cH62kL481lj/OoRco2zx+KHmcwSj8DxDL8LMfnRfZV+uXAOPRBzCDJ9
Za2S+VyJ/cDClrvhRBkxKw3a57+9LrI9KvUZViusv9ZCdHzexdTrLg4g9U22DKafHbIZ3FIg7f72
kpZmSj+bR3qABwblqirTbLKRYoshXmQQ+YonTns6GJRbacI6rYd/1FNWZWzKG/PBlJsNy5EL2Gek
OjQ3wCPRoLKXgSbBMv4ZhRUT1DKFz17trf69JUSXSzYzh1p4SiE6UmERn/nBcmAa/eZ5aSRJw9I6
Xll5LI+7z/uglBJt+/ThySbGRkUZcdceDgLkhwhnFEk1lep/3CD3MBSCqVbY6TOU/Gml2/DQTd/4
CfnlQpUvN8OxJtm5dzsvico+ltQLxNWCvA72/ZKt0/sVKhvqDnTCOboRseUfidZLf7pQfOnuz/eH
KF3e0ZQlAByiP0QAywc0vIZSSglUs14bfyq2ED/EGwcrZM6pdS3OTeFpSLXXnL5m69xkU9leA9FU
eq+ZoVDZdO+l4il5ylT0hfmTsb4w3V4c8p9yfZB8PwuCqw2vNfC+1ODv5wQU1AKT2MyaAnTm378M
Emr1V9QsP7HsoCHNF/3J9h2cl4uUgYLcrkhPp6JVndaUrOUBTkZ3KgEcjaN8VCxBb2iYRspWpWPN
Gej3NxmVfNrAK3p0+GtDgI0oqejKzcQdNEPcgIeM0smu2+gtAbxVT7zDGOX+WpY6T4CQS8sf+x+N
bQH4u8E7v10CWPo2slIWlLGGzhfJbLkWpqrk5tLv28S3KzgRjAAErDCobYCSO6uJ51Py6p2nM1HK
HYGFTi+NCgSYl8RrrOuudcmH/Zb/Z6lYx6H8qimYSb5TGaryHOQ5VdewJ2eao42H7pdagteiANMY
ic/AvPxtITKt2WxViJH34TTE4FdTV7DkSZzEtCPSWJn0C9Ol1/5EgRUu5UFtXfQ4tr3r02d3QLwt
vjep59xd2RmTlUvOX0ZaOaqGsBktCS17BhctB3UmFD3u5gR2tt996tocBzjKpMCDETZi1UHQsMOT
kBaCrjyf+y2ymwxUIfs51WngY9OEF8E0NKABv9UqRKL9XMpcnM58WMpapduynGzhOgs/TjVxrg/U
1X6EdNil8mk3O+ER6ICeEMS6WOnxdo3IbYGm5szifFB9JbfYmu70dWBGJVOkXbWPk5c46pVRVb8Q
IO1x47uyV7jAZt0APRrtgRdyxafNRboDn3PAw4qGqTL7RWrtSaDpMxkpgxb8yQLdFDa90BUL4C0I
AzJq2woA+IJ8qURm+yMmQ19UDJ67gRfnkHH1UTonlb2ZxdbBv4Q9sxUsaCg6+yeXuMvUvQY0RcrE
qIiCJSozWipVcuUjLvskCwlpUvDpgVleqVyUZPFL0S7lhYpbY8zt4x2CC27D9n4DdgybWcCAzq/d
jrab68axLSN8iknxEwSvYy4DK7/UEu7I5BhyIqZyzT+ab5xG40ys684VJqn3gJ9Op4HkNTFy7ckZ
Y4OtjA6mugBwpmdNkPNsYOapz4Q2JoBcrb3SaOpVVCKG4tJTgUBc4C2BT0x5cIDTTaQrjeVuHq5c
g1ws/w91rFv/Ted81IvgFVoiepY7gRs2XoCavhtg1MZyU9tPaTMDAH6lQDvt8fbAZ0YDVMff7kpY
erFm8Xqu07NxIbNCqA+6gGNJB1vj/AONW/7gjB3bGWJGbpaTskL6f1Foz8oynSdm+WsgIXDNBrTm
XS4YP8QT3OKzO/wFGYhAyTpXB+F1tjj5oF/bEPn8pNo5BT48Po7yMfhCvyQKByfKFoB8pWp8RjRH
OpW1n9kkIOZ7kdHMJ+YQyTvS5D89GJpiGoRp4zuR9BTE2b3Q9QNkbpW6tQ8xs/xq3PqDIyQ1NRXB
/pTSmG/IyqMHhNSez/QmIiq043CocT63nx2svGOa9MIsQxquVYl4WrwHr4l68sF2RLVnxfDugSSa
UXiMXQnxeqgpMUrMOM9+bz3bjQL7Bkb7VgPe51RIzZuYj6jOmCz6UWMKjYek6NH4LOKtBiFtiL9Q
dqkPjj8wnYvNvR7ijGrOuZpMqDQiEpfdkS2BshfvW/YmrTNJdA8DwygJxAwQ2LYW5uuQBN1nhbM5
4+qLD1TsjOal7TKgyFacEl12PDJbL7PAp8n6d+w8FlglhkKIspdenhoqlV8v2T9L8FVQT3KeuzPk
aIckAe90Q3RCN32MghacwBL50XKOc4gFCOjLVVcg/JNnzVyErMj6GrWeod4uoBPmRzS4Ml6dQdxP
1IMUZlPYXzTCxN61GDjzRjylr0USzIWVmWIgFthsSuqTxT83HhW2r8bYJKdRqU4Dj29jjHyb9i02
5usL1T70+jRMNUbRWW7SU1ptGKiEP5e00emVz/pma7BxkDhhOwN0qIZu8OJkIUhsoAe0TvuCgdmg
puv092b8ohYEzW64VuJvw2L6hVk72OSCC6IbCKRTqxAD/Y0ffzY9zuJjwj/k3fImwoKByh4nE/Ld
lxUks7YnC51sIKBKZ5oT6PnZx1DzdRI4D0YZPb7udc7Uul8CXlHDIkyVcVIqNVIhU+e5TeVZV5Et
litS8egEVSGBQ47vqvsd08ylWKPBksgogNEdxj3usx5F6g9kPExosUVCM8OoTHdjr+dFQ2fcnHhL
TR+9i6/cWrcVwzWwWwYKJBJRA5cr/vmYbZ4D8Y+vyg8zLNMm8juMVn+1O7YeC0jVjl4SP6OXRnoG
SCS1Tuh5bUCZkOhNmll6ai16UlXLnrinLmrz3bTJGlX1kuwyhTfchkVWtkTod6jlQ5VLYMx79KK3
i8eXw6VSwbcH7aLb84txCT5LA0eNI2UOSEBVlhOyC15KEYzgbWQFkjeEGwwgr9hjdH8QheRLMg34
ZTGkwXw0iPZoCQ/8sm0wcJmaqsZu0fo35k88Rl6EeBF8ZhjbLoyLDSp6k18WK0jDY26sz7Rh5FnX
Va4FnrvZmgr7MiByTuQcSi//XonkpEfLPEUa6S0zISFMTJzSe9RiSzXPDN3QB3+n5A5+03klV9Jn
HeUbBlcxP5aUc7Nd+1AOExPfpJIcRscza/yEzMuqVle+DmisNvon38sORyPfMU4ocwC+cqEet7sh
etBiLxAhYiBYaOawG8pIc45NHUze86w8Wub359Zw+LnAfoBT9Ux1P7VDukh2OXeb0CT3b1/EtqhK
4G74d9XBxC8YSjhjFR1FHv0kCtU5btLbgkZA+yUK9+nrVkdnldcq0rjVwp1rPxrQ7b1g6qKBFl/i
eTdQGuM8onIzvW1t64lW0jmo1HZR6b+t/w0Ckasq54rrn5vHQfi46D29v2srSm9mcV0i7lW5YSHd
DHUEX9qAgNpYmQ7xQO+iDF6YfK/qnjDHEklj6psWDvbkWlrC95sKIdYBto3fm5sBNB3CnrqDSG2o
RhfkprkAohyYHKwi8r/u6yxDoIi2VerJdYFoESEmL8tYxWwcQAnf38x2tzQRP6HLnCt+C4S+j0LC
F0TIh9bHew6ZEKZQrVnQQgVG5pSHdxj/3eZFTh5E8sR3JSo2NNxDunODy2IV3f+/ow8lv+fnuHeD
mXSRoyfUVyY9wj/xKrhPG7SzfAxvZtIZ8A+4L0yZRBUukmGnrPto3Kc8nPrRaC9itT1dP7q9QyRu
sRFShX2hytthA7vF0IOaA69KukU0cIRG3EtmNB/WGM19gymFsaPkLI1Riv79ePjsbrseE6WmSAwl
FvP4bNCxvzqCxK0ZUseiCaE6Oe2UQ4zDfvPkyxrGWqXIBqLWD5CxYlG3K4lQyClfPJKOQLm2elfx
jdxIqGhFoUWag4izfG19B8GNnVmSH0tMIWDfY2d5jDDLWjoQJQsslreIt8aoFZ3cHNvz+NxFJPFA
llRdjyENsk4AGRkI3q0VPQNcnJv0dN1WDqyix0MyCz/aB8FPoKPPMnT2OI/FLJC+6SaY/jxDBhG/
wbRIxQ2lho8Se1g0J8EUwOL7Q2UpSHUHKMTVrWAeBBh4yjkFBVXOgBLpqOAvtRGjVGwA1lVbrAD+
pUQfFwhKmJ/4mBVggKS45BTr1snvOPpjcW9FeqbXz0LZcOfkPUnPeTQ1Me+I81xmAxO9B+krz4uC
4l4uUo4eJpC51t/NKeMOKbB53FEbNJuwR3YEKOjtzWjEnFF80ujw4Ny/wN+8dsHNxPMlCM7pWoY7
5ffe1R11JARK6EnAlMZVIUy2DSE6uhSIYmRuaipGs2SzZ6C8RVY11x7JQahL4dqdFPXsXzF9fI4c
kRRoGEG9/jbh1Y3D8fIT94DBpqFSj5EV7bQgrt6swSbmrRCdvHhlnVxACgJULEm25P2Sb5QWF33V
aitp5aifum93dtLfuLH9iNX0kIQppegC4u3Q1K/gSM7r02lmc2oilMY5qLeFsx677HFtnx/wp9np
58UckvSdmiqLYM+ct3K1/vNiGa7xUet5kjFHEoACWpl91gLvo8CmheX0hKHRF9fZs3k3jyzHBhUG
D7DGLNeORZ4NZ77EVCnJgOnzfJRNEfrJp+djPX1fA6LwzEr/Ty9DYOi/7OrWBoQpSpSXOj6pz2fy
w/0waeTL6I7KoYTuwAxtVe1N9RzVFEXIdVJoBdmMoghKYm1aAUqGsBMfKrQtFqa88XZFlti37Qi4
7qwjT2zV8nRfHJZzeOuasq/Dk8nUel/Sl74Q+GXvDt1lfv7tYF8UcND31G4U/4WcoZFwEgydu5Wl
cShdXye49LRb+hXGA8kvU/qtdmDcI0XhlV3eMPpZCFpB4H0qHUkRnn99+EWllB8qEhf7LuqyysXC
54J66Vw3A1U+sTKZsz7S4ED1/H0qmPn0Lry0oaWVU7UVzIMiRnS/GQ4gEZ1Z5f71V0PpnWMyPSGS
N8FY6MiWjXFOUoqf0InkRfcPOQSZc1rSVw4f3VMkdZjQq+5lng6P/TWfkA4nMwzimwzwkrTKtIuP
5MUzsR+HlJDQdJNO8YqLPclBCz5rmhJ1tPv/EdgHaHvpJLHCJdO07tbLnIRaPi6wIGKqZZgkgaIf
9bUIN48WjCdUjzRDx2S4xtFFnesmArCXI5wlQoK6OgAXTHdA+jkMmbNLdWJKSvFbkFOWas/3AgHK
hKZ98Ce1fRDWEn4WrCx2NBVUhpNKXdtjqAnttdmQ4aWyfnnnSEeNj600nA41tC7VFEnV11ZMXM5C
sehV9AhIGjAzqfX1el4gCiS9dlUq5WueEbKiY3Te6YPvHCso1Ms5qKStss9FfYIdjnVcTgPYxDOm
DNODGILofXT8bIHht/gDkQRr34Y7oZiVHi3jAw42vTrOmeWP9c5Gf5y2Mk+6ndcPRX8jY0DC+pOM
z1gdSaVTSeVnZT7z9DUKUn6g2+zE6vilFPWR7gV54a6LnCgO01Kxs2CC7BkuqFDzb0Q6cc5jkhNk
f6rtV2n1dIHwcxFDW6Kp86StroT7cIuvNoYrOr7O2L9N/CpDUSsDEbrJc0Hew9YyCfsGVZplnPo5
SyAbGiRsv/AdXiodtfeQyaaCnage0YYoAYg3SnMjfuD3BKz7URW3HBKn9lB8Iy72Vt2xirsx2qkE
1oDJS+bd7+5UH1gqccvzuU71R/H8XVpAhQvdBxWHeFXVDbvr2+C1g83TfUq8fVCaaxbzqjMla/2W
YS33xR+R0THyt4bWtoW6E+7LQgiGV6LsOd2XgQyK9YVylK7KpU+5VYFo/1IwH4RmmRG6D8BAumnZ
0dWovbiOup9EIXqWaenKDfVldtKeltrdqRAntI8B/Qr7DgLPJS7a0/VX2cKyh26GwFkU4afH8W6v
7Sj2dneh2MGVRNRfW9PbDyXotSyNYbxxo980fO2zX2qlYe0qQN03xSFR1mK5emlZ2ahPU3hpjE7f
OVhcpzcd9LUYJ+l1o/RjDrzpOnvtCs5Lsejfe/U53ax8AW6JaLCKeXTuscdUKQ7oO7zazTf58isp
Hw4oNgOu9TVNX30CurTNloyBx0sN9G7tuerMf/+/aRhDxdpXMFvrBodNFZr+SvnOYPsmXqwOYrSU
UyMZSkAzO/KGYD1tr3YsurOv/8/b8sYjV9iU5nMqkF5vwNaU70xZ9gMk4WIp1EC+CZSNIirg3bkh
IOZMfgAg56Y0w1d2gWiAErJKFUknKxS+VkTTlAzAcNzAyXmvBCv0RR6YO8f8S/EoSCX1xpRXGGOy
Ttsn3YUQRKORHvn6is8mBjDjiB86ha+Vr03B6ut19CXdYZBXamFLYIPeOiCvTeItnvdRLb+49Qgf
kebWeZS+vAW4MCFB4XLO9mmcmI18ZCLpgyGI5pUdGu/Lif+9ra58NOX+XZmZ2HOQGV+C5RlSt9M3
ab+hfASByBDbh58hoSc0fsqZtEEn6XpTi1g0cSfREqYkMzpphA2OSQ+y5Ug68DH2eFxS8DIqTDf8
ArQ7PMojuugMqfwmxuAzpRU2x7cNwyWFsBmECXEyVIHjC5IMHUCrVM0pOPVAg84+9CdTXRZBeKes
UviiI+q3gnM+6kvxbUiLNDpYM0JgdW7R3F5xc2VrWBUtLXzHhTzSscJ0qEfYTU9MVnJSLfEcn2eB
KqxSfpCsYKdX4SfR3RWXxzi1jxbK1bPnnJstlb6KZjVCOnuJj3LiPqlxfCueBnFVTsuLX0kyzwR1
ia1mYqAzi9HWHPRhyTf8WzUwHoY/uA5c6dZd1/iXWSm3juiYAQAljzcVXbmQkJJpVrCdBz08KhZH
FTv5oqinYd+iDP4XkV6eFu7Tg1v0EmKmzmdyYZjME7VeFtxr9irtY14SYvawu6OM5psofNIUQ/9N
np6ABfWzCUm8b6pch6QR9PrlXv96wvmhYWVOWsAIBVe+N09+WRLzksE1qz+Zq1UrOzowytp8x+TS
Y1Jc/zGc2mM0rSRdSQfke6fqVESSuClGlxM2YgZLidHOnVTst5a9J4Fz1MLQIt0D8QQ/TANqJL3h
my28/CBfXqu/idMu/rqlxk6Mf6SfSDcm1JEemXjxhR1V2Rb563L3fRWspQpIjgmxoYGEH7zBP/DS
gPb1y1iD5yKO1frvvi8j9sWdr3I1yQCwob3o38R+7exmJncEIqSfJWMun23dCGYqPtXLC2V0s38U
8sBDIGQNzMa9zwQGpY5NGtUfKGdYU1EpZd8eDxWhL43kltbBoLWEVQWZwy3eepNbPkZCFtHwueAg
x7ha3EAOLGQ9kAdUhbO1lSkdmogYFm6ZnhWcAwWADghdHFPkejwVXurEo9LA3Z9jrB9VfVey4GVX
osdtDPFEQ5ZYqhD2Ylsb2HfeKuWepKRen+axknmSkztV8PZVKzT+hf/wz+3o70p1l8d4p30qSEvc
hzBgfPj/jLl1J8omLrCHDeC3Rg+lX1922VXItBZs/Tvah3NpShctT90OEl3+653aSPrfpGqRkjMw
zpxc0m6KytlhzV6OERiZMdT1LhcDKAzDn+TyMVBCXtIQyxMN6bD0nCSryNTHirnfpA5z2D7nLQZI
ysA51mKAYLSFiLgGF22AZl17MwI8TIfdV6aFVIMyftaiJ0n8S4pgIFtsAQR+/X9VGlZZMlFgBkVx
4oS5f6I+jgA/xVkgEOy3kuOaDTJ9YO0MhizVkuCl+zelliOJ2C/qY8z4MHcPrzdqnUmXOUovsaXv
59bZzsm2VMR/z6Pl50bonB8oDQBszmn5pqS802GA4EwvZN5ErSLnN0xPuvFmjkRR5i4XFPMn5DjM
GMXHYf+5gor0pNQuEj/2FhADO3Bm22y/osq269R6W8uxhhO55gTnDQvfS+y1HuHDlA2tG0KiZwde
c8WNRCl+d7/vtcstmtYJSr4Aqu0BSE8cCjMXZdATSo8ZW79c+vsqiNg62VeAoQnX4gHFxRR9lFfL
sFqWqnPg8dpav26TUg/nmFMEl7ndcu77z/OFgk+WKCUv3GEeqkGyiTnmlMo/nmT+asMZJutGKO5t
1UhG4scqwrrMAzGv7/Hw1Frp2DluhniVfmjIDE1KTF0BXkoIHVy8rA59gGB0x4aCHIHhNXlSPLz7
uNDoXkDlb1pPGrECwLrU0+UBulgNca7VVgVzp/jVIH6uvxYehX3O8SpMZ1aqUHgVKDwqNnO06edK
MAQLJwSBU6LAxRdZMwAbeH6Sm8i9HASDTpiX/ju37STaXtE14m72SBP2oHwNYVd8KHQMtuemwaw/
2weUqGB0wZjevQP3CI0tpndi3UN3FBIvkxrYYV1Dn6HKcw1lMvpBI03AY7RFpJleBE+Y/MNy2mWX
BV/ZSdLw1wYZEAlDdTSjFTdMtN7WjtLvdKPfOxYhDf90zvYb3F2SrJ0evtoEjti3bw3SgpftO2xv
fkoRoNY6rDaa/nKms8sb8iuN/cp0YsMT7qX2B49MrZGfg74miQ+MCHx/RL0Xfo2I36spkbyk/CyX
H7/MESOEBG+F0xnpGbjryPJFQA0aICBTk5MHVc0vWeLf8dGSiNIDQqtd8lgQw1EaHXfEl+pyGCV3
iNSP46nM6jDJQHfX4Wk1fBlzH1HkFMVd3xd0dxp/+Syfv5fnmR7wgnPtIuWUC7cxhnCqYWTxG020
/B3gzVkMGm2zxlf4xfuO6IxpQvOr+9e510PAU4sUTaUBqeiO/qqa4HaS3L7bLkQJplVv4cT+D/wu
r7ZyWMNDRICnaoZICCgW8mha7wdPNwFQMQDcvpCgIbdUTQJbz9Bc/5tOHJMaNKUSgS1KraRTDPEc
33SCLeQuQogwAQbIruXDjsGOP8c9aMc9KbPN+AwD4dR8H8iXwu1FnsjhvHfjereGO+MLx1x9/PfA
IRMvBR9jQBOCwtXxTgYuKwSpHcmtGasiNr+foc/Mj+fYEpB1yAp0OkMxuGSPMGtPLcwVegrFwvem
viQ7hyaW1ov2zHuGBd9dW7hH/LPmBd4iozbznkNkbms9vJBbRrbWuT5LwvUUwhaXHPcQNR4agAGy
QJbKGyqQrrboWw6P60LgFFAaN9+tGDvfqhGfbBPN9ZIjLr3dEeZ7F6Aamxxw8jrKUDAUVPjnHE6t
VXuajHE1Plhccfe30bOpSYFK9AtvAuZNDbRUMhHK2XHXCaOXsnKUf0BJVz721CwXVd5EaYHn717f
1eWaQWgb4kCQBwot0Lo1jjX4QXLwVuVC/IUmxQZYA5B9TgM7+oIOqdkGERrevm8II6KzqZt3XCPH
rUae+GbQInXpjndyT/F4Q/ReW8bhCAyDAiuLHCFqFVHB2wAVd+EZT7L6dqkmM7zPGGMSzQKfYd2L
Mk+vQw0MUZKMjK+W0myF9ALqV4du3skQtO3+LGfa1wo6QP2z9B6mhzmIo8CXRZQRo+QNsvmRg6hc
5pFlo7/1BmtuQZGVfoWrhLKjg1RuI4rSvYqKe7Clk+ndnhWg2V1o6dUwJqxlnHx1w5KFWeFAbht9
McfBMzUG1zzdfbrIaMrIfjsiN9VbQ0aNUpbAA9k3Qd0nzCj5GKCM/2Ju1Qun4cgyBNNqXh3j6U/k
t23SQxFZUTOVHXuXfG67cvgs6cxzT/LzlJCLo6aRTmwPZbj8qjbfCwwrePSolCt6+s41TmhmM/Rr
d0axwpSbt1prwAUABQfWfz/2KI6PVyzFJzplb/r5WjruTFJ/8Vdt55QEU3K6sW2WWVjVYPYmdOO+
L27fRq0QDpxCxjJKc+omUx7vU+4jlexMQFqic3if4JqnNQLrYYddESgPfwellWeb6BmMvWYOXXpJ
JE8XcBwtjjMVZwpdy1KEyqO5A/w6r7REb6sWq1pp7ZZ4jKLKcEFTBy9MaAG4+2rY1UpD/oGxetqr
MwlhsFC/T9qGNxJcPwiACSgLwJ169ZYhxEzradzBzbPeZrX/NnZv9HcuFR7NOW821i+P/DABwpys
StZ03dNNEcXfQ+EODKijekJhAMAaDEcLxHmKiIbjSUS+RzMzmoT1sQnYQoOwlKqiXJkdahk4xTzh
2I1EPzJbC86xUcVMwUYKoTjhyRVMk/ipARA/W8/3QToeoKP7S65wD3Usx3PLBq9X6v8Rz3evfZHd
9GxO1mSDx9G0u5jw0tTRb2jFCjb611B1VyM6Tzm+SXuRKsmtHQWm6wc4qiJYR23F5jyP3b4NwY9e
DZOOuwuOsr9VHTy5oahYcCWMH8r0Fjt+EOG61/tRTN5ielUho/InzpMLwkGFCezMN2TvM0TDd+nh
qiK/NLbSxQDSGtW4eQ/YtJQMq31Ope+h809ORxgtOy4vhQlXSsl9S4ExAwNaEPW9vZ9a6hXproZ+
yh9SoCxRfDoztugLT4z1A803fDrk3se7jKFMIWP9gOD4iCYi464AbnlVYMQbQAZk1ewMJK7g0BL6
EPpdYfcQa9tL3Grnn+wnIAZbz+W+K9Y7FIIz+YlMoYHvMlw1myihzAOJQe3jxkONLQ7dH9b407do
KHgQH17Lr3e3Ug/BXwwqqlLQNQXazMX9o9w54PShOgd2jOto+6GpI0Y742PNyc19FIdHeZy5pcQn
XJYmYoJ/hYkelLdHG6xwDGHnwohiGVghVzfrzxqf1PWBNeRFcaacfZSaiE7miNDXI3QJ/7vQeo8y
hKcPw4wuix+Il2brhIJ6jmPoPOKRzJ7+GBnClWX6m8ISp4DbUmqv2f3QltBYv9dAYGrvZd31qHqU
mQ263zhJybCwcf4iDfARE8N/de00BWG9edJQv58PcqXlQOWPK0QYAG4z8pJm70aeQLeOW1+U36Af
irUuFKyEE/kfncSQZNoslp5WjMW+KdDVl1684h3adZlU9sYVvWkZcmBtKZuNqm5bHuJC1lGVgLyI
1CdmMey5d5J33bPTrMyY4cLrhtbHHqVeXQk40ljmPgVLb3N/kfxTfeSfjNCK+BViD5wqIllVT0XV
6u942cTOaMbJH4Umt9zCgrYex1La7oBLisO1Wy5HMPz0l+lFUurrcATGNC2I8JrNmqHH4UwhU3yE
wbv8JLV4PbXiRPXr79fs+qrWlfHElZotJyPpDJGBCUntW7eNWwBQaUH6x0SQlL73WRqAigB99gCX
hv/eluO9MrxF8mvGl3i6gUV1rpOZBqD1YMI0nRW9eQtJz8ag/N7hniqLR+cXnw5BJAJ9o9GnMupK
O9FblTo/8LQhiOMALUKkGZtevmP/hNCissHXOObO6AhnZAT3kiu8VNtS4DcE1+fvZXzx1mMoxBXb
eRzG1i6Mgm87Inn9iHYeoqdfusCBjCTTIibLhBfrkLNnpA3d7MxtRUV4RE+SSIbvHfBEifp/nZSM
qRhKKJ5WuU1lmkHvV/XZ/b4vS4KI8pqv/KkyeUITsoQC0rrDiid8UfiRvj46HL2+qwELSoQhtNTS
CiW1pXsSdmtPGqP8wznORnsw6UnMKYd3ud4aXibrpLQ8/GVibVptL0YtfmR7QnsN5wYKlBQs0RjE
SzuTOWnTijcg+khudptyp4KBn7lwntoKTzuvCtX+7uzEXqhi3dOBGga+C2AX9HYCU4Oc8T0L3R7z
2+dV8r3fqBw4o2JwsV6G363a3rZMr9JuKmHzil72EkhXTfu25d/T0Sj4jbg/G2GnPAVQXV7nJvr5
piRK4CyGjLYptlBGOpTnUQ6k2X12CE6jtbs+ZvwpjNgtIuclk2EZjMiHS6Se
`protect end_protected
