`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W9ikAzfkNAB9r6UjwYkkLbO7xSa6Pa5uk+WdU1HnuyZEhmVth9jtplxOjM44FNqSQvXccO8yxQi/
NOIWOqyRuQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hEuem1/oUd4/OEXkW2OvYqIxpyUbHGfY7GOC6MYHG11DUK95IJjyjs7VGLCJVTSk7aMQu8m0Up8B
V7A2i5Ur1C/MGpffEfJZxWT9TmFVFogk48CVrfRqfUf+EY/RnTok8AxbPM/CybW1sngqZ0CjEdAR
WFwF2WmA9kANp7DyS9Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YvMHbfeLoNrrdjK8MzZ3wyAsEds/aUUU1qihbPDmGwW2kx85UhHj3XK9rxLVtguq6gNEFC6HhSRq
ElvLoh05rPkMnw6WFsbKYG4H4bGxyS47kd8q3QuXnE6sCz6iwiKIv3dpxTb7XlMwEgrVo5qwxGVL
s9GGRvYTehzL7krjc0uS4aFXrE0IozDVS75JoLN8e6buKPj0LqKxI7eJDZG7nEfNSuwPJgV9jjsn
hBN7sE/TpmRuBxik41OE9HAXgcn8nnK+V1lhlH0VRFNNoFpqAT/MO7xuOSQjqp+eRafuukS3cAC0
2Sj1JyG5X2zzvgGRtR4WAzC70VggYtvYSDr4fA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
odYDbVugJa4zsNoidrU3zfx00EVw1f1F4ZM7PMiUD5vBKIyGujE3/2kpootoEODrHYYL5BLfkUxF
BOQX5PSqpPgaDdiSWs2KCidYq7PHZN3L6Rfg3lupSDrgIHrKR+n/0uxrr/QGDaV+/KOkCbB4EmF3
NyOLBbCEbB/cyic67Z4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eIzvt2wVqO3FcBIgfe/d1GrO8xAJyZ1wgW6um6UoZcItt2tjAa8e4PowdMaz78drHioWBIt7t7sB
imWtFcP0XMZDfFZ2wKw3JJinSToIdJDnmZ+SigbxdzjvPvdZmXqc/soqccpjzaBwx0DzDM+jpCRD
sdcRaQP44+rEYmGdQzUtkX5LMZ/ySPHZt7L2ejRcX1NR7tjsbb6iftGBFtOOKIolJXES4o+D0lFM
w4plD0zfXEeIpYzOx/B+7FZQ8lYPkEeG3Q4nhVL4OPIVDrnnmCTdbedEddsMjHf/oddTYPxyD/Ra
iW41N9W4EeySOPEdcOEovPgHrZ+ZDykNGAE4tg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11024)
`protect data_block
wCi1EGWEcepbgW5uOEPN0evgYS9XZMSzJsF/EcLsBFhCvSD1oOzqmP8fJeDLmEdNQF/7YfTTGwOG
s/wOi78uIdGAW8EknbP1v8GZ5t6AckJ+EAbHX2Fw5Pv9eiMTrctGH8sk1YlZDCuPnfV55Q2O0zud
+0ZgXnZlrc7F/yyZf/0sL5RdhKarwiOYPkVaXJQy9vCiCznzitdbynS2yKkF1aLC3vIZhryEd2L6
6bsXkgm7ee4SOk169T8++p+1X37L+DO43l3b6H/OI1+62kC4OMfxcvL1jRl+vSBIkdl3HUEXQrCw
BmWHZcuGnpe/iwZc1V6oVxIxWi4cGY3ejnO6+VJ5a4rzjl4OlufiZr9qpgclLk1fxBa6TbGihHi9
RDMs4KeyGEvpcjzh6tGhCG/gvV3VK3M7wp9uT7YEPNHxQO3EM7PlrsX/DYSZ9PzM4RJjzCocSe/3
XiNKaR345NJXRC+Wex8XcPYAGljr9J9w5GUwlC2iu4yMn3fsLiDyiN15qNEGr0Tl4Xth4CG1sfYc
glnF3CpxdEWH4FnY86Et46HYGX+ezVvSVjzWPfQII4x4TuqPCdxM4hq53UY9L8QnDPjkJidKkAYJ
A9SVIQVaSdUJb/fJsTc5rdQBFybAaNUc3RWW//Q/aegz6j9UZTB4EY+Fq0UzFmtB/D263K+5m5R2
k1jVDCHI37Mw5Q3mIzezR7HEVX5NJGQP30WUpwf5n0QmslBWheGmAaBdXi1VQAj2oDgSvzK4Roj1
oqpd3mMkX30De+pToc2HoY/rZUV73JMlIMw0KCIskkPCTA7ip+VF1+MO5EsiF0xIZ8p/FkZhkGPo
Gi5RbLu1rEg2F05pIat444Nyyr3Pej93fE8aJc67F+/NYr9AVk21O3C5g7oFX+l2Nce1AuajhKwK
0zB93kklzSo7mCDRBC8q7PEMADV7fFxZucBy3aK8WU++rS6aGKvHQYo+2p75y3i4EMMBkH1Rcqoz
CBDgAyuUqGwrEfY65q2fL/2jRGPjSuml/rXDYuZlu0e8j0ReNOjghdJSehSVOXHCyHM/xw1qBYIo
uu0QnGqCpTsM4q4RdHu9HlYeb7yCMqSkjYeM1+X3xYu8J8+p5KKY2mUE4eWgHtP8CE1KaM/Tb0Ow
M2P2+liiXliBjWMtM85usfHCJ7fmmm1r3P8jk9iuggYxmEjXFC63ULsDz6owyUT1VfVXpAIp9/ZJ
u7uajzC8LEbqWkwqWgryamL21YBZNwlyNfVdbSiclHupKmo3pNGFhYwOmYlqS352zcow2F7u9+xi
hUqZH7C4inw9SAFF63DmJqxhVE1mQjcWzRkw85tY1KWM6B7udsNpoKEM1WTqI7qQ+53iDoEu5xYX
4TWSLv2MSWK+djqLm37+GWvOwVSDkIkJhLGlxOienriYDND0QfWDwNcyTjeD15JdJMZTVEYtmU8y
IQISw1STkXPechQz3a1Rh5jWVUyLi0HTzdHo52FenD9MVRpYD0qxoBH+H2Sj536fFfKbTI2ikQPG
z8jiimt1UA4pRXwRZ2SdUFdLHp++REwX+6F3gnZbDjjJfhP1j1akVyqDtJiJOsDEaC1xx6PwaQWV
1lFxpoiRpTgQGBwDj4H6zqpUJELMM9xoQdNcVawIlV8H4xSQNp0KFquOdMjw7gk43HAvEoV52Ucx
T8G0SOKKXyQmn+d6RoF4TZiPzLsGLI9JQ3fDOnU+ONTmPwIa97TF2/1jt5rEC3BoZlZl5J3iLjym
+HwPiDdyxWmDVN8eh8YTbIUbx23sWRkXdO2OxFnLn7wNQKPAtPw2rVHbDty/enJJ05RyJrrLrsDT
cucwoxxeBYKjwEAfjRZqkCDGUioTv3uC9+7XJvxjI1GNCyFTtLwCCL5ERtiC25hSec/rtw4U1PyC
LFRTHU5FERCf0Uha12OzrTndcISwL0Q9nb5McAttt44W9asyyeSQXJmtjxx8vZhBBv3KDFEJVZYd
NLNr3+KqXxd5e5EsUXiXu6JDrjgmjVcg4CY0fyKZ6AzWLIO23g+fLrmTjEjkaqg93g2rcxdibiC2
waVnqlSwtmaBJdGxdDlVJpgmHKE62H9wO9fM9/uDkEfQQtfIlXIA+9k8PDVKueAwexRIhgb3mIFN
uptop6MXrrb4kSu4iuxMzbCT6fl+/NgFz1AXVItp8SH1h/Trer8XpdiXcvO778r+66DugCLXYS/s
OIRR25AD48R1w2GP0649sZpXLfBz7F0HqCLmdgVn8gMNQ5eKsWdXOnpcQIiP6hX/l1FOLdMdceNP
gaatnO4SVC+162i9QswQXO7OlN+epuzGKmPSiTLYygv85pACrYF/KnSZm/x2tlWh+wVZkReOksgQ
2N+D0z0RXeDWwtyHcsOM61s5kuGRbNgEf8K1bhCo2G9Gfv31XQMTLNupQOTuFm3oVLClNt5WhDm/
mrV8YpxXM9JhQP8wV2zVAO45sV6/pqZGkqOOB4nSI4nsbD2ISQn2325dzZ25uZMmUGVvlbQ19cAz
LLV+EzYlV9c8Br9KeG8BGUrxR8dFCunXrnTGyVRQeszGYBJaBtJm69UpBBxF3Jh5mGvmr0n0sJFo
F7Mgz5IglCO4mIUfOPRMsWmb8JPB6yUX9MaCvjILyawpazflhCDi8aAjE07GCW7VaERKnY1hAVIA
Re6UzqWdTIOWz8miNNWoJWor/+ScvfzOwPaGhPVALiP4pZVERb7JIDgUDeR/6EBJ6grJjM8Bu3Ll
9m7bsjxFoSJfwkkrkjkgjKlOL3fl1/FLFoL+aPfk9H87k9cQ6Bv9RFUGNLF/taOw+n8UT90Zlh3a
/HmP4OyxGohsCGcc9FDhLDhdwKVIg4otoyF8/ZE0B6O8DE4K+o+CKG6MC8GPyEbnCgcQ8P21P/b1
wvydvR1ISUCwoSZmkgDtXFfnaL3UPnWHm/xsOWX+/MJLNsoXslawTgVjT25e8J8Yyflj5vyKiHNI
5lpNEPTvrBzidpYSoQ9+v62kKOyKwT9V00ne8rXZxXK5/Ei9h0wc0DJAzRVX5C9/CL53uulh/Xvu
Q8yU76t3lpZGujaqWf3XCHi+TEqjxkrVubny3pUuBw9GoclaqlYCeV8OAdkce7C535FnNXlfZfn6
vqF1Kbti+iAFI2TGU8NDv1O1+2ns05P9++TRXeyKJUYBVnhUswAg5xZ6nkar8fcORx98ziNa6fwZ
1uuPktpyjrXFSq64UbVTERIA6TwHImc3el1+hKsFQRS+nWfZDvKLqngq31yEjkFttrJBfI+hCaDl
JnQNOpuFklfg4bYw5L3P46b97uKq9uNmAHy0ezNU9BSoVI4xvVG8thF+tC/UnN353/LZ/u/2nr7T
VFX4x9doWaEtMnpADsz6lxQZNSKjh2DEIA4GztQ9ix6GamPsINzITUnvzGBzpScLm5VseBy2PMQi
SSDhcsdX2aymtT8K0SOkIIT0ImnjqK6nuq4qx89cCQqIIXMlmESMbhcJjA+iinWl9iy1f8uF2Z7l
dVk3fVcJtcPlnVjOCYj2Rc9cspPF9v+Nt7csYxadnwcAkr2LHGzme4309qjdh4Af847tlVAbuid8
CYV4eMBbTaBkI6WpVeU0vBd53e4j2L4e/i2AwhY/o9BdtONqeLM8QjbYOGN8H+Hhuj3Qm+8Qs9EX
emAmIvxoh8nFtlOxwCOVtRNuj7sMWjAZdt3x6+MLm6NOas7DYqopXWOrpT2oOtZvHQ5p/GuEgDSe
6Uw6Jju9Zq3Q7WrP+++YfW/Rg4F+M2f8EPRLBPXQ3ofmID2MNsBOrOTPT9lP0P6/LO0/lVfnTRnf
UODpU4GJtAqQ0Zb5Ckwa/7idPRN716prGurD8uY8lxZuoKcXPZ4sRnt21SGZvXSZAneSnLHkrFfP
Q2XwfJI/ilsUgxf7cwQF3IJq/xpvVUzYguPYt9UHGukSNgxiECvXWdWxVJS/UHX0s+RPz8Cxrrxm
6GUQQZ2VHelxubUgbVemoZVBSr/50f+GDFmYocgabwl3XFQna4WZVtmx0j2Djr0ZMvlghtlFCDbH
26xgqSUWD0lF4rs2yDcfpJMuK7p6NBC8yTqo7PJ+wi4JaypSPQrUv8AsuqYO2mS2BD5wN3gM55MR
uJGpM5PoRnNDYCe5okDEzh+vfVBtd1vmewSCfzqbtKrQvw0AN/2b3iSF2wKsd6elS/JBbvDJeXR0
vcaLurJt73FtjHzMvDVWwBjs2XZVAkRy2g/6ax3EJel+aSsxrCLdVwUg//cF+dNP8O57BZ4taE7y
LClTQL0stTDosvi8b4DMpWvMEU/y+/EAf7Gooh55Bth3hcWzU+Z++HciBWGJVnZA3w041qkK7F7k
nrcpXABgxCSW05l0Am2jQOHdm9gqrsG0jOHBSWvpIeQZ/6cgotjsCH2T6a0cAFG+D0FyJ1h3pY/w
QEc4gvHNhj1vUxt4LHVcEXZ7d9PUdjLY80iZNaT6XAq2OvwGoBkGZ0EIA+jaTFbMwc5M++i5MHxw
AtbcGVZ/DvSV2A6ZfjMB0BJ910HgMsHkFPk8gpx09xssqKyoickNmqbOTRzKkApmOtpCKkV4XYxL
OjvRP7hQIcHhmu9808MLz4C7gYfHiMl79EhttiWyB3PrPvxavHXmfa1dnEJLVOIGncRBk50GIIGg
HrO+kb3YjNpx46IT2NY+/VCTXNJ3mBRkkUGyUMD/LxnONccqZ/D0+eVoVT4wL+cmeCsUTMt3HbLI
yLAGCdPejK16Jw9Q1FR4JhYK8pgHUvJyHi8zEkKe1g2ajfMWGBgTLk1I6uuSvnXJLLxbddK2gJfK
JDMgtlc8E+h4laKrZA2jBiTH2mweBeZNzsaBtO95Vg8jqXNI4BgwovJzk4O3Zcg0UYiuyq9E+iCM
8MVkTxPuWYPh8tuVMSY3TrwQmGJt50A7CjAKalLx44K8UN3L4zZtpzNJRuOuKU5dg1ssAUaCiVjj
zhtIhRJh8MphYXXxi35HSuWRlQ12KRrpsXefBadtqgrfoNpmBtFxwZR8vrBc1uaS9NwPWnbBk63M
daE2DGX07+agz5imV+o3DM60yc2/40St3Fp0EuGGYBF/RiHJyhRfENOrQf1Zlk5xNCqyhR+RmXOF
EDdWJYA5+eLQICqMCN/ZK+ImITU4xnsdpr2lLhCS1q9I4ivLjGy6VY/8CoVwpScON+33WdsOHqU+
HiQl4sAd2n05aFi/kCKfnGBY9Dwo7+MuVH3/A3SwyPcIYHMEdAngKYbdq7+OETPEAvPnukxPeQo8
WvjZsG+kvu1ngllQBwYYjnEAF5HhiZP0MnadKUS6o0C2t13rOEPB0qaBsYB9ELEcy+KRWX0Y4k0Y
CKch2/HMoaSNrgolSVp9Uj78ko+cpf2hO/7Ap4CedHfgv/qo9TNjNBbBicnW6pqgvMZgLmEjzBGg
J7WOrMNNDvIrA8gBP3FHAbAXOr8Gs699EQPkQCi4+1P+j3tvsZ7z3gBCyUPHXvkD+StxtnA3BZq5
dlA0EKVU5E3QNPqHTqDFiJgnrGKz1uvgOp/MLkPwbAnfv+k+Cb3P+4Blg0qHdKaLX1okmpODaSa8
JvKQoLJbgl8gGklvGrlORf+OAdO6wEs0mA681HnRhFvkzHCB8CtpZnMkj+XtBexkeEUYZHvOh3pL
yOfBF1a6qizc/RNu2+FannoWoR96t1fPF8eklFf+cedAWEfaPK3nWGej8ukaMXjIKbg9fVT6KyDf
wLQrQL4LdRFWB6Y/9kBiMxDuWdP0gE397ePL+HOLP6bsGjqN9zWsntcqkBRmqO2CMVVGS3Y8148S
gU4iPECb6FwXbwc3yjcu4DxPuJ6YETrlybH/nb+kZsFNms0XKO6ND2xTUixnwzyr1N3vv6F0CWe1
1UacUML6Dk2ndWa+E3zqOBVwFSpRIHGZwb9syoT9PMvJXmNM11cc6WEzzhZpbQJB8SW4rNqe4f0L
n1fRwmvHyQefdv1eZKvQr0EL2i4CEGAdh+8pKR5QgI04d57PCoJQJjvXiR2JfYNd89BWMtGK6zd2
+UWaNp9uXCurzNVgXb7Q5XctS1Bl7fqnhGkifP9GBi0sOaLzlYrOWUreezuC/Wm/i80zm3HIxrbh
CphcYYEUwf+scO/1cCTYZWeOt64nPlNZC/I+ONWyG1/iUfpT4pLH6NLZysqRDlZRDML3VUQNUxDr
XOujCaTRinuglfapVDRf7ZVegPTnWssuG+QXNuur50QuDW3K6WkBWx7bDiKH2h9rvNc7ktkERk38
heGQygaO0qeo+uB4twoVBNfyNKfO2Nd5pwVIaLKHxTmNNb3NvaJZ3dctvoC4viNP4WaaK4Q2cmTD
aym+cyLi3OUq7Pd3kQQPWaxZXbAIojzcBRS0HAryuzXScnsbL9493fqEe7di3jS+qWizMjlx9aGD
3+8RQEb50X34FqOjMHFadbS0Smz9vqgi88BXX1tA1m0cBYYdZ97ZIBEj06txiK+MTHDQdxhxNWAg
3orony6RMm+lKifnHDZZWReSVW4x4aHjASJMMCSVAmk6sjjmrzAdL/QO7Bx9+UgElmvLlpmMZPpD
m0X1c7KJJ7VqDsT5QmKXCnwd5X8BDxE2155esUsxOsx8q+rDw0MzXZwCf1U2Jb6Dw8xEbwOZ40jz
ttetB2fjsJIbDrJZe4ZwWhtTPwIFI5A4w21PmugJtsBDNw6M73CEoy4+PgYYxT+VLBuzc0VSG+gN
qYJ4lwrkBzxFmgU5kYhvkkLV5o7UXPHq+Dn2BwVK6J3Kbd2pGu8Dzhc4Cpit5kDLuwWfA3gt4TGD
rykl0ClqIG0HYJZynx8FUtv5DfHrwLhaJZ33418ifEQqrJuGR27CkXR5v3zsElLqcpM6y5jglrxN
JP4k1npi+7jM6E0i8wEU71eOm95QD6BUd4aZij7R7vjD/02R9l/7L3j/HHpgjPFi78CfpwLhfuyB
H5OPlCC1tPAbtWVsNtcXN8Ab0HWNuPsPIiDtLwvIe5F0SzXnX1tjbXzJuKUOZwPqTeCJJWOELJdk
wdvUfjCTcB1FcGoLeUfdmuIFE+RKyS7zbt2FqcRIUzgzRzB2bDZ/uL8A1diLwS/IRfEo07STqm5v
NFdVn/tcWfWws8udUK+rDuF8r60p+oeUEoj7LsrOpT0dIkIISxjGpuPjh4Pr4RfDnFyIsGK6o1YG
GGI7bo0D486P0n1B+zNqE/Y0t54PzRLzgNeDYmLPRSoXWQsVMNkuHQRQrlCEYY5y/FwoHy4yc+/o
T/mBxinOwAM+S8jDUnG18R9HmgohJk5o+s8+L5v3GxxKkSkpXFZAmUrVEOfoqnKMwxsiwsiyDE4z
ogdndONAvMG7y2pWm/kdTpLY+tYkdoatms8zlAZMPX2N8wWD/GhYzIwd27BaEdmeeFDhzY7bB/I5
LTo5U9yM3sYxUOCqSuUf/VG7yiNIvmRVehgNk/s1G1ewwZCEr8gi9gOLTePLF9aQUhNMJS+VU6AW
qrh6xlsbGVUYk2oHtGWBlw40/Wqe1okdkZUKvlMxUUMxkHBMCphMyuCjhF3uwRkdH3nD0cKJI6cd
MzAADauO/m9767UuQvlgltNUk9HJbpvnt/67xQA5vu67/GTyZGu60uToCuEMImMsBzZaiUo1NGIS
vdpfVnGfM0nAe0EM+kGVQSdP1QLgkqCW/5UYzPtibyMA+A0KAr3T8dEHBnkO1JMntrE8arM8VP6P
M9klHAIXIb4Pnzt5IunE5leV7dy6WPepP+F9uyv4O2oPDA1PTL6BWj61uKlUg0xPO8KCtWEW2lAT
IRLjFdJJvXslKd84Tne5jvwRQAQMg2WocmHiwk7TYyWihN0odqKNtmSdqYcauD2QDzTT3ihBnBjJ
6ltHjrCfFwe5NeWOnqUMypMPtZXxjH17d1nIPpdm+zqa79/nSB95FS4FG9vAprWvmwr5X8RcJojD
5vkOmoQtpYaKgWYJz28RekldLSfNPb4H8mYjUxOmizCSgbfo45l+6b/hTwFCCgPG1W89qgOhlrYf
HECCi9tEPk5XYM/WHVBty3A8vxcms7TF4e5f5u0rxRnM8JnwYuosVCmJpfjo7myfsexQkF/BhyLx
ewQbT1k0UWHWV3B6a7yO8G+DLz+kOt71BICmvR3AeQFVwyaX4ldNbsaJeUZu4jOkyx7IpDFpSLa7
z90EvaHOShqu4nlPI95Ke8kgKOaQ3GukwILrFwz4w+0NvWcGNFH37ozx3QxCsQlKpdgt+Ib0iBBg
h7iL7B5oYOeHm1Lc0fKIspVm0GvHXamYCK1xaqQKpuC1qd/sHrc33ACYzcDxNDeaVS89wgDfh2vc
3R3sO4PsurtD8zXuIUcptEfgUpJnUTRWgKmD0P7H8pg5PPHlvoq0B0xXOZj2lhAvr0pSwputKXLb
Wv4M8F/+aWXf7HL7bonuqT2EHCOe+qWEOdGOr6e7YYOkUULd+c54YnAtaPBkI5pWIWSzy5U3b9nJ
/p8+zVgoXXBkUo36PMqQjoppaKHP8xGwMY9IjndFt4XtXwpbAHxExUQCyLRRcvPDJnswjxNGD8Cx
c3kJa74PjFdAzbejqNdOFviT/EFkwyO1pLxLs5BoK6dRgiqQbc1ZphImlMG5wiB3DU1d2QQSTMn3
fVkF2YXM4/i9WO7bFT+jDzCPPD2INmiF2wjzr2d1cOGoKU/ROPAxk6ZFyhCJ74czt/CIdy9oUWPm
ZIALnrzH/+RdOMKIk7NO1XHj2xU855YLuPUBu7GJgfdCNsSdKuCQgWaeUINi2YLbiXtRKZqSkKB9
o7h463WBwWTKeX2hiYlr0c1BnMW6kgqSbEFx75kLUaTUMm2+UI/+lw+1x2BHBP9TB+jvx112YtyW
udDOW7g/7aAlDYIyYZQAqYZUWI2n5SKHrZH+aMUz6oz0jy7yTczjEHocXFu9s1uzEu9/awHX4161
qlL97LWPVkGWhLx2cTevjlDrpoukUEBE+RHXXfm+XP9jkd0QA3+1rUoGGoabbWpmhkUl1yeDWm/2
iUa4y9s931hkHMfw7/DeqyX+H0WjGthxkHOvBLEIuv1bd02/1vXlZcKAtgK+yApXUvn/XqqWEZI1
jGzM9Rugp+rMb4Vca042m2SrTg+k0ip+8NbQGbHFK98uEjPBb2NqWw30qxEIvxYlcirlImi8osGq
QKigQVTuoiJz1z4MS9C6nZmj+6bWZUuzZm8b44kJMuyF3YFgXjWRE2VjYUGSWDb4Zlr6830oflJb
FvmFbe3ZPaJiXqTQETeXuI6fSSkDZpTw+XJbdMLOD62UHG06clgTHF9NZwR4yyHPB0jWQ5TLPDjf
I57V8jTs0lYVDnHL34BguNJJXtkU1a48C5BbuOlwheBO6Ir5E1Jo7HEaShY0wA77rMAgWqg9MV1k
doND6yGLaoudGXQll9HmIROFWe4NG//FKhdqGOqv20sm5/Gts9vhjdulxNfOw9mepUUamVYl7olU
XpwPjoWjBx7zYiOTrirUqH96iTccpCIb7ickww6IbM6QQjOgbX3Rz5sTqTa9xAVx/IPxBAS7FXOq
GuSPD4sXIjXpZIQ98cQLdQnnrGGl/lltEa5B6B1wjrf4JHb+07V+K0kX4qf1rzMaxcY3QIuc+V7B
XV4GrgBD/97DWOFOV22elPnURolVFxUr7AV1QVdcAwklf9h9Br4gHxQ9Wf0u05AfKT6EQMpkJwwa
P47sjB5PWc4/NWzuMxyFv5X3mGnugwrpGt7nbD59Nbv0r2P2FENy8zjXXZ80KMK87YKyn3LXPmb2
q6dOWAgaWrEZrFR50Qev5aS5Pnf36DgKNvU5E+J0/BwjjShVU8XwgAI9G4Ur3/GRez0Pe8izzQG6
xQV5+nn5WgdnvnxJvKyYvUfcqtqXLv/OZ+EK0dmadT0eKPoCPyQUzywwlI7FNjn319Di4YIcdxXq
K7q2IdPuXb76sT2MjAEJArApz1hGIYIYkVwPxAFrwzMCDbyl8EIuG3oIeUqyDjPZTK6+kLxt47ba
8G2R0/udH+CHwRW8JZ7ap15J0LCVLVa/n+gamRuaNCO86/BAObtCNuixubfs8vQImjkefo1SMY5Q
B6fB0iVbcdbxEc0bQ72a9RKFnMJzkICcdiNv4Qpty8ShgBcTGEkvuMLDARtmOjBRIoMuKwcPYmLn
JvsfGm5Re5EAAJYFC3FviXp+6ps4bdWu2t2NyvWXZ1ajaV4uwXLe9lgSgyTY+MKDY3US3b6+8HM0
BVkvIpSkeaDwua4C9nlm7JoOIEoDL2Ll3V+ABi0ki3BPa3Ye+s0iXZVbMgLPhBrDgQwdTeNWY2iZ
9kydxvCQpPagovce5+KpCINv1RaYyWqzep7grGyfVccfitrc3vC6NPpJnPuLwfudK/4+OM6/J+PG
rXkhzDxVq9/NmqvRCR3Bh8Tv3BmxiZmLJKlvADm86eI7sYs0QF0Cq+PG7SI221Z8aWx08vo0RYLJ
5Shm1keaQFbDw+1jS+1Bvamj+L4K407vmquZwMfK2dM0zQrkgCWq4Yfed0lurnkb7mej17T46+vO
uSI9luoSWTWZCYymqz+hKcEzOrIQS5yvn9HrXXbveQhUxyROqHtxRpJqnbl0wZ3DJgVYmbXCSS7W
k7lDnduuW4kyvzKoL+6/UNTRED/rVGJnqwBB+NMCg1wJTdZ2Xi3GIVucxZRx2hzWZXkQ1YF6TxA9
lymDZjAh9psFClQxxpWOmfL0F7e5viWzjSKFim+aRUwdaPWHIdYSbBSkv4faJEbmC2QToilLjNkM
+icgBYlr34gshG/BhzLW00QTvhA+UdvLMRC24SPGPVsokbrMVSWSAM60gjljTdBUFbJDm50wkm6s
HMg6t4IHvdsXH8TvyInwyZ8JN2aVyOwab5jx7Byf0mjgQx6ZzKlo4XDCffHTWiSfOhYc58C7e6JK
QHxD/QAJGit0pCrdy6LA00ZynR6tfTiUpd2x0OcXYIg82ChjvQ2TbtxSFx8EAd+/yPwnn83fJd5W
fvZp8MWz098AMUWTUPo4helY+FA9tYpczfEgTIqCs4ptE+WE4gA/rneEEPwqkoOgWzgMYO43F6lf
f4TD4M0AK5uWR/lxD89GTjQYnHILNoG9ci4E1kQsxVtXyGZlIr12gSpdDKWXexuJ42YPaqddbyNi
ymODEWI6bxyQCAAsF83994oadmIyxeAg2RjqXpN37mhroY6FHN8SkLIS9FOTZl8VTSgv1fp9vjiA
Jx/h0b303s7xNZ7hHMwwOgMwGYxYTHJzxnbAMf8GTXtcirnBEHvH+HGawnsC6quCcVpapJBSwH3Q
1SSFJThAkI5R+eLRK0nstV/nzKLcAqFlH3XujpVZ8+jNTBqlK4GxBRFLt4Aw7S4V7F+6ujg+dZ53
SCMMt2KA1AMK0CRiv/G3phXD0atibwKb0wSjaHVnfGa3idHdIxGI1Fog981FdLEcTBer1rs4zymB
Z14gb7YkIFI8aYUBz7CtECXwOcBw+jABdqGmQuMPoNJnGkXV431I14MZRJpuqfcD0b5jbHkp14DN
wzbom/0YYjAJPzAwXr/58oQWpPCczxq8ZC09sztQw00hmgMErYIEysWFjpNTqCMRLjuY9tmrceWM
PJa/qWDr6yCSOduTZ/gEenngtXm2orzroHdOPGKKzHz490U36HVEKNr3Pt/XQU6AUVvQ3GLs88y5
cTDrZ4SgmiNf0UfEQDYFzwG3wHL4p8Tnl2nmuxrAVRQ0nNSst+3ydz19l/QN7x/fZmoC4YLyB6J4
ndKKDCgwb94G1LR6PCLZYh9olBov2fv3h8H2rtQMBZdBVLPMj6E2a2KHr9NahH/amAQNL/ZBgUqI
z7K2myNcHxZ8ABBf9yKc0c/Shb+xrhI+ysMFLE/3qOKFc9qrMOylDYZcvaq5z07Fgl+9WpHpNnGB
D49l2Un42iL4EeofMpBuYYEZ7/++bYP6o96ldaxcehGkbb1F+NtMXwVQW/XgYVqFY9J2SF5BujnE
g6SuA26MsVpksJuD7vbxOzPtjPicuw1Fm+DD6IL+Bq90tgfrTAZMQW1IxCqcGKH4nSyqVHhKpTjs
Ron4T9adljJYR7DsFNH6bjXm3ePk/snq7/D4WcWVkmY6Zsb88h5jZOV4Mp/QRnx2zaO0BoXebgAs
HBCw/RqcD65HY8+/uGOqtudNS/tYd6hr/8llyel3dTB/xv5T3PXKIP2IuPLs33xKkJHRN7F4aJs4
Qt/dWv3iRG9cqvX8NyZMArBxAnDbD2ywVTGk6ZwRbzb4riv5frsaSnuO2Cbajiw7677Bxup0pd5V
5Io5QoTAkmIOd5uJ5FbziKKo+bghTpBE+4RXrq46GIC7iEVtAqEaursEsfNIWu0XecFEyHurmnwA
T2z3iSMqF2WT00US5fdoE7oBAfCaCEJZqF3M2ywIvWHf3Bw1Ce3H8CZVdIKERaP/zWu+VN8a+D5A
S/MfehnY3jfnvS+G2WA2jSHVyeWwjTxo7nCfQWPIbJDucHdJySiyiYQh1+15NhEwi5mRVR+bJ6Y4
eX2ndPdswspVL5y0+H0RsXZkoXmLodbG1mI7b/BL3DdEWg45Kp68QF3yuGw6iwvd1Q2fWce8/+IJ
p7473UwrOkEvRWzP6aVC76E/hpJobCuXIASIlPfJIOoIt4R6WwCXNB4ZIIN3N5a5go5YfAANWYky
tU5jxCxLyR/J0nF1eG47Krp0cTZ8Xnazpr3n/wbq1Y8hNUuGcdsel1RWleITOy0OWtQVctghqftx
0PFzNp/Vidh+/YHwUYA49cPon79VEjLEfQLS7lTt/jBDESAWnwEaLaK2TzQlknPHK/NiGqQRAVrU
v13x33eL4ep0ZLtfQPNipieZ8qNnn3xmBt/+t1i4eVPhqKwTkw9rrU5pI1Q5Gsrz4ruaUvZq8A+f
QpLBhoMnB3blMpzxQeqakg8X4WV5XQXT+KjqPEvyIovYcBNg1f970NRiJo7+AB/uMUpi0o0qlSOU
Gz4cjwe4WEQ1YVgKDFpZlJimkuroij6Tm+avlzoxDqD3m/gpEhGbfyEddFfDBM5iCJ/3fF2i9BHw
PX1ZIibfjGwFDbv62/FZjHBJuyQdEObKiWzY83GOOWy0chAqSfLf0NG0dmaHmKU08Fxf+TetX4O4
/AfLBiALQVWsyDm5ME01cmG/F0wGoIMJh3v8p2FyFLcxbuR/2wKD1Ki0fpHV54xw9yXhwDc1pwve
T7mmWQ2uoqmVnCtn0WKsMu2dT2D4ShX4wzxEyg5y1mUQ/jbhUQ8tqpTp0YLW4RBu3pmSG82IpK4E
lBrX2yZMFLy+5P1DC/hFvzS4qVLgXxVrqebDA/D3/oLt5nZ/Y4+Y0OtS8TlhFeVHlJyPSpAfbR7u
wpPu/uMxl4BhF9CxwSlRsz1Zj3R7CfUvrbKqbnvIx6jRf/VUgEj0jHTKl5c7nZAWCmsQNoqU18V0
lE0hmaqSchE6dfhFV3OEDisMmT2UD3byoy76CavG5LbMjQyfpqFA/zcvCH4jogR3UybCKtXGd3zu
JWjOAyCZ2EsISs9uVxqi6H9W4iZhnJS94o4+FkwUt9wtP5H4McFninSONxAz/P+H9EKIqt54ddce
W3NxZ2g741cfWMXrTxT96NHVzuPqaCx8o0k5ACUiJEktWcaY3zgySVJYl78EC7UYbUAc6ugBCVdy
k1+bImun3EC0iSvy7QJMo2iR0fJTdSNwWoCIlPXyChMZjazGrGdNYs+RBRoScNr1si7zsNNiyowh
pTjVDUCHnaR+D0EpynL4gGGQVKovn8zRm5JcVMpJl+9/dNph0Cxr1ESdMpmk2FKrZKRdVYGj6fQ2
nG52LBZWAG2owBc16RlTG4naILE5Tbo6omsQ6u6xuT8nEqlvJctkzNiwbWOAiayZIMKWTFHr123Q
hzzevdPgq+PLETWVpuqWVwABs2Zry5Cn8/1bY1ycLn979JIAWPZ+CWFYFNlN25pN+EsX/RHG6R5S
KJiTZkoSVqcMgA0DpqLox75PBFPyJ7i1cvjK8YtTujok8e4VVhXsI/lNXWMTC/UbijxZwtH267Ce
I4fMGbQQIMESXMd6WE9C3YnZ5MH6x2UpDFIkzWsQJQA7KZolxExV1s5ks4RNysoYkXVDzvo/mCmX
k4oR9apqKxMCecmDlaBiNOoZiwzn5hqEyIJKPLKsH9nSDyj+JnoZMyQQvyMZlh+vPrf8rCFqY6hi
RkbrD+u1Mq9vMeE7pidNai1Srz9yGef2OGgIq/L53Utc6vbDnICqYFW5f1xEB75dcUvzqG4rdo+T
5CggBverDRcHd0mfv6/cuCDA50UKoXchT7um7hrHO8Bpg+5LcmfN/Ih2pHLF3ljBEhcB0vXfOlcK
Iy4D241vvk6g27GzhLpE8ygbJd5gdgAf46O7SwseHXBhsP9j8KWZt5BXtsTED+LI3kePgYlW+5RF
uE2dDRAmi02Ick7uqMtVEvW0iPsXfaZBD4uIyTkVxJEl4PuvxkRMzxk9UpXqxzBED4LKQu9Xx0mO
TDZWT/WXqCembv4/MjB+VKBed6NZzUIVa5hoa/RHKhjwueQLtiOCFeBXMECrtjcv66lhe7vfb9z6
+5/p/1CVftcsyrdAPnK0cRwNJDf1EAaYh7BPwK6H30ueXZtm0tsVo7VdSz/sYtSzIdG72vXqeyCt
kntpF3Ak8hJmnt883z/0Lav6YRbzEKfW90EuPMm4AiewTM/zdWNHdUN23cJOcLrF77qEGEYDe8Sb
Ridq1vEgTVRnwCYMu4+7sDFYg6jXRfk=
`protect end_protected
