`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jrgcvB6NpgzNJdRVHlSeDwQMVl7aDQyabgapGh7rqmEjznKI1NCLrR9ImJTcdoeLOH3xBtfWWaGw
yILZZ+w5TQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ag4YkSmodLksNyI//vguhKIb+29r48eSSBnSekONPTiY5KDvwEVk7FPHt2IwDIgp/+lHIEVNuvl9
mSG5KZ9jPHSPZPyN/4vfwOqsa1suwTYwLnCPSwuQv7t2wLyPCu/QCBXqrtpbIj5KiydhleAx1/yo
23YHJk0egLp0iDQ3TsM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVCy0uaMTpqXTvUIzq3E49Qh5tjtPCjUtR5Z0GJzxDQt4fBZLtMlbWao8zrxVXXuPptlCW0nZPN7
Pb1wZL2OJBvZdpUOT8g8t8cHZrubY/a17tJAMTFLjFUd2Cu36GIseWCHNz+iflFRrkSn4RfZu/Qj
2DFLLhHmK6zPRYo48n6QUALR7JLe2Ls3gt6U+JhzuK+AMijToKTiejQK2QXcgoz7swaa3FZ0FeLH
ykamoUQWtwHWo2XRnvRfbr44YvPS67/sOTlSxJ9wISSVlWulUVdLnbgt+BQkbR8iZL7Gkgh7Jf+o
F5J74x3vJ7lb1i1WkuSsGrJZl+WjFODRBuW1hg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2CNH0zDSx/qy/S4Wzv0Ghu9L67oywnGBNit8FqDzTy7nb++SXXwHCNc2D/9N5LhjapQZrwlrbfgn
OcbLtgGWd0I5hDexG92TQhNUS6RBfFrIGcZtHla78CUuV2C+p07h+9XVeCTNAHcy0msrkbxXSlkn
rB8273SulEPyiFiT658=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R0RGo4b09yf7xrNRZdxn1IK5E0Ta+4gdve/4VDSCQ68Y+u8TBciR3+qCAWIdzXJezD5JvN6Y6ecv
zOfXJsdxyQb+mcGNqbN/OMeAHTzNiEwwhjfobMrn4SBSEIcg2Tw6Om0FRF+Ibu4a7C/UUE7zsL7j
TcT+QCn4Aw0JXsglEuMq3U0nyE1ZYHK5dym33Zmvlwt1mm0pWZlexHoVJxybfH3/gDwfuvSbKxOy
lHJcet/xY7TUyuFHD1IceBoktuKyRQ24koj8AatheSSbLCOOGQsiQNqvE2CEQN/oHsPg8Fy8Sfs0
1gpTuG4liLXH7SYtNDO3iPLq91fmFtMZeSH0Lw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51456)
`protect data_block
H5QoqV0rheFNVhteN6HdgpOoaA4XLf8h5t8/Iu+b67XYyZdggzkTCFvHPzNb7XEywV+qt320bxGf
QHdw8OK8ZgW1yvOGBOZwTjniMPQfElt5Uq7vkxXfnsvAegNURH4aoVwekr1gNgZM2r0PApxRzlhD
JDVn5avxh25Dw3Ukv8NxNR45eAS0r0AxqFuRn91q5nNFNOAl2najooWcdpq/uHnRplDaI3vzvKRP
py4wrn6NVmwaTjaPzg7frt1YMnROPDguU/Quuy+wH8ji6jOo+C0S7jFV2wqNgLu51j8JSam1Mdyj
BbUpz4f031eJ0PpWhcZS8SkmHXXfAdgTrStlXE1yjokV4L1Tx3jhIHkCQcB/zAx/EIe0ORU8O4kS
oIVnwSgaIZULRyuJhJ7FLLD7Uo+a/vvEIPWR/FW3ZD9sG4upMv/bTRpnuymOJ25PDJf983F/0Dnj
uCqaqilr0knZPXgG5Er1aLNfRbw5KVuORVbFx1eALve5+6GpxDFt//I5MLpoRfrUv6O4FQ/EqPsP
qrr7UcQqONcD8nPDN1CqCaEukCmpXEIfijltoukEjLgm0bkTcL75PhDxMFdr28+8a2qWCfgN7IL2
K9QuMF1ggD7FZJkdOOYN7SukMACAi+Be6bJ/uQv+4mSfDUL7cLupQu6EcvnnbVOFhmOcG+S1EwZf
4roSeUxFrz0qjfNoE6sfdJL9RHkq1Z8vwI3gdHJy0IkJyEFszvUks5mTZjDbhYbdZoyIONRBYXTL
33KySOcyg62Y4gpmEz8xjqBjJwfsZu4gmo8lcwW3eTSUdSjk06IzQS8ef9rjhCm6DkAg/gY8tTNR
dPy/c4V5zi/MmTw2O+4NNSY5wJe5H+kSJDG1Gh0oIHm7S/l2o5HQvFhV9itPUUN54K+VJs6Jfg4f
zGoWjbtKe8ksQ4uD8qi1yJDw1PuUZb5OuhwW+nM3Bo73efynlATAbL2Un5pEjTRxrbST89mjmeTD
HLxIEp9M6oQhtPXnvSpU7yuNaknvSs4lmQoOhHzFfGdDYqE7exY2J+5454icVTOH48H6OMeRwKyb
FJrzmEEqwojMNothHMJY3VqoklZleUgVKDcI8mhZ3MdCZDNg90GyUGL99sA1AILLMxNN9zNKXfde
aU72GZHAHve/IDGhkmPbVGvRPDMtT15PcG4eLjqj4j/5kL2bnbIv+oNOFNpHcjaFNb7lNnqxbaZK
fj9uZoHUK1DHVGrnefSWSs9eqOLa8ACSD2Uh6FBqcbiSma2NEwUiOnZrkivr/wHRsY7GreYDZFbK
qvXw6IIFpymy0EWZ9P4v7NssCC5TEIv10dOKKHcatmN/P3gE3mDaPsupg8oZQeO+pF6WoL+LEOPP
P4iJ4OsZofmL01nB24c2nEJZtarS+iz2puEEfjZwEdkKhsITbt0XbROVNegXT5E6m0woXWaaQ6RT
C4Ev8YX7+mGCyMi7gsjfzE54C/qkW6XfdESSdurF7sHoMxsIIXg0MfYmFBZIhZfzkHTSpoLXzqiW
QZiNo69vT7vEynrxT+9GjTjUcjOSEn6XubV23scdBW3+GFHpG4fEvV8eMsvs7gNobV00j+C5bgjH
hkxKd9kmt1DnLWxgQyZkAiSlpbiBkGczix//vFF4TwCN8y68X31N6ms+7Qz0LbHLSpc5hbLePUUD
s1C06iGfXqMvRT1HpmQnV8hS6fteiCkKG0ThYRKIpJ7COFXqTRj1hyF2/19yYvwnXCvw5Yn6o4IG
t3I1VXWdnxg4QejStjyXCjTqRiJJFwolaHSx9YDpZPCswKCJC7N8tou/MXTW/B10mkQ1Xip2b/8V
xe3blbxhhl8AjfTQ46EAjSJNG5ZZ4KY0lbKUfhiAoL9WRonE0tiyz4R7gedVsT71TkUnVpYjoNRu
ObiiWw06HitRCR8MfA47cChFDP2slBPzFJV4GqgLjsQI3Cjs7+TPU/tC05atztD7TmqdatP8oCaC
Wmes35aEdSnqiZP1exJ3v3kShSx6LRiyQGfexBxpC55c6F/DpDP3Gthi201KkdFf7kvqkWoVtegb
mjKXjs8TeT8X9AliSCVPai5IgLzgmGX/JB1ArTvqD+KcUhu1lDn0Qpe4fdvxz6fJ1dq78m9dCMjo
ygvvTvBmicaKCqwiBvazCua+bMNiXOfl3xEwQGR+aX3TXsZKaqj6TeivfYLWkYSHKvC1WOD80vDY
u2T7OKlbMTBWkflLXzcEJJzV+/nJWxiGx8IpCwBY7BxZ7WiYBYb6MFKPQ+pTu9jhG2vG9+mZmTK4
OfF3YWKVethRaitI/2BLUB+ARGK1BpILHxafYa53UcZsvhaZ/RIwlgjLqbp4AV47g+vowqqTk6hj
nih/jwSy4GAHwOHu1EvSjY8NokA6U1YiMz+1HnKD9or55+0ZYWxD511bqBZoku8o4IhEg4IE/Bbr
r56aZ830N7GE9m7wOyJ8joSpZFHCed0U3q9ZAG7ivqrBf7G16YjZa1BzLXBUTEaaRbytP2eGPzbR
zfwB+nqgop1uSiQi9LzThUxZaJuOJaUOo41gVv6x1jh88GGspPIy0fvt33sh5hqmBwHKd2FLROOM
5cywRhtK8/6IBipJmYLup26Nb77D7WFW7omVQlZMsrx4HUJhn9lmhexr10jgrm52Lkw9Biq04HhF
MKU6oNzIEpxcSHw+SRAjfKAEUcaeaAiJkWxz+A9zPFGZn1UKrTy4YtQMgKzLStw6yisVBXW1X41Q
hTsowtUKjii0/pmP9BLWECjos8qIFEq6c4ZsGbAOZ80vuysC59p39HFLA4WY6eI81U3/exVMPJYI
u5sqIDmu86AABOj3WJs4jyh9GPJf/R3Wf+7IWj01Vk1BfFZ/z2OHZ4ZX+QM2i8Z0THee4bM5xaWv
iVUD5YJHtZxxVorVL8PnHvGqA4h5T2VJoF5tVKE82kHBgjhUb0iLG4cweI8sqNq11/0uvq1dcWsD
agvtDF/1oKq136iRqS5zbxOfCRiP86tISM03KK499EYB3w5/OB4mbXQ5jHPjKNR9NFYhDUOllqzm
vTBr/7oi7qNP7sOi5rCj9JMol12uAX3wl/W+qhsGAZzcw1gteyX8rX2IbIE5AW+B5kf4+lyu2pQ/
WsoJd/Dc1pz9sbjILAmHwcFUaCXumID11Z13/i+IQY9Z1JhfUyh7ievjw2oeTNqTxAGKc9XKg5KY
b7iT3KlutAssvCrttdj3kiZ2Dgbilz98kRdiNzYn/B/ClDHFAK0EJHz8QJarJ/rE4iDa4dgEmga4
/lj2Ki8DvoppnrBstL/5vCFne+B/mObj37NfQbJtVZ04pPupjL5drK+uUiWt4MnCB9R4bzr/6e39
SQcsGOd/qjWR7VC3N5/nMQoB4vknQHyD0HU9d+sEB4gFduU4jC75gPBOXFpEAltMTmTBIartHopW
fQGRb9k0pXvWwOuMk86+yJRN4G/3+ORZGrrMfEn5J//HatD3ROSzYX5LiYmx2Z3jdSJsOD4ZrpCq
J5cMQwuSTv77Sd77zxjDt/YmIBqjawouprI52B8Lws93DlSftJJzPZJPreeo0K7NTKIkj7RHHhSS
nsbN4o9O6xtA4QcF/6+snyvPqCuOerCdVZZ3AWWGV7B+u7r8zXbN6IxT4MQ2WVNS5QKjTPVYql9F
PHjGpyqwfB6MVRrlsGisspYs0uv/RjxmpUHuVnNuZntsfdiNGkRhUisdIwxXdnofEplej/cJnGdZ
Oo/6Afk3Kl8Ju3nB3UZT+O03cqG0nmKRsCKOspHAftvqlPE7qgL73qonW3G3oZOppO6m95AjJCK7
Ss4nbwpgam5SfXtj95uvlslm/cVJe5IOWcmIT/IDp+7SCx7xiQaMg9GhBxikrDopji8tlNZ5bJMj
n/492BLSwxeQvaSXoU4deUa0Ek8hbACZ3ouCPFAsetsFsu7djtp9OIW0nsuYOx1IrxEgoJnRGd5V
4shr4Q2l6iYK/C/bxZGbnHELtFQZThaKqkCH07QERe9K2Ryoa5FY0mrXP9TGJqCCSw7P7ZsmSsi4
gewFBzdP95rbSb9Cqcd2w6jmmaYnw5uZcwiJc7EtXILrnznuaxnOuBSXMySCNmv35FA0W2ifny6K
q8OPGFDBqWJTBTQVr9fd4AN1h28JAq7zWL3CtMMxdl3bF6d2qjcNWkBc94iJuk7+MPU8DCSnnlGl
EmzkfI9S6SUsIJAwiGW5wmHu/XCmedgZFOBUH8YCwuncqW+n00CT4FRtWL25ulYvC56zkjvLDUeo
lsVj65Odzi8tGyQMDVR0zJh/8DvKyAynK0jhegIvMLD2B2wLjtIduEJg8r3oFvMnPlwI+e7CSVv3
Q3rYD/xs7kMaN/b2JD2CqaeM5wwsN5UdZMmSNvzRhny/M2nxTeF2B/I+bYYh3d0NWccx8vPMCH9A
dyugHOyXnOkeoZpsq51eMUyVI3AnjvUiNR9mccRfmOvTKl369Fa95GLGVErGRvun6fIZe5s7sqGL
ausGiwwEqzEuzZUys0/lSiaVSoqENf2K8bXo/L9cNpbS2g/Cp0//LqgdNFDPn/CafHTcEto86AJj
S335VPX7kK3kuLjGwTB8gzOtpa/+r4uHxZP5DuZYO3ebkJcFxzu0oacMUH66fUvB/+PMMdfC4bBI
O+jUmU5lcKyR/kajSZxAK1iPwvHW5ZSTOmJ6GjAImJx2qMdECOHQQ49gidLLzcewAjhOtzoURu++
QnfM4Gnm+i7vhIaCCUm4YO1zAtCjgc8ufzBtpIEN1v0mo0nWbpx6tcSEjbxVKwACFsm0kHykrEby
U5UqxBSs10dk2p9FVV/aw1+K6dgb0/2Kgpfw67iWuHVTcz01bD2YPg6IbwpKaLBFplL0y7N2OveU
63cW1zYNTnW9SAJUXSgJHgjKIwK5qgyD+QlDqBJ7HTjb2aTJ2479/ZpFjbOQFe4MI3cSCNEBQToA
dORo0mpAXXXiErr+Zc233h++vc9ZKu/OAwHe2z66CgevK/hJemGYrq8ns+xlL0boC+gvpIJ97g6B
GSHuatjZHVoiYSzoV1TBn2yPa1g1yw8tx+N1lMHVigTS2GjqvA3yyvVbwOHqXnudX0mrYKDssRWC
O56iJt9NEQ5dW2DPbvEoCDaMAsX15Ak+y4tQ1FAlxTJjjqv/FHljhDheTogz2DdOX5e355yzQi1C
9sP90qSD/aeJ5GHruq5IQpuemR+Dbsk2Uyj5exGDCRKMfCgKZvBmp6uX0523JGZeBZYKWqzGJ/qV
HE1du7sxUxJnG5RK7pKUm44K4V3r3X2DIRqmwy7Bt+Cfoyk57ssq6iTWS9H+rPTC6KvWF1tno0ye
/PoYLP/2BCIxCGENmT1L56eel2YTMcrZorhGJ45tHdAJiPjeJk6aM1dp+6HhMxFXpD44X4ysjnce
87EvCW1f3ZJ+QStykJLnDFi2eWk5pOO4kV0zTHFWaF3gMQiu7lZQbBb+PyAdXA4twjMSQl7bRzN0
oOg+VS2q0Up5uWG2blmCiveWzeRXkQSQ54o7wiZgfAIsCiyuF7Udt8wAmHP/9G9FvUTilRimMexU
Hvnu3YTZHsFlZJgKo6O2b4wLV87gc6OnH7pDPgHV5U463ctFM4DIOqawa9a+q9m5V6RzFEf9Ygi+
/BLwsUe7fh6JJWlg7PIUDG8Z5ECas/w1bVWf7ULzj5u/wBVSvqDV08shcP1jARPXDk+Qgj++L6iS
2lPacG5ldbdk1RD+fB71HuFkGhDOrueh5DVbnPstX9SX0Hf5B2MPmVF9iD1LYBwH+6RzP7oMitcH
r9i5ojRQiDiE4gV3d+YF+dpZX2hq9PqbOdgiGHRof70lhAgvMLIOYBD0574nkRHHhNle8IdfdHzX
BsG0JH0HxT17V7cOkDhgynkxl4GL4wONw2+DDrfmDDpF808iUMMXhK28MwSvW/1LVgJSfYsZMwMV
fRTHVXh58f0jSe5o1k/vfpHaE5Aq0fJ/MrJ2WMwIF2G9gtUbQjNN0y0sPpIRnktL68ksNMK3dW+R
00jAT5i6LPbf8mWLM7z4uARaaffACAMI4DDHUs2DkSEq3YHaV3MborfOdNXwhheUlmEFHhZC5041
kX8j5teaGPU8rpQV7/1C/WB5zuIz4+tXGcPnSgcWo2JFI3PrhqG2fyFp6vf/1Qb7BVcSraOfLHXK
7yxIY2Aax6JWQ6K79sq+KjyxPf7u1OB5RPQ61iaWPbEF2B1I+JubkaljrAGVm+KRD1cJM5hA5Aor
xlE8wLc/YcKO2MubXtkJHXxcBxI+qmzZNjTVGIjqSl03iARQrg8HkLyPWLxwPggMSNdKifzX8lKe
t0K5hhjGn2xlv3T2wckP3f2GDLo8gtABfm0Ol+tGdBQYxpLeY5gOezP1CtOCUi5EanoskoyKp/SI
YKE3d+aNjVk5Y+pNl//U2t4KnpZI6SZUSJ9hQoMgpOXo+E1fU7Ba75AIhZPVL3430Vxgy1w3JJfb
kUetSUxwYf9MaOUlUjnb8nOTj0N/AgijBdU68TEjIyibCWzs3Ok69VtsaOgjBRQ+M/nL8GHPzerI
wAS1A9HtUqRgGFqz7Ms0Me2iBNfeDH+u/VipDD1Uwq4AzU/seLxrrYVffdff2tSRXaUdQv+OULjz
2rMioy6xD3PlBwu3j96UqtIwCQPhqdgVk0mk3yBadzCnJNFYET3z3t6ipdu1kEG6YIwvOm4Rc85S
A7mVoIDJ6wO6rkfYRUID4aVLJPfWgjyIiDGUQcmhKPp7Xy5tmwhLrOGL3VB+yc2pdmZ1kq5+3JRV
PPauFZsSk5380aU2uDjO9pjtsHP+pyHhAhkzGNvN/Yu7Z0939XPtp2Bor1NtxPrcj9tGC5OgRFOL
na+yxoInuE+ssHJ4BNASsvWfxWMkOr+9cbgPYVc01uhtLiay8/EW/+32Vww7n5ndkwftA0B7kWJV
ZBZu/HTrS0JyiomDlR61ZKut/I0AfRYnN4f0uHQAv4zDFVIYlqVuQL7cbaAB/DZm8pdnrEq8KtSi
nLGZsfO3ItyN34SJspjsDPypNn+H0IwWSmthOLCGtEWMMpYT1wUBfx+m3raf+wrM/S2IqlVjuGW0
dsdGytmHaY7i2z0/HgLaL/O+Td/ZWaPtm+9jnT2gKAzxhKil2FUTCDR5nHdm+VttDD0c518SaI3o
SkeQMBHpGTCew3Kwl3QM7ku55fDy0LrhkwkjGWMwgoK9y5meQdShDCPBeCjEWfF457JtU85grocJ
vUvbdjP+Ou7qRu2LMxj1m3xdmNOSjifY8oBa0fU6xSkuN1mLOIooQ+fkpaur6aAG3onRSuE6BrKY
NV9wSELGHznGd4SH13KvXeLK80iuMXJA11g+RVtDs9RSiuu1eIb3QJmV2y9zOcBMWUVIsJVR7Qqy
gZB5fqUEb5QMJWFmk/zTOJGibgLp5ojP7nH2XkyRyxacON9fYrZR27hn/XOpkbe1nKDLiQ7f+QSs
QoegshGKuEiz0Jcq/CUyrHwMuIcr96PBr6t9jZaM3KT3lev2sNIR+RR+DxGPRYHNqOmz3+/R+xE8
PnJJx6r4htdWc8Ba7U3O8taWA8SskYp9IeiTnGzRfyO3ggP/vnnpKarjZf1kDKgdj4aRBTr1qjol
00OO9VdnpqJJsLMv9oKVfiO8xlM+dLAC6RsBwFwchY24y4Ly5AA+tVfMI+f4KKKeJjIPpu6KVcMZ
LaA2rpBYzNdZ0iO59jpr/woxfgN6DR8BSqHQZhs8h5Byc1tEzzlw0NaTm7NU1TVu+uDxMopfBvdT
w8Qsjcz7/gV5JoJnzdjhdoI3Fiu/qK/INEnGkk6SU9zkZJzCyL5zm8G+Dd3Y6MsceTmamu3Grcmp
HoUnSnymDTh1ivirH4x7lsY0S/f6ZYgdNDAq3cvpecehl7Ke9iGyAXfsyttOYHfNAUo8juROzLFk
HyVoIgazQTSAm3qib+DBNbAx8wgNYaOdrx9gYYD3giC7I0n5ipfxdZmCVcK/Bjsq+rNY/IxLwjyz
Fj0pBAdGOmfBTwfNRCatW9+Wtq1fhG/F4Cgwx+htiYpubDv7IAfc78pp3uOQCp7NoxMOJZA/tfLM
hC3IHJIOH87OM8TMNjVAjjsItkfJ80QlOgjwr7KUgDtl9FoDL2iJd/fv4/LazIUstWSO0rgQcQC5
+LDGa57F2rSgwcZ9auuYYlVPgzMU1RQGXVAM5YKmFW0OzhItlGCLbKYUB0tjTb4vJizXx0BGX8sw
GjzfOFWB1LmKRRg6Gz9AmF/8W2JCXRP3T0VmcJ8ke8254msVmqOpIVaIkAn9TzshaBktNavNt0xa
yc8CzcWxWC1SFKr+xD3LXgaQCyLjCp4+mB/VTPkf/8iHhgViMPXzizXMPz+9dJZKJpjhSjTY1mQM
owUsvhSAEL/eugwP5M14KCHUvin1F7ij9HDQp2hKt3UU8qt1El2RiB1z1pO3qm4GAFiE/8SJ2H4a
ucGWWMW6U0pMQWebmTxAjl7m9F7hu6GarUza7nxxtJifUnTf8Blj4+O3Sm+LxXRPuasGoTwhIeq9
M6iCXDwoA+vzT8LU46L5a8sonOEOjYOBGRHnkUyqF+zDsYQTo3PdlVVwK+GfxIzx8HjGPJffLU/D
AFg0hYgqzJwlERtp05jUqDEo5U6H/OP7ffaMqDQ/CaFMLxtwLaAG88aG8OXtKtQoRwtmY975t4Lf
DMJdzv0uDs9+xeIyPNWdeF/hP5Nr1xfIGcJlaUA022HNrfKt7TA2EDKn1wtyp+DJ9MjOOcRBgox7
NMfIZlafEm0qIt9rKDnReULnCTzKQqa7ItjOhoo3OD1+A6UzT4fbAZTKW5az6ByEowbKov219o05
6qwbpCuYEEEVVuhGppUqGL/H9Lvz9NT1wF1hFj4OaqL3Ugu2hO01khGGn1X3O1omGcvJx25pnaaZ
VG4mA1rGiH9AfDfPbK7bn8K157qiXvkzytbyTOwZpcNeZ+bqJ9TXOhWA+Mx4+aTvOmbOYwL/Nhf9
WnoOZfbVQ4G7dIhL5z9TPdrA9edkARO/Im7Jxb99eqLg3Cb6yR3g0UUcUdeGrFkLRcLT6kg0nRv0
VfhU5t1M1I6VXlujn5EM9Lu7s9dI2t1Az8ZAmq4PbYsqc/5DRel7BY1VA214oQPkaVyTEdlKpQCC
mzMrYGOO3MhGtnhNKJ03BUG9xe0Sdk1I4A6odW9o4Q2FlisF3ViWS3PDZXIKAB7Flkln58vkn9Lp
l55UJNVF/MPojiXlL36f6O8a0KaAw39TTeYCCpov/DSam/ZlpPbfLk4cd7o0pVwAGWRNOzw0lq/2
34B05PcOXfe8rdV584QdyFzaVqq+bDOnGE537sBlcXJFxeMXqQeSNEd16/D+jvIna2gw4UayFihK
CaibJUawnVFeqhej6F7H0qbyIT8FITtezdO8FB4LcwL1rJh+tI5ynlfDntHwCjej3AhIuJ2Nf8bZ
al36Cx2mUt/p0POuFsajt32Q+ifd85qXRV7vybw4oGWCX+3SF7mOZ1pPzmGAEXEKYLZvgKE4a+ON
XcCjTXcywTflBM44vlBOHYvUjKBHBgBzOeXR/Ut+yXCGLUBy3CiFghaGGGFtHAbq0qZXmetmR0TK
FVA34WMSbV0mIA89EIwgBrbq9pgefpVZVuyAsERe8LWoLETcjcr7KLr3mvE+LJ8WV8wiqq3lc20n
jGREYVdGPkONNPm5b/VirVnA2P8YdkZ6/W/OporJuuh4V6SOM2Sgw1mMcBnJ/Qa4jdRMBAabHOrq
ZCZfMMWp3j0xVrE7Hm+sOXtHN6NCNORV4nnAf8vUepfmXe29IOKEpXDnKtFdcOsUpob5Sx/d/l+a
AJQXgxI37oPNMACn5XuylOmVSTNciiJjPRT2sFGk7mj4HcLh2xvY1R/NDX2317FqJX3BY0zINZ0V
YC15zfpOeHkaVK5nXWYvyQ/nGVBWaKzHaa2X7lDbG4TCBReWjOkE2ZdsuwZp8C/CDJyXlDfbk/jU
aaZRUbNh9Nt9Voa9SH90UOZJErkIaLpjZBhuNwyhSTl1rkTbEdz9yUF6UFg6XgGwYZwbqtddlrOS
ZQ+ti4VE5F8RGvP71GgdwOdMrxltHZGLdmUebjn1V92i7cI+N26L+hzfcKQv4ZESahJ0diQskreo
FLUxRwyxGdnwFWI8XCpenh7vn1XKk0lY5bndZwvCBDGS0xR/7TDr7IPFSdDJOMksecFTPqzO2j/0
7woSiz/i69VpOO0u13yzuZRcFnEn+fS2yfkmtRl67o/0R1GiLYmpVcPlC1LIZ3Chm1q97/b8N0vc
84S00N1m4C5dhMdZXvNx66BLEHvBDT+I6Bq7nSlbA8mocaH57cPGhjw7eCOSWrnIRi7vvfjIDWjt
SrTupLd7bgJ0mNdwatEmzRjm0OKNAxFq9tP3o0o0zKf6CNJGRjk9WtKrP4Efw2LcUvbfEczji6eW
zCv2wCkxCli8tPI22LBrpR5X+0Mv9Tm+rdMuUhJIu/t1Bt12fEx8fuydcqAgNC+9cG8YD5mbYKSO
b6AON4nLg9ZIXLeP37ON3Qvx6byzXLHmLgfSZZili7DhqEFJiINlBbunMCmG/2CI8ZRtdrG7LdFh
kBmlYdqcc/gMQZcJKnBue4zFBBeQnlN3xeyRapkAgEqntVfksBzWMqdkPpukucLKfCvPag90TfVO
Jofy9NoXav0Cwk8JdHKz1m6W5qoWaJY/ruhz+tHGzLPrUu+1w7hj0RFUI0hl1fV7tOnrwdMOquRX
Jnzxw8JPzKex0+f15vk0Ce9agJTl4AYXT7ihZYdJGsiAauhF9gBLhkIcUhCXEfWHW5Tp3VbElG6r
bktkLwoAWjqiYqo6j21zW70VKR1v6my543bOLTtLOONdzejsrdeVOAwQyPhoMyq+XY1jMiFUzlhR
Q0LTqVi+bx2IGgeRg98GYRiE2ZqNOQTNgj3pPdcC5T7eOKfm4Z0FbtdO76dXSBxGopZmaFu28NMc
z3CjknVBHueWU4A/goKaBE1BOF3fAFYg4Qz9pFd/jkeUa0LWBW8hHZzGObPU+35WyICxdVcd4Y6p
cStZAK8lrcXZGW7nNSq5EV/Ef5BwManpRkZK8J3x5Y2iBAA8KMvSjIKjhRg8TjKjZGaOJnKAlQKk
ZodEyEMNFFUsZRjBZW2OhCrNX7o5m+cxwpwuuMi1c4bV2nVddzdiGbve2fzZ6p/4Ab9enkSwDh9Y
ux/je8Fes2s6P5+6nBGu2Iw2mxUQ+QP5z7Ll58VNJVbe2jPkOCQrVDVH4CB9d4DCJdeEr+ZHw/kg
x1mH3zffCavwqpNo1sUBnOedCkIhvuDUzP+m1heoy8qyGO0EQ3Sv1xBR+680OVHTwXeKgt03RA6+
OTvM9QcKczsdp7leb96yYqWk4tF1HCt1jbjGMAdIK9dD/sKp1rWMlfdZ0+VusUieNfKk3jFyhBpo
h4nxvrwl2ByQHq6S83xJZjANNlkW2ntTugvBVQhIdbj7RYUc3O6Y7U+t/ulr5TFDMiB7UBK/C69I
kjJ8a3gP5cAxE/OoUttu1WJX9rsDlGk6Ty3KOscQK6ct41PkKzfNNY3XLdkHi8cVlv8znGoO5B1U
lAAFVhjac8II1/c0Dce0WMFr0sH/GY6YcDmieDXlRehLAVPaSqG/pjvPQdMaxcbdEAGMdYE07hEi
s/0NrURuyIbgwA8n3ZzZeT6McfrKdTeut6UtGu8X0pBQMzfuVqy5Ql+bya507d+P7kz3B/YnNM9b
jWNNDWk21DTDYzhfXEtjNOPbeLhjHHwqj+afdwTihb5PdhCZDNbF1NTtdqg6saa7+M+fWhpFLo2Y
V/j/5OCQ1LaS8hY+cXDYDUeeorzbpfs/utYiUUNWLXIrkpVGerfMsbWqyOUpODaWJAewHtgcbyUF
S79zeZaOjEAm/Xh4Cl+5ntD4r0jqQObLLP86t/6KpZuHGQ1RBJGYy0DFo1W6BU/DyvDoShDEmNjg
1EfnEuAk+m6aad536xhEE3n69MAElorKt6jmRJe0ggePofSqAYlXJ6fRpA9c5Kuj7kXp5WxfDZpj
zVpreNZBgK6lyulaOgtl0hWqxtEb8dGwyr0/ieNtnYCWOTlxhSZVC+DxasNM2aadKmLWz2ArhNy3
b5wZBEIKpBjL7o9EFptJvo/j34292p1B+dY4yy9qsOWsEP1e1kWUvW3VCEKYCgaN9wAogcOOi989
bpU39uKB2T0f85gWr7UIKIWWG8NR0GoTvaIg0Qd1YHk97CY/G8Q6Fe1RXFF+nRKDhXJiH+l39urL
MzEyp+S6C4bhrSX3dvgtrhxcsV0f7yerGUDofeyU3Z4V2xa0DFKH11JIN4wX5Jtrv5ZIMNpYTGQp
BVhpL+AbwGaqb2JkmD0E5LfRAJV55PkywUrNn2Vcc5/G7nOJ5/op5eodRgdGs3tRunOMsugJ2k15
tUMRYpnrlm0ThtuzT0+IH9zCItmz7Yytg9tPiMhsY3LDOzhkhrroylsdySGC/1qvdUq2DRXqPAxO
KpD5AyQbYrFJy4aF2ykXPow2wRf3aB763GMzQ/4JkgwSWspQoALmfcIKs/xjWMPp77f/yMwGb5f5
egYSVOKNSuRcdfaXN5hB6rymqL0Sfu9zMJj3hfPhNPwdUOVXU1UxENIOx2ISl4uTPr0rXanLTAvE
8fVAT4LdPJIFTUheS5TzyJSWkNX2x43P+An2hEqrRwazj4gV73/2Q24MyJCCoZbT0exBOdm+zLg+
JZDwYQKO5BiXDujpGXFlidAPh17wqWD3G+DVJ3yDc1Z97d/4mIYhE1+5JoPWrA2S4xEaZKs3kd8B
yeuglTHB/FmZDa9Wc+f9e39VhW1OVzL8/oqofu85og9XKMUBTWclkE+J9x183vrN7rnKwD8USg3g
uKGAKVZSOq8qpAy5mR02cVBaTOU28EJu95b19fZKru7WcNUz0oDd6mFW3l8HBs/AUH//s3+j2OfL
KpmGWq/a1q6rjdzVIueb08r+uDj2KazEXqGxs8Z8jff72MEjN9CtpqKU/NXrs5uSPf799BFeMxGL
Fy9nS65f13FvZuhjnfE8bRY5QJ23ewG8ezQHg1ngLiU7UmiJqPhTTYVhknU0tQhftZX8vhn3xQqQ
0CsKebjYcko7EUw/ZgaaiMglNZtZDqkRZ2Yoc9/DAzZLDeMp02LEJLkInMnPBJC8q5BHk2KGp57y
61M1OKG/PujZl54cGgA47DLpXDH/RgHfQDmAF2ZXztkKuRcHchb0rxHScpxzPxQCgSD9PP+yvRS6
yjngbGLqiZeJJv0JwABwu4JleqWCrH0OA3L0zLuooOCOF8IlKCLe2fePsI/Hah47eys9D9B6g1g7
ZnSZCi8IY+eWX7IZlKwdF1x7Ku/xPaDZ54p9FBXBYes7oOjcQH3h/icht5otjBM0JB1ASPXYXalN
drKpHPqmNeTl0FTByOhFOuPH9uMYBGeqdW8JUyUPhIrHTfG+47/dg6bZwEH/gZ0QmvMbv6Pt/J/q
hqCMDGKgNm6hdElAMRpI3HfVZPybG3+J/kQUq8D3mQrLTS73TVxQr7TmRabuEKlYZUARkq4H/a4W
UwzCXd3h3/Ho5cKrVIOLG4sluEpxgnftld5DfQcm9ZZf7OlvI/U/Wpf+Pe9zB7kuiGe0IwGal926
TVD/r0uIOsMMlybON9mn5DlgVXkrby4GhB3EhWQUutAGEivpojf8iCZfEpOtOsCjP1l+EuljcPVo
/sa/zNp04dr2cqCuF7ZgPLGNg+hZI5EbOPZdU36sWUc+iCzouwS0ARlWCBqii/krga4wPnYRmfpC
fOPrWj9Zx0lgVSypRrVsdcHxEvCXVbfViEe9C7cui+RFQwPlKkXSZ5/PqZ/HaSjw2tJvEMnH2q9e
l2FfrMN0i2Dc47ZKLH/YfQdCrCoBFnHl1sk8oZMC6M8DQFHUmiY+rve4MT/nlaOsx2orK5oDwMVY
6mpBB+B8sXQbLzNJuelNHTXD/P0HglVGwGxsztA8DrmKGIuzCazbuyBNS2aTyfB6XrFbTGa49nPw
kJqB/nNoQQjWg+n81yszvT6Ayshq0xchKCaZZZ1UlOzOmArrUMYY0Loi9qRWVJgsCzgwF1wzLqKl
+9mFOiflRKeuwwMlraHYL79c+e2rWGAwtpm6bBfaFJ0dXI8JmUtGe8PqrIA7jRkqGp2i5ZEyDdRg
I6TjjACeKetdF2oze/hW2LlqMYibrrS0qWMaONjv5qtq02+2+B8axcWYUulJLw4YRiW0wUt9frpX
gRBj+1gfXdh+Txw+n9a+X2PWAN2j0JUNWLwenOj/NT/k4EwoYoMcIHwH87zUANadDV9udrMTyZUr
pNpwIB2xg47wOgBr4fpHwi5LFEhzEvZ5aAaWqZhORK543wdWU4GG6iS7B1Vb4IV3gf33knYf2+YM
08sl5aCAIGhY9eOmAjXKsZJnt1xomYlXTvjaHWytIDOcllcOh2Yq2Etw+eVnpFo4xDFi8/xLrb19
WwuaPFSyHrp0r7KF7BfzXtM8etiBoh8vP8CcjBvtaMv12U4BAvhUQ/izelVPb7CtmG+XImNKPhtO
Me8BZAYWIkFPRCejQKm5s3ruam9ERaY2RMlNuqqdp3C9rge5XbZalLmxkUAIo96DJByoTDKL1fkJ
Rg4SgO8L3xVyrGmiM2BBBmfGVBkLdDKXGOG0meTxBHZKKrbyD+VbSTtQ4GhDDZAmCgL/HKk3nRBO
L9+dVWioeUMh/PzixgJTzo5JuYjXCXzmApnDtOkC4ZaApP6jMWiScittCXYDkKZyqH8/GRtmp9n6
ahmZ3SQBOplaq6k78ytN4feNavgis1lWglbE8pskSjZYfHnx2koXQk5buNxxWDTw5/3U+kIDaIn/
8PxkL5vZlzUAFJrJ7oo/6saME3jFuvd7LcL/unyuC0GExK2sfSQHrQtnlnz5OV9WZxoUkZo2aQka
zUDR5jrvzEJJn6ejU17rHNtqpqj5jWZ3sNTgrWG3fAFxs+uypezwZ4qYEbOaQKdf2oVy0zEN4z5e
x7+lGu0SZRQH40IUbuDZKnuIuy3wkKEGJUUlOWOHyBozpwnCddzBkZDKecWmqzd46ZLOQWyZec9+
6DKeCV7NfwGMa58bHBmrA40f2Dup8N+xK6kmE2/RgFpVJug04zbw/IywqqP17dKP/4r3CgbRKC1h
1XR5qMcWOTazCkfix8wVtyWoXjSk/MsLS9KPOSEolY8SGxcPNKHhXnbYzAzCTyZqC4YsjccQJgn0
RT8XmcS0gPFKZDq1iLbR+JgzHL5ehtuX/u5PQ89/d2DAq8iPtB/hj4spIVxNuBugzKljKCyZex3t
AfPIO7kqEBbCMqwt3u7zJZWP1tX3yArPcWKGnem0tYYor2kWzOT+meShTpEL8jtdcy0ZACaj0f4a
RGfADhnmUUmMa0Jema/4QS+oYRP2rB4Vjq9I5uGmftg0Ap+rABgMLHQuGLop5OY0NUPago5c+sLD
hjz2gr/ZhiFzgUMMsb/0+mK7tcNtt3B5dqbCBgTNwEhNMCWu8FqR+LnwmjkODU1YgtzbA92twVB7
7m7yVl5dRbKeXtH6au8DLN9LiSRFBJ2shLVdS4svH05bCwW8+vbejMwhypYojH3Ne2yRDKFq1mk8
4Yfn0rbdldYgiEdWoEzclq8EkvKnwh0cqFLY2EEpyBxo2uSTOYbsUpUQYTfzX2Cmn891pkYrAVh4
lCRQExd6wATzZ/nVYCI0xJWh2upaaAEthmvuUAsjmrL3Wd9bnj+hikXf4fSxqeh+cmIW8lF7lhnt
7ADwcc3P5xykKsJZvZXGkhm3uaON/UvQN1dJuiT+qTx/Xgw62SI/zwzGTVp2Ps5xOJZ2G5gLstLW
4mRmAJheynfAnWnTlHcoYckhdHZ2qFsvgFaeHP6c7HvfzWAqg8Rbym0MzLhFebMhQHYI8Xl01gV/
6Cz7Yj+Ym2g03OurgGB5NOy5WqmEFbeRLPJMxI9NPCqTkRJe6vHsIm9Vy+01THTSpRBqQTS3KXOf
UGqk9j5K15pBCdQlsxuOYyIfbVyNty8rW/5GctSXwEk7JKcFgEwjtOLv6eZ3Zv937T9tJqTQEzCU
84+GVNQJAHAFu8FQajpk6ANmotvFQv+wDD0Cdbl24nWenl28GF2nucxon6suhvSREWuE6rzgIQA+
OpABAqU//xaJGZMRZ2nVGQW/n7XxD5HcJs1Q9dUlpkmMYozxU3aE1WDM06B3w/ItT5n0D2Y+mFrJ
aOuXMFkt+A/rT+qEBbcSOEjTlK6/AGY08XL91fE4inVH3rH+PAX7ZJkCrxy41jfzqH+aofskhGZU
DTEYWSDeg9o1LO70ga1X7CMWJEVu8e73CQg1RcTtO2CRBW+q4yorcgXrXv5mwx7sHd627c9xbb9s
IeE1gl9zjHYj/MNCpwVwsWfARdgrNbQs7a8mV2L6CvDl9rdgiwqTU3JMbrGqNUpsvePa17450eMB
dGeLf3O8uEoE+vQeN5LYTqMpDx1jNaJVTeppXU+wNuzAnm0V75Idrs3EuDSfQjGBZ/St5yQW2IcB
hbxrrBN1AqO62rwebs2KaVH+eQdAUolDod+AQMGhfgYFrPtIvoU6JzfzPcYY6uXOaaB6dHZCU2gg
ZQl6uH7eYt2k0023JS5ITirdvDDWmZ3Bnw1Z/54QUGX5vbJTkLjVGqflVNa69QPkf5Dumq1nYJ3c
/L3ihvzD4ifIhqZUeAm3+w775Yo3tTd02WkmT69OTXEpsvqwiTnoTM2IoGhe2Tg8sCVHPUFiz9EA
fIsKDvpv8MRY72SxD27bXDpzLUoO1a8LoAId4smao9VCz6IBCEcf0/tRdrL8DI2YPTxH/8oXTKf7
SrU4l0qei//+dGLzALy3SOGFnyaHacPQsmK1HdR+n9BoaRZwgB5xgkzn4s7qLHmnPRbpcsuz1hMm
WNdyne5jDC18WuXi4rRyT40IIn9rH25w4JuIB8tVpTuQudUEnkzUoWAXUd4RCRA8iqtCJ66pL6bK
Dc6ag+sRd0P8rmBlo3P7IvFqKCuijiHQjLOodfxoJnkYkBaWR4x5W7AEnLM9udF9P7t8k6TI9yh+
f2yIbMf+38Dkbb4XciLiT2Xbc3N/hyHWZLctyHDL6i8hcR8opHae6WHjAb5WUUzAUBRVBKUdqyFc
xW5hIMg31NpCoCQRKVzKsJBUZz/z+XuWWPG8nujantbkti1qe/hqrosAHQshVB7w5FCxNeJReUHr
DF+HVmY0JeUm9E0jnng6w2lX747Eim4S/DxEbWAuOFpm2eN71Ax2asfvNZtAJoAaGgWKnmVUy+UH
FmQnboDH5tyMj/0BR7gbIMG2sdY5y7ye68fqhjkJCvr/ahrnA7xBGFCrWE5x7PuwqqCMk1j4nfv9
u2FEsnSKrENVvq6Sm4sfUv8L9KwXOl0E0iyzwsAvnQivd9H5uHbiUeLMRv8ryUP41kHLEqOXzP4d
VIVZHVf1UB7kW6PuTGLfSwQMS63vcdTqvaX3SaMty0EX5pMTZ+ILdDnHNYEoYnDP+2TLHEUK7KwP
QWBE4Qq9e64dgITdLLe8iuxKLUFVorSG/xxpyiYMzE591GEQJW9cOwEFal0hYUpzPOw4j8qMMRr/
itA1XKABb9AM5OTDTJcJiiK203WVHQcO3OHf7edW2p//CNO7hX2XT0IYTbm9u0lo/oNZyobMyhlq
vTtNEblMsk/OPBjG7UQnlxuJzJWpAQptMKpQMRrqs9ipCHXoWHiVjyMLXENRwWrsRCG2XfHrlQZS
dCcKmlhh/MmSmJxVm8EibQMkzBptjuvzdc3OMOTQrdDKnLSoh7xh5GDmCBr0c6Y3cXHmp9447UkW
NN1+5NrP631zRU0VhIB2B0xOTPm8UoABKk2pCtQgcERtMjkBkmtA/XaWFkf6uUlhlcqipTwGyw09
YGfkSuj0J2yiZxODm9hSVe+nOdi8HAwqYRzTzkUr2Wu/I6y8VKyACpUXNFi//aMXvW8IdCZHs8q2
FAg2evASFa8bU3fnQAE2HibhQNLiDKegEQ6xu6yAdmxDo0MPxn593ZCzGekPQKbsLfBlr6DL1xQn
D1NTTCXGqWkXqANCSsLts54MWI+ilSfL99sLcH1MmxMklQBwifcc04V6GPEqIGdy2X5YS/AEnFFA
KU4Hs63i4mk8YUKf8CYH6D2Tol9zm4685rLAp84piE6RACVS34vqAYKgVt3SACsFz0SeX748X0yp
XHzJ9wCaluZ8+XUAnV2G1p99FoLfVqOt37NNE9ZFTYJkReLsAONJ+u8DUfjd6eWJCFpIeqE+AEkU
II8bJ6ecZQWhh4rZNBseWJo5vw/DuESsF+y3DHvwIHHvHc+VeXUbOSa1yPYZ4j6P8c3C2Plx/VRE
8QFNNlRAC59B5vdHubFWMH9w6e3BliCbPKUTPADLTZlSa432gMrC6mkBpY6h9+PQlTCInulOkkz9
0WPNPNEbDrk+9Zme9obhp78wM8I3rkFB2TEwCwTxJ0cDw2PVG/aq1DHRF1Ez6d0mPMSAQ11mmovP
78I1XEkQiT8ehd+PBEnsKw0xHrUIvsMZqRQgo/p5VZIqMsUYZyDy+lXBx/yXrjbJsDw3Yj/S+HFJ
WnAXIfObgQYrNv4TKWes9fI8rfOg7yOtsVEx1s5r5neIyAI/Twd/SjdKPo42OT8hRBDrYR+Q/LRb
QJiFTlb385UerzJnyTShZjh7apqwzj1sBtxk/LA1HgLG9/08z2f56yuNmJ9i9Ugj4Gd7TfD34v5f
Nky0VL5I/wM3wPcUloN9RfsoSmKfp2xSG5QAKSe5mxn0Ek7Ewi7up80m/GvIPtGHk33AmXYkvoX0
jBtEHDx0PwzT598sY5sUmnUY2E0OQH6BHQZlfEwHGmoh4gr5n2mYq21gAvPiZidWOjCm7vzwNFkQ
Zid4Jhs++TmhBpRrAWLkche+t9xm5trFxqGdJzzvhUsZCYAGpTyFge+r1eebwIJysyK5qFybGt+L
2aZsb7qViGbmgsZ/k3o+peeX9wu0m5L1fyvv4HDNZs2eqpLu53ArrrgkNsKC3wfOjvHGPUlb4hlQ
451RxG5Oi08pk/krzvPY8271ZsDs2bOIU+VC/nToJDJdPyo6bCq9GTifW3T9vOuygzb6bApALWhO
Bw+pLSG5zF+eDIcQ07xUg45PNu/I1Irue6wDx95HRxv6W3Moo8tpm9kGQuYAfOnevkG7Jx2Va2Tq
lb+N8FWawyuRESIR5xr+g3gqmefYDiThVtvOxRlH9x7unhSoKubTiH0BYdN9zoAHjWswPzKQXVLf
uSWlxv1BfsIpEQ8Qtiahn7hkXjiBp3MeFIMq4yKdMNdn+iT10rl0feajQVpaeIQQ01GedYRwyITx
dX15rN83vSIqX/rabF3Lp8tcIiNWtpXpjDFU9mo3XHGBFybmd5hxZTEP+xZUMDtLs7g7eJu5a6HP
qUluXn3FNLvFU60jARRrz9zW1opMImhqvgiI4uik2EpuqbnkSLW8JAaWjyLS4GF7fpGQiO9Lf451
z+yvVQ7Ws5iJq1hIVVu9virqf1nXkfuHHEdGfcqyWWn3LmyDP6DtnZNf7pB/8f18u9F5AAom0s1+
n5MirmHHB4L1gJuJeTso0y0TquUVyLmNS6SOci2mwaRCsTobqfnS5T1q6cIwV8ERuH8oK/1AnoPt
Bk4BgYZut37oY7kptX83nCPz2oag1fxTE/NXyAGtQdElwNFjr0RE0F6e/eKXFWr+4jGDny78/VA6
4w6FNFg37DjG7kJtajpLP/p8aKCoJGJ4Bdp5TmB36hFf1I/dI+2xEU9uTwSVmailEn59fbPOy2dc
QLT2cxNMj1ZblrmXD4l81r5WuHEiPXXGjg9RU43ASw72SOnMWfAheZvoq4+7GJGMNoIEah8r3CCY
EhqH5z6GUS3XHgc48uzBHcHtoMgP/SmFlqs1YRw1cAjDZvJeFJ0M2nl/KDt6eIn282cWzDnF2Ly+
X0LDtidWp6col8dSkPbMasJTS1rZmlXO4OggZNRGZ6aFhrkSoHQdUGvcv96gugCY9l1kOyEUCtdw
3OX4nyvElySwWzixCHmUG3OF6LVYPMGjSrbX4fZsoKctJIgjcEdrJPmAXeNatbvOJH8iFXg3nQEt
6gPJbQY2sG991ibcGdnVIYEbT4qy7pdnPREe5m9GVZyyZx0Y8Lmp3qMlib0aHOZkVkjRAooN2tB1
M3ZVUsaZCsq/mPvk4WLx36CnP1slB8eeqLJWZpLjfIBlSnU6qs1ea/1w+tayCiR8d3sv7o7UeCoe
0FyY2RP0HzeSNnETZdl5yb/ChETcH7gbmC+UGR9d3bXAs8fhQ1VIta2NCDXdmFQcIDbhCSVCuPmS
iayV+EWOIv4vzt3FsfAp3rJsgqDltgejMMZYbqyuGtcI7l/EHXAI5dc2Zwl2wAZ1sJLjXRPKWKBy
NdR7DDedODaVcYVNFvDRibJt2BpD3giHdKk19bEXII4Z63s/E0otgtnio99hqNUR5ZFrUvfUIasD
Ww93G4RooeTGjPfNeSrhV68et80BisII6FcYJaax6IR+ZE/51AQIoZhNoEGk7jOlBbqrAUlwyO9y
nrWMpTI+01YHPaTsDENxMywhicCsyE9zt0JE1e11zNtML1cxKrUW8oZgIf4Yso99ZPs2bUJ8b1Tx
1kfzJkudiNBGgGkm42BVYvbba8enbRL2TtFDndpz4tE3wx9UiI0IXZLbfQ2fmq+5JNJ8SqTCx3iK
rY2IDalqjucrOp0bJi8TzSmas7gl0YR4ApX3ioLsdDpwbxifv7f9JTPVD8dCW+IDJmmtq6oSatSy
wjBgmX0eyoVKTriAYvV4Kp6dI3QX/WpnY6Pal/THx5sssS2lC+eHHQltego3gUT6HVBBT+GukEj3
xtgZkTnYNVB/37SedBU+dnjqagD1jtuRS2SLTEDo0zD3PICl98eQoqxQxxGeI+0qDoEhCflF1lzH
mb3q6opucd8Z7oaplXL3qQqFu3cqVB9tvge17sTHroX6+bh6DZp/cWOpwm5QhvHV+ZtRHnDfGxD1
0cd++MSJyPidLecRk2616Wa23FOuJF/a7xLIW0T7snGDew6thZM8IcB4aQ7nOTTiSVQZ/NtvJ+fQ
1970/xeMpY1IVT4rslfDF+RBlA2XZrOLsfHgt1Os0KcSOfrEyobaf37HkN7eIR2YoOhukfyMH0pm
1WtQsq+R6fNa8+AcC2Cuo1ABJq3zNQLkk30txCvS38t2EPvlkUEsptkcG+4uKkzKmsoTGdgYe3+K
TEzkFu901SVsUdprntMxdNwLdFFz0XVvm7NP45OVoKULEj06rB+ve0BFdNhFz7KmNNT5QuLttIg1
xRtTzGivsruioEAb5JassamPLKR10MFiP4iJUiksxXP1VdOJ/nSksVkfO779TLJ3KJXdYtInSEhC
0HsrU6iqYePdMno+AJv/zc8eTypkFS7jICuGN+td77mESaPY6HFARZ3/BEVlZuR1Z+pVRgrLREbF
Wze17CLlTtJAmDrvjsxb3OS/GW4/9hIuLt3WgtEgJQRJWT2Zf/2EXe9yeGvxpF26APDtWXPogoST
p8zAE1MFiX2gEYM1uxPSNu/Z5IpjGmZbmj0jZfOnKVtJQ16mWdP4HDg2sIPMVfzDwo4ubzB6iLqP
NFQc8FrA7aONuelRJOZxV3wYpF99iZjA/meORkWymDR78JUHSbnFz49F3e0QwW1qP4ZK3EZZ1IlQ
Lxk2UlIiuPsztu85bkSVEV4Jwn2BqDqWBOiSSPdCiB9vxoMcEIX8+AU254LrOLKAxSBfOCtmmBHi
Ea1gwbm94nwtG+d36dbLpgf0uhKBlGROz/QzxltW8z+Lo8K4u492I/aTET7xHk7I7b9wWIR/7nVn
WKZJVlOwVPjg+IjtNFd380A6n9zu7QBr4dozrG5lLvDI2BXm/nkmQ2hUj20yhVz/fb8vu5vxEzMq
RuqfnCbSBa602Eu91WQS/TSkSOuIasu2JNGq3o4HkMvpwWfsSpmz12lSCamTmyUEfzxtmvWszajx
IkXsA0zFlT8llL32owbqT9Z2c9zhaCii5nLghDqCf0GstGTIFPteE8+cE6o1v4Wd1iV3tHnU1HaA
LMyL0STXpjK4vsybDBFz58B62ISDvAgRadNkGYRtZz1RkNIMw+wFsKzuDmaKDEjiePcYLHau3sDj
9sgEpI6NH0Ghbdd+C9C/hho51HvL5F2sxXnZEpsdYyR0Lnnwkz6Odu6e5NB0j1/9NDWkRik9B+3E
KsFJb8I7wNOO/zlYV1y8xYXEaOZ6MPjkciuo1Ti/pgNSphcMP6LlXyoHGI6D9p4c452uuoTdpkMt
C+qqQmDFYbtOfTkXpAQh4ltL0PLnyq+tjKJPPqOit6GL317dV90V3sXSmzxKZChUa7njlraqKu/V
qKz0GoTRach4i4R7qwbGxWhB+pqcU0An2PFeq71hivhb2F4tDo3WdIgMgYGVopbZ0bbezCZd//DY
1l5JJyUu53/kRTIbK3KzGtjE1bxBcLVHuQeEPLlCX8pBByiqabFo7oqIHA13+zbPGNwvDDIGjN3u
UUyI/8MOwWJ3NFzWSRlqXd9OxmdftvfGKCCEMD3u+S+EBtMYpnFQiNUjVvlk7s2sU1ttWhxFFE/x
9XEOyVbBMZrSWHUkdT6MY2f2VMXqwnWdPB+ZJndUK8WklxA+fqpAGI7B127hn00h1i4gzO/hH9MC
tQC8LcoJtgXCO4ehrOKWfu2gEH97yoYdEYqoDPxZwV1KceXt8cltwnM/Yl9/eop655+kMp59Plvo
oFqW9F24bTH3mMN9bG71uIS1wsftTLry/mIZnbGa2GdmsXAVQCjm5xm0LCiICqc4Udr/oX+RM6Jl
0r1bfvU6+Gc7HOz/1QXX815z1qdyipaUqZ2G7dsBryZnfHgqu65mrkHG/Uu0lT/a9Q5nSLx9BULQ
Erye0Os+Gjc99rOFUlHsY1/BYad/GjpsfzOgBTk6sTqmW8rMu5ZlUh1/JHd9APiHAqbkCKUzayhc
hoAXvMpRL/B8khJl6Bf9KLi4Y8gMSMrtXxWI4BWVxt3M5GB4OkRdbmfkJspkmie67whIpPR5J1/m
Wwh5vQm5g6+LIKavfv1+3nFBr3SmKpToQxo4A69yMZ9ccz2HW3PKsP4kUKoConIVx3veOhvl3hzk
ghytQc3ILG/hQWTkPOUWmpbgzw8cwQRx0+z/5Z6zJrNKuxb+2GGDkQN+u7Y+k3JktUDPVnmJfWvP
mvz+qNnzQFxO6SC/7HjOkt0AresUIt8V2If9vvDGVZh1hhVlkytQJreQ9mH89GlVm3171W0U7VaA
lgSQ4erOMrw5MXVOSQNTggB20x6vYBAx3Rn/8RFK2hNCoWjmeT9pw83YvwefJI7PpbzD/PrpbAyD
0T4/boVk2EF846DWEuRo30BW+hPicEtEyfNKIGUkIXPOl7JZ69gyJwdla33gyGcXnTII9T7Us1py
e0b3NZRVewqG8g61NX+hCOXRwXTCE1bDRulc0FdVcoe/PIUGenwQjbSJ+f2xfPJt1OMPPqsAA7n6
om1+8uUufGJTU+9S/0tIME6NNZUCy0HZ7BG3uNF9f4UmHm3GP5oT55kkweGYB1GLPTsBsXP1d6qp
OC1fpuWLomiYtiDiXdxRbkhOepfLqKspCBzkAVyOdrCmJh2Lnb4kAwnzMRKtH7dekSD6fprOt4y0
xRcCV+tQ5lZZws5MgTlyPfgo7bVwO0J1blndrGtGo1VIlg+Z2XFtbG5ExHQKMkr/aB7CtvnUt8ar
WwlO1bs0hvZ+hv42BRYFDrpwVYhGjiB8Hhu48tCqZp8mxeOWfa9F3Fikr4L7LMDbimy8+R7kWvjP
a92lL5A6QmuW6rgl4dyxOyrZgddkIn51+lS1UCkAZ5XT7yctuo65H0kmORXD7Z3sH2sH478lA1sn
ssjS2O4qc70rsF+7kiehyyabvM42wQXoiKn1rPNf7g0ESOgWERLFbmp2XRUl+sKuTeHk4Kb9doZr
7vsX2mEY6fpU1V0Tm4jI9zFq5ImIqo7SicRAxMAuBKOBBBGTb9bW4W7cgQJsEP2zfNsDeSLQYVW1
u70+zNf6ymn+3qbGVDddoUGDkDwYpoG4KwOShBJ+gM2MoQMh51Sh+oJyOtOPLtbJs15i8vjQ7G0J
afHvwMRUxo36o3KrrzKd5q/J4x6pSzWZmDZZbOockyscJe7k39XFMCjgK4u3qEq/CRMNY45drcy7
G8HwqoYDZk/7YZtUlY56ZtKE9gljhcAto213n6oVHaHa+jr9qcE/cKD6T2v7LJoXcTbZXASUioj0
l3oTHWQ3KOTyxnkczgzqYJCzvCTTMvh19jdTYWTdPmrlKT5qQn/7Xt2xk12BB4CZbFpeC8K71cL6
k57IKeitvTBVwC1/Cpl2h5cnQpwbOeVyu03WZaABC5oTXHkaAw4Iq2KQaOu9HHxJYRCliVOHIsLK
vEmhure0sV/SQ3oG3MX2Ly9Q1Ju5ilgZrduM8EcKSDKu9/cfCJHAr9aZ+4z5hxKc4aMi+ebdfSZ4
MqcQKJw4nalfk2zKm6IxhLKwJbOisWOH14D4BU7ijb4Ud/go4Cs6ao+icO7p/beMELmmFCgIh2GI
WS0jXesvgwI+P4cw8294wXuILzbsCqwcFFA2IK1cginu0rz6dc/gjqV7HbYDaKFAtRnixXu9FccJ
UiIc69iZA28unWeMq504oBo1oe7+pvixbfiYWljAb/loAalLCNdYQrOxog8UaCoRDt74pxsg0RZe
qTTxtRBe8IknGKScV5669CCMKA9KYc26tW3a51dn+PB08zgmTaYrzc3GLK6hMeJyimQfLmmPAg4j
nFamyLD3lO8WnMoZ0KHpiAcLF7V1jRwM8tIZivWpla9N5K2FJhW4O21XVcEUl8pUASFIeYD6zuiJ
kuPgN3IMrwq1MrgVd39nrt84NGClbpJp0y7SMikvOZ/bh4e9UytaJKConOo1uGAoew0MpKLiM725
6GNs0KrRzqQrHuWFTbOc7kvV1zTnx+aiDEGQkcYlPBx7RKyNo+hUatJvmG+5sADJD8MRPe/OALhi
FBSLwV+Dg1IHz6eaBMy7S+ERlJkFVghcnu3Qm89Yua567bfURajgnckDiIGEw0ba0EzFQaA7UXXB
dXbwoWryPJcU1VazSnyCznfAKOfj1PgKizz8O8q0dRaqgsu5HQD0tScNT1UYr9mzBG4kPyeIEMam
buk8VLk5vh5uEXDHxcFlu9s1CBr9dOxdaHxuuMzHwIOwfZE6RXiW0osFTNppKcCKj+qEdr/wVF+q
jpM0dXVGh8bN3FGeeqiE6lDuAchjDykQcm/u5/pyRxYwAzWCOHxZT7XsH648pHjEq4NbCKm4x4L+
JK4uXB9B1gQI1K7UxPKWVIU5CbllUQ4qjnFLHkszvHHoyCdchEoFtohlEchmpdm0RD16JD3HFnMP
1Ywwu6oacLy4+CqLIEaGN0Iyk8fJWoEuMWp1zUqc2vTYCg+Bv1ULfvVzyrl6oaRG7p91PzWjgm04
Ab+y/UaNd16noYH7sOrNzHVffzxpO/umg/4DO2WGldoVzbi/Zrv0GOib1A/KTyn0vIJCGOn0bA3J
4Omw8T3gDx6GY2tgzbEHr8RkRMFYO2SMoULHzePDFdZybK6xiK0RfNtC0XDr3g2o4UO+8HD1GsWn
sVHd+UkTpn2ibohaVCN1opG6+VOc+YuE2es/xAz044WCHjiq9pOfpLBgWw1Q0b6xzOFkdUxe1vqn
TRiB0xX/c0BrkPpSl7m+Y4xDYxTOSG/mgWnkpshC4szLbFubgUOL/YkE4qEo/JlbGKZOXrG00JiO
bdhodbrNVB/2k1yzA8is4ZoVk/oq1svfXUHl35fO2kCf3QW5jiFUGq76wnnuhY37yQvCDeJZ8bSn
8QmYcWAQMr9A/Ay2mxwugVbV+wjJnjpa1xFtaRbGTBQ4+VjPSAqmaq3GaW5jgU0bM3M1Wf4I2wS6
Sg02K5vuKTBCjD8mO/kk9CCPNw19xB3mrhKMYaSfvm8oih+3T6nTkz51LXvHNNB2N3Vtxi/b2UkO
EdLmZWaErRYi3h8rPCmBmzlbfeEC6IMsWzfNqqs74A2E0Mz/orD0shGt6Mwer5VjNPjiMThfdr1G
2lw3xdXDmkcyooaLN6BXdGhTLTdlIJLhUB5qwNJ4FLKdOSkfvZlQmsLgVVpoQbcg15+kDszLLjyT
OuzMjk6k/oej8A8pK9uaWqT04EPqg3QdePxEFf0+OeGcPI1rKyNcipuHRmk2mPeUTnp3t20NbCyY
nS6GR5P/omg24r6dreRFWmAWiylXK8Dws+NYyycb2dw/He6usg6P5SJc5GOdI3SRAtJ2tKosLtwv
HEgAmo/QZG8q0qjxcZ6v86ACre+aenL5cTiXI8/rJJ9QcDDbb1+ZFJ+oz5BkG0mwuyL80w3XwEYM
AJpLuSNMvTpKYGQ+Faqn4SWJHZFLR+c4lrdao2aLuHzFMF6I/u/efOS6mRz2EpNEgFw6uraZLEOp
eBitPJJSBz1JKZMXcnqz5VX+9Xd2KYSQbMZv7p86MI2SceDuQfEcfNjQaoPf47AiN9J9AWRoNQ5u
g1IalM8PiK5qLCeLnLMuYo0rAl5Qe5ygOKd4eJSLEHrcS6Z1jMopCFHxiVTftOYQA2VVYXARa7Yv
Jc4wkdF5qDQXDlqSzTUBz+rZMRw8rj+3uEND/GSyPbEKVk4Y0XcRB/Rc0vIkNINcgX+pdWDSudNN
XeYMyKKSDhAVYahtq3dLQ6z01S48lE8If3b2vLVF42qaI3d3hUp5lsTF/obMbdj8SDXe8HXFfXB7
SdeuiGHiUMUREpDjaLvbfl3cR8dNd2NVtL7uYZdn5BRt1VExA+qCyvo6Ju7McdQbQwofY9aPRn/Z
h9iqtlzf0SxomWTRwfN4znkj5EH4ybBP+o/V2111Z7d2AN7Il4H0XxmbXrDEViygpP2cgboNYn0Y
XmLliVW8k6uzkQ35n8KdP5T2PsHH6up3IshsEUSu/Ieica4eVVu8FhKL33YJYqNOdLO8AWKd7Cis
rKdUJMf3dM/UxKULPy3LcW17I5IEKck2ZFpqfjG9DIBQJWwYuBq1pvKo0KE8EKrB8Cvpgqji0S0I
gcRI6/c9h8BNAT0RCUip4rurxrgI72SO3UEyhBwEJSX4vobg6usTrPOOssq3jXt8WdiVrj4az3bT
a2M8WZwsLBa7imYhuOU7L+qmZfqTs2J3jvKkAIl4xUfvBb1G5VFJoJe5R113bF4kPTYM8C/+zQPN
olr7xqe1/egvZ90yMATiAYMnGiTYa3JtZNPhCwbB0EPa2fsSSQRe2H2HC1nuiYXB1dNSIJuihPNt
6XP9GbDvkWJZ9tas2L032qrw4hrJKNnejOKFuFS2eQoRySXJW/637iPvBV7t7cuGiWzaM1bYjdwE
8AD3kqY6YjIO7coRH+r/FX2Zn9riXqMwAZBKfHIYWyPWsAmoKVS4DL65Way1dzsaD1tJiR4ckrX+
cuP2sVllOQy//bjcgNAXexADNhrGiieRzLU6j6btp9juCtaMbgdXk3fdOQLMhrQHNKicj3hIKPPC
D1n7huY/Jrg49PGP8snTrPFZugkQL7kFrXFq8wPKWssFVBpXI9vE5qXZvMaF84QEFtk7dwNBs13o
PA9M7M8b+V7lz5VgMWDUJvDU+dHZFvwXKIPH9f6dP56bxqlQUkTA5wMldEXRAJY39pYtSjqowFTm
BzV1Qr6jjwzk2G/AX+a95NcHaoc1cEKJf6enQ2YeLWueHknC2/lR0zIS40bkZomlsxDGc6s1T7Yx
s67pRcnsJ8WNvXEqpbA3mJGOig9WH3pPDY1IECf++5VsAg1VPMQFfdQKExmvBzfhlw/nh0cY6TGi
ZUsOx5dgZJWT/Nue6tUYs40CV1LUbvyl81WkecNbHi69ludoqzr7AuRhnE2wBY1v+rBeewurfsjg
hFqO/+3nKsv7D/I0qNuxNXIU9Bso0lkP3cuPm2QMeRPvd5/ygSVZdyE0f5NccexdSMaUP9FAA48N
BjV+++sVEpFeAHWCrMj4J0zZBN0dWOjjy47pR5dic0U1DgAoDbe0HUnCP6cqzNcbceqCFNpMOtWw
NHqD9EriqyA0Tsd6UWHppu47XnLHp7lGuadX7J2UnKO3qcfz4vMbwX9LBH5vGmiPfU0PdrKY+LLP
HEfVgtXJHQ5Y0Ne8kJU4B3sFg1BFHz4/ddcztP8XqnDSlpMUoc8FwIlXXdUpmHQRzSPDNIaL2s76
BHG/Dgj+JQckLWGam9dbf3Aiw8uZ/uBGQU9hTDF2djzIhJxxyf/BwlBMUHTUJt668exC9iBNK/wc
s36kvPXJhCZZxsBPv1IZQw0L4n9CfPFG2hsZRWLnlauhUYLyEmbXkQESZ/Qr7c0lRQltwAAjdtDp
+ep6Yuwr7nZ7MStbHRMrnidaVODZClid3tF7kctpWuiiPEIEvBvIGrDztUQwlfFiROXaax26dwIJ
jBJ8chyeDzXtZHrL+262qhTg5+le0AMbI6G4SxV4Bd9uOl7qpFMwDZ9tXlaHzbMSSmzr6lztX5qT
SlMAwyincbwlzwUwgeGfx7GiQQ8zP0mcKXscgLcKO8eufVGTYwQ4SjlMxkeSbTSt14o/kAVDbyZn
tC18teLZ/X99Cgi0PNEf1hVkzIxiI1NakmRt8LI6GLBcIX9dsCpLnbFx/jHyeFdDmV/PedCFV6Qj
wea6IML4K8IlKWmxueXXSOvGAuCUb6005utr5ozxxikcLESKs1+lYqXH8MqY7tObvI0FfYeIcyoW
43Ch33YNitKVHYQDxoMsqAF7REb3/goTLKv2pUnORn32V+L+KTVCcGvNlBIavyjDtjS98AqXeUTk
kc1Fo2eNIm7nBj3sljbYrp9mhZlxLQaZitqkSB++Fg7iqxU0Afh1zXHv0U04UoLlpnDBJx+Ny04k
MNl6HUvG52oLVtE0i2EDMeOU/pt9FRUkv328wYQWCYgAWv93fhX0DNw0011vIADqzpitfpdWEl2K
+GDYIyYzmaa89+Zdc+lY+3duDojPiWfHWnxFKCfXJ9Tx/wNAN44vVRzFScbWlMKuHO3pofMkhNqB
NMkXXa3hmPx8WnB9Rci5HH7uJWpwxHh2Q9UKN2M2CHjkynhhTVozsUMFhHim3rtCYQenW/lj14lH
qW9bH1HbxKQxB88mi6iz00wdTqYhyft29k9uhi6zRhoy9M4OUyhZ5n0qJmDVwenJZPEStQ/LpP3X
rD/2uUdlbDTOORtxhYCERZrgfiblaUOX9GAWlaCISMOrsqDaSXNuK9pUBs/71/Da9SF1JZ1/GYwP
uv3SAEnvlYaQTSEO+jrtdnhBS1bkEBmY+JoSg/6obbHH48faHGcooX87Gi/QbZASLjq1/kc3n/ie
1qcX8hdxPu9A/VXr6U28wa8wmiZBdDdpdTM3rKOSAo6ePkZqNOUKd0gtM5JTZTMz4VanAdGRqz9u
7N+nDG3SOSK4r6yr4QLs4SutRA/gOYhqisUQIMPf+T+lzpLTSb/q1F8VRk3bsyr4Ft/GWf1Rl3/b
K6DYoST3ucXKSCyHkrHCjNWxWCiLqAh3JFUKWs3X+gFvJgdIp1MzltehUDi1dYtJtMpL2KUyw7ox
hbEkZNaR9dOLSqAjO2JSp+wkhAL9dzEQ7xUAJb3cMrsUZ+HL9GXSoruujeXa2d1T3j2elBWm1xfW
NLl7QejE3k7whfoPXgfIEhPHD5bf3iutJgKmSick2fA46YID9FbcLqknp7hf1NgKYX8qdBFGfCRM
ocoJNvriNWNbGiMt06a+vsi3LTTqVElgbWwKaOYwWcCIppRWz+qs2D3F85k+m2jsFv9cMDi5I83H
6LX65/lqNr6VBXnGC8rD68w2YLYml+Zb1Br+B4Q8kWOxmFLRtGK77yVN+KbYq9zvS842KmHT2uFF
G1kBIJaKEuiJ6mOQFv1XjAl0JZkCqG+viiZ8DY7zd8kt2/C4D7Hg/XaApVYmgYjw1bJDFUN7tdny
wqfDBG7rhBCjcRMobHO+UOVP0nJOHfE3ja0Uo+8tZFwyBvkKRnAfaIIUpikirOF3o/ft4g2nuSyv
5A6ClpfbzNpIjt1tjQeqKgdAYmiW4cqgKTfGAPodZYIqft8YJdvVYyQgMqjdb4Qm+LQ+1j4huQw4
bXMxuRZ0AYv5EGArCNlbYPp8xpMVsB9olyn8zgigMN6LLu1RgBWY7ZsbaDt8PJDosNVDQGlyqHW+
d+YPOOQs/khQU6J4MczAZDxGZzo8Gmnlhg6b4OlYTGud/vqIiwAhXjGFCAGa3Ymohqqk6lFMBGOb
bcY9BbK/gDYqhORsaIGZk1I30UzI7uHg4kg6+7G0ICba4FMZwKfuPjI8gkfK3suzRlGyoTUt8Ere
3P4tIpzWmDzfyiUjV1y71L7K8fSG8MSWR9KwByydb2wZIeRI2FYYL09QHy3d+s2GJPqePXQAoCr/
nwUyJx+Fukj7UAu6k0/IlI6fLkCMzlX15ElF5Nfo6bXu0bSzr7A0Q8CLFL3heFEXGJg7ALdtCvV7
hnGo5ruu2l8q15Mq0TgYXNBJKi+UNktdxtciR50jzXIrcOuqnOGkAnfwQDvOsV9qBEUs4n3CNMqL
NTSHMNqNENf1cqun+BKSbhziTshev8LIMHNX8Hw+wNTX7IqUfHoP4M2lb3u3//oH0iSZsjvO+vqS
fhLcVrXCLE03g9L/0Wcyygd3wgi+UjMhKixaihsD78DuzYWlc0Mo6Lplqq82VTF+3XZeJHPnaNCH
p4ekKbFbjNXmEcRq3bbMZk1x1ta9U8CwtaXryhONK1oknn84Wb3PFc5XVJUAqfXQXmmHEn3VXQMr
6DWqXW3gF70XREv8atCvvtCfzfsmG6RR5R1oUlHbR2l7Boht43kQepqcA7YQNQOszyhz4o/A/2eV
V9nrm/DeFX7O2tLkdmsR9WfzeDZEm3pOVmX4S4T13r5CnFlHTix6RyjxBme7rY98diSAJS8SpRop
te4+vk+95EW+F0OqIbdm0Ql58wBbF4e3vmx/Xw9OROVjDvqW9MvOpNE/Itb+ukOj21DiLIxX8KIZ
99mDcBKhGir1hoLsTSwiZ1p0wtk4m3do4hSPwxJnbcm4V4yXA+im1sv18YFLNUBfJA780ecbvXoV
LSakcbGLvn2PAUkkjmi0EkefRL3FEHTn3BueWzyiQ30QIYmPvP54KWkfI8HslOXiDKYYpdhKXVhR
UrLY+j2PrEZk8qvEtd+8+nDWwafBT1ZUB/ILtaqgn+uwM531S0zQ1t6Q8H6FkeY1es3KT9rR8RVL
PkDwnWTbhYVh1IeHa1XvLmX0Qsq1EYgnHwbBXv44+mhcoOlHs0l+Oz0i89rs6UZIq+32uSbt1mxh
DQXicEnWAnsMjW66PxlkKTP095XLmwC1v5QXvw/bqQY/6CaXv7RsZyh0UTBwYIi94Y6AdXYHDy5a
3OUQ/m56mAYXFeDU2t1WSO+ZG04DLXHXLgu9W1w2xhiCoKcxhtaVF7kQlkSFqfF0oyT+XdjOmEyu
CYKkoTuO8P5C10uS8w6/hWAWmGfa5C6KTO6pfgfRbuHqPHKYUNHdgf7m5ZgSZxW76XRctsG49FJr
a8sVz/R/RKzSRclGEmcK4Qi9VJtLNe1x2LkSxImK6XGZ+IKEhIh8iO1N0m4CnOBiUi5nYpuFhGbo
mtf5chFVtoiIXX7oLbpkMfm8KK824RV8t68ieuz0moPMy9rkudPcNIJTLw87Qe/xKQjKNgU+CAHn
TWbMLDWNR+8GJFod5tWTdrTVBjgnclzMYvQnywptSO63xZtza5qBnrAH1vzEBv8CmaTjX6N4c80/
YCzFZpzVxJ4qSNjEWVa4P2dfZ15EYfMB7MX38WmXV9pMKvgwlBPTyE8lVpVmhyAib/Iz9r7Rfw69
4UPjCelLrM557QB7N3f+hWDXm+VmB+xZZnJd0+XjsJUVskw4eSq++LEkEj96ll29Whf0OScwhlrr
FBbOv/osBFtz8lf6w+Y0Z0yBrPRgcU/vQtDTF0NhYMTw/EfITI+z8uzZ8stc9MkkNY1GUwilktCc
5o5kNItPwZ8jdiTcZzT6LHZlum0St0SYv5b8jbe2PjvRG2Ttw93qWOrN5nnFqWalSgJZ+0v6kpo3
uo4nZ3jLIlsMFU3AoLKUYntlaxQv5YfkEjYoFvb29Nh9ONaVsOMGJI9CEQcYcNqPrP0QiRwLjmgP
kZCwjqeOdvvX0b2Tr93qPynS9EzcaMO0k0EGmBwz5zLITukD9Nu88hy72B7p+WrY5E7cKss1kr3U
wTNLeitBjgt9ktppDT2R3kygJKoUxRksMVbo95HQNq8jYJ+tuSlujrRltXfKkHsFcCi8+C2oM6rF
xD1sf4FcYHybi4FJGs6ZLO/Oc2Av5OZW8hbitbAUwoH7ZQdwo029LvBXqrHOB/YPTISpnGk/IVlp
tUKK6m/e6cM18fhVrowbUu6Usiaq8PfsYUIeVhaLQvrhvNkwQpBD1H1JdqpzC6EmGb5zN/1w9Ugq
unmsZ6hU6U4BdHOkpkAkH5govaNW76qLsXxCokquPwFUpyi74jL0MoAfgWiC/wjbD0px5WBsY47J
6cFQihcuuHORHtQBywxnH5xEIkagnmRfIcA+SSOhUlPBOEkP+poUWoDEpIyVmekP2JfTk4MQ7wVu
qhA/UVony9NzwVRRs7mr5R3ih2EQUJ69Y5GcKOviyuORnlT7itHDuWZMhdBKeHwuJnImnC1POgit
6HYE6VP/l4Hh/aJ4DyDEQGxOMg/KLiIcIj6Tavu8XhRmNxzvvC8odlltY30K8zTnDMDXOfeIyu8Q
M2cX8/iLmHjNRNKeByJTwSWApFifWxezNIFUuUtwiIu/zbSubn0ZNyo7uYD/01q6snyd8LjF2wWW
B9Ls4QV3OhLRzrc0WcFyNysTqkUWDm4orL0zjIsGsCjGH52gtMkQrkSLq0vdRpP5smKFjEc8I3pt
0pW6H7F0qFypXAQrNs/lxiu3o+RUZnqb6L+Ox1gS047aqAK5HR42UiCxKGS83Fd3/Poz5nNc+aMu
DwqMdRg/YzSDPKszuRa+8IasEfFq0IsaGjh1nVn2USxoUasC3brTNwI0Xe9pzw3R5zbSAw37KS/p
82Qm6Bpz3xNp6VAsaDGqOajGSvqnpzVWy6rtu7xyTA2poKBgFyT8HYDyyeeMqYe6IAdWxsbq3o18
97m3eBRt4iTDKc1Yb6elCvWWo4rAOp6b8j4Joi2Zr1vkacvFih9iGLk5v3QgWwknTiW+CjIqBwYP
ul2KXPsMywchHsrbyCVMhOMcmwLquNYq+y2c1cLPBiSyqIFL3te6U+ZNXmmi02PFvlXtYNGNXcXR
EhOPUR127So9HbeHIAeh/3yzWemtbShgeLjcx+sAHjc6+3VjV01Jg66EiBhi18oOXRtLUztI9ZWI
xdP3Cq7qvFOG6wRF+/Q6JSJjnamJy5xHBt+o7sXwZCspoAlbUexXjg6kIpCax1isROxQr/i6vqzf
qERGGm3pP4obEUgr+IyMyhCsqFdq0IFxA1zew7j6v6SUt+rAQ+hUuIYQ3wd9P1TRf7KYVyQrTLkr
4RWc7xVppyowGZKs4R8pN2SVTg0O7zg+BUnlN0f0gOVjGQLCJ3vHmb2uEOY7pJ/vjal4UpYQCUii
lK+pFvy3/s3ykdAfSRd+qWp5D9enAss8M2ytw/vt/x+nrQ4rsK+ZBIr5XV1vx1qcarJdHNp78exZ
REIKEPTe0/h7kezQGFF7r46P74kzppGC9VdsCdDaUnz7dJwBFt7H8NnpcBVb+Ccb22pixr3mRUjM
6M3j2cQpIpRWd9JB8h4VgJZ7hi2+duFef7j/HgUSBw1x47vcj9E+xkXZlUgKLmex/6sYGfpWK3v3
Jzq9Ri0QcB1zpQJrbyDI61yQIVUPcfKQcoAQU+kK/Ue6CkjfZsHw03UjNOBbJWSSMjmyHqAFE+Dk
Rz/DgJjpgakWGpnJe6AgYYHkhuOL6/F0UCUzVYpD92PjTu7lXi4a6xdL8T2z+M5+KXz0uANdXaR4
9ujT6lyNlnYDxPk9WX805eTb+Vi3wOO020xwJK9ivyIyuXNTu4FZdPJcjFA+EZPpmxwlAV0DcTF9
mIfAB4Dbmns2Xcsl9PAdMjO888OugPNkMlOpVa6TCRxV9uuZY1UcrVFg2Xov4B/xf1XGi24GaIkt
jlBoe+DzBldhRsONkkecAZUlqDGVWqrqMptjHxhiUv8gwUHcOGGPeNlrXjTijCuhhqEhBBuj3CH0
CXwn0hSIK4JBmRWzGo+i10syq+Nf9H6sxD8H+E/asKKQr/EceO5OwPnC+vdSMcyTsvcXH3KpKSj6
AzxMF9RCRdXIG/TDn9e0TMIW1HI3o9FvQnytQsRUKbZhY0LKEyS/Fxnb75re//Aw4mxC/RjPRszP
Se5hG6KmfAP3l+xPwIsDF8NyS+ubb1xvHwyxQV0ffErsfnse18PU90EYyXgMtDxIWnRtl6VOpHpV
GfQ0r7MQkBhXceVzeygsUSyi5N7bPfJfAUnLQUGdGLdtVYMLN3CmzX71rAx5Tw1ijallG0etlFAS
wppD2dWHMHO8vXfx3F6jq23c27oQt7RM/V/V5nCd7Y/5+QirDlccevUKcXJmztFuTaASsaCBt3H5
xtdtcp23+RWMV7Kh6NTKOCFlELKS+5795CFDJt5+kz8Q1eL9it+ewYlJhtgoazW4Ue5CUZMRqMg6
/ud0+jBKb0J7rOmEuknTDWUmg9FMCXXo+cpirHjahCeudk2CN/HsHl2mYztlHoV2ghLsNeH4kAhW
35j5HLrzYM7x7bYJD4QwFDrv8cjiGgGL+WcHjy5Mo9MJ3/OXd2W+Ln925+T3bBAA5OWXZympQpqY
cCQrgM86INJs6b4p1n39ltN80NkoSIiWPqN9hx4o4JK7HXbqoGz4fUqV9tO0wQPeNFVA2cO8p+0Y
3AiqsBo7YNVCfGRqjz3BoQRDhuu9j2GJ1AgikMs9XdPx4VOjDOYJ2iwngvvLf0JGIkcIBngLnT16
4RElqFTj4mwDNmh1OqFACNETZp5HtKr/Esvqvtj5aKCBd+v8ZZyIDX0oXzq+oJdZp6PntRZv9RQa
B/EppK1tv8WraARmb/prTTIDRpEtoq9+xDgyWn2L3KoCZ9Y6VLmZrNiCGLKNoAD08fhwy0YYRHm7
D03CKx+kMI0tiAtPlb7e52Ql16FXmiKQr5ByB+vfjLA0wuS7LZjjbTaMLJtD8Uvloj6bYJNp+wJJ
XOchwaldoZluHfLZH84MPtooF9h2Xlxs8aP5v8KOu1fT9jX0r2NlVLKsCnZWiDz6GYiV+HtPzEag
S/ISArHmNwwBXGhQtW2XJ2tmixb4k2JWEgII2uQrMlA3vQPsHqRdlnnAKhNS8cbPyE+xKx3qxiQ4
djMzuH3O6mRRsWOccGjVFr8sx5QyRSe45Eyy/++FUUZtsuIj+42Wm1hyqcxgEBizd4P/7o2dE2ea
gJtoyU4Iktu75DyPy8JpPZgUSRn+dtaoAdmNuw+0IxhvWAKED4UA6zFebCbNBh8D0mHaJcatJnF4
s5RqwHNHW45d90HoluO2mbkef0DlkSJI5TvfJOxYmI1UzrDfSfv7XV5pbncp2wPipoomBdOB0uiD
ElWuEMXzZh0ExKXcIzZH1tvwAgOT45KNvLpJ5/l2CisrXoVOOMuKKAmLcPA2WFkHl2CK6dHX1iZC
FPA0lZXi/AMyHrgIM/jk4fyYbvT6QaM7KJdrTFi3b2Brojb86rjM8Z4yt96OV6EfALnTSh5++Wqy
wIyD+5OyZ1rKxuWQQ8GMQT1UuF0D+sXKvx0hUJuKQVDXLffAXlHcrBvLaxHD9MOYUvTRQGNYXQ9A
TmeWoXA9veQg2+vL6UnzrfCLwUt1u5PaudCPzR/SpTrYJnRsd2pH40tbsCCDNhFo3CVRkF8joySx
/TZAg7fgFELbaG6Cv2jj2tzX3yNQDiOvHPOmLBuW+VVa88hzswGCTvgoYtMS1Gu3GO+nfnRLhqKX
+LefDrX3C7pSn+4cD2LFtOaC/OVf/QDF2c8+TZSE2XEFfNIf09kDXrWYLeB8l7V/tO1l1iSEFlvH
NMfJ/TkxBwibTDwgbP3T5U6oJRpPdNGw0SNtH6U1taVBXbwn4Eo+CBHwsLll6cIr/G8z3VebLMKv
gXsGtC/FppDguP8iMfx/eTwGa/8bi/sOR/pTLmGO8JQ8wDD3XuQWHJF/HBToYTdfc88ykb6pLauW
L+lvibtFZ1oGE9YcWPRtyQh439o8WWVoiK9ZtFu0AOjBiUETc6yEsZ51AroBjFOKSNCaAzo2xWlb
PslRtiPhatS2dQtdcN2UIZWSQLzgfcz/C3qRQEmveqA/l7Hgx4PbaOGZCc5ORMl6gP166uN5oZrP
a/VqmL1TpsefbYoU8jRotZ2kwmNgRhGBGfLzcaNdnNU2gBzb55dX/dMBMPhOrApwOVPtx6y60exo
hSTkHge9bgG68y/16+eYw5UBncRcI50nCXX/qSdEQirVEW61AbQ8CswtTwBIDLM5OIMizklIvf/9
3hkkRpsAKLPyKtFSuhgCgitm7G+dRyp5BKSyQa4hlxIq6ynLPinQnFaMAC5cpU6jjEVdZvKa0d7G
Kpbkxiace+RK1rU0+2G4YbQIjNCxlq2vjZFJ9GHgQEb3W0SyD+6/vIPJjNxpQU4Nyvnw3gnpGnoe
H3YioX/X3bzH+81YVdZhLcpCNGmTaFA0mkrFuX8cQarNztMORSsP8x5DA2lcDjAU34OpU1wVp7G+
+pd1w3P5UQeTCFECIoEoR3ZyFh9NUk3jKtE9iGRutTiNTpShRrNE8wgJeRsfn5JyXKfFku237MgV
6HRASQBsi1vMtXg1wy8c/v25ioNLKp1EdSGyYLzu0R0QO4tZZkdXL18A6qgZGZJE0o6zOBYHHC1X
zk+a221wEuiLas5W7a1YEMpKtoY3yrrTf+7TI2sGjGdoiFwet0sldaVbfl//aGG68SI35ETmN93M
i+6Vlhz76vB7mQxhH276Rfzjt9J0CV1MsMpC03cokq9pYdFB037NQ1JuIIlzu6iNx2psQCdEpYcs
xlOduhp4+euwSLKd86U/H6uo5RUUHno58Xx5OaLa9SJgsJ0BA1st/nnoQpIFcN/feUjZ6Z/RfOwk
MLk8ZEbLnc08XLXVeeoOuJgCbRyH1RQHrM4Q75QeedETXRtaTUZjPgWcyjt0cA8Ua0ihmm9b5/S5
Umboo5WCdg/Xvhp2qzlVHy5OUjBfoxaowDAY9Swnb4r6Zt0vXodSJayLgoEFfjDDmHT3doCWtULy
16jvY1c4MOlm834HzcSumWNNNwXElSAm1UCHoZOCz4F4PH9cpto3B8vfEfqgt0twOQc5IMGpD44t
bDrJLjJiAhYOlUhItbQcmDkSDqzQJ/tdO92gBeibNeopLO2MktLmb5DKfDb/dKWKjQ+0yCX1rxIK
pV4LenPIJzf5aVY+YMpfUg84vTcO2iguXnLuzSUhCKERMsIg57L7pYbMetNyey3iSddGpeiEacMX
We8V9t1XVsEqwfy+TNwxCkJ2G9ulppIE4YyS0vpZmke0VpaFHtLBA+6DVFMXUd6HrnAo6UfGHGDb
h5nqFOE7yhGtBvYJS05yjBC5wp18C5DfTXMbgKwAlvaDku61dZUQNDvhHBWWERFDS+9gwgZTFrnV
T5+97zrG+msuVqzMyN8vyQeSe3p0no+4BC8iMXNdFG6vPuA9wbtys1k51MyEsUNhDOvED23MD3fF
6acjX4zfQwQ65M40CnGKmw+ono1F0GtsIc3bCIVXVhWHHEchzod9zXK/EleD4gEgckqFLHP0vrjB
Y6XiELCTT+C4u/5qMQZ01NWSso0BFz76T61nTNxTCIbQjcHLvdcZuLyhx7w5izr7Hqr8LPAfaA6r
cN+qRkom/SwK4TP61zgfC1/11Aa58QSz5ky6AJ2oYM/kxdu6eTsU6eZfYlzopXHOhtZGlj8zPWEM
YyeL2ljd1SxACKreFjP35LhI/ilup3510mSUMfQzXuvEhpwxfDrukb0tZDkG5VM0ask0qXhmQ/rC
YlAqAI8DxMl0oNIY9GCeKFq2p6fNxQVnYA3nwB4kW5dhKooKCz0GBeErPV3YXc1tXXtaQ/SU/nnU
Mc+/TMPxiD6XmN++neJdVo+Zexqg7kqm82Djcg9lPEFWzp3uqcDjDAD/OqaO5Oxeu4IowuzK+kNt
IocZ12rRpXwYsHLeLgDKKYsdX55s+VDk+dhERAllXsX7pOX2LsHcRvZcbgCPSfszMpy6uRAFW1+H
E+DNGOtXeIl/siaAmJqaPgKxRo7PHDCcXLKuFEqkG8pAKCNLh/5jaeIV9yLBZHtBS6Y5Iy0c085u
1dhu2Al8B20HksDudlQrANfHwgNs+Z22v8Gt+gaHzBXX2vScuap54IVX/91Z3SBQyvBKFH/l5rrD
dnRLPXGcN9um5uMX7pDwu6NTDfDkcYlPb+milQXd6oNpm2pWtJzO4atZQ1Re9fDuKhfYkVwR0Nu/
GdJu671bBOoePbaebxPBo2ApZrnMAI87Df+C56PzXJOJ1qP79n1UJWVlF3IU7i90Zc2S8aR4DSk0
jWk+y4ysWtMSu+DXL+EyphDtBOI3U45Er579WP0lHB6Lp31p/mP4wgizEkNhuq/vr+whFdbqTBut
dMtrYxZ4hoEF9XxFVfUWnW41f/jUFEg41spmZJTA4+zttPoz4Tziovsb2B77Bru/p8UFqyi+e/ye
l0r+KCGr9vNxbxpytdOJnL1sGNxnJsq81GXVem7uC8wCOgRTzg1CRNmXbc7RsX1AIhB9UzqdEseN
b4QNtG7Pi/uTk+XY9S1tJ0NM7J8AsiP5cJT5TQs/5ak8GBfv6n23IDuT7h57HcE2o7OzXbpGT9CZ
dKo1EL67lwExWNY5TqHgl/LageUrj+qCuZd8/tRnN5dhuRaiD14f4BgloJIxazbLyLr4lHh1W5bT
4ur0G847vQDkfOhw63w2Q+jdIQTttYg8LEMTANRzh4Qod8BqylEysSyS7LDZpbcXBF/Fs8wExrJ0
GCLlFPmYK+r0G45TWMVZqdEB4TcbPdVLAml7qo+DialyCnzGKTQvcqMS/EanLu2g0DkmWawwSZGF
WIjbyTZMdjRMNfHuVoYgJCB58aaHA9w14EN2ntRdyDaLR/0p9+LclzYdqvRM3Cd+ZtHQIBJ9/wyo
kfV/TRcn6kJaMXip+Wc5/wDYYjFS5/yYWI0sCsmxW9ljgBhiEDTELPdBoVF2K5/deOTcmFW5fqK6
QdurmPusJ6iW0LqvmIAHTs5x1+vyNv0iKyBYv11j2CLE+WzdNnMlIT5qsp2FYLbZMDuCnNdBtFeW
AJcmu2GrdbHkLx8vfV9v+DOv9ALbJWDafSXi/lWujwSS1L4JHlaz+wDLlo+zrO0r8kt0gfBHjL5G
kjggSYRMXHDo8yBeoNmLD4jolwvO4DHfDsFnL+C4TLqQpN5VTWnUmggJ/M69qDp/fHGniqRxuZYp
6PGs2Rx8EKoueRowIjX0+CRxFoe8w1GeTFHBFN/yOGnB58KYnrTRJXWvSglPTcmBjbfB6b+et11/
8PKJILhUxewjVToyJq8av54slS2XVwJeJRLFjOI/aAJLWoc93ibfYEofTo1mCC4tYYl/Q3FvkKBh
uXpduT9i9KpnLgZGQC7AoPKAGNqBYTRn0XXGi6jUfG1sUt3MkS2+GKPUWr7eZK45YdGDwLTdhdKk
zcwLDEvnPgAZ3ABAvIPCyjhA+dKtmVoYF8dgZpzSTiHEDyDMWVPpZSDiwQpC0ON+ktFyVqb5Bef/
oA/nzlw/UbrUnc7YyPpjIp2Nx9QyZ5dxjyxoQCER4Wuzdpm7iEu+BKSrIn56zmhFqiEpZAih7wS8
MqgJfHZCrNa/5/kmh2S5vuOU8CbExoeDLISIRnfSLrStW9PRx1zUcpgFU4OC2HK1EOlB7cTVnpuk
GlNGKuxdpGCzRxfE35Dp/JyxzU+fwnOPIJgjlTI/8OiQIHtsXTR57SwASkOrUfe/SOIBrj3WQjWM
0kzw5hoTB8+5SQByXOFVYvP/9xSzudr5pJ4WbVlXV8rMHh4Uj3pqcO0fytV1+Jt+k8CywxBehfum
d9527ni90FljgyVf9RF2bTVZzlZCLRPAYrUA37C0moKvJF8wCHZ+rc8cPf7jznbg0RR2Khtl+eCN
0Vv54TcfKwyMdnjl+YYmjfNIsdMgQ1VdUKhtemjX4twHUSbSxepXAN51AdKB1f0Obo8io180eT1/
fEugty7pkDFL5sOR9MJUZG995kYe7JV4abZqeQfVLDLytNKsW4H83hwLZrkPlMbaKPkQpW2vwzFp
DRFuMhNoSZ0acZ3fFvYwmfM/vZdIUQNUcereKWq5o1fgxPr5+Iqq8w5WDKHAq5tDJl+2vO4/m4wV
CNLm+oF9OuuCktdsAOJhlQ2d1IOYzlZWZPHUjsQud8259/V8iyeMUNR/p9wxMAEqTvUvbNMApbeC
qzp1KKFSmBSooHbvv3lEhKevwZ/vOSzT8UTn8L2we+mAeRsAi0XosqpJekLj+HPmj1V47CJL7s+4
2DCRnnLhC6UKK6YD2cTwm6nSrVB0rgaH9NBcni8HaLcglDJq9bvJmshO6fU7Gwj3fTRohBPDQbq0
T5kEMS/HZevRhf//WFzUVceYvXvp/o7KRaSFvw5DzvsxEJIl2Y35Tnqen1f8og/auXOHWux53RPr
LjxSbgb42/ScfZBW7Nd10Y3ilmqNOGpael/eFSYtcPnz0jyPerdGVUp8i3BRgzisQyy96V3r91tA
agtMBY7oiypby+qZUQ9SNPdg7kQJ/e3GqUnhf123lYl/9jA2JhxEOJJZvrA2dUz/7PaG037zZAFC
WEJs7GCPtcCUimM27LICQv1VuTKQPE6DYpYx6caX7oKd8khh4Nu340EO8tL2lPtbP8cp60pnGyai
4BzzS4Niv1Cc6EQPYR3XwbPYFv9VpDnSTbc79nUGst3oObQe8pDmJEn1dgzcVdzO2G01L0GUWis1
WFIkYvGIrhANN8mhkIS8oLtRefSgPrM0IWt6vDi2iDkpL/C7T4wKlM++2BliYljf0uVM5CqP7R+C
8cf5t1l6/0uZPtlcyJuGEDfmgSMObaOozwGamK4fiotdqAnsRydc2hATd4laIcTTxxjhMZIPcM+f
Hwre7p3DOB5BVXBIem/iYeyn0C1HIKMl0TJveWsKy3mPcBIohULMBKW8+X6PPyFFNj0TcnGRXQ4k
6oFqT9WTuXe0MplRNC5or1yyQnOtzWT5uRdOIv1tS/j6dQH5sA0PyOk++uAyqINQ5HECY+1bvyii
vuLckho2Xe9ZK9b0zuVFRZUHtMF+X65ioMFYpxqG2XBlfM90NMD2VE+MXr0YY5GNEMFeJGrQT5ft
37hL5ywvFWFgzfvnD1dosc7sPvXKHi6tvUuIc45zskiexSGbpVT/JCeDt+FkG7E7ajr0pxo2vSls
/j6gW31pzAm/eAoKII2ETYvfIEkNF3pyilRsbElHEviOOFIOxozrwJ4RSo6KR3LBaiuopgGy77IX
wlMn8TT2/wHcKV1wGq+QxxeRhVMhPK3092WixVBZn0yyDecS6F93XMwqXfSSyLNwxvMY9W8dK1nT
vqh6qWUB5bJlHEurf5/SFEQKkEQ09dybV6tF9tkK0m6Xv7ahBmczzMPRfPonyT6/TV671YhSWWzQ
Ks/ioE776eD4WWWdiHDGcSn/SQPT3SjQyrVnnIayRgAeFjXE5ANZWzLOHnWAma/RkoXMgpeYxlrp
NTRw9fBvT72QofM5vTqKzKmvulrR7a1x89dx6JP4OyDm+UyqTV0FfHpHaTwGGZOPfA/e9M+jPe3d
O7mnXr62UfvdOuW5t8vm3Xuvqz0kGdHwsho1odr/OjxJPIT+Mn5hHXJooRIWgJahfWpj+b57/Qpf
avEScwRPr2Mw6p9smSZMWPOKcTr88heYeiOM4N0RfVz3Ev5rIFaeiS7g1PiMUKBPsSbWjy+rvE9u
lkudjwxbB6Dp+qWfo642aRk6UyzkSrP3OTxHY3CQzENfbV+GnZKKSu3ZGVZ/YIfmD+zaWJZfL+E2
Jq3PgofxeVzDXTOGlwzmXjiMza4Pw8vr39O68GGBufhOer0P/UArjT2xw+eNfWPSNT4oT8ccv6xH
7JA+ffMy35W7IY2i9VBVtB3LN71GKKr1WjAD7RBhwXH4D+FJAWJhBzOE/jLVFq2+GnnC4XrBCOkn
tTt6GtT5oaoim26msa5B3kuwM7Lyg9WNpm1DzS1fMZvVumtSrkV2egByNjjbHt/uxQ64v4HghfKc
izToqQiO5tZDMh0zc5slcqpkPSdA9/C2YrGhmpz9BVyu1eyQLkx7wkxcKW95QI9MW4liJ4hyDMDX
WooIUjm/Kk5179d+9e7huyDw59OUV14zWT2fFy3kSQvhYCXK5zrhcWuOTxarF4cnZCYbTs99uDRB
7CsE04OhZ1rErxV+st7hngLqbx9xz72Q2Gj+6zRZ4ES19FxYFfBN8/dtAAuYIvH5CWwVmQeQRYyF
7udlyxi6rmGABjanZSI3FFBXDDkkkMuN1GbHaQkMY9iUOsoSnDIbNuLIL+kIzjGMQjjn1b1VuhzC
Ok/sBDOccVRgOEkWOJ8nEXkbh1tfT5/N6ZWUhUjJu4ZSMRYCWE5cQGWCeBy/HrmUhkVu2mJokcek
vK9tFALqYDwPBfs9wDv8EC9HsZHCocJoCPUIzqOHvqiZ2O+d2ivsWVNm5SnYPfSDu1Z2IUHB2NJu
LqRC4UOLoDv8y7bTdybuw11Vet452HkWjWBO9hM3V2y1qrboz90vgMHMXSYMTIwxgo7cYyRGewMC
2Xqq324YfhrnAuCc6AD1EWLznOiFIsbu2AgxVICFIxUOkYejFu+bx6l9FeM/M4yAgfAazNCwJqjn
2frlag33rgkwCOzANBbYONkKaMtNq7HltbMMxEqfwCQ3FlOon5P3LLEnV0FFpaKcdjcQZ7ZqWKwf
GIVArdpvlR0aaK+OMq0a5Zxr1PdkS8pT8fhzZ67loDBnFnVUsIiWDIe0lVrKQvaO77RrEMa1rgOt
bG8MuLQXCw8ESIuVl4g6EZTFiJK1nki511Iu2zhkz/HbMIecgm2mun6ykvY0UkMSLa1ArWllXpod
pCGBJqqkG2B4MhaVYeEhd4x62oMKjaX7zKD4tvWgLFF4VDq4IlJu9BZrYQTnRWtpHMq/m9w2fymZ
lZOrPDL6DRtewSwnoi6J0DTCaFIMD6OKiRWWtfZzQSbpc8DiAs+9Ry5rPswJqYOFyOKwDCw44qNN
8ABZQbInAGNlRMGJ0obu2C6A4sVnYys8B+uFShLNcNCCNaChOTHvFq0zHbIFob7ub12JQRll8OjL
ldF/Cya0wrdfpPIu31qKp6MYhU4nQUZ/Jsbq5hUJmQZbDA0NTSnnlpa7oK1vRGxoztyDxKpUfoNs
oQ8mmdqdA0lp9FZ2OLmHBL+V9NV3DzqrwDtWHcvY0NutE8t2XhbNaqtrlNiOY4Ezo7YTZaGPYDUY
sluyfbppMQLXBBguKduLMl6uR6YsiDDyLPgl6HIpNqOf7Peox9hIVpVLO4SOrjmWRLziTZTJb5gG
xm+2ZGduPpPEPcRZkX/FRqPTcrAkM1hmzMdOIub8Yvbpvg2GMULo34hECEYjC8FzLJnZj2bxz98k
50kTfzY1FTKPMCZre62iCNSdeYEw2PZsdZjX8nhhMAfb1m2th1GQKgAysxQiu5Wt93h6L3t9nm12
D5q9h9yef1FVWmUetf+z7kznCEPEAsd1EtzMqqDyGeeLFaV05tNTbVpFtgFJ2p93yCLhpl0Zy6vO
hfgVDgQfXsKlHfa2kqiwlXtDJNsh5Z8IdyQo9Tqq5xlYGJbjJZgnrOFLH+mMJ6Ec6/TU6CWNTwj6
L5MQoexrfRLAK+djugisMAK3vvxkDGwHKUSLBPNlOeMZIBy7UuVMh4D1K7r7wSwpdXngIoW9ErVp
eCyNkuhhbbLSwh5MQ1Y3opJ8EqWP7HVVegfcCEAzVS2i9aTpiH5y2jbF0ZIY57eM7U7zete4e51d
nsJwXTQVTXLJOHZfU8xdQD43O3oioJN84R0mkmlH+WZuJ1gmL/OU/MJW/jtRfnXx3OcD939ijnH1
kGoTkoo5MDiEC5XJLZ28n7DD0SzMK8VE6fVGEf1CwzzXpUtvxhUDAlFhmaHPX2wcakfI02BQIeSq
dUx/5M20lug4ChtKNZy3KuvlHhtbc2hgmQm0rurD1D8x0muIViK2Fy7/zxYSan0YNd6ceJN9xMIc
W2Ikd0aPTszV61Rkh2Ulc7/E0YHgj93WzJ7mZIlbcbZd+5WtL5yWWlMvl/W1hPX+k/gFGyc5h7Lp
n7clNThmEkrQwX225ypT37fmIZbxfWeQjV/8Pzrn9mIQktBq/t1NvCJBWuYuAQ2VWu+C5Uq4EFNL
R6M/78nHMg9JuArpbnxbgVvd8fyLCSjWT1H3Sg0gdmoSTT6Kn8mwTVVRk2pIwszzSbNB4HFMCxQ9
p+cENST20AlDKIxs8OVRwZMHoyCAE0K787wOeT+7YkCoD9tiTLqQZ0WtUfL1HhGwjAlZ6dXP3xpa
xcVImrlO4XKa0YOCgYOvdcvhc2KT9mZTLUpk3kGzqV/XiskdvQBOjnhGJlE66R2UxY++yZBj54Lq
uG3W7hH+PpwQFNGB7sXTkBrkVHKYe6n2+Actnvtt89+gbStJATASZhyzBvseW216M28CY5lDAnLp
RhXZPF3JSwIn/vdn0MAu6+Tz/VU+KOw3Z/GPiFh9E8k/wb7h5O0xRueU7D8BgbqtqSoYwB6GCM0/
NJ1KyIfazkxZGfXN+y8E93IoPM3uCWk6ClcXtuRwwY7x8abGs2gmTbysMChFYYZHo3hNYfulFvCf
qm+iRA2ovfPAFAFsHsqVTmNRHxzV2msThmO3MkZrccbuxK+B3jWpbNp5jYaKBPqVVGad37IOQ6UR
w+tdq89paKizLkY6qhNDVKfcaWom4VfFnm9W3Jf5ayxG1i8DdU7IdbpEaUbYrign9xorVJz8D/9S
n8DK3rUGhBfVsht3WXkspukLwnNdFwSfGE766T+M+pbF+pp9IP9KzLN3HEgslh5LEM/ZKKoIFtyg
gwvLHPQAtnHItWxoctWDCurjNfaF/5AxmaQdB7sclaqZ+N4DKZJgG26K3YoFWIlREcvtPgGvLhTF
Hy5ewicP+hVm8ChtEV7Hpf/jkFSYHlahloFj0nHBo7nKlljFsGmHSMKYfPGuTRQFHr4BlwNpAj4Z
/0IHH4ISCVour/bSJtQTmWv74tfMyrxtKfbPW6uwWTSgK6UL4o0zb8M0+f1AY/RC4g4/Pso6vR49
EDbJ7jK8ZQTefGIQUqFFiua0k+yH8iyZPAUjX+w7yGKLFSP6yEZDLJ5XRwPTDa8vNhhj0RCwEuKI
UlN6v87xasFHvageCRLPRN3cQMkik4fya3JZ/tB2MHNbYF6YYPbRyXiky3TE8nCKe5B7cCFSAjIy
kzG6k54rrf7PLAUCOFNvMOjnHlmzgj+gm//q/AvvJoEtOSVmxJJwZypsMehGRu9yqLaEXcL1+oC5
GsYRXvGnP2f1tB18bVem+D6bMG+RIcUTTaATbWJkRwQPbLSF1AORIXvpekrlJrZI11khNHDvsr0m
vxd4oaEbXwd8zxlQdTgXw6J82ZrF4fInGgBUsEDmKnTdoIXmKpTbdeBQnC5JLbJuxzzleZc4mCcz
nU5H6+xgOpkRqWqhCNxQoHJsjevhh7aEcIaa+T6TErjnZ9M4p0KCr7N3SAivCyHF7mfX3l66ZCmT
PV4nwmuN0dRguXAa3qspfWX1gJbav2oedwRSWgBjDt2Ou+2flmzWHBEE3a8rVpsNlABAyCyXFXk6
IWG0UPr5qEiggp+IDQS/LDfmW7/xFV42y8gQQuqzORdSjxjQwrR7eygmIBfvFDus5jdNwwoPUyC7
OGGMZs4bIfTS+GOuAKbIrFhboyTkyXUAu8baBedeZ6gwBiaKLZlfQanrkX0TLB0myK/DXONGsQN4
imB3qr6hM1WbETMnuSo4r7s0FL3Ato67GcT0Ud4oLKtfMmPKc/kay8JoFoRIA+4ca8HycZfghDFR
wISfaDiTEzqDvoOUc8I/GTca4S7SkKZtN0K5/4aWz4P/U1a3ogAiaml9QISJisUzeYRYeSXMg1qk
nG4+FyObkTN2joXP5WkPSrL85uDSKbd1GwObRlbI97Maoj6/MRPGeHKXnDlCxllBk91X0fFBgwez
IjiXkLH4bZ2by+57iIc+iTRZQbYuKLIWibeQmGxYxXQVZtk9SSCur5tBAMA72jsSAtsILBSr6uyT
0tSZ+k2lVTeZEDG5loTYePQB0tDTJy3SX3TZcI6EaIvQDQh22eMbzbuY41kZBeT7QpHlmFOrmLQ7
6l8Etp2ViFXlm3NHtH8nbAR+YhB+cQ9/6aDQtLUriRa5qdEtiJ0a6yUi0Kk0Q8icaIcpGcdgM7Gu
kgcKpPHrtM8zDQTFbB+3D+TVnVHjoemN+qmJay+4d18DS/ohFp/fzsYgCDc+zWrTqwAbrpn6ZdSW
iAzTP5bfam6RdYBZODv366n/W0/sYV6niFSK6PA9v40UH2xUrEzvZWqQhkGYbwneaCZRQs5NNrqD
vCHZa6JRP9rd/RyPGpVQrJYSKdD0K1wAygfiycUKd4FYngr0rbiihR8g2a26UR/gqVB4/txS0ZQ4
/zTIn1AOlPEhfXwYuJgCHqFAwGOVUQ5ioSUzCprNboh9/EBu3jnTEAyiZuwhBXMjSXDT/R7+lO6b
mvHEjKQjDZTApipaMnQU6sBEDKXsMfTzlt6QjMDSUe98+2jGNx0kPn0U15tkmhw9eRIyGHyNzRCD
J5QQfySUShy16CPDFsMEiC4CoFeWuPf5n68I7GjznIrezfvwd3Y28jBgJD8jEo3yNBkm/2a8QRMO
M+6Sjf82FI8e8blb5DUg0IMv3zjPxea+KjcnwophxcXWuiwm2tXB9sQUvPeq7jOBOBUNbn+htlgi
Ode9PaobWEnStspsZLSvYEsO1rZE427uniHL70Y1P2ORyjfrLZFZWqMWiDm5Ha4HmES2ud6FDqxa
JVlMjvXdQSKpkAZVAAg+uugCXpqQjx5M/UWYRSTiq8PqYDyJ4ymH8ho9NVIqAqkOto5vyCTy8DvT
VD4bsNSakYa8BRKl2/qENQYlCqwnV8Z5KS4UNLnQCJorjXwovucGPbnWzSDuP77OvHfArUuUfB/o
h8b2tQkNRYPMWC5GrWELDA2rfEyfBMlXfjx9hklCL2mqcAWZ2gRhuTF22i3JsjLPuAgJ39QpY6NX
sRthgC1xNLqoRsXJzp3EmRhdY13rTSJTeBatNUChglQOxZ/oNAiWtQBtuOhKYZHzgz6q1lry9v5q
7leDwr8AY16D8IAfFYHpdfyVJIkg65oSckUyP7BFm2Lnsj4JZ/tjYttvjJwlgdiclQvT/TGsjAVB
mBzmu3gOD1xrS5JdUksu5J4ObUdtrW8BbMPOFRQk+IR2Eh59MXUAvoGYAZW+ER5bfF4/DZ1iLJVT
K5Tiv6bmjm94VXs32RXTZOcFErfOKTka6O+Z+7brNSW14Kt1QjD8hjspkCdrkbXUuGxToOdAfDji
VzlJZn+oiTSddUOCek1rmI+ZIS2GP6H49iGO8x9r4mHDxrqt05Z+E3vj99H3MXSj9efBmO2mZYBS
ZfAyoJhUWILAlPG+N1gzg0ohLhnwyv77yrlv8lBeEVvbLwKXieCwINjEg0LuqpjUhhUwLwarCZqO
VG9iBMjXflC+wOCPQrdP5tyFqXDoW+wRl9BU8V4ZjdxtjnTdB1RBFjs2RNag4CGXfmchLD0k94k0
47wvHTad8y7AoHQSysYTlUmTt7iBGSsLlHniMNZylnKDZwkyiSwE1kfOVKC/g9efR27aWqq2QkXp
DB0w8VmfH1db1J0hLd3Zr7tScjoDUTyn+fsugyvt7+vE73sQOMpGAPVAnOY7rz8kdhTZDqkRm424
SKK5xo8cVIWeMNP8gaUI00Tdt7pVp0g+7zXWbq2DaRiNj3Elct8a/5JNoRZheYNSeMvUwr8f6A6j
Uk1nJlFA8Okt/Ww6nyJL8WCdWWCCDqSPYiSFS+pAO1Erk7srFPbWolbc6B/9eFCMBfPv+TvQJOku
4Auhxh0dF8HFakuWfTNJNGpwSjmhpIW9f8NkbRo+mCFPu4V9TpTa4YMkvAo9nv4sKbToN42X2R+i
skTCIOj45nfMsG3SkzgWCS7/E+jgf4ZAPEOBKqFoQpDKxA9RUsnsS3ntGzdPlPgw0F8kIsxaPjwd
wvXIZ4uprjuR7WZX5JB3sb4EFI14bEpm6uSzKUoghMLT5esURTc4lZ0Tekhrm+xX9ka6uRvBmKS0
gB4gVteJwCsqEooafdV2Bni6HMDRWj2IgXgQYC8gmbt13/20viM9qr8S0yjzHfp4RqDeWq1DC+wa
yl1GtN/XhMOdLVwtIYmlS0bwKC6XnZFHXijPOA9YD4l7JDd93khZBDmtiRErv30zuPrE6J1g4Vsy
vNnjFsRp7LY3GiYw8jZFNxk+nCsXEoIqDNEpx3GFpzeY//kyYRvIf4fo9hm0MMxjYQtwOTd93dRu
N2mRiu+eaEfBuJM+O4Up3wF9QcNtu7b+o8htsZszxBHe7tIWqeK7wTBzySpbgFd7sRmRpQI1iLFq
xZr6kebZW1CBPlWd6wZLF5EpzgjBOIZuKvZANT5Yt6DW2NQ43o193Iuvs4UQg7kmI59c6YfEPGjz
kH7MBd4zrKmDP9SHNvFJfE95pNji0nMrUEGFmSnUXBIOwgBL2r03aoqx9b1P6MVH0UXI7l6Hkhcg
0Gb9xwkDrlFY7ScMk3yGT4qMPVxmnOxsVglaN+Ha79qw6dEBorZIaXRayknIOObi0UTwVFx7M98f
X89dz4LkHSAn0JEvuX5rPsHZ9dMEbwgytFOTueG7I85KqXinwERPvmLFgtr409YdiqnwDTn6+BmE
jXPYoNTQ0ryO4rPeFT54qAh7a6Y3zdSm5xORb2wrMvRaxo3NIZJU6aG/dF6Cn/DMyaFJU+E1MngC
Vu5cfFKdD1WzQGniDXMuXf5wtI1rO0vMjBivlOv5XT41L8QSyJeEJpqwpzXmdB6BPa6c58JxUc0T
/rmWEQpavZVEtes6SW0ExUbnyvrQOCQOLMuhpFU4J37FZT00478Ir7mr7E3W6pBcG9hlnQpE2RCw
Iny1GXu6G0JGiVXWj9tbCAcVZbPonR53L9ptuANI8eLtysIFZmxgTALByYhUVfGjRCyOHbxaTWrQ
gTN8KPy+WqtOVu/UKOP57PiKGTVZmUmgcbTnVMVTttTeooJFkWyfTAauUyHfXl4FAueDK2Xjxj+A
8MhkOQE4pyy7BclL0sCXAVHGrzGP39D/TXnqrfumpeISwB69xLmW+7VH2WSYeGbWYLrhPSTm8PQs
xUaAzRVRljKzYBZ+TUmukiZ+o/WCOJ1LIVj6sp1EmzEHg0rBpL9fY90JtkCySNJUCyvAuOSGdw6E
51EqvIv580Atm2zIShaNHsXlhcSKFFepThXcLuew+RUdBEXVbsAbHOy51mt+FK+waeAcKt8TJoGo
ht3cm9CVhO28OLprmIBMStjPVQDUyBdv0TyK24XXWHaFb9G0L91KePM/PXgZXxRPPlkOjpzut7UK
v7tU8lW7GwUHtOrtvbbhzAfizFLpDf2CO1tgLIWTTtX+iWU9sKolp1gyb8eXdyHPjOuk2uLzuEaj
B6ngtVgCVQtWChrOvAgSksQSbWdH/q9JrourZuBdGIbmNvqVNqTdM8fdH3CTlWmxh59Qp6hdC9Q2
yCUGhQIU6GiAEE4Hk4F3TMtHwX1ERPU50v9qbPWC2A9tleE5F3I6Z+3lLjzMstqUJpu6SiuhCuoB
5oNt1YpVRtCLXYZwpXMOoOTZYpC8hXMH4ophKli9jm3pGnUA4rM0C5cE9WPWCgAPIFQD3HdalUik
eQxJqakPSoJMJ1JppakHEm2sYMSfjC1tkgm6w+qnc5u4KIodoRhKjaQQsI7b2qfztPCu6mdJ1sqH
OtaHo6wWeaCIaNtxBky696ndmPPaIZoQaopAT5jHf0UizrzrsOPnc2noVSXxzxP+JbzoVem2OAlJ
Peqz74yW85jS5oL0+qb0+FfQ9f19fmWxM9rK/B9E1eVAYmAmorMP5KdOzbks8WzCDaX3koXVa/Hn
/cYG2OOWmvIa9hC0CyHibXDC2q1TiEQmmTt0a6/Z0vPSKs3rMpbzqccbLHL3zjYUNzArUslo6x1D
qALvPhqu2ApuzkthtLltiRgJHzeCSj4NdegQ6RP2J+Dd2ExDom7N41QeGLCEtJwHjeFjfGuVQh9K
1gIZC/TMIunCoKkjV54zx585ihXSE3zzLYMBgXBvXfnDOmXXHOnvHQTlQ1Q43I8LQoGvlkPdYPqG
yMy0fDZMd9saG+sNHFJci4FAF4LmV9cCKDOuS8SZa2yquZjo1ZAPgq4OWKqf/1Mz0Mo0uHx1EMOH
s8Cf+biOCwh601Y+tTNbNDE2/i2VKxOlEiPtmjZgNYz2P13FdS28/trLj8QDQko4dxErPzlEHosx
yQ8ZmCsP9bsPrnyDHrmhwl0UCLe+Wvkbs3W1UorWll91FmcIBaBH/un1Fpfsf3gpXSs7y76oCPlM
9vM5Eb784vMgIm+dRTQI13yq28FjD9dei1XArk1R2bLcgKiID4snK7sK4vyKEYKh/Ch+ryN80Lxw
UyWs0CTOc3GpPrb+fzOMwkB6+/ZXI2f1iIRfJ+iLa+M6pC5WKwv+7Jf+4Fz8DlOc1V2jiPkNueU9
K2i0tvWPv6DPPZEvdoqkB5R/WxEvjovIVEB5JKCY6CG5Dlg7fAw0YGKEixXRdHtT55Yzmch37Ugy
C+WXEeqJKsASYzPmljwiQlokboeT8Gy0yTjxR03JwNBSCCP7G920hoftoOyS6vQEwJ1njYKQBJCc
dD1gjoYg5dCmz3NsygGGRjnfBqdJmmTUiii0wE9P7b04CuGCsgyB1aamYyodiXy/2l5pKSxO6CN0
d/MvG4DX7esIpm/9kA+MOdMqRsDjrBt/lS+0w7Rnb5EOe6iUR2qt3YWCtO4DsAlb6s8dv8ryA4f6
jQ7yNXd7DicXrQbwJjG7jFXAhWz5hU+rtfutI+BgLuzc4n+ncbetPBuzBbbnd9SsGB+AuH/ypbjE
8YniDOyvJNHRZFXJWOWU2UhuW0EXGNg3ygDbLPYEgA+yvECIHf/YGV8yo/SNmAqWbu+bwgEhgaNF
NIxUs/fba0JWR/cNVt58a9rQBdinpYglst+ar/+FOzRzkkWJT5bQbjpZ+eQiRbsDEKFYrUJrB9lb
QdFtBktqVxPn5OvZSOTqPmNsInwbY7luKcrRpIBAOB700e7eHZpX0sMi8QcHDCUTMTNiXV3HsY/7
sWx+nKS0n7Pj+RC9kuUd+/57P8RWoJnNQvxTRkP/oKpzlnFmo4OjkK9odUfnOr5EgnV7SuHzPG5G
YHKHUI/6MATR8t8SAtu9YFxSHT3kHshMK7q7FA2aa+uZYysDMyNW2AAX0sM6iKiM4SHrTAZamnh3
6J35PIfMyNLaMDinH6dGoz+b7Hwbqwxzids4yR6z3i7bXJ/a4mrV6dK10v6eDNmHYhptt6m4fNta
Lu8OqvOdYh8suRKVBlJnYm+jGcrQzozVDfGMZQrxrPYB4u4+OwbUB9BneYzllDZ6jkX3hfGRSMQG
5qOXNf9hlAF3Yhsszq5bHEyFyZ6z6tdIU5k+VrgLNPmJn48M3+Cm+RR9AycwbEQP5ZneAoGwS0Fq
V4/hs7hAmEAZjNsYvW3z75cDm9Y86N14lDKN3XvQzkaOLAeI6NZtsGLGXfYBCUKW+eB7HlovC8kZ
QY7BkSVeALRl40MboQtddFn4bRKwVMhuITVuOpewTuVX5u/oiqzfqERIC298kVmPXLWIH7pT7wIt
tRMeYCWtu8QgY45wtru0PRgEZPYmeQiWRfVZzxjEsbfe1HybUSr5laJpmtduQoX1xM+QDbgs/ovA
bZU55GJfbuKU+d2uv1kyB/F2hLoeCJnub6oWryez7if/TRRYOoSy8A0pggtYQZWeM6simQxmRU7J
hy6xqYwB6MZP/YEkmDU4gqUn1nhpjzYapThupLj6ibAk3pUyu7QjanqsiWem3lfg3k9Xx13F708E
eSK2+J3FQERXkwxaBria/WA4dwTtcDb55tjiDC1X5V7ylW+ULjX0tZ1FbxjP8vFm5nJvzFJoYCed
Dn1tWr/tjsuLhcdSg7Llt0jKCe3D8KQfIvJtV6iGzZK6ODYNzrUpgC2gzCV7U+srWRuxiPkSWtxx
MSCVxASrjek97EluhDQ0L5s0EPfonBpult1ZnnhUX3TpoGa++CuV6e/DdmuWI2pbpVunrHgy/yz7
0lJ9LJWYDk9jZFrB29cyxKSt77OdtEg2yJ9pZIuZju3ZFezHxSEbUZJIRmRWpeztCDNv+kAg2w7U
NJolMCmL27YJTxuJfTTkT/o8yQRXc4ufBlwmrg9q/xr7+CcTFkDWZK+OPp/92yfOog5Gtg6Xw7Ru
qY0+/uOJFe3VTN+Wpv9xH9tLaU/b80zHJDaEyr6ZXE/pKHqwKVTprShUHJw16qLAu5lztngH8N8j
4jp3VRaOlZX64e/R4jUKkfkz3A+3aIoXmM4TcFtg3GnWC0XZ4yJeRo1Zz8ucknnAVJA2920fUlWx
qa3+SDxwXidqNQQlCwBYGaMh/6ZEOg5yiBCyvboG/hUJTgJr78019OgU8TFc/WoKL1rFoErAX0Op
XISepzFy8mkQHlKxUI9mnTADYungTuLRi9Hak87y5Zkog/1kGVYMWJJJrvNisMBWW4WocLDQinGL
sIQcsW3nYfQz0TIgYN4CgpCulI9GZEFozA8bpO1VsXxpm4tP+gZstytiaTSzt49dLXfxnpCVScsz
Sj3bN5VpsEuewT+2fPsbUDjDl0IV0ku7HYuigiu61kWiZyU4i9gdzFjuR3mXSYiMdrj8XUVHd5y6
Pe+SWm+XXK78We7zZtjhwV6VbjVEZBIF1ePywmYVpNcqB4Txn8Z2voZ6J+M8CmCt0XGfvVRG5KFL
UamLIF/HMEPf+aBoNwux754946DWGJZLp/HK1kVkQYe7PsVvVjwXJ7m6ZFm3ElbU6wlTuttMtgb0
6OIbiI1iss/JzTo7I9fF/m8C1ILlRP1h1avnxxaS2mMpgU/LNNwl9DCqZSACtLUPTO3GdgAnPPne
6UrhX0JYVachi1u3a6zcBGmoRNlpJZnQ09U1drpyK/oRnBsYXC4joADz2vxlPT058t85GrX3kcIT
iu4QvnCsf8qcCYH9LssJTX2jBBySvUEXo3O2ujr0VuYsVVeV3pahOm4K3eKTpT+vR6KxTS+JnHl9
Xd5c7wGnUYSFxutO/DktraJggYtAfEMaVrpBwQxFHeb0GNrnBiLTiACvUhdCvpm+svmnQ7iFwRjT
tD+aKV5iVNeDOlukuLM9t9itVPPaeex2zt5MtKb3Ga0tIzZmscYs72ooS9Cg200RNsY3JSA46ZJX
HiJYpWM8fQtsBEFhZjeo1ynsIGJxovx/0ffv/p4IiolUzPdO17ogwx6lvWlplbm+z+WFCFGVjlOr
K+YFUv22quIEW9K97UJatL2Juh53jMZfVJT6kxIIZvyjL++bigWb0EUJFe5P2E8BdqIJdL3YWTMK
2S1gO+rQEmerqH2zRcTNr7OsKUp1wDIlcUuW8nfwpl7vktns170/po/U4k6PAWujURVF+GKefupY
mrUUEY4JVFk8y8xqzNYXkfuHLfusVM8fDpt8XGBEgjv8x7O9scqDbhjlryBWnH74nDuzvVF3dctk
V9E9jNF1XlbNdgFcQOPrUBmsx0f3cY3Upqh7f+B9SAf+AjQfwSdKe/olMzVO2wuyASY2nQjCsyjz
Bym6qfruxlQSEq3TM1gSuhSmm69c9i7zSGHtIOaFWXJLRjOgiiOgjhQKNx9SfppgX/G4GnK/wIES
LAmgjMSPyU2uj6obH1zWkaYuPFqe7/0UraaX3IfdxJrRN2vDvsgxV/xdIHqgYUEPzmFd49o4Vl5F
0mLYCvTFA0MA+65BoRxhEEKRhBk/p8n+oNOknB/u4a2GOuxH6u6OzKb04TxRaSqBjCYajR0wRXCs
9KgLsZ+N5/shr3WvEllTuuW7arwBSYAWLV0r3Bd2QmyF4tiw8voBwoT6tdkV+WCM9VXOHrejJCBI
z8uyeZgYB0GpcnOQZPgli+EB1mNVWMPqLJHsGPBrqKufIGc21/34rZbnhmplfVMA8Ch7JduSqzu3
i9GU+e6o01BPuJqsvwQZkEUgC67heDvE2IDwyXhHWJrjIFWfBuVg1nZdKOy/hzicOzlPBaxqWapY
YjuCPaAKrO34RmL3EoXM4EPvvjtcbef5Ok8bjkUW3PscVLd3+sAk2yVGJzmfl3kALJZkOiA+cu4k
U1OFohCBhMKDqkD1ds8UI3E21GHH3LXLas9Tt01oXgwrvdhEwREgdq1vVV64/dAFOgDa0fMw0EK5
hy59/IEgHGpKT457NolNBcmYHlgVQNYrw/AMqoldVnhJZnUpozXRbGbNaK4Q4Sf/jEiBMoRIXeJm
31DTYwOYS6o6FZJ70wX3kErkC9h2qnF3PD7iBIL3T0wmgsu5IVWCTOJ2TdyXXqrHt47eWULxKNct
zrkpOSmHv2d6zzO3LOseuqt8d66NA9X7lhtB1m1OW212SdIFLR3GZSJBJn08TUVFZacxO1cy5VKF
Y4Ip82MplPs4UZZ94XcoUrUepcSUhFv8nZbAEWuYAvCNvx4GjaAU4/U59rOdRPfZT7dFysbXzhA4
ZDMa89a89lug38AnDrbDc96ednuRapn6DZGdfcTsUOa/DWPxvzVxafGqx+sPg6Valf5Krr44lK7R
9glisa4USnY5wodcYisZ+uU5Q3m4a207183FPlwGqU3ekWQMq1nlG5mS7B8Yq0wbSjkRDfSs42zB
Zo3AMwP4Ket2UYnwLteQxSY3KWEWbdbPY7Vu9Wt6m2LtGw2OpsF1Opq+yXybcWWrdBfSiLl4F3IB
wiYeHDmuLpbX5bjJkGULQ2qz3V+0nwdrXax3puuzCySjTH+pXafNGWB2A/o3oHvovlqAtE9m98jC
kG88zRPYH4jN9LP5djvZj36GoHxgcXzPgE1TRpOTQXsduNhrQIm0W6cB/mvisGqGxdWPb8r5xVGK
GYEQok9CvwTus6+mpWcnGxFD1TsbtBbAJtsKkTkQdhjqdWMiUR4dwDYUqJ3f+jqVyw7KohqQPIPX
qJ9le5IE39QRVhVXAb33uFuGBu+WWtrzi6FbrBQNyLiyGPZbN9diRlrGNuy/b9/CWslh1bPmiLqv
FSjiYu4KHG5HwO1kSfEkAj8zeeADoHIdVWcen+qUVRGx6ufAGVdenvcFPtb6ORr5Z60JVKgS6Tre
De7C6zhpQQhvUs1Pba42Vmd93XmorRqrLjewts8slZ6U0maVuxSTdaSzMIwjMV1MF9uNM/ryMmJL
uSfv0tvjMhsuynpgZ8cfw9QsKw9v2PafQsnF6OCjKK61BCDpXcs2hGW4AQoKfybshnB8H0q0/LmY
UkQnbmKPHMGJJSaw3QUfjkCTV/fzBs+w0r5LX9Nj+kP9tg7H7jQEnUH79nCg1HdY6uiOAPrjqjva
O/oCAXZtE5a2BFIIBUFHR8AkolVMk6DK4Q89kXRF5rzTekXoTirZI7V+LON+wpcBG3eGWc0bg9xU
11cvq7hFN5BeRxLFxQEcELut7/sP1BBLB9mNi9Sqk3mvcT3VEZmywQWZPYfVh0r/vYij5IH1NXeX
TONiqaG1sggI9t8zEbYxcYoThFYB3kHPFu5U/8O5D/TfCaEb1puufJeTM/gSh2igGk40lJCZHrZC
nX86f4NispwQurrn4trq6clNC1gHAvF+behOVnsT4ccfFWdLIz0EPxBUWCKqko7LsTabu3kEOe9r
woGEzrwmaOq3Nwo6vmDvGOoWZvt4JfG/A7g5ZdxPxNtFRtY2nyrWTQbrmbUwdYE8OAJ/F8Yy0HOP
yfzRU7P2aB+kAn/F86AyPnL07FjwDnTMIMyWcJz9H179w7VeHElJfnMSID0BWxD0bSSo3QjB/zm2
u3DZ/bC/DEwMC8OOCceVBG44NPY+1j6fNejAfGVHsGZyjSGrVkYwwIk5YzyvRl2a3BapKTPeqqUx
X9iHLBE0qt+jaRn/VZ977pSZ1c1atLNcVJNptD3LLr+GSzk0+W2n2mwRShcDEzf2aR3TiVFvC3rE
nAbXfMNdA+iquW4kGsn7UmXKy4YUsjC9h7gpyP8P5V4V5hTT0CgurMUG7cGoHsNgcd3LOWnFZ3Vs
QJtrz7B4vEpraeTQrG+gaEg4qV/5guVWOht/BiaWfcMX2Y7BJfvQXJrfuv8zdjkzzxURVF6JO9uY
YiiIdRMNuQcE89W8ZmoxylBVODilFWtHIqNbrolwF2NgFjp1oV4tCPKgKwIqKXk0qgRf2+LI7uHS
IJRyhFnY3f27zEdM5XV0R8BYmf21e957db+kEJKfOo3WgK1YWhFX8V0j/7r/2xF7zXU8NrXWscLk
CbkL6ECaVgCMkO1rIO2yWlahHEbD9uufdNZBCwrLbJRvOfMx9NMc/trmpLXd+5iDsKRwIAvtsWi1
w3CWGo12LbDq54XLRJFdLwl1+jMYt4ptILMPcH3V30gp1S4kyMyVm8DTFF5MzQwJfxOlMblQgxpF
qbLiXlTthn+aVBxxzulONecKt7HoOnIcov86e9XkgY6x9qEazbS0gdc0+SAGOUH+hdHyvRUu7qrT
495aeb5LMaEHN7H0SqhaPTwyGJuLmZMWc343MCxpUvR659/4vOTDnboYdvDU55w6fH1vUyhzqzJQ
YtTxhP4+yEs1lIijJp8QQ+pqVc+3lRSnEoEusJ5cte1669T+H1fB3vFVopzVPMwY5B0GUTnpaa69
fS8glvt24g1rA3TH8eDke6EAw+CEoejahVy8b3xavjx5GRcidI0T5VQwVjxNceSGfn575t6BdUaR
KnACmMKYvEBd4U91eUQvlpfZXCEUEmW7g9DNHjWllLrhwq5nvxq4iUpKT8N1uOq/QrCB1U4NmdH0
E4r874ogeIK0+h/t5PZDsywr4fvIkehx68Z5uhcN+7hgqu+jOSBU/5hZgq78/MBgF1ThUZx34MlO
azZRwbAbx80b1Gu0CmtalG4BEgil6P7CKh343VXyiVO+4VcJzL6LGw/Gk/oxmzjMgPQr6PxUldhv
heSk1vXjVIOTUnDalsyzNt58MCRoYJVNcuc+fmqLdXClqPzDaqtTkEqsZa53vOxs5eQ8S3oWE4iI
or36Gb2kksIAqNawkAbbcu5IM19AohaByy2P1X19Icfz9JwllPzovtNiRxw3oTR26K8fYrr8DquY
7nhPlg3UgyWJLyniqAzR3k/7XAfLp9mEzA66s+KzRqYCLyIGizDsQ/CktWpsEzaWkrppbrGCN6jf
wzqZg7xdFHKKRSldDMViO8nLhT3xHAM2z9Lsnwnvik327ZlJTwMOlEPiSWQIP+el7DXJP+5arnpK
/HbqYVvKHvhgFGaOgaoEQmKaxG/zPl37iYLpJcj5gpUSzDw91BSgjUnLz+g90RFHEcRJnqjANoRv
P+9xdF7axEfjpnnadwLqGOQ0O8jKKEfqUycIe6VmzS98zZ7YTAlbf/CHFd8kR6RzySMKRYmcLwOf
LlbrrbWyU1RkbMeSTMQLsoEFi9/SI4ZFC4rgglAaCy2xBOEJaNPq9WIouSeLjaQ0DK8RWxZF9kRv
9ZoV49KPauVi1knpFZCRd6ZJUNSOk1Z+Ss5dJZll+uqFiDPC8cgT0eT7CHb94kwQnZOT6pAL/Dpe
dj9d3ZCBcN4v8/tSOQ1lbcZyvn+r7jg2XbOGxFqkVmbJL75isFJmi/yV9SvWK+2kWyRX5xJmnxHt
L4l6QHNwQ/Gvvk2x/dTiZYcF24SZ8/vsuOIvSgeEPOsZaOeuRlWAnOq3qDs+y/R3ue0V5SvkA4JD
VzYzJcY3yw49/pSYqB1FZbNHYA1xmRJPLu+0WNFoaSVYvnsHcVSXX8kF1bk3eGxrUW3u/b7A4Oqq
j3HZwOwLRVuPAsTrubyK29fjh1JlzR2iNY84dG2SVpUCj6/1ASfoKB/YF5fBw62om82cdVF3masb
6sEMf1NEvsy9tDfVxRscft3rj3YhmjAMX5KxsTazlhvAbDD1rtvR3ijYJ3L1H0ZQcbcG3cAqbanp
6+qKxoODsWD7kEAX2Q+JSk7Hl/GPhn0kJDERWm6S6SI/cmbMapmky9xJEINf1nxqAim76Td2gFhk
wgPTNl1A8fMKOrME2fCWfg4mAfQ1PnEL6FDR0zCXeP7lwQ4eFzKfOVujQGSgxvQS7VYT7c8ahqW3
NUeKLG+6niFirNiO2eEh6obMTisIp5yakMy0UJuwO25Getj3aWn37aIiHBccXiLuMJXE/K4T4dTJ
NvePtK4GQf4+aQa/oub/qPrpViUwMjjEGd6s2eb28mcMkbtZCuj71CQMLA75WwNm+KTS+qySDTZA
y6MT4cP3ZdPMCd1I5T+nSK/oBhKu11HdAyv61eScGogE1j0e+uIx15F9JiXqOK9EwlcPAZVSCh7q
3bzioRStJd4FIWY+foOFqM0v/yGgS0m+ZSDaGW08RV+kf6ubgZ8AkTaarz/Wo9/P5rfYTZKSy20T
cyA2ycBodj5nPun4MhEcvJMciJ9d+oTgGJ4PE8RtB8WdeIwZEnBnLUGZCy1d093iYHq3wgviDn15
r5SGtCcsjUgwOhPau0ogRe3V5wDw1oqU2cOtfGdB58XMLIUjaUHau+k/EiPcE5R2ulxOpcCoPRq2
iogtII+qmEUhm2dBorqQcTN6+kOkO0F8lFqUo7GS0P/gCJosyHSSlr4P8iIwy4XJdVChubSwNrnc
5sV9QGJLBy0wnHi1qljc6q+Ebqsl940uxD4I0YZoCJx2HsZMG4GFn4IBngm+nZ8OJJuSV/LqiZXh
zKhW2Zkg/e2DHk7KkRL+h+RIPLSwG+SfjB2sQIDaNKvqc6MTT5Yr/e2a7ztIF9vXpzh5GGzPIVpu
pPfj41OCiPve/H5VLVhLnin9FyYT9dMfAR1/8mIwqTAdEj4wzlLbhLMgC6us0mExR6la9rK97muG
5e8g95x1RHqEpnNpX+K3MpUZDheKTUdUOll9o+uvdMqZpXAGqvxpqbQegSHatZWwp3MLTpQed1XS
LFezL9qYtLo8qvogGioc1HOPzbZViGvKxjBB4ZXgbQgfBpixVQxRfePS5RF+79iQ8XrKg428Pzs1
IS8FpACZYqavuTHRkqoJfI30WgyknLju92GOD8LKM5hY0Qhhe/94SchaeHvWZuH9BCZrfn+pttQq
mF/utjK5WNJh+R1X612rIuxANmgXipPdEJyXPF4tVPkUWAHXL2VCEQC+I/xgZqVlVGAgMtenbxRj
gNeKnFVlJftM4n9boLYUaEaHLlyYwDx7/cIlyJg0cHvrO22YOLXcVvZUYuac2eWgGlme14bhM4QT
O9v/YouWJPA6W8c8JBA7epe0OC06YzBvXOqRSir7tyFH+R1+ej4VhJ+2IgGfzGe1cqixowNcLwXP
8w7kde6vQzwTZ7l8Xh5CiY2scWowoCQ2infXzeeIv+FOXGlV3d8jgSf4kYKKEIDYkBhs6IgFrQ+s
F1nbxTzCECfNrAO/E/t4t8dUD1b7ej+VvKn6gl0wGxQTauZbrWhjGEPv5RsHo5kmZIZN2IxhIqzG
RfN0oxj+sNdmTiVV+s43nq/17DkU351LWA0FwZe8qkULXeh2IdfVLNSHy4g96Vpmzm5U4p/ClhL9
pSZNmggodowes0J5E3BunYuJ+kmFWXO+qPsoeeB+gfKuKWzavsQBX6QpWSz7FGngiIegeMT8jB7J
xf524LB85jO2tmwKi5nsBh1J608GoKwKsKFrCt0ndJ9A7XUSXZN+acZ9KIpQzSdcyNQqzQl827Dv
ELUTrrl7+S+ynRrRxB2AxMWjuncoxIFHmTo1BUFHBq3mO4hE0tADcx5oZv2BIerWy6nYmUHLm+v+
BqIuWUlkuASww2g0NjmJ2ZnZSuVNV55U8z3zBubtlbJRWX6vJuvLLjaTU8gqmcUL+CX8lCg3NjFb
43LUHkdBswe+Ew1unc1/yH/IpMR2OkzKpoukbdEskdxRDovS0CxrzeNL/Lw2+MS3/uRs+09SkVr+
95yPJPcNnCZp7165gBiy4HZ2yOvuDj2gEClL8G7YxAnMxSSuzINx8A6GnCrPoSb5WGX7zDYmKd77
SAwRLy8EWuyK+sKbKEIc1gy75rpyVt/T2sBkzBukOQknRy0FQIZcIcLj2fagfXa6Q31yes05EhlY
/MfIEUB8mb/GxMcOrknMdIw480nIzBXA5xHxN7wS4y8g1HqLIZXlmr+CAOKTw32AE1H1iP1mesy/
wTuHdFAx7FlQynYM+OiZY5nykMJdF8/EV63S0hFUzsnv6aIhrPeVuYwJs23ESotMWuRyPdVt476W
vI+8XDhEvA65PBPMIAR8Eg2mCrBxkhP8pdh0/Ok62U3g27QMqKc6D25KUvBMHmxDYqtlRhimjpNh
pLJ92HPOscJM+iz5l50xGIK6iqpnDpMwHnR4wh9lFFHruDxWhUgg03jVEqF2eGWxfK70jA+BtC/z
L1TfSNgU3IHKyf2tYBv9PVjHLzcfMSY+EqkHupKBhKNpHwXx9Q0mwX1SbuN6Ig1/0Ucty0kaUsvh
4YTws40we6820s/DASyzvulWXvYa1XVdNs9E1feFkGA+6lAvriarcb6kCD+J9pTcBlCkR8bwZp4C
aB17wBaJBafajAEIoEWub6i6b9OocvRWa/+DpvMjRkiTvUu8JXGFNZ1z130kSk7LDxO4Kq7xGU4M
eskC5wtly1mvyb+VzfyomWE6DhxC+CpSkSUKLlwqiLsYH/ibmzR1IZKFDhlrADEPseEFO9ZvVV/X
z9LFnAmuv86CnAv0BTPpLFyDg2vAgsn8tiQxqZkTOQlitsH8mXvrLaAo/MlVDtQrmwaevlQYswox
ravXWfjC8DxU7JpzTCOVEMDJpDRKIZuhpHdaC1OCKMqTQWXDEu+woSMWJM4DACRlM6Fxx/E/uPWX
c/GW6iz2MkZGNSKo6g2+fJqi+q6EbTFrfn39q5LvzpPAvPTq+T3RH2kobWkm4vLa0rmDrpItmJq5
fr0jBm1gIqrKzL3IJM9ul5wFuQdioAJJCBwJAESeSly5dvh7Vdh30kb78vKXXVdKEGKLw23sIfWR
bE4/QBY/esFCnsFFFmJdZlZgnSQZanTtMTp5yqHdpmkvf6k2UlGiRds7wrGOI+J5NTJjo/3ReJYM
sRWiY8p3N/JjjLzIH2iR9n5P3pr1+Z3nfsSM+KnfvFSqRGGjmiyvnNpt8oz+ywEhfe3dQiEDt4px
I9rg6ZAPvhU2h+lFMqGF75edl+cyKxwldtUVi1P6yRfy56BiGEzh6yWb5fFMiXG4JbCvr0DcG5k+
gzIWQ8dvFP0YBKGrxb8fxQJF+mxmcyLd0i88GhT4MwfAd2qY9rw8zJxakdORDc05jj1QvKE8QRKo
GgsCXgW2Yf/jRS3+UcgbkvMRh2GKK6Wjbytu6mlIz3WKLMHt460MJBMJIG9hpFS572IZjm/0+ndq
ImBSAVbPG3CcgqcZ03s6sEA4cGh9xZmpuGZgB89Sy0ZN7YjKd2plMEuupC7B5s1rGjbSbNzjMSUk
DW/52vQ29BHlLY59jesi0KuaVkQHE/YQjCcN8oisUNBfrIun4z870zhuajVvMg1Tjy0VdVbABrvE
PE52sVx3YEjXsxFXXomwTd4K7soOTTyJpbJ+TXGSw46JAzq6xFOLo94YakP2G/H1ngxwGL0UAyxe
03wh1avVaqWlEsmYAQSj+whw2jCBNjFCe+N9TEtvIJiB7efi01upLTVqarfV+rCUo53p2DXWa7Zj
xWgpJ/bb6+LkiCgmv4L28iOMmA8hCkxo4SSksFuZGgth2yMUlfnsL/DHZnaw3stFF86Qj+Ua341s
x3EiFLq7MkAYjcrA95MmU85X+zr8JhWU5/emqbeRTKhW5vF6dm9VhCSA19a+T5MBEUoo9in37yBk
C860rDWEFv5Ou5vJ0Ny5yqH5X/RS8OAyesLKyWLfqAgSHUoFviyQAd/khbbA1scORYm6hPKQ6/V3
5lPma1+CsMtpHprtz43/Qj05/Wxu0CIktF6Eb/cSmC9i3odQptcbjHR98VDNVN/M+W8wbp4kOUd+
xKrrK8B/MKzR2rlXDQhzVyKw/ZepFkerULT8BTPd1k8PeOnLtyugY0My3xGoKrpchBWCHOa1YhYn
Rjo3tTnedg5ud7eX1Wf23sGZ8ED1ub234Zn1kk0mdS9/+ChMZAPA9/QVZCfZAzsem4I+75TuO6XM
YUnn+4cnkXDROnLI6jSr424Zs/ePZKbx1ciUAMjmR4L3vFCn6HcERyMiWb9R8p0iEShJePE2UCxb
2twrFolQeFHh59m2ymhnmsxj8WE7H6bJ4IlXT6LBPgxkBChYytTFcyJ5CrRRLjw8qDeob6/efqV8
nh186mgp3himu6ChoS2opWQm5J8f/XoMjSPqcaO5RzM3sMjyjwzk6AOB1cnaS4QldyHuyXpTrNvO
v/mW6c1+QChf9m71tHbj9xDf+cR7LoTjxQ/i7IxioGdId5Lr6TBJ6lU90v9Ldvdc3lCLTyYVoi+A
aXmgUL5z5R8Cr5yMhEU3lt4GBmdxm7bbSFfE9FN/+cWM7RS0El7hZM8AJOHQGn2jOsPf9e09yTQ/
ETm52XtLw5nZsTVucW8mAFAU9D/Rqyp1R/a1FUqgsxsUqOo8uvLP8XrOIime/tnC4eSqNNybNeJs
Fs2ldm0vs1nSxUR/DXAMNxwD1zrAK+2gvuTRK9kw48TpX0eV/WX7jPPpdCUyBQ+BehmrxnJ1R9mD
IRQP+8vC584FvxbQ09pQsEJ92lhAlCH9dKLROcx2TXu5f+oLHZOdHP3UDrcJ+77V0om9EsWe5YI4
26umQFCscn95gEi52Uw2FoEQzilHpc4TbOW1JRmZ139apcrTmpZe8LoujWg/LxJfY9ApSnLglDcl
/1p2UnNNiMnc1ZotoEdOUvIOMu4SugSVKRVVeSVUzQe+aaS6bcuBaAD9fmm3TWDBr5JTn4aakzrQ
JNFnCr5r7SV8xltfd9rvY9Ugt+nmPk32NyWVBqRYGzssWqOiF+d38wJcAk+tuvkteOGGMO8Cjkix
5ZzATlgU0Lh0G5As8hc7UMYChJiuX9VEb9wzP44mIIYkYOdbbr9FJ+3HLfmRO7tju/WYtwKalfAw
rLuxt7lJ0yV9hjYKxvUiMlRftAmSUe2N0MJhiYlgaIKna+eA/KTVrummr0hoRoTHuudz4iHGiphb
EABinHwgmnBlVwryZFgJB/exvQkeRZTwidV1jGrD5uZ1dMPbHSCQRtLFtE3mUm2M0A5kENFdrnSh
FVKaF8uS4oSs37a+oiWUgr17nJkxo5s8puTQmyFLgonY+6nbSMFEcEKnn50bx8liwNpowNOr8vIR
OEEMAz54FFZs4Fg7PjsdkQ/lJWZN+H1lRAk723Do4uB7kry8r9XYk1EA0/2QBxVmfxMmH3kMsqL/
o96eld9VyePipPfTYa8N4n5cGQVuZBbKH9R5M2VNYpgaWLK2Vl+ia56LzI9xdmNHngBNe9bCzZef
7Yebc8LujivTva55bd75ScfDDjqHFMsMQRtEhOWGrvQ9OGSmi0lQfPrrswa3QF/fNIRniU17jqwl
s6Ys0Iu/7O8bCwwKYtqRLvaTQedxqjHeSyDimLXt/gfXiWY28qikHcPagTDcfMj4D/qotVFptvgM
x6KGYdYGo0ApqBeddOm5VXKRmGXTMqitoaFjdEEgS/kFmOX42wb3a7bAGX+RFepEm4im4zVzu5zX
AvvcWYBEMW2MFN3nVfWC7+a9eCHsaDofMAzBKCrHhgHqdJKqrb5On5x8KIcv9tUuBw5ILyCjaM0P
Ra/pQrdlcSWnI+yEujGKTY6pPgUWGjT4kJfV4eriUku/ExQDmjTbeKy5Q7vxrleqbDw2KIpMZ59I
j0q7MSB8S5e2luPRBMuWEJhIR8/ghmj9/Nu6pVLYfMxuwwFgD7rEiOtv+/obzq5XrHZjeypizsUt
qmDKDG7+ipWm6WvX8b0FfzLzrxZIJMw+dZmOTnvcXqZI139azbyX1ezfsNY1DQ+UnTrJ8eGRfWcT
kFdn391bdzfRE2tdRT4DLuxbBlQuwKNkgCs8njsrqiN7/cCn+L5hwhx35anbDOzODTU3OKd+Tj03
WZlSGpsMB93Z0lIrBoBCMCTVlCoz1Sv/xX8yz2t9YqV3pdEP6+rU0wrMPcLjPkUjxl8+gxQnfZRL
sIr0zN4evO2pJH5vuC/Tqlq0UrkYgfAv3Y8D2G07hE11NJgRoT1NMG817dn4ndC/DMVRCj/XyQSY
Y9uDvJQMbJ/Mq09cSp2DNLutTh+DqdjesicEHMrwxx72aqD77OfVkgM0hmybwLZV8QqmVDJvl1nK
TFXSNWu9KJPLXZpl7J7JnHhYBRhdRBd9hvboc2ox+ru3L4jBCKf8veVfc1C7PF1V9+9Kl+0yiNEO
j1CtYiFV00IriWE0eNpKZTxGXv09/kIoXGrey20ZhjuDuMw+Dx6yxCQ1r4rWXFhtNiuZjejgHQE3
FBwGSYcO+eYU0IL67lQrYs19cwN5d51qe7dT3SbNxB8y3q+TnmeLWpNyP8dyfk7sdWyM4htMqSS9
BQAHFaXlom1ACby7vzLx5+3vM6UyRsWo2WrRy3pE10RwGbcN9Wacm27PqyPvLTlhtPPF3UdrsK/e
XjuJROnpgUJzLOqETCbEq8i1lSxF9k12qkelejcWIpfjQrajmiC6G2qvmrSiK5E3Cli8+V6Wm9Bn
0lhtvve+lfukm5aR/c57MZ38+rMjLxup6gqHsHdiCD6EWoqP9tSEtvA3KSNdJjrQ0PbqvT/6dyAc
Ofri/CpNE7qEWkGaZ11YzgxOoexanQfJFbTp4fkhpzXVyAi1brOsJkYbHjTgVTJdckuGtt46Kg2i
n+ERUWcqyKflpoWJjiB/VWR5tHc7iXUSXyuXMsQtReSOLXitc+UMkq3pjiO/tj5RjCvgVaQGlk0q
UhLfNX/h9vpb1hzZwHD7UYoGSEwdbrgNUc2bJwu/SNNGcK0SfTchP/7IKGj3bvssLIQ7z7bGDuEr
pEx+aL7qwhEBNQb13Me2uG1o/qi3hPh4tasdfrAM+UBpsTDwVOg9hTT454QC99AfpNbAOMRxf8Zt
9keUo02YgkeaSezD1FlNNK7NlOkZ+KU6XwdgW33kbOcrINhtCPa8Te4S5+79uURoYN/iXQx6oSba
1TgWjLdviWiNV1qmGgXjtnQSX0tSfJydhytgQihLlygzAe2oHE8uNk+g5sL6N89QpvdlaPBpgJDx
Wbiwm9YBnlnvHfruF4nv/toq1km+WgI52RSy7aOh9Vgp1FaZzzqyzHof1LgH/ZOD9vCGTrsuhb9O
0kyggruF0b/buumJrxvYaKaT9ozSWhisEY3gEVIXhnJdS6Ei5ZgCJ+xDkJHxevSufatvjePnOtpI
mzCByEFi2lPEEbPeB4bDfKa7lNXUrUIAO3rut2UfbaGJEAURNN4BJpPpi2wgm+ztJ6Th28PO91/3
lhC7crGaqB0ycQS/x/FEk7HW0FkBnPtNmc3DSxTjXwcy2Hn3ASuvDM9N3s4Hw5t3OUU94VScXdqX
VeD7sT1dEyP2oqCBEt1pHLBb6tagTdHR9xNSlCS03pIqFfT7/k3EW/Us3Pa+5JjhUIyTGAum56am
/V8Fu3FQiFR4C+fRqj87YD7MkXAYPh3kSZdA+XdiQgqOdNeOaUtj0Gh8YDu3CDUp0kBJ4yg84fj7
GxBrwdYGuDBsyEoYDcUAURFl3IBNNvdmCDXlTFdMAAGAoHYJ3iKY779yUliHQGeswYlcC7nHYm8x
Vr9GJNGMlBEsT7cP0iqaD/1n1wl3XHZ8EcCOGBE+Ds39Me7D4OXe3gRCDOYoMKGHzKS+Vy9HVOaP
P5Rx6zzuQdlOq6oiRHjFMI/dB6tpwOEIHmrrHEuZxE3xXHbzdHHRMfJzXHCOD8TuYqcZrReGbPDX
avduR75Np6fbsXezKYGy9cbVAV8nPNebmT6Zye/UPe1lNkFwUTZKgqkUMuakFsEZlYIFll/i8Xsf
9pUcvqa+GeyYIncYoNUUbs8LPSgdbx4bhuNgxwxy9LuquNEhoSwKh8moUuoXEQAE0+1dpfO4kE30
X+V+EoYE1oGqmEgprL8A8n7TAlhdaLRdU+p94pjHrtj20oOrf5OyX1nkcwiecYj6TObVEOf46V+/
fugIn6PEKFzidJI0RkfP19AX/BHWhTO/2M8KFYNOASGSUbALPB1aDHaoRtKC2/OEx4P1QOJoPPIt
Ny9WuCf0H73B6/GhRcNn2apfTRSeqsIeHHDsKDtuesbqJOQwFYNVQKaYCHU5p3CoISpNT4MZ6Yrc
ZDh9v8+9VpByRdwAKJ/7gRvvyE4YmZqQnf1Wug/trubkrJDCFx8VoYQC5Xs0vbA/fXeT95DDRyUz
2MR1ma/hSYF0hZmEL+gOBHvAuKnM3/A7abbB72Fxat7FEYuQKFz33ZQdAMCNftgRfsZC79slc3NJ
5Nbv+2cUeU3cgKf61y5oPvz6Q1kmdEK/ZD8NMIrMU6qLhsZNHlv1sG9QUgR4ICD2TqO2gfs/ziLO
0us8byPov0UovCbxnp7JjzjMii/mHPtKL/PIvN9bacwN+Wg5y/gTrYK/VIa533/ly/06Z2dcmYL7
kY9jbB9WOzdUMoWCa/6uEc1Sx85hT2Zru+d1shczLuXA8684wA3LBfupXot2b8tylTu0jSbNwa9M
Db5fsePXf9M0+AnUzEyeae6hKPP62WAXSCbdOUH1liwUSu6jRET8c80Q4ZR/k2w8CObkUWi0GTdq
TL/ruAhq7YGMHEaKGk9UXFeH7/eXPcRC72OI4Sfh17Lha2ARjt71aJaFAa2MQW9Dd3GilFa55/OL
izy11BZudItxIy+ONSxOKN8CdsLToBOszefYZP61cSvtnAs0sOSQo+q4KbrEbJcJw2D6uMaghRFQ
NLTXKvZRrly/RUmP1DPfil2CTaTfQca0vr8EwQ4L1N58i0JdqEuDeXi+NdZZdJ5jXy23tp9DVeqS
hHfB3GtJoPkpY68toxfR84LRQvt9+sZP56CnwU2pT5kjOCNC6WRqGpGyGudMOwX+wvFo+ZKLthw7
/F7E6B+qYwNw8k3uwpM+0irqN7MesuC+PqjmNHdeo2i0wcx/9SP7TSL1v2kQozfP6jVv/j90cSWF
o4ACgwt7ouTHpvuByTMonFH6pZNsH28XaNoD7xLPoQehnAFNZOA6EjbR/3ddf5Z6WLiZOn1R6awl
GLYlCvs53dA5CROpjCtzV7KE74Qez5Nhp4WLhJ27n1n8shIlE15Qsojj1wrNW4Th6+yI4Yl/WOdG
mKgoXHXQnoflIP6auaisRPA19EZVub3O9aI15eS873xv/1Qxn1NzuxbBV/E/xknoUZUBGs9OBQAe
8AmgYCNpEu4FWJeUfG7wY2b36wPTxFmxItnDy3vuJDoAes8A/rfm0gkLNmcGB+Gs3vYgbet4+ETm
qnugcPcjlNHmzbOqgGQprOiEQoaf216+puczJzzqxqQEaoNmygIYQOlE0gs+a8zNY0KySmzZvhJ8
8iS7i7fK6Crer0PfwmHU0tm17CzQK/LPbHPZkGi85EsCER/E0p9RJUwvrg5P+BRbBaVHlt8+TJ3H
TzRcQKL/fvcWBrlpKzyYDBWoYfzyEv6jEEKrQaq3s8pF4C+gEjKZmTluxfiQraT7RYeTQs5SUsTz
9D3OIID/6GCgIi6xlgp6QfMNgaa2lo+jGyhMZr7/LbIuxYtruwH7ZCPnV+PyWieIVBsTMNnV4KEV
52H8UQ/Q2ct6vRUPU+q1jr4vtF6Whzb6NXEIxTebggE8sPrwVc+BfAYb3j+VC9xW3zJDgXmAJ4Rg
Lnau/4k/wc7JiVYcUP3cegqTEH63D9nZNB9jR4lKQAQwz2LFWFgkHLOmtHFVlLrT7RRZD6S1PW8b
6TZdZWRWvu744MfhYwqczb3ybP2H8Bs+4DEOljA4Gd9uihHFuUazJfh0tg3V6pgvkT3r6g05uOfE
h38feKFKrs6g/T2ve86Zl3JO96hwBmr6NdHIUXz27fVxRjpnZWRYcGnLXCnmJez923FFi6W3tvJK
p68Vpaqnb/ZIXtXdJDHmd/92UvnyL9Woo1DvQuRHOapsg9nZbOd5v8Sf9Hg2QjhCH7iWRkCpz8Ut
3MbhDU96KecW/weMb3Yf/hVLzRCkd6RO+ggtZeKWdszq1VQv4jAff4VXkFYT1jvyLSS6l8Vyl1Te
CsXW8wkMR5B+LbeleC3bSihkLcVXlD4Kh2WSav7T6KF9tU4ZaFwWdaHD+EIZs5Efywa6S36ZDNkt
gs/Yx0qmDyTJ1ZWACwdw/i6+u9ilPedRJ+CWWGji0wCfT3Ba4Qe1Hvo9P1Qf6hve+Q7ufmltlm48
QG6rE0Prn251qxdTxaURTmQl5wU1kKpQ/bczSKYHFoZaHhhheMm/PxU9
`protect end_protected
