`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PGHFNiR3BP7XGoNdt+sZaTmGZWIHImrHr96onkZN6M2wSWG6MSzLnz3xTdAOzrEb6GdU/I3SQ1/j
1+lecrUFNA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MM5jU9TWbR6/PtrLhERYQFUfWh1JDYUP7wzhyRLgamuHE/Wi2r2uXHiNpYGCrSz45T74W41GsUgm
9j3mMtKtZA888jKVdsKre9IS7ln3Qjrse/HwU/HOuRjQCYTzBCThVnxR8/oeSAPnT9pJZpEHuD+A
zpyCvRauvZTEG5j+scE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fi4nhbaxpRjqCDd0M+9OyfKserp7DStZWpnATpp9K5HcMKXXPcKQuvXtuOUfLNkJ6/72ODDZUv5s
NLXbc2oGGClaRwTUlPy/zDhhyGD0SdKZjg/1wKTIvwt9SYjLQTIlj2hFAI3n0xZcsDXA0pbuM/xl
XH7YQLcEUH3YH5qoLkmgkhPbmTXc2KPGjbYYIHaNZWuGZJU7o1uI+ek2P6xx8ctzEu3HsAo45nFC
pkPS5QOdITs6At2bp9c4hPHKgdIHxE03FP7exaI8HjOQVl+vQxzTTPGcmbRSjfgA6+Iqp4cM46I5
iHmVPY6nZXLj5z0oMk8+Q+8ka0admCYkTIFJLA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SMBn+Jq11bmR7KsSKMN/Ncfxt59glEf5XDov78erxANfLvk5rp8O4KeSybmVABHVHGwnaOCbjI9X
Go3+bpOcVcgtlajNGY9HSWVVqsxS48RWPpRm/0DlUcNwjcdHSHyMUaYgDVlc/hlppbOgHJaPrbNz
1tAeewMQfrB3dx/2BXQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YXz4WZBI+ZuRrCi4Gfpmj9u007zhUaapkKLeEvEugtpisG9TvoG+IdugsLUxk3/cVor1HoPm/QO1
wluJVsz3KGJAXTtuWA/G3rEwGRbTLvAkwUR1D3GEekAYWWpx8qYGzYk9iVldd5qkpPJp+utczsVY
VXlhLuQvsaUI3g5IXrW9/nD7tPCJrFG222qhCnuZoBaGj6PQtJ1XoyHpkOLjiV/ewV6NJqNp4m6O
59u+GtK+7P5m6nnmbSdhQDFMZt2N46N8Heecoc552V+SNhU042QleG1xn8JYmm+tIO0ppZ3lWhM7
q37Xm623uEmvkgQvIBgd1+0N//XilBipT3JQvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18352)
`protect data_block
BGbGyJA49ilw/PQso0auWhuK+BEQ6+KJHHeHuBaC41ydAaPUKQNbIMfnJ+qEF/pLo4Q8BUglhRph
iujA+9DKW7EK572eomDh3XMKEylnuW0MMAkQoPAYZX3Zv0zj42gF9KdTMXU4VIZEmoPUDjyVeCNi
zSn8w7eQa9EquOfnr5V9xgZWgjd3ltIgVFnZWtQ8hiMma2GYtzQJId+4ZKHkpySmRDT9bgGB7ag0
BFEscy+2JImNu6jPAdJ7W++PHg+9ivApXnD4JHJFbmD6xoUJ1QkBS2hS/WTKRgLa58V/VlO46TMM
xEqUceaQyNXI5x+NGlVFZwbI1oEtGfxVmsIXusfvUPj2GRnEZ+Gk5Jo+ekyymNTKCCeic6lFzlBC
SibqDWs5f3jR0DTnHzvy/6WajFEkWBqDS+cbCrkSz04yzI6LNqzn/Uf3/v3BcYFutO9cd/D7sbWf
gxORqw7PLBmL1jdpoSHO2XCv0g96anqP0UROQfQYVzzuBldkxb/OnkjuSR8599JWoVWEn5Gw7SJu
KE2lB3Ng0yIYoPSwPAD2HZ7aacWtIFw9d+OZFCnu9SpR5f3G5oxSeOQ+3+GH4YHzcgeG9m/6pqDi
NZkbEJ2yU0JsJxZyjKo+V6NaTlo7/F+tjU8L3T+p+J1mEvMXoS+MNXcGCD+KzKqq7DHJO695trWJ
mdzgByumVT5xOxCsZ3y0w6FbcZ4CE7sJhvDnWzLhCc6QedXNlv8qI8rSMfCou/tllbbCP3qVKjXX
56kj7hUWPEoA9ulghkZZwS1rCkejhuvwQ5IKxYq2pU8csJKYdGhjgLwCLoPNG8QaKB/ElbXbg+lU
M1U/SjuentKsD18aqy073aJZZ6+lP48R65EO2BoHv2FKKm1kDi2gOa3zcg+2TmT8/83x2iFjuQGQ
TAGulKNj2JCbGqMUopXDPsRX7Oy7EJj2j+RadajTabJMQu5YdiGaPGbaL5NC1pl2bfGHdKyV6eLP
biLPO7gTBT3lB9MpJZzsc5qJFffQEZyvmvYvnL7dNCYKSr/MRI4e/owu2FhPRrNZ52BBO778NiXM
LI6QLK/Oxe/ZmkP5IBdrBLBmKRcia9kgekIGOhe2ZV8WUPE+RPXNCSiv5ueW0Z5OEsKzZkthx/7Q
dJn9WHXyo/ByyCCbA8+iGaDx1aDWuRRy/GTvk5/OGjc0prT0i/WlbnhWpkZhvxxfJiC6Df4LdpC1
OoNDzD5sVH3mQqogjvGZxz66US6yPqsi8h8jYapmusIJ1Vdv0e8M9hu06v0X2QOZz8TOPE0S2bas
OSZDqh4/nL7ybDQSc2sPSZXR4RcP35LLmxoNN4ZvXdlIuyjYtLis3pJz2xLq3Mfp5c5QEe+X1OXb
+ZN6B3ALQrzbuBJX2KKHB96aq6lKUuRnigYLg8eNniWHNeV7ihTilBRiLKFWwEMnISUiYYH/qRwh
ddp+yqEgx+gEToUFBLDAO5psyBbExiJTcpo+kYozhkFmntWMz5ktyugXS0/6xh91LUzMgTy5vn74
cSmE7UX3VDgXN3nRJqum3C8rSkYjGGnVQP14zId1vI5Ag7JFW6B8KLtSbqUq71uTZx312A1aUpU+
OmWanqdNde0/TomJ9riuJtD/FL5yoa6tAHFe3y/c8JNDJRDlSZussYcYGNUF75sK+Qd3y3tfQrMv
gzkAeLo7aJj+sHPp8HFAEJz4EaoxjemAin6/S+BVaOz/MEzttH8DO/j997P32BiiSElR6N1gekYO
x+Qp8YXTCb7XK1ao7QhV7V2Bn33uKwny1dPdQl55Dll3TwINybauLTbnyzmYO6Tl2X8TmGdLDo1M
1Nx4WCLr8v2bOLE1wRBqH+PPcHo8rS88Qh2Gtc/+ffF80Pg65z5nugQ+Aa44z+sjMcSiIbkrJi85
zrdlsEeA/IABVCrtli/ge+Gx21n5YIHBSaL4IV6gQL2+pCbjLoYFWILgSlfZAkO6uK2Dk/wUfdLT
8oOUwsJxjhZnRjK0y5Cgb/1sWWz8JGD+aQ+M0MAsEkKA9V5gBF/+IauNf7jrRkO+/HcEJrBDE3NS
avRzmItxX4P8lUYCVAV5Vg43WuNtPQRXgWzKM+7vycDTvFHsajF9B4PFoumOXhFYVMiccvxmqizd
GKI/ec8/37zyDYD7TfHq5JA0YSm2UGptlVEzuWgeJk+9SNdSJ6WWyYXc6Oh6r/oXO3POn8BE+bGY
BBm1gBJVUNHM/XYKni3y7+Au79QSIaO5Kh8l9Xlcm+v+BL7sam8uR3nsX35Oc2TvX50txfMsB3wV
IPlVHxLHMj4zQox9fs1G2CMXWdtWceVfup6+Q3vh/6/9fx7bSzpa8heUntsVzFPmffafy9nFEUQT
th46JP9qWiHaxYS/jjwP13GS7N2WsMVzHKifPV8IjbWB05aC26+Am0CaX03FwTFSMqLzIZjBYacS
Hk/JDEIQwH/ZQ4mqB+F3XUP0hyeap5Riu0og79bBUPYMvlP9euQjPvjq5HJmwDMYDg76AQOaqP2s
3UZohUCY68gbr0GsSRLOooCwzCnkoESzEZvgLMJBAsvPi/o2Ki3ZRKdt5dmwDrmFzrppmu8Tmf4d
NkOvPB+abWOMe0chi9A+R8KeiAU7x8jdLtmLxJHhpJcE5yWjn4mplQSPOSfh8TmAgd2jRdLj/23A
CahDd94F0XsHcyx/nqKY17bjRTYe27nujnM+j/EZ+2VBbT+cQz8qdBP/lr70XlGZHke/O8RxE2WW
kCaIxLmHMzXvZCc16NC91/i6h0t8xB0gp6SDfpO5vPrvcAb+Oj9jqaxyAzgR9i73ZHmqzur+WCvI
GFtP/6sF64so3e3CX7IQR8uAj8ZIQNfUvQncoXWyaKNz2YSxIo0DYQorrO9710gVQzgq0BInYEuN
qCh9QtOUZhh/DtuJLAOwY3FtKqqbVD8/hlgdzj/8jOKR4zm2Z+htrB3loLPntBH9gFqw4WFoKdL3
wQYI5LVR+3NxqO6Z68tpSbvdLm8ZkGQGlySijYT+zuimjZd8fgZmbKaQvrC33eTJqmonaROVEvAt
3rU/sK2I24mV+DncENj7sERA1jkMFzI9NidcgUohIfDXJOr2GnVQUN++TzULNUGATS8uIyiiOM1Q
6JtjXDLSXRPhEOCdeZlqm4t+4TnQO/HOvSUElyaPywSiHZ1qasScrPWAgd/4UudACF8notyzdrIN
zRlgQFeet+L7pgviqkMyrNT5rhxicCuzCSdtz1W8q0UXGfb6WyHOsOltgE8mqpk8LyTuhJXgJKX2
16LPI03SwAxb4YXfHCY4Eav0xGkZeqi40IhfeY5WZpoDurVKFI02qxUE/IPOih/dI5uYoY6QjwQT
n6TGxV7P0qMG2bDFwq/hNIO9MqkUaeGPjXe96rtGxtvJPkJzJIDRwTQviiotVTjdc7wVUKiXWtW8
gu0GZMNs6aTnb9m6hjCglC+tmD56D40j7Gg6wouRgdUdtjsV4thsC09a+TFwgZ9hKdHHcx6lknhD
kZsURXfjr2K8iQLKi+E9tiq9hj1004GRY/g+/DyuQ62DyLz2XVPNYqkHESJ0hOlQNAUlj7/xI88K
1T7/sanLTlXXd8szmRgCsKuQmVMMA24HJsotcBT+kdGTKWktpgpLVze8qU9uMqFbWL8qxpc1/3J9
l0/Ooo10QRQe+fg77nUThJvyrnwES1j75XqsWpJi3jF+9x0lG93pGTawLI/t4ztvrxqylfaRzFtj
Kw48idWDAbXsoSsvFb846kRFSU+PrF282taEafQRjdmEqr8bMJX7Vsd6WJvRA4jViTjdp6tl/fcQ
ESQ04oOOmxmq0vKl+JOjzz75NsgZ2ELm2DV8qECOlLW5ztNogFFqTi9zRorwqsyDRGHCLkbWbMJY
R+krP5jLWACgRphYdATeV3g/QIxChcA4t1deIJIg0Iqj+d6v/EZdcMeEjrZ9z8kyF16IGI1azmeM
gVO1Swja7XA0rbTs1/a3/C5Fw5ktPOhr7ZHad/MafajqW7TReYq/dG1eyEEhZ+PcP3McHqCpNK+r
P/W8MoCXolj+uZLGK19MBYPA/U3zbsMrd+qQ/VrNJMJnJ9Vf5N+C+37ZmdAYoFchWqlkn+8Hs5yk
PmARg6YRVr1m97JVaqYlgzqlVDEjlf9469gD4uKJSXlswPGWCEPczsp8sUuWox8OCydRzxI47iwL
qRYbvvwEIB0mjqANcO2AwY/gRZjIIbxbH7w0sFoxm7IBr27xKhJL/IglkhpMMud/O8eFc37Ezo4u
hAVcVgmdst35S3q9wj4F6kYfOg17gW89XIOxr/7WYjM/2O1kcV+cqmlB+vjeo9VKZEGFw/DeaHLd
/cZHP8TPdj2uZwTxDaYWw+SSverdUKE0gKr7xnsSGoj16opqICrUIbtGMJMavXfzvz/CgVvQ1Qce
Qx5T+4iWwcp+8S0Rx+aJS6tzKmo+kH5sD8ToGdFx5kOCSER8ZLtPTv6p9NeDFg4Y3WlOQxezA0xT
9FUukOqTi+CqxUr/BA0wX+bdIYjDvRXm4PQfU8j/o2o4s1YfhWBZfShmsISTZ1gyirBg79Yhs8Zg
Jw+GsMEvTmq/6d6DCrvAtJc80UfVtyfMPbAklOW/aAxl4qevCwIvEOcQ9uKAvm2r768kF6rjJODh
/MRyV1V/LVhzcQCSJR0jxi6nruPJ1shr59+bFxkZ4kcg8sOhoMMeRPKbdxnypHE6euypZagpLyjw
nDLrTEftIRsq2FBoU4iSOWZjjrhqWjMKL5K+8d2GmEviTVuXcSpPBPRVYKfUroY7R3O9A/pzMPvx
pSN4t06caoedU65ogSkMd2Y3sDDlGzFFah3c4MW7qRNIUtZZ4REXH/O0zg37lpAFm7PoXnAHGHPW
jkufmOq7XCCI/Mbp8X8CBirtY9F8e6yZLcAq/LQ13Bweo3zKjuQT+UG7Bf9NzH7BqOaNYtsCI0a3
3cUJEqsYZ6ITd5tP6hjtvlRiO74aHwP71ImpezwqWPyZUepTjYjTE14EtNJ+Z+ap0EdXMJtYnocL
oXSw6TM9sbmEMDGFqcEOrOj5Z5RwECAJnn/PCUXWidwzvJdTFwK7BG3gFUnMYSaDdNWs6o7PMknV
wS+t3kbgudvZ8ZC+DxJsAq4wvGG21PYHXrYFIjU5XlX3utE73snN4YONX1vYpog/RAoQBVlyT+Oz
wrMtCygr/sd9IgGJzUqdqiXhdwAHBRc/vJj1Eejqm1VRhkMHdKNxYMbnb8Y9BH1MBCc1AxQUj3lw
KxlBPFk3n/ACMnSThm9ia7jTP15MElx8PyLQwrx+BmNg3WRz9ExgZdb6uAhcaXv7cQNRkIxD2FyO
SS6kX71Fc+nS0odTRWrlOqEO8u9wS98vPZdfd4jr++8jfKUrxm0g99h0AXoTbmCk16dygF47F2zt
kwf5XsmHlYpebdSxZ2vEBIyGJ0kGYL8E93gGaRQQaF1qAWbnIH4JrjMIFpZrC9d3URQMK+K3wfYk
shwrZmdOM+bc7T4D3l+s/HheaP7rmuu/hA4HpSsNEu19/CSOkBk8y25Kbje6FuTSraKQKYaDHVSz
qtIT/ACPa1EiUBs4Yidv/KC9oiJUCg7+ToaiyCNkabRHc7BVm5eN2PRSnMdEsTlH438qTPlDnSkU
s9q3s73cCojDVrgtyGmPZYC2ZuvBm24+LBSCan3g9SRNUw9LxeCnJGMAC5PEQoc/0BFYU0513YTR
wU5paVIkZ4krFUoB8yiQAx3BsmwTOVqWSqBKCmuNSuPOrk+c2kyeBj6gQCfNK6TUi2MRjVjYxVr6
5k7huim3Gty/AC6hD9MSWF1SWLazSjiu2Atmnb3gRCH94r4sDUIna/708+pOtDy6EAK/G6NnpJ9s
gl6ph1D2qup1Sc1L9x118+GFBPbF2sL1IAvk/G+pimTbvIZ2XW9Wj8WTsXSYBA0aAsH2QXzVlmZx
pL62JJo46pPcMEblafkp+Bs+zzGLJyh+oq/uxE/esZKbkALOUpoO7OjeU18YTdXSRpyinOJRpNrD
M8tIHdoKpsh65CPqnRcV2y//b5Mai/B3ZEN64s5j2dkQMjDc5MtqbnYpJqY/p635Vv0+Rp58PAjX
uslRyP6ySp/w8wd5R6ZnaRhCsQiQ1PQHLubLBOArx4H1aM6YtHxJLcV1N4x4cq5m97a6DY26oJzO
0kHfa/q3t3a8EaefugmLn4tzvfltwhlFrxObI3M4LPm/Mrc0USor7h1d7gdI4BZLpIJafkVzrVXf
d3k2VGSvLVWoRF5QkbLt4Nnzq/ob/n/2kCNGMMoZ5Qewzt+RsH7CabyFgMVylRbKWw44XtS3P1nX
A9QGQIOJFRL5prnPS8PxmxLKV15XwsMi/IHbaPFMG7GlOY2lbicqgWQ5uu9kwkmiSK8M+M3ra0CT
sS0ZWnXzqmWvRLI2lug9Gm2muhV9LKt3wafo1OQyMjAOvgg4Qo34A3FLgsanH33sURsLBV6P9p6L
ISH8dVdZhJTeWzMhQ7GP4EChzuL3mybT5xgxHwZXV5lNgmALXZ8lS2sZS2QC9L7VTYGzrk4RSDkb
C8Uag/2jEIpTGrFvBMeAZd/di37712UgXFfuMuP+T5gHhCzre+dCkYJkhbuaxlN1TA7ZBdayAbzM
Rh6zVRua/jOCJsvaJMSkJvL5kWDeD1/4DyDfL67miOyutmUTaMYy81ury8NZbORYbYXWcas4LM7y
zmN6aiABIy1t35VDcNuI6Is4vmjWn5uQqr/ZoguPj5eaE1k6lC1EGKay4XSIwmURiYCP7vltlFSx
FBkhpG8Wgk746BbgQM/LaFwPKXqN6sWFNMpo5/z5KiGKdVQs5XJ+xWgRLNgti7ilX6xkmOvtSRMO
+qk1MnA65nBUAOol0LKb/qAafOQKP3WgyN4cxg/SdpPun3Fx0WhIJQO2TVrmETG7eo5NC7/03R8n
jcAw5FLcW3gGNPPodEE1N9IKByMsjun5CK47vcTcZtKxk9exUAZGWfLyXZ43H5T6CKVqLr351BEt
JE5vuf6ugii+OfVv8YFxkugxsQLGqmuPaihme5QIksBGONdi06oSKujoYsj0RN/psQu/DnK9pB9E
4dSIndX8gBURNFEteJaOz0t7cFes4deFXfFhDQXW3QGubf1fsu6ecuZlslwuwnFd4+uKaE0pZrBZ
psu/N2Kf9FWXDZZZeEorPjsicL7MgMUhpF23jGTZhj6DiPKdgZCEHjlz2agI/rgTHUA/QJgQwLzc
+4XfKBHG3xPaeK8vz048H74/1y108GNd7xh/HZFWAvgc/YLZ0Ko3LlOwhBXPhTBn/ktByMAI/sIc
xcUSyifmLxJD2xxR9dK0fpRPLbVISUC6vzwtjAUj+4eXhb2f3JsZNfrl1CI2RK0wuwn+7IjxV1ZJ
yWWH1SsqC18/AZsODdnBpdY7mpY/r7VKSOt+Pr9Y9No9Xpe+B8QnvdrlZaHaUIiBHwki1lJEdaG5
A7zSFEG7D/I3pvUENL61Q+FA623WlrhdfIhXA8r4UMWnb38+4cNV3aY9N498+8jBH9SEOZXZfWoH
uQesJ3BNgjJIg+rKCzvRMAr1MGOmJDT0Na4L3yzUx1aDn7lQ9uL6a1IgLHkeZbJdSnDgg9TqRuMj
zZ+aEYmki+ID0kDpZI1j6LMEdihnqDv6AEecPFJOldQmqgNtQVXhK7girTCidp1wAB8djQDtTIZ5
JBsBlGYGoYg+Xi6SWESMxkDeFVSbFw3oKYqyS17b/jzpJ0jX9fLINfSeoOnSmXdX9wFiuNLI71B6
0xFKb9we7OaJU6aK7NMcXQIVueKiLQKwPo3SL8J5NIEkGdZFDTorYT2rm6GacJyDp+NhjMR2WLUV
YX2HmyduVVl2+8uvrmo0D18o4hPAzmNax2wTrSLEbEwW6XS/SCQWRh0MQTE82/1aL770d4h8ogdB
UrXlQp2vmdQtFRxjt6EzKCOgAyiR+B+O9wReiQ7zYR+ZSOZkeT36tqWYj1pTmiEOUWdTVlSLURCW
oZc1wKkOFAooULIh56J/KVzq5ml0kUXi1bFk3NsBthaB00hMa7gOVZrcLLlTEMvdYyloYKiR1DJk
wroCzD1VvFW8Ofh/DIoB8cvxGyQXTrzlSdLAaEIdtsTa+3R4zSIL38+Vc5IGH6+/ISz+y8/wX2ak
nA4U+nYvHGLWyBgWP1kavTJkonPOB8S86kcKlC6lu1G9uL6/dclOpvmcA9Ksz+ZyQtGeW6BySZM2
5ZdIlXeS+ljdtu2aBwrB4LFGNj6wCG8Gg4+oj+hCIF+woj62Ek3HJQ3k683D/WoqiSuNuB1qHttw
o2eK91sqf0nkesa/7WDWK+YcOWY27exes0UXdzDa1wi+dBEnjPk2N9k+Xr+HBvcRKTg/06vfWYUT
zfGmpJfCqGzpiREnO54QCqMdXoYUeSFpKZPyUlm1UhsKwo6LQEN6/NlT7iQdoPoZcL35bFOLm8mX
iMe8S3AAAAm0+yDkO9AD9VMdxQ9Fr1s3ufOCvbH3Rh/8k56evHIMprqNapvSE8cN6xDXd/WdktqM
+ay3OmNKUxvT7kuZbXdenDfzX830QEqdklFJIjScG1xewEm/VjhXxI7cIKk7y00kfDndL311Hz+s
r+ZcPdWFUWzGO0x7g+EngioxJ7NzDbS55VE7KeTBvCn341+oZaN0npt2lpwxTpb8UeKEt5XO05hS
SlUBpp3LA7sETq4cev34MaqT3AtZnAeUkywySUJEuuv4JSsXAZ1CMDQ4emFn1lQDO9PvgpwUNMRn
soGLCioL5cgCzILLUVqECEZ+xOa3y4I5lxY4yU+t+HnrX5QoMwV6JJSMZIXC2ipMxvhBxYEecBsA
G0hZavHy0RgZGhk3ErTp2qgqQ8r4pDR/UlN5L1whoHA6+xTxSQm0mPwKO+Csp5hGLied0ZzWXoXw
OQK3fBMDPg07q1web0Uj0gEE5OSvdfCuA4/Fqj09bxSNZCoML4jBHoz5YMH94cwJfTUdXfhBV480
u24juguOL+c2XRPnF7thX71LT3xZtDF5CDzg5Ed0ngMZSz4NK31DtSmmlSRYYC5+vPEboVM23+1z
RgSK+lEQgUrM10WYFyDJCwBB3h43Vvw2Gtnd5T2Mh5HUcTfZuIepvY02vwvEfB28JjoDIpIRka+U
1BYKdy1thIcYYOVBy8XSUYJOGri/VB7n+WpBaspWUiX2Fbpq++f2VI8HIxhAvi+sMcDvNQnbOQMy
XEixL4bHvfdQuqOUw/0a7ISC4pob5RiZtnpFalIF/u/a2TtzPCi3l1pVBPYvMVqYdJfRcF/iy13C
nhi9JiMtxl8sfUBVhis3ieCTz1iagCQres5cUqJYB5immIeXZ01RFNA5sWyN3xeXFmbht86C91Ub
Z5NUyu3oXu9Qnanky5esbphXGO2RCZsRRHGiMxSZiDD8KOWu8vGC9Vj+h1BbMcDD9Axhs/44JjQI
yZERa1e5i471DZBthrrQIeqboIjArv2flsKalZ6TXG5LlZP4diGZscvKrzTvYoax/EWW22owS85b
Z2V3bbyyZ2A/GggMgmZuaYyGdF6NZ19H5R3KF7PFm+WbOvNI8XW6XuScBO8GkXtSpZE+c8T00nOd
PrNc8VAkUOlNWJs7VGCgYvbwbvVYNj2ErORm2Uk41qwk37QF+yH2VXmjOs1jnVOuA24j2mX3qeAH
lqE76jLANiAoiVl+CERP4Jq5yySO9GfiTkH9xsEuK8cVM6Y1I8tmvxKs6NHBu7GwtkajpIcVuhMh
DdkiJ4IucxiTykystEqYy8MxSViRGb1Y98IqXK1n1e9+GqRFe187Wli+DLzb12PH6cqfUo3hd3gj
BP+RfQCXy6+6NL0wtrEWR11f7IvkRO5Y+T6syN/1g1CObu8JDrzhiN6v6LinYYLMtyocF+wvdkwj
r1gPiXKUBNhrzWwHXDgYBZUe9ZRVtmt9zGnUCvo2/po/CzlzOTUlqeCkvsTg+zlL2XIVMXy9F272
yhwrLyErbFT8gb11BkQZP2ue8sHoA8Jie8oFjRaqnvCwemgRS1+z0cjRKVHTgIObS24zKh0Z+/km
MfX58EUBHPyQhOEWWcdkb0SDYWKO8ovr5t0sJ8P9ftl2uLkR/Zm3tvkLALvB0G/CK6R9u/Nx/V6g
z3d5GJRsq7WBAONbKi7ZLwRRvY5cVlODMI4s/OVp54VigJCCGoLrVKxWw7JXe8+JdgS0R9dciP74
0JCY774jb8IBP3+IbUGb/xysE5PjAFR7XE2kp0OZpMatPJ0VPnbtLZujB4H1n8dKMbrMw8FqC7oa
nEjuj7sLxzbKBRz5J1rVX3tulVjOL0bdYLtVldiVgmsAeIlr1dvf/4ycQVX8aJbMrcrpE4/1wqAd
dMt9lMvUiVn7PyiBxFUIfeN24MQLa3r71itNrRhEg3jPuqfkc1MDTSeZ2zVhdN2pSCSuykV3gasY
6fjXSv2Uz3EesMVWxOkxLzIDpvVVnQNmqpSfTJJ3pP1+qUcgmZtSqJq1Lj3voyLPJay82LwkHzJT
qQHBwUCTCqaZ4qXODvNVQwy9YgwtV5erJx9F6khG53RnBnlua3yfTf4W3w6aWnIJnMDStNrfRYhY
J4cYfpHIxmBC7yVnbZa3NJBID1op0DHVZz6VQWyFbcFAet3zwHbZB8ibwVCnvHyOedkkGpEtdM3J
1aj3DKTplRryxjmwIPVGx4EsRpJc1bu84Vszz0xTIq0GuEVNRltxipuuYYn9soQazhB398j3e/Zg
CW6plhCYzyypZ3ypa3/Zghm2hfFMrvU9DkXc3L6bbELmw8sn/jdkXFKHV5Bzjazc/Rt+z6YrOQy9
s7aq6athyY+y/Eh6Zbo+WL+4wZVVEIJmmfZyp4yED300+MEl5T+Sb6NrrQJxgzTx7KcB1UoqOjur
ZLMqFfDra3JGyna1MVkij1pkLBkzHbsrgQaAnOwCacLMmdY5bOPD8WCED3fss8iBoX+Cj5KRCcty
qZbu4qrT3w+ikhQyB2gGtyUMEQZyYzEBqo+l2/uHq7lWZqB9LBx4+Cr6h6g0JbazTO34FrPMOY2G
nvK3aCbqOtKbEdfDxhCJZoAhZbWITGq6nHKSV4Av11syOO762BlRiqANpDk8pk4U6VbxfRetO/D+
3D8M6Ld5VM2uF30gqN8hJRXw4AMSAnrnIh4P30xzGi9ZgdLKnLzQw5IIq9d5PnspvkkTVuLo8nen
A5uaBFz/0SobG4THR8jRQBv2tBPTciQGxTijbbbmTQAp7ILnk2sEQ+z1654rvpOGa9pJCzuDsNkF
NAo3EmdO14ZkYTKeUTWVrqC8u1uPMF2cmKqDkCLZUr11thH7B1khItkEucJiZbH2a0j2oU7UiAgP
iAg1wHO0cuQboWDjxeP4VD3HXNdEnHnRoumpgITkhgiPQgNbacAvYGNJv3nZjS/ttuNFPz4WvwWh
azNJVIbp1TlynXoHTjpojCiz9m53h0bQfzy+77i1VZeMypDidqJRIuXCcU5v50AM9QA/NAu7cty9
0WAStmCltdgSDaPrVYeuV6QswyutCjR5DKGVtCAs3LMs3jZ4BiHOLLvOfXvS/0zERlZY8oPYY/l7
sh8kjyemcvGWfM/aSsLh78KWfy1huf0uVNUdb+T3W8D8YKxwp9sR3RWuLqRsESve0tI7wwfHuIOF
bncBpRkmBHfcV9g3C+Ox+4wpI5KUXKJrRL+gXK4G7wC7eqhk8BbHD/nVH1wB+4qijgllanbpsD/r
ieMatfYyYl4XrpEYULybGQirTzePV04+gR8PRe+hLDGVP5op9KdKRXhKfE8bUl/Q8x+g8r1IN+vO
YtiGrIhKI92V4gJlUAI5Cr2oikyH3Xt6iqGN/ti1c8UvHEkPGvKZeDCfpxI4GYpFDRKeDh3uklhL
G81msgS9B/WhDdZz6i4Pe/JZcVyyFgmbXPBDkrIfbPt6Gep+LQHyR4z/XfxA4r3kdx2gSEVI8Lm0
YYWYuj+h6qRwytN3RlPzo2EeaA2WiUMMm/4vyO7SDbZkYHAfrWVDKCme2tEm8cxnYvJDwikQTRAu
9cqQqEflHXccZLU34BVUkXByMPFCM+MDCc4sqLc78yhnFEHdlTIv0afSIxZmIk/3A5gsGFasi1CL
cCFNo1wsvzObnswnO5mq5jkVFteGc3M2ywIpJjGMuu3Q3PMkuItsFHO3/vJ5IqGzS4E3hsOlKUfF
B+R0H08QMcN+YBAQkvK6MmkPcI+lR8bVzcOlq8C4LoW6nihi3UdogyYJ37p0/Et6M96U1zDUefiS
NZDcbrDax7Ul5aeklA1u7WaaBQBdhGB8f1pPIXAkl/1/TnV6U+KUC4LeM8+9C4VXTFNdoSOCX79r
nS8M59Tp6iHXFEXlPIqJO720q43a+xjvhQ59uWC/t0ncddlfn2D3h60BST1R/Mm3al+UKXV51hqI
Z/zsj21RW/Ahl3YqIecAyRkhc+rj+9JYZ7p6UQvTbjs0eUQGloCv9+NdiBeYsNv+GBVm9cRiUTxd
xj3lxwiWA2FJENlCjupGlwMITbgNV8cdQnOFHqfcZSDUvqgofL3s3BJNl86zFGM0HaCbkcatbzBv
IGtUcxmg7kLNyFpJ/cWpc4fytIpYVnZl8URT/9Gfj0hHZfvVj8OVHP9FLkFj2d2u6dtaK2BPwX3y
CiHEsNPQb2YdtKOJph2EaF2p9kxdsTamYUF9hC22xGP2nRV2Nr3mz06pvlgn+jryqE9UhVz9Fq6D
00j8HbIIzPMA9IJSE4vV3LUDqDtB1KCYEMAnjrtF0sV5yFS0XCfVy8beDfyoEHgt+ePU06MQq3g1
ruxqJi/1JDLDn+hSqo4lua792FSp3bzlDUVltaNKDqWlWDzAp4RittUQp9wc7fORxJQozEoSMmKZ
zxfnJ10bLO+hFwC1vXPUcZ2z6bgou6S2tQFKhYj8BubqbXe9qwzGan9Q+4g8lcMfYBYAaWXQEPaX
Xfi0iZmY9dUMdA6MKNin77r3zRZHx5aUbIHpi/zi9GaEe2vjf+WXSArRcrX7ugTHncm4QUy6HcFO
ROPuy7mXakzMJAzcNTogOxRNulShKKPqXVQnT2PA6uMvLF5VuJbQZVb5qLSypyE37+jcu3QawzMu
LOqcnWwhMwLPQt0sQYB+8G52S4mXVgb0wH5S9a6YRQ59F2KCmspA6hvQI9VhnUAdgNq9IQuZwRz2
gbH99wT+kjRxZzOMPxrLvd8qsxJ/MwuKnN4MMiW/gEjxWnoOC3H3ntS5K3+uxYvE88wKaL1nQPXO
B61+KecY7hjuVXx/u/jsnwTz/IOSLvR58mX3H85eK7TCRQdyvb/W+7f9x8uYbyyONpWzfqgbXDTZ
v253TkgJDEL4cCmEZcaFvOMMff0nZktT8MFzxJTOjYk3OHC0KzYMxJ0U8RxIMRWKyNrczY0k0UnX
iLkeU9MzPugYt4TfVzL3Sv3JKj6Zk2xSricwsxIGWhi4aJLzhWIcphRbf3JPFZbDFrOBRXR6uiyv
necPxWSOF2i0Ovi99S2Co2CeA6RPCay/BrMSrNit9x68sC31gj9gntjQCEpNsqgKf8bK+aRk++At
PyDBSC0HNYufgJL8TwL5na7yCcN5l+GxLSuV1n78tiPZIiQWTiJoRo+YeAxs33z0k1TiWCpSR984
o5Ya5kUl0WdL9Pex4OzepWmD6SpfY1IcddgY5f4tXR7JRQQO13XS6WSq4FL4YLzOP8yoF2exMG+E
/RFVORbxr8LtPZcl1LE8+n7tKU4aPwUcPp6RXajuQYKJdDFqwt2W1GYOKgEJ9Y705pOdoge1f3Z0
qd92VM3v9/HIJPCUgkASu5pACXqqt0aBUxltnVwe7zDn8hJ2A8KSMJXOBrVwT4WZQMPPl4xQFPJC
KHffhnoKvxthBedJHAWgtJC28DbZqPjNn5WcYICKyTZWMDgFqpNQ0WxzUP9T6WzJOnI1+1+wniV0
6xM9yslcyXXWk1SdjvKyjVKzSDnEvrTXdl8GKD88FAYFB5b2vgfBUpsNxkLJddE17NOioWMNEiY5
sCIrWqy+amyfSC2obbL6UePr1vDVz3Ofwq2NRnKLSMqd+hWbBCGOw534mGmi5b/TRivzuhybFdF1
RYoSFaOTGybfTw7L9JaCCa4Fet0B8iC7EoVWxK6HAeVcmO0XiIr1g02A7w13VJO7Q01igIWFMucA
PjaflyCkglWhVFxiiY8gwR9VUtHseeeBflpl9fbxccg5CzOM1g5d21m9XvUaW7xftt82HwXO9Tpa
5RRp/HpmIwgBG99L0DqElWz0MgzFt8TlPbDQ9tGHxNx/9OuK6G6DpzXYpoUfK4OYw9vniCkgmPq+
j8Dug5gtTxEJIBGD2ck1RUWY5UPwsAnzemurHxc8b5TmIxfQe1gV/v/qip8rqF5Yb0LNRPEu/rKY
T+G/+0bNABTPfehjt+bwI3Wdj09bTPQL8S8cyj+BSM41odlW8eO4NvMpk8gM3/KwAigQrdZsYtQ8
1oYBcUZJvAb9TdRf45FLKhtrI96zmOupxwMQveiHEZQa3Dm3/qIQaTeN7vo+DhpxP1CwYfY8d1B/
BsWjRRQ0PHIZgS2k0tiRLyGLYdAOErPYXsDeg+6VGRJGaZGMBOQ9vBH1ZOIlRXxAvQ6tkiYRHwpo
olvY/F1JN2aF+rWh/hyPF6gSooO571h16m8kgaX3wg8Az/wrZOCgRgh+4HOG+382orBymywzFo5D
QlBuVydizgY1EGviQu/zB+m0m0aTJ4d175tJiOCNVKIENfZFKTSqFzDZCmUwDBqnPt12kNVcYsRw
VWYZMvfAKJBzGkhVxCrM8J9hTSu9fjIb/9FT/ulCEYomtyr7pNrb/BZRnUDHiqIdWBtQdwpVyKw7
jvbRceiZPkqiH9dKLkXfjC1uL8F0/PJu1qjPRF0dIBMhmDTfFk9/UGCW72BAhysoiL2rxWT+c7sT
93KedXQ5Lcvt+2/MjqUGyUh/lM5NI0Iyo2sYzqznEB5jR7xdzFbe/4PHvRusENK28KAK6mGpPmvU
5AXngUjiuX8j/Zpr/5fMzi5r4iA9g+87pVzAS5krcZ/Hv8GfEFtjUmVsqdsrzW9u2xvCDKidqVq/
T01uBEIcfUB9/0oNaxOjD/fvMIeaQXQqyFuof6qBo7nEPGMDD1pxLAEHWu2BCTE6bLMilaVpmw0t
2kMueCq9WldIaCng+xRANwupuVXaXSNy7clC82WK0hOsRm4zBvK4EcD+HhZeNaOFjivDrT2ReNmD
6r9WmokjEFM6giEJjWyt0T6EckYPBcW69mVDrAgWffOuEaEZbpaanG5eIyerfe+6/Qh8blMDfmgs
J4YqXEWIhpZpwVp677V7hWBwlZiitDN4gDVM5DRiI2BvDoOz51iLhqitWC0tmy9d61lCaDI+zfJt
LPWsw96PsScZEyGtwWvyU7F3omObI7MWtvtckm+ENY9Otz1iupjwPW1bqwahRVkyRsa1+gu/dGEv
QsVlO8c2gqDqufH9FaROZnjbXub1rLKXGPIkB2LijtOBmCf+4cREUaUvdrGnqjlMiMovKQeijDWy
rZHJKqw7/+v2MeMSVeMe7sP1yrb37Z51ylRSM9vTLhYj0FRP5Q0AKFe3dEsE4/GEbVBMljkPUfXj
owMYW+5Rgx5P8lBDOKytKzW6Xt7A5noLbVwvcoPOAvNVb3xcxMLUSA/2NNun1wPI9fNyYke57won
VoqRRiz9MpVkYQMCa3LqbrFaKIgwCT7u1U2fBZiTQ2MezkrzPoNdGZKA24J9AEg3oFUc0avCCWIO
CmkvGr/oLucJ4q5Ef0N2PkroxBJ+8c+nMeV1lk6vIjAl3V/940L+2tFP8Ob6S/c3nLq1UwtDibPD
7MNrNAZx5j7gceEJYCpXxI9EFVBTaYunS1XrBaOQTO/k6yeMYB4Xjx8nHPwoVz0vRisdX5Y6uu67
GEXwr2NuBMjU1b46eQkVXgA1vmX1c4oBSswO9fA21aQnSwJ0asRDVKbSzR0RCcRyg5Tpz1ORjRo8
E6aDBHVtHTWTE6Z4QQlxbWBj/NlM29Ep/ccUebvOrSYuKFoaexkIVfWpCqgMWxlAn8V6CJPViVKQ
Qq78QjBCPacM8QvWHCw5jPV4pfrh2q1ghofINhMI6rQfzwf7/qo2dOh6FKJKG0Tfg4QnorvH5Ll5
0teBYv0011MKXE0tl1EAEI53qKpgeru0/Q2E0YzJcYj/r7fY8k5XjNiiOOhwqQ7h1Xqx5/vYRxo7
2HvKydL931v/avQmBc/PcFsD0gltIc/4DxRhC1PL3RUw7eTwob0W0ZXudp3y7Ca4Bc0fxLo+jofV
E9oUVWB1lXqSGW1fyDqhhxKHPd6lWlPdsINdtmIZpG6s0Xbhr6HwOVc8ruEZo1FckStKR2P62eY0
843b04bWSP2hN5bos4Xd9Th77Kd1tRpEkG6WeZg5UmnQatDun54iEGBgC8XJIX4AKZxr+bmuIY6X
axJWXiNxnMPdmhII5JV718Sc24L4zLsCpx9ryAmG1IAAyLI2hK1CLITa9ZqBTa2rIeNTfWK9m9Z6
fLGAAhYE/OmBvNc9t9K/rfkRUXtirve6vFlgTMcWd1mtOtSwZK4npQZenMuEWGmt0gRbPF1C5qHz
Wz10Y94UHf63g4NsMVO/PQnyK6OkccJaFYL+EVT+0X3b+O6vAbD+vcOZbaSQA37X7aGUGMB9jEdm
NEZgTXH2ldgfdDkd4DV4WFY+GGSRs2rxoWH6tDbyJiVYPCU3yR6BweuwsOzYh3nbNm2o0dtBnUzC
UwIUPOmhCszvjdDsPj6fHjM+WqTsq6aNqZrD60cjYpGVeLALBlopID8oOXFso5l0psw3rcIMpB5p
IhNxAokNyyCT1T34L4M/kbPdhMh39lfscsmuYSHJy4ajuHPZ7/M06VLuu2zueGq9F6RR9hDGcArR
Utr+7Ql+UviZNrfpyBD8RbpDisYMt7+qVo9IJvpuKKc+nIC7HlR1YxpuGRbAFoeiCKksYNNL/6tN
NBV5TDJWrU4U6Lhk3V+7GY+WFneljIvGFYRHXAuu/smTR3Xn4RRSrgpw0RQLO0ebCQLMAenHVzVl
VF7SVfd+utXwq990YEHxdzyBfsr8KYIW6uI0y0h0tpCc8Wl0P19sSQSEw4OymPr7d6Ma7J6Ia4IQ
6sMPQF08QeesdBKBv/HKA2rwXXFl6wdyWQqC64lqFXw1G4m6vO+0vo7IoKr9+nY+hRtKQMYSVH1l
+SS/hEwmlp335SSdGxz1BNGrL4TFuufGhVCWzUWY+Wef8sxM3GwlibpEsDsVmlpVxRnMmNdCqk3Z
WSpPomy4CaKWMxIF1Pg2zs2dBY6eEiiNySSnq2PrQ8p5iO6k0JyfXWJrGNGrWyqawwwCuTVDUSYV
2CVqx82IoGYrgEp7xqMx1db893z/xpRTMmTTzQdM0VHgByWTGtVB/oumGjJXngEwVNLrT43g8+Oq
coIQqzuVaQkS1KjcyS5o4FXN9KM0reyomRfyHDyvPixVsxveHBko/tAt9DF2KTZHsrrHRMhhzYPg
RWQUQdNyQ39hZ0buACgu/ZQWXGOiKuaPAQJwdIqIWntO6/d6NNBtezgqa6KGMSsXxj2LmTiGSovI
wkY4Ogh8P3I6jwb1UZpUxvP9PZqU81GxnlfaTCixPqkqNMKSUaMqPyKhyFqKFMufBv15X/CzHcpk
88ipu2fdeH1xhtnUG+i6SuRTRTqvHuFnwF37k8zYEa0Ngt0lT7yKXo7ICcBlR+mEY3/wpEv5aWX5
b3jNIAxMCOgFxw0WYwhjQsmOIV0MCjcHgptoLwCr4/mU/eBN6rGRntAMwqGcGNY0odNTFt9qSp3A
pQFvfNc2Qp7Ju00Zz1b6J+dtIKuj62SWU7f0NMHC/asXuyALGoefrmYPBuFykYkJFdSLncn0Ywfd
N+G3/vgldiNdZ2qG46On2p9m1lsLcyPmlokwbJ97XwBKQqZyUEXZtMCV6qGtY22iyZxoFUtIHVQy
ft07lWmfu6NkjlV+LJNmlCcPveppThc72QJh8L+VA3M5+1aRg3IUBXXZKUjn5owfHXV4cjVMzk6L
rqaWG/Oz10CfU+Ae+WjgkjVu+t9oAtuzyS8TNA0SPDUDqNYf/ghrnWKz6OtViKLl+6naHoH/mErR
crGLf7Y10Q7YHchcFHRMbPA3KJl6gu7xuRUMmXIG6H+bBvXTmpOJSN//jmkscBuHjtJlVQuv/hrp
cyLbefFUbpRkU+kfLAtD41bfQ1S8uFZRwl17rhLvJw9hOm7S0ooE6+JmUETqz8oC4+JDbuhOhvvo
7ihucO2hmkMdwbBmHQr6iZvyWDvlhVoVOGkuK8/mZ5Ace6BEYoqX/Pk9TsJdLtYG47YygsgrJ9Sl
24dUdKmEu/4ncIANPyiQL3xZR31cBhaoc/kD6uLuNYAJhky0yNLuN4PIZG5D49OG4T9IWZxNv1OT
Bkark/+pjQWZ6Cycn0Pfv/aLz1zX+o4yPO8Iaws71Wymb6jBSeErhNf/HufxPnZCqaBnZWva1iMW
xJMB94PNSGNAN8/5bx3FtMdCAQ5S66zw1fOEGai3Z0YPR2dETlui8faHgAqdEy2kY0yZgMLk+wyX
KOK7LQqDM9uTvnORDkF46a22cK5AoG4zTEIxi79Hw9qEcK4SkvqTtcVb3t5OU8cgJMgxAnALqGi3
0hp7b742pduKfiSmYs5qoTzeTWhKEctC3pz2mFw2nG9ielRZuL4yNa8dkgudrwSwKVBx4JF852w8
9vLw97Kw4m1Jzeu63lusbuRGNFg89Tk0WEuGVdUDlzUOMMUy/CS2mIF20bLxDc72YfeOpAFEEwmm
7FKIbeKnTQtHc1lOWgrBbnY1IpLZtvzF5mKSCU2TwKhHQKg8suN5E2RyreBfcTTXDWpMF41YakNb
5SjbcWldFHYR5Gt5slX8C7HWxJsyGp6Jrio+NXJk8/xLBcQuheb1k6WgUTXOpgeLtbBUf8DmWZg+
c3h5vHnWES5Z6OfhPVLKNcaC0oaMiMjQQgez+KTsFVUnLVKhW7d0bBEkvqfGOsU0tgh9jJGTF9N8
N69yzjy0voGGn8oH8JkUub2UmMKxXHqFi/5Dbn3/OxpbqL9p0pkYEpRUOJJjAyNzp9sccuvkXex2
18QnGqk554lZmvbAjbVGf+5L7SHE0kid8u4CVob0toJAIj+O/VWN8WBaWRNrKLSe15YtkGaPe5Xv
aQWAsZbAZHFP4DywTl2Cu/A1JeFFGszhSIVqMNgp7/66xRfP1UDMNWgIj6WfcnddEXZCN/o69AX0
xjFe/OFx/6n4QUYQuIF8LHtRMdCvEOycsbBh+AEIV45ywKnng76Lk4s0YzWOMSx/dl1NJO+2PSPw
LEW2pNhLX3FAXRN6rbyPrww2VAxyJNDWEJVwINpnQIv1wF7jVSvFdzgBBHPSgRTYJtBaxjMoMs1B
e8Ly2saVOXvSkpJlGSbJcoQWanLS4XV8TTCKs6HdGgvumFF74hrYrayQKgfbvypilQmm9/o/LLeh
5zXcPR9OPgcqrRpiB0kdBwZwR30tWugWODTKYaTvTj8AQxIFhwZh9qdVENokd3CoUfU/cZL0VTCr
SZOdbRvQicX1ZVsNFETcJWnh9k5c8LPbgTywgGvUMy7TrLmiLP4+KFHsiMVzeUvTtnXr9fwOmmOQ
yZeFCK6/F8FIrMNp1Y61pMZy0yIUE2Ahotnj2l1KP6JM8bvADp6yiqndTdaFdnnsUwAYvQJcOC5C
X9gXRXeHC9i22eeg0i4qBtOz82Fhs8Vndvvfiqkz26R9xx0gQ7j+PjT3w1i6kTeLo3eehK3IkEzZ
DcU/2sw9ht8xKKyMaXMxCC54YMWBFfRLkpOFvRrv6debowchzHyoNNqArT3Jl0qlduyD3dTdxTCk
Js+H2X2h0AajBoPcVjuyPCLOcA4kTWRMAfRhQmBqaJWvyvHF/lFSk7ndP1AHf+3xEYnPBmz13RnJ
EmbDCcAJm3hSvMTJr0GJvwxkx1n9hLgOCKZk9oYBl+ZW4eXPAOC2QSll874K6N12KY9/fK8WpDTe
86KRaxDRuaXHu8I0zn9PYDTG9JU1mHesT1kebFHNjLIv44jmP7w3Vu7nERILIocUWlSd9SgJt2wx
84uMCzVGrj5cQIS7c26FgDrmMN0zee8V1xPvmLORLdQ8s+GNned+NjzgT9jJnW0VVWjEJSs+9JI5
xuKuaVMP4jPySMjBiFMsnJzVs477/DfZqFZLxAzDB35NW44yOXNp0bVUv+XHBgoCtPn93TDUHQ8X
fiHQOa+kJ/D85YtYnTVSWGddLBtaAzIOhrO5RkEACL32CTe5oceOVBbsEPPWhtLdeeJoJZwLjVvn
lz55/f6WW9ibe9LtZOjRRSgb7eDKriegSYTMqdGws4c73RcPcwa3Kv0WSa8NZ3f0w6mHNBYNQ9ij
4edfnm5xJd+5pT/jMo/dEPs9wlCssB3qokhLuFV3ibYI0ejbSLYMapTIcMAQyncWVnndv1YlPBPC
LU7kBCb3K7GV0+OYIMGJASXCEXr4NeyZDz+q4woSD4J1SUuPSJ8iS655U9PbYLJOl9HwbAB5Ardx
6Ie6fvSoPzmDqOl1KpzPN4UWXqe+ajhwuYY2rfnBgEyak/QaNlknJR6B6IG6/p6YrnK26EUa1sUS
1v7BlkeTScpt6zFBZ1QS0fWTzJWEXVlbnkH5qzFZ8EjvuZbPAzwyZonu8ep98jtXb4LjAC7ogy2H
Aim8o/p3v1VAS69vgepfat5AzKmr1wQbtCmUS+FpHu61zjjY9nfrEKVI/nqTDb0/xtZ2PcIlvVEG
R6v1s4M+S12HwrW0YfWkqq0TbWL0ZBIxT1QNflXTdvCTMHkrEBzYsaPjAXoYUrFbjiSkLOhfBBvX
PrxV/qjMPhSACaZFFryXEFzEHSGyw6TgHy+SUwdzulz88Lf/uA26GAAgjc5K0j4IENTixQNNs03Y
rFJuQZX3BXTAjfMiH2iAozmYrXA8duHS+d/3XQGnIDKrdPAkohmglVfoyJnxRqUm+nznv3oQqJvR
KUcRsYTJAndOUswZ/O7wuTlFUKdJwx6Ed+KGjipnP4R+VAD3xOv/Wzbtd6FS75Gnoq380juV7q/g
Xipvk0b64uJvGcV2bH8F3wGZFU4OaHnLFct9DlTUu8rXuh3hPjWpStmwzcFsh1f9TtaIMKT1I6Up
Dhd1kFPyLPZ9EnGgm5qevJ3lQoFrGuM7rx1LR/2Ua7WHlRI8oOsAr9VdM3khP2UqINOpZAwhgpB9
P6VZiYBJazGw2IirQWqrd7Y0OVn+R6d6qI4VPZE/8FZ2lEvCI+SrIoBKH65v8/HYgDfeA33X9gru
r9oZsqvJRBEhOtg1izmLqDo4ZKnviZEViXfnzi3QKZHd5ssCpH6OwHPdhxCRwslmecp4CEzqgCDL
7TOm1aiGRYlWiSJaGp4rJf6xXT+7nBktGKDB9vYTHlXW0NXOUwlKzNsepHasHehSxTcTwvA9d7wu
et3gdhf3ngGNSGDDr/7DXTXvZ23tZQVLIJK6HoJ9ZMUobFJ9JoY1HVgbmYsK5CoSj6xKGb/oCyC9
63ja3hXjgGyxGUCwQYbHxL25JVp0m8puDkTdFP0LiuqerER3QY5HEZoJfCb7P+ehdmlm2YxgO/+p
Gio7OdiT1nalTj55RZQKAB+CgBZotCWwa+80DB/Tmv2YWlPmPd4AidVgaS5xIPRuJaa6t7rtTqoG
fsRQRT+l/EEQSaV80clGhxDDPIMVTSGXl83+1QSq4UYSN5a7ShO5+T2DFiXE9TYEY0B82s43Ysdg
gb2w8/Uy9CLnICTEemLuPw3DH3Rd+MuSeJgp1k9q6GtJfPdTg/LlywM/pPzutqB6x+CYcHcaVoA+
RjXNU4XEMJW7QnULj0Py0vZwW2A44AMqWv2WqGsbmTuwBdsYubJxuzBKORhxGTYahGgbMS9qMj1j
bLFVdsfObkhHQsit9ZLCoqCvYo4NxJCLV4yyrKJnGEQbBnJ7nt8D6be6NIH/IPQ160o0cmCzg8br
DhnFfduTaGOOLaB1hjBipHroemn1T+Qz6OhH9/D872z/mFTJNGgCI+SRmrBYelrDT/HGFAgDrA2q
D55tQ/LtKGCeFtq2cMXpZgzHSail6EtsxGEZRqUEiBT0kcAV6CbK6HaD0P2gYmiGRxtJuUK3+iIt
s35QF8Fjy+MCaWoK0a8H3Z2DI6uKBts8Ex0nj9xI6pWOdEpDxe/iP9ZVQLEYRKU0jHaKaeb6RSs0
ieRDuH9DpM15AZLXPxNLQ3vPt4RgX/RJShVruy2kgMujIla09chFpXrGI/ko6m3S8+YK03Tptj6y
cDKdPVMVndwJwypljOAUhsaq5R/fnkhEAXkg2JliJq9DbVZ1ouIvUAzsw9Rcy+kPuDW59PvOkRLR
lun7eTPRwHh8ujJqni1mU3yEpR0o8K1KMEVqdg8GICFe1y6Xzl8xLULPK2Q+H3/RmbhjeDmlW/dl
rOe/I5XUy/nHHycBbDBN6c/44TO0pPcTgP5/GG9YxK2IgPrOk+2RS4AL8z3JAk4obPolP4D6pb7l
JLdK5wG1kT7pvBXu6GL6barN6H1cPTkmnfSjwiinMuYq5XorMCnLBjhpnYUNWb6dEi4J0IfPC+3e
ysHyN/RiF2c5fo/ebPFF/MqwHzB5cDqBuv/Q8PYxgfgaY96gIj7yxUJUofQ3p0PKbKJpzHT5u5Dp
MUMtHNShfWv1molEOAc0AHQWwxK6vG/GfoOMg/1skDeLDXjYJRRqk+83e13sSZIq4jHtICG1vGG7
utJQkyUwo+/zHaFfJwrzuzAjxiDoPg1ZmiH6u6jfpp411Qdl8HOSWB9Nz3M4Ldu5bx/exXOEGfjF
79UK+Tk5E3GYwgUi/8A4TStxIUQufByk5NHFEwKIEwe6mc7V/BGAaLPN2Zvtw2qfPjzgi80DbPH8
S/GrQrFzyZA2nlRnE/RYhhOlA2K+3NtKzpu0GZ8pnZncW95ORm8pKHFBsge9IRKkvkRX0h7CChIO
tAfZrJmdlgDqZk5j9ofbZRFZlp0PxVose9HK994vni0wXbrQ5XPTFPWA2FUR8fMZfW6igTxgCR6b
OmQghTJx7/RjVoX7tPqFIkmNsnJc7yHyiQo/xLhBLZl3jjd3jvYVb5UgwVJVNvaqIg4g3FM7f2dw
vnwPCYekFG0K+ouq0Ldvq+SPGuB4M+IC1b7yVNuCcAPuQDOLcH9oc7P4wnbB0UiFYIiTL2TmzJos
06I4+170pAYSXkDJTC83KPn1Nb26Ixw1iV2AhIhQTPoGQvV7LJTy77ZB72l2X/41lGzB0kopbcQF
PjBMXhfLmq5zKObhraYKbbJLTX+MRpas1F1qK3Xz0RuqV6xIgeAu6sCqEUHWNQsJEqiGxNnMl61+
//w9GKLMwD0/BUNdWKDU5S2KL36iT3VJ6S1EBqoq8tClqPiFZam0FCY97ktSS/jUwIUcjuQ4q5yz
NErCjTVuC96TTZAQiVTqjtCgQPFykchk40Kyb8uGWIezjRgFpTvgeN4i9UMO0UDkk9gRAAjzXfm6
rb6v+fZ/suQXuYBn5wVI2uro+3ZJxy4aW5ioPu2rTdmiT6nTprJJPGXr1OsUU2Gmg9FOx8BKboXY
+sq703uNogW1EfeaGaEh6z3UR+/zIvp/m0qUxQRV7ZO4/f/6VMfEV7oeZJS7YR4vBzGMkCwceiLJ
0pCV++j52v7ofbjK3AVnjKUWpjOGil+NnW+v3RAujyBrNw6R7dGegwxtP7Qi6dMrrcOB9I14hURX
L7vCqHpHbJQVhY8+K+drEsq7Hn3BxE9tYpPMmLH8Iim9VMQ+D6HYCsdD1vkokcJBvfaCAKL39AIn
T/Jik4VuPpo6DB1NRz+v4gh20wohOMPUy2/2SSJWv9JDlAn+WXgiQv0qHm9A72EbDBGx+BOz3KdB
CKfDTLlnyGbudOOtrxOtLh6cv0A9bAtvZmV/h2EqtCUVDzSq0ZZHVWNTaqUW9eDyP4lImxV4Vflf
F3w/oj0dlhCnFx3FeVucTohxXAPqX0/FFVXPXUvpph35KAzD9fB6d6n6vSI6IzTbhqxDIgDsJHlx
QWgC9XPSctOO/u3tMnu3lwu/f6oP9g37wbLqosw02AFzyI0kLdYZTuYULCX9qgsc6BhQFVeoDT8q
8dwHnMrWCiwwQNr6qIyjmFaCu9rF0RxS1y4uZSBo8YK5kidaumsWtaxtEU+fKEf7vnNrhandoESX
Mkt3uKrhZEaRMXTA75QQyq4qwNatvrPYYw3KfffF8o5quny/yBsPKtumtDvYW4QUxz7mocf1l1uC
5EbHgroNgiSSJCGI33O3ggFH0VtpNOZAcbVZ7bovW+oEk4WU4R1DnETaVBOZMV//OXDEbFdTrBnU
1MAu+3YNG/stMY7brbBi/b/h/xd2AwO/QUfqagM6OCWgld20iUph5VXvgGjSOeY7CJVXbLXXAMs8
Ml7C0C8msEaUHzyJQjPhxH4TtudqfJDbc34udTeAXgn0W4mYDlqP6kBgltUN8N7u+97IbNLbfA==
`protect end_protected
