`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OcvYd5i0BcKeWB/Jp7nnNElW4m5b6NeYExc0Bwhjzp0FEC1Bh5YNMJ/JK1EKaBwH7+Ish06Dsccs
JkSXdGML1A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/UjyAM0GBjGiZFYR89t4uZo9uyf8umitBYRNI2RNuveuiL6SoMIrSXFVzCPTq1wz3UIKZHuMDcn
t9K4nwVnfoojlNoIB8QzPBfcfs07YR0tOMWu1zNwi2SNyTGPbqbbBlnoPf9QxUV5KFZWWP3AaQ4u
A2Hsf08+3sBH3itm480=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nlFFAJaPniMh72vyWFgO+S+GMy707MUAvORFUP8hgAblTDJq4v3E+DBxlyzYCKJq+CQtrOUn4asq
dydlBNdOo//bNpjGacC4H/lO3WbIs5qBbdYgFmXOWuPaQDZKa1zAnLgFo6gwTZYux0Eyce1qpO8Q
e3N9M3PIASrkRYE8lZIcghBs0DRsqSCkdX07zmogKIoSNzeZocfr3q6REi2TvjyAPN+pveeltSWZ
b5QFuBO43G5CO5S2oYzaXTt9fsLs/iHJKHGoF82HWx19M5fDajQJGrnssrcSB9Dv2/UAnSd7UwFM
HSHhCHR5BPJLXNZ8OW4cHpnr3XMSIlXn7f33Ow==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qIff327NTNs08x5xtfB4R7EYUcKpPpkHncae9xEsfgWhQ+Lg2CEV09OZXvIa9XDwWBtWmdxd+WdN
aIFjt5FRUGLcXr3K9k9EYpbDftjhwuN+v8cbZW5TVJFVy8Lq40bL5Hi+TBCJcRgUJx/r6UGP+Zhq
1iRegRw9P3oFsr2j6vE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qRUL7l1F7/yBshvPneLXPL+TQcMvMDzs15L3qdQ1ylp07VeTLJspX8TapU+nI0+WlDf17rMDysSe
yJweoxo8GMGEMTBv+DsEpEPX3uxzV6OCAdofPdnxycff7CJXo+t1mHteo0YSIUJiuTG2iT9rmCgd
TE31vL4Va7NANbP6CCDCSZcNsho62mWXco7u1qy2H5sxa14xH51EAFaCUbma9fd50KU9JCFdCRcK
j6ngw3TD8nqdb4/ZJ9kJ6iitmDayuv/umjz+yGXnV/VjHczkxlc02C/gObytf7vYFdsohzpy8kbz
EGdRxPGgVZTJOBa8c3mSMpv4fWVIH+WcxgyH2w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`protect data_block
cQ/94dxCXVWcV+humrKVAscEajdM3xL0w3xtQLzqMo268AU4vU0esJTjeDRx/n5iM5ZCmZQK9E/p
yMAt39FgRmsctO3h5zugg4CC7GI5hpqwaiV1lK3z3RlRMQTFuU7BzH5k++EU87+v6d86rUDYqg6U
75VLQxPzDjNAKH6XCdxbeEy75a9KCcrsW+YVUW4KG9DparbZ0PtojjaZ6dya+X+Lb2EBMQvhD7Sd
3IqE6XKPGwMD7AISblL/UpxlQgruae9lSQiT/8E98Xc+9Bww6oQCzPx1yK3N0UAb87LaMIdgAWpE
ah+wy56Z3WpmmU2BywtIDfDCRjabb24vgeGqyOpx90BI1+qkMUm0AKqOcgxZQGTqOWPYhoUlVdTI
5o9PpErR7HpJj+URJpviDs1U9ZGakvpY9h91RHJWJTrg1VS77NsjMNUKmESWUTVFnKwwiwOxfH9n
sIeHGCInNWKhVEyv78EOcaBALt3f7fkKArf9MmRFz01ur/2NzYjoZWP4VuCuA6eUPEZaY7skFO31
IaK/HV/7krsTXYleq4wvFTkth30EanSPoG2Xa8oogT1xrKKynCr+KSS1LB7D+ql+98huWhbX8q9k
AB67hDtwaEciEYyf+bgdbSNDQ7kEpJoIcFCW4YOeMhsF8JZQpz8T+9P6dYkAkdt5Jj3OC4i1hrNR
NFM2ZDOa6BmwwiDseD+ecI/d9TkJy9B5QwhcLBsepzAV13RBiBsR5lttDQzKCODWeVaeAn6jJGwP
W+YFzRGha4cberOL8jG/gCFAye/1FR052R2uG5luNB8myiQWegCI3QRxfNpNHNS1GYFhEwPOD29C
XHxc5hY7UG/5j+kdgZubk0bB/qVAQG8NxDzP9G626EmESQ9JRT6eL9p0nzsRXUvpqKb+GUq4DH75
+YualUaWYxcLnSDAGbRNqk+xSD4e10KG2NdcuqZY6hN8iBtY2mv0hQkTTAYIaS4vxRWg1neHrLAg
gkhSZMsTCr52Lv2WJ9K5rbwbjLC+vAKY7ysp1I0jrzgA6ftOZOtf9VtSE2WSanlBK/7xFJN5emj3
PPNK0oF8XloIjoQ4bsDlUBccCgY9bWTaf3aYqLwMgqt6YR7uprnXuaWkR03HBeA/HEq1tTgUQZcX
nWQIzCWUnlEp1Q4KmqbvZK1IGBu1BowlxfYD2eN0+y0IaTPF9SoylDxN59JHPEBB58xXo1HQMvkL
bA7ds6qeX998EBMu2SwD9e4+YDQVbhI1jU90e5oRTC04IAYJO6kJUL333NvqKXtk7KKJF2Y9MMBY
APK2swt1BGUxPXG1scj65PNClDucugjevE23eagAoqdkwDP4HMj7146w45w1AbFkg5aDIBvJs7XV
Ll4dOEl7BlvsXRu0wML7ADl1cvJBMpkSYCSxak6a26nSuw6SnistRsxRRrBrVkPsgLGyJAvkuSec
tavXDaO/iUQHeVvvNARCTZzTVhVntnTBnc9FTeDyuME45fjetvmL8WwjuISfqcDmK6HxSvELzyuG
YwcHToEvnua8wbQQ7kB8fbRFhbSytjUqEASAdmXrGJb7tP+hV4/NB8aeh1/3tl+LLtmLgeM91sdh
H23BMaaAZ6LsyZBE46/8CEN1+6eGA7ByXV8g/bSScrs5nuj6plXYCvmT5m528D+fsTGW+giiT7gT
bR8Bqa/wIoyvEAMEZqrodl56KaW+uPcYvg1uulB1PwEmxGM++6sN8Dm1Yzgzyl4QvVuS5LcwtNCI
yEnPwz/J7NvpzMb+4tEgBBex0PQ3MauYOH4xPqR+31XHIx3FkGqFTwnU8hZD+3XIdHCkaa1u1TVO
mIvzhF3pHtLaGp0WeflsPg6zGlJhT7mIg0Fnlc470gK1Te2gtnjEh9RWNxxBgcEsMot9fc2UQ32/
vcNz4lCA/kV76mHazIAwBvX6nzsEfFsGlqPzrf4CflQLBRUInLw/uLwP/3T8KEkRDVKfKQmXut0X
HlrHdWvbIZ0t3yGIaaSVP6Z648CsBFPwXxjaSWuPd3kGqppg1D9JqbxkE6mzUOdVbyhOWM6hH77i
9tnLN+Q+4QSVNOVeCgd/1uctc5fi/4oc1wUq1XKOqcDHBp4WKotWnCJvlvRKC124dKmsPGJcaWG5
VgawvHbwy3OqckSoPH3qnvsszK5pbxvaR0XtMJVQojShJavdBEInzvDDkA1erlrCgc/YKv8UEA2r
iotb4zCbwKj+LlAI5RoVhJtHfN1ne0rZXJDv3l33eZU3WTZZf4+ukHzT/SbzEIvSo3eyvfgQliaQ
SsyOXLExFOtr0eJKZDZD2hlq9ELOdn6bp9OEsEapyNP9iRxRzuEIibkFGyjmGEnYZ7O+oEg6xlb3
7wMqViWLchmlyABWun4Fx6QFdFovl+ZXY4900OouMtr46xjCJLK3NauNLOclamZY2ILA7hHzD36H
CbARM+9oFA0wu2lix4Z3p4UVlCD5BAFvjkkBn0eUgNKQviE64LQiQMJyz0rHLHt93Bt1uxEWvDD2
S1CEAtcHH3jfYxVtKvXJguH3Yqk5UU3bxRxe9YHvQO7xX98OLokj9vcFUd1/4mMSTJU0McfkcoD3
1q/Q6QwXVuVWABV4cNNF0lLZFJrHxf0R0vhMLiLNGHe8e/hf+mrMvY6cS5H1dFIR02HV8CaqXh9I
xsHRjD6hEcNPT8zo3kGwAzn7Ly/NGEZB2QI0LSJGHMI2ME7h+pMc/iQ1nxsBLJRynWlaGs+cxyli
Bb9Uab/MHL7KxythPAEv3tR0o3g6AbzArYZWD8sZRnq8opUOQLQ1h8rBMlCf5NsDpDikJjdJ7BQH
5V8JCUAvu0mzAKWn4nSLgzy1fz4lK8phSFmFRNOGVu+OF1DO1bJpeD71niddcstzFzcYp+vescYk
zwHTLu25CcomD/LTXuwvujsHXksDTVJcNyj7L66xx8ymV6CsCUuck37XZx+6NjCL8LMXfl6oa9ct
eHwREJvyGtQVDH88ymKYnNPhEzUmBxpXzDx0AH5kEBlFhm0X+2g3Lbx7JnDaq/miR0o04F7nva5f
h00uodwPurpOI6EolSHQLuh/oePrG3BFRdtIzkFbNVmjZqjBGwWMWZpHmS4OCHK7YNQcfAZ7BFyH
mPBPJ92LLR6byrGTGUX0OdReNORU8FXuMbKI5v6ooYkGnMRjVvBP43nA1vaE/aRsJjJl0rZ7EYHN
1f7waqJ7e8w6kV3M2aENzO3poEB4L/P6HjRIPphzw51fhuk7AftNy0gVoKmyLVoaWcIU+2fPbRwy
Sq25i0liNgHC1/lXN0EPwlWbeaN+YP/evu66LdIFJ5J4YXRWxQb/RtN/aY9r1y1p6sqMvn8xXF+M
LFKA4dvOCaDMWKmBC3CZ6m3y+1S7FTK5ltlsKfxQI5g9sLtnlSpXVS+oUI1C6fKvdSA2qatQ2bYq
BGnqZiB61EuCwZjOKjM+WMsiwg4qT5ra/mWuTSu0H2qUKHpkJqZ8eVyCtpORHPTgJ6uuRs1Cl+gF
VZvJpUr1oleCJJ+zjkfh9aKNQE4o0h/tbUpqg1RUtbQjTTxnixiuDxnWBkFuRniCwsdZOXkqxxKY
uUD0AGXaVJeleEPzjNvppLnaZgRpAu1+D3Y0QcdqIuECOdroj4sqynmS3Gdnrn6kYGRKwlyOnLhM
Pm+J40YgAbICTNn7gbME74r8kwky/WSlzxR4eMyXNt3F8g32dqh/K70SBehGnaMedZbWbzFwpcEW
WPzxu7J5nUgy0XlYpMEbjUBkETjg+vGlfd0ZhgKP0eNuYY5oBH7keH4N50kkruRX9EEqWf4Iwzij
4eZGfR2h9irDuiSMveh44UXsGrpELF4jiUzT2ZbWZ6gLPqpEfi/C+ZOlxXTtE0UYn56Waxj/qUgh
HTwoVSD83p4VlH+QCd/ioEczbfAe6qSaEZpaakbqy8t/IY3dfpJiLQ96F1G0suM9nP0xyrFBnl1o
1f+PRwqRDqgAdYgx0xf1D1vcRYMp5uTRKQ6sfprESX+w2yVOIhoJJ+tDAPQF9cebRIx9cjmwO+hA
JIgAKVefIvsE+pEZzq/6cDt0M/eqTkvIOziQEzzlfbpR0Dp81VCsOUafptQ5YmDFf50FF/pPyS9L
dN1mPNoO98R4pazIs1qVn6paGKGQAX2EZY7Df4Lu6lMehJDedylEpRsLj0buK2CNNUOmNSRuGTkY
SA9zxiiYMGE1kXctw7kNC4J6kMOJ5hzUklT+hCoxfpQa+hq6TwJ0Qw8f/17+9vmRgtl/wxBGFUcp
SFW67CB7q/xnQSPi54QSpqutIYP4/iW7/LGYlgpEZpYJKkNJKGIeyqDpjl4vCd1nInGaXFKZLhpl
tRqKAbZPKIuq/9WX3jMHJVHNbi5mUYWJHclBLiVPT3J+qABNZRDCyHSZe1vCuZxN2BUL9c6GJgQ1
I+vJhi7IvM5khX5aOJAk+uJgDGWBS62Amj/5BlmNF9CCYPhjr+kwgJQm3KD/yMixdPRGcl/tqXLE
fcqiiOQMCOQ5DpbF+d1dGsPh1xzzPPEvMyzAqwbD5qB6cN92RmH9kEFidRyOtmjekOoIHfTMcrdl
StEcjJusbUnP4AE9K4ASAs3vcuzahdt2rhTTdiUgFOgYB+QtpGichdTwwe9ECjSaGfP0YySK7qUz
x9PXrC/aPiN9IXPcRbFvDGEWLNnJTyobSTQPcvXBQOtpP5RZOZo0OfH6P4jBtXfrZejcWYcuOtAz
w/w3fBDEek3rlbaJK0WpzKlYO0+DK6HS0XLYfpKmVBZSzP/wq36I2HL8FIZtsT6w68H6NpaGstET
Xy+cyZ0IDNhVVrVShWbqOjNGdrOOd5IlXiQuDsEh2TQD9gJoFPMtBRkF/R0DFMCH7Q06zBk2iosI
y3p1gqGpG6GI6Y/klHD/zYqTDKEi/Qv3M7ZRXI1HPjJ8v4iQJPei1FX/4eneiiKmy0Ykll6vfu6H
QfA+zljI24J/SpiXjuk4XemWmh8ARQSfB1dHMoh8Wau4+0lFRoBDL82p6XjCoE86rdMPRO3Ddyj1
IMN7LGjUVAJq3nfERjq5kzd75aXPLxwZMXNkbgakVVJl2h0a/EEffXBie5bywT8re7zHN62IoCi0
Ult1ugWc9OxsmhR7DIe0rUl8MvFhxmRJ9Q7u/L1EtEPHUydLt8KGsTv0HmUCEk5FdwxYl0c+rAt/
6V4IHK2sqvy5M5cxWrzbjfnMqJ7SPIy46HWnqRxCqOah5T5nivdN66R1zm0Y8sqOEewld7wjatMN
ZfHyXyvpS6vhnnF+8jov1wKOyoRbH7RBtmrkyso6MTOVjG2x09VMb8581pdc+Qqq/7A/v1PLapdM
3UgncfPgievP0GO5DfjMmKac13QpDDmjO4M4Zkmz2P/KdGw4d5pBnv7xUZI50dfv9RGyKrYKT18Z
pE3Eyk2SqOeU9Qdv1XwM22wLfqS8pKHxITMgdX4a2b0G9TWwnaS6hdrzmvUW2PjYKWOuDDS3Vk9a
DX7ZIvCU3IKPLXxCdOh/KS3KwnROo5d1EBaPvqs0yC8+IXDxEqaepIjs5Lf7unVUIf5mQQs3GTjp
snT7hi6tiiE8HxtLxg4f2gzKFRAV0+AfIWFZv6MxDCtc2jV5abKk5PD9ebUjFxbtmDo+cEBL87fK
N/Y8hcpCNQ0QIQ4MO6zGYk+Lv0q2yKbPSKsbcvUa7KWZAizi1paqptzR4DGZZkrPhmtkrzvxLZ8r
i2Y2LzBr9WmVr/2gYCvcDRMRQphNbZIYQKeFMeiuEVme6a/526XPs8P2I3VCfXRWKVTb1CFKmxoe
86RytYAtCvmbgbia/n1LzubVILpw/ujhe5uEv49ah7pXA+NPr1SdtnUBVxJpMu2W4MBBjrLHs5zS
Y9ARRoB2x2QV5xYHkVoChAUyPe9dwcfJHb5QXlBi4Ty6F7r+httzhwR9Q/OqOPVyfwHRfXHhgDLa
IvdpEY+n+YqwOIjJk3pCm5voaMvKnji630bS1xvN2QbEg3hQq4cUrgKgPONbHNQl10kHlwOO1b7u
UfOvqqWkW5ZEpiuk2rzUxbl5yqbyYHB/vDlTC1FR0Km5tKHWbJNHojRkdzlhHIsRRXgQCXaH/TxK
l2+BPxQ7YRs4B+SpgTmOFQ7i/1/Vzde+XrW6YAJ5ESw5aKudPloRh+D2lJzothbbp/XvvplKXAAk
RrYvbc0GPkFGoViv2E/c4aMgWsEosAYFPqPkiZs+0IgvnNpCVok4mGqV3wMVQjj3daAge1n9+WWB
yhSAbGds0GmFBDQ+RTNvxWO+pw5Z3HwYCWkta+B0PonjY1hnuq8gZWjpcMxb/35a1lpYMZyMhVRp
8uXbK7W0M8QfuLUFKmoz2hBhsaxkMT7qTp6uBGvBDOQM8hpA3D/kGnJqafYLEpK0nPjoAajBUlLc
KAMIpEdpXnR+6groQIAMviQ6UpJPBAeYJgmrcJ1TxnrzbxEknXJ+wU01+no2svywXOqgV0ieGbrq
xdIvuN9hX1jPx2fIiYvQAuf4SSsifObJNpmT4Bft17hdjrcRsTNedxm3X8B3fL3hRyvPRyXhs22b
CWYCkmocISnSNvx3XWlBtveznLNxlW5lfFaOF5QaMdPeMei0swSuwMwy1V+f/ZLv5xgkq3VB+otI
+1Jx/al+F3ZrXn2n3pPpjGiq/qHv21p2cDvT5dmFwJZ1fGmXmV4enlT92Zinu0f4T6n78JegqXaR
nhvlJvsPL4aSB18VxQA0BsWE5fWurkqCUE50pl9oMXL6PSt0jVWrh1GQYGtXkNQkwfCNxfEDU/eA
hc2HQMfauAR4IUUDVDmxZwUf6aPuofOaM4qEFuRcS3gusWoMBA3SNfYGFVYJAJorp72jj/Ac6SS9
dvYwswh/MQiAoPoHqvf3YO2spZKUn4NTRdnn2bVMnsSFFyDAD0SImHQhZYYFKqIEXH7Iqh9TkPag
8oCt60aWRIqOeBa305lUA4LZ7OfXiCQwlD5aZGx7OhDfzS5gNCnQ5hKmrlAIHexjBXIZDbkAVz3+
j9KrUJLGd3lYYHfXoCWrOW06A1ukoMsl5ss5peis6/ZeTWZy5eJ+b8+xJmvrVZz7/T2a+GfYh+a3
/4RuGGxOSLgKOZ0Gv8cPD6v8kbarFSR2z6MRw+eft+Y889a1J7Olo/WDZdBkdexFfVjM3hunzTYQ
0pvZM/bnNK7Pw9HfdlfY3LA0Hi3R6cE2FJ78WnzZFo26XDP/PrP2SqSPczIeVauPImlfTdGbwnDr
K7Z3YmL+3qgcYROiSUdYIhRWMbsCmEKpBos8Uo48NLgUC2+aeCERO+RkvXcxv/Ou+lS5CDUkgN32
lbFucx7vO/h71ZU7p8f9Ud/eDq3EvxXGt9DMwWBOHCqU1dLK0ZLu08ytYbmE3EEF0y1/aYT5co0g
oDnBIclgEEWmvniddP2RvCeNfIFiz1SwcjSYZ57P79jfF9E9wMYDMY5EM7wh5toEcnlqREI+jt2I
PK0tcotZwlRec8KahrBrkHJW5grp4u8ud0Qn01AnMgddrUoGQRe1PSQtg/+PeVcqNUp/dftp0O/H
25CosH19pttIY8fLtKM5Vj9VAN0q8sT5NFxV9DrqYFAbGhXMWr8mgAKm/adZisj1ofp7NGJeY4DG
61H/ZbSCmRaBsbQX8+NRZbF1pXUMOYiuxjXycbIFwaCeijqzEONjgrqOFzlGeaoZ8LZXg6MIayof
GVGedWA+7M8KgJKNbeCVJ+/Pn3pTLIEzgdvpq+z8pww7pdr7qD74key4q+rG1CxjFCLi9oLxqwYV
f34Hzvys/A2LAqgMBTMrJhl9gI7fD/QVFUrm9FG/tNvzIpjOo4/V/IRigbirurs/b2HzrKJA/2TK
YUe6gKK3uEd6uc407BAvPuulcpUBHkroPKbfLkxeg8flFKA6kZc5Kflh2B8iUVC7dJKduY5po7nM
vGih4vl+VLa/CdoSZuv7uF2fpi2mnODte5bQUC1D0xoIw2sFPtXoHo5GV8uu0wZuJR9NNLrhLLhH
oQwWdE+gmR/SyJ6rR1Pn4OOmCpD/g4S6ZcGniPK3P4GgJRGcEZhKmX1yDJAEc1BQEAfadZDk7FyI
rocUyDaVSWDM8lhksqyz/2XwwRNaKwpRrE+7rTjcEBnAwro8bD+V+NjrYbDd8MVX472x7keCdPqv
8fFQo78Ybo0eIM4q1OTJYzmNHYl9H1s/cBEmeeSwxMij5iut/KVDSNxjq47Bzq7KhRBNwbn7Itkq
ducZth2uoQYKmZnqzi3z2v8zsx0E8CZjnQblwlEm1+KVtetPDVrXlkH3AYjwfBQp0oayKykBXx59
w/pyAYyixscUB7izmjkCgOOujbVlt6SZffb/EjvKgDMXYy+G4cjWtigrPKR2gMm1Yl925oqha0mg
+r+Fvh5Iy2W1W66LGyvsPr9hQqOxExHzYmx2/mekqyODKQ==
`protect end_protected
