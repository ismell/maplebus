`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
X9tqRM1Ldp3veD5JR6nib/Yah7rNuzujWVoEJ/KsnuK+H3a3VbjPwpRdvRjGEEncOkQuCMKvc1Rz
qN/qA11OFw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PoeesUIChM6pr56WGy27Ub94whBuJL8D1tA0f7JuZwGYyEMs06k5StsVd0EoEKG7z1AGJ+tg0B2T
kzQ0c7+n+ZJ2P/bRGyu514RCetYFq3UF8Mv6vrJYj/Pgk+aaYtPaz1H5+KNAOGQOCQuoanvrrXDy
JUg5vbMZL4tpy3r5n5g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lqTssHZksaYsGTxPtHCnsfkKAf/ogIUdNmDA6xEB3w5vibYgk0/dSpi6IDDPdvjkRXP/u+1yrm16
+YPK3caH67BdQxujJde/5wqOxELwT03TerxDcl/90UZeVOr8OhM+hKu49ond9B4/iSmu3s1tXXnL
ti+c3hkm0k8aNzuxPYM90Q55P105XIeSzaajLMinx9SpmAXG4q+Ejh+WwVK10qmLtb0jWMFZjRw7
RJZeiiZ/ZEm/jewKU3km+vZlNVyJQqvP6atgv8diGGekUTTfOSuDYD9SERNxR62a7r0TgN63tVrf
ihRf13doegqFKtUuOfO+L1z14sO0VdlFzyCohw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3n0mKG+c8a5rAfH38kljmv0sHJu9mH4qK1bFANq+x3cPePHohsazGbxedmTfsLxvQv66PmA/LvIh
4Dr01v/9QM3+zV4pWHls3DfTgpqMPa6kTqLB77SOqEVCZm3lKvNzrCMTRfxX9/24zyPOLCwcZz9K
Fdg7fJ853OwdI6iwuv0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dLJfzkou4RwNfYaZ96WPGKCHnbE04rtkw0l85srAPggz9EJ7X/Y9m77gcc/iUVsRyhXfDLiNjY/u
kozxXMDckZLER3RPrWtjxORYqQnFO5HbnV3CZYhcpiRjVjeqhQ1t7kJ2/usNJB32TiNK6Nh+j4W2
M62jJ4dgv8umIAnbLE86vgZslFXArNfnSiEVTG4zyeFP0VpBygLFcBg2A6u/nCoijDbQOGfweFAy
kkef0Z/fdGYMKyFWaQtf8/3cImNDYqmsd/NcK1bXmFzbHGhDsyrv7/4Qdtz7hT0TLCLFHvbc0NUK
6tflOAhoxymvEwHsCmTVcQWaKKGeAJeN9wp3jA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
xwoM7ayotW43xesP6+RU14Nmc58AUvvbInUQY5zu5Fuee07fAYPlDu/uZW++gVsYFSEjyTe2agM+
nUT2rLXeNMMfJvbyM1Hizf/x6iudcDzqin/4FSCc6U6Fl1RTyfPiu1TN6J9XKCgsMnc8KxdJS3ps
c3eXfsTBLKvXNX2HSbkHtBF3NfEKdDh5xavueihC/PumZRS63EEQSJ79HXxlzF6cU6w2jeDJnv/R
FGsm5NpxS86Do2/7eSCYWLY6gXORIRXYdil10fwtGh6cCNTMuHP2v+J5WuAusmt1v5cxQS3eJgUh
jxxL5DRHK6xSW8IRN6bgCJIZxES+9l8d2A/OfDApumCCYZBW5at0o6Z/qN+Mf/S/YONjQtuBR0ws
5sBOPodmTVnuvq3cGM+QHnKZX1dV/bdSHhrMLwUNQzYzXgVlMuBYhTigc0xvpcFAzFWrYMOT6JuD
4XoUIGYD9ZAhfe3I1BCUDld7AT+UQ6OLNmIYWgefyufsqe9VrTePcQigHnHz0ej0is/5sGnnfGpR
pcE2ELe4sWalWMnsQFpR+DI1wcWi8Z4E561l7af6OB5laaaC21HW6oJxRa4+qKd//PIg2mLJGzQ1
pr85MzA6TcPKFVpVULHvweWup/BU5brz4j8ldj0Jmqu6mxKFcP6RRj3NpVTe7ha6oZinhI4In32K
vKBErNT9PbQPaWT9bkJtiBG9NHwLGRFEXyVjH8tY4mCkUfYg6uPqskzv+J2xVHPpmpiVyhQhO5hj
GcByWGDoe7/AkwowCpj6qKanLWWeXYugZ/2BMycoI9ZH0J9b3MegrDLwUCl+1xU+ghbcLzjpD8bf
Tz+zxJrSY6bvKsCPTe4JfmJCCIY7Xw5m9yP/+jIv84YKRG9fx6xSkZMo4Hmw1432pVm4D0KJCcRP
HhW83xnUiFQ9Ei8esxpddVhmYjccIJ8yayb4PV5r4u/Ndp9lGQMiU1W3ieqGS61BgfbAMAJw14ov
h3ZRqBxxBb7PhWly3xrjIWwMI2AlpiOkFLm04o/rAgfWLEdXtGg+eitLNnU8TYiX5v2i8PrVH9Fo
BMUKS9vqPQl9LssB9nqGC8mmfoONm/74/UKHNtE6o8JE47Edj7eIEj5P6zOCHvFoNbIUcqqvIBbk
wnFavxgme3bVjR3KNWRZnUcHnEV2e5O989zPVNEyQl+KA86RGJgvODbDhd/5gp4sVAFoDt+MIeWZ
nfY4MTfsBHAxXhOopocWNlWy6PKPHaxOFHNjFjVlb1pVxTZRv4f51knxsSJEvS8A5kU9Vp7DM9NA
FYlBQiTYdVT0J0Q8bgbZPerSQxFX9uUfHIsusrP53W61BnnSivbg/lCR49lQsWctCV5vY7+3/zje
puuXmUrvjUAOR6QTzez3VeTn2a1aeuZHOqbfKuxbBS1sfyyl1El7a7tBaBqdu+Jjoq+m13n5BoZB
Z9iHotP5gXoWtMp/Kl5+OtFXS6dxryRAvjplWikrDejQhDsQuauFmVPeowsFcBu3QqGdj7I1g7e9
hTAZDvHjR/qXScUGhfzzSKkA6uGRiYdl8tZ98iM+CCi5BjebSLd8WYcCF/2I4eRyY4bz7u08Ivl7
LGjx8PjLfSYecjwuzCJr+OIekwoCqMwaOLqDsKjW1/O5msBzyt318+xYE0mZxNCOxM1SSPSZrHnu
qmeHIi+2o0Oi5+TzrX/yYX7x7R6ixJDwwP2l1fRtPbt2tJA87DtzuLcFlrFvOJY+9gpRUtA1AkGh
eLs7ZKHHn5+Y/HVg1GvRe4L5XuKFTJLmKXjddLZOtmCKZmdY0S52NNkbdV8jrquQLD7LBeAJxzJy
xTZilgHbXCQM1zFSSkdnrZxfZyu6laVFRPHx66GZR04iwLRnC4bj4vO/3wzO1MILuI1wcHBe7iIp
cT6W320qlC+ytazAsLqfXezNsN0gUzxZGjSURnCg1qRVaXlxR6GZQeb3Q2rf0+3dcxf2ERHMbNxA
Y1ysWFVd56WrIMhtlE3PYligeTS40V92KehFiBpnoiLNl31W6oPABE9ehB07sOWAIWYPAPDGsFX4
e7/ZSPo2dy5ncB2zX/Aw0zNSHBnlS8wOqIBn5PhX3dfWF7/9CUEdnpTKwYno3lxyNP6dFFuw+aOP
/OqIC86InH6pRHg/y0nzJ+OskMSFaCdDAGoyduXKtPGpeDJuED3Wz6jhehLBb1x0QOXnXcxhBqTi
/5Mjm3l3enuSqtninmRWR7DezOfFBH2EbDpx3iKQEbR4JIEpcV3WhdDpTz5IEffixu7FohPr9jV4
gGug7S7vxmTXQJ0MxydgbsjBRxANmLAmYM54u7E5qievaLWn9dkTiPViwrAiPvv/3yJZzhEtQ8Oi
5SamZ2Ug/HiM9oHIcq+q+p2qMFPLZSc5boehoU58ohak2tyJAtItLGTP2efA0GZ765TSWKVUWZdG
F6hZGkkO4N8Ulvsv5xCUlNIE6WiCerXB1l4M/QJ5jfSV+gWKP+T2bHEuTvrkfkDHhNH9IdDIi4G6
8PAjKhEluosJH23bIP9Ba1gnZMbP30ZBbXBHQ0SsxNDQLMouXJxO/PPJ+iWO1ddfBqpxXMxpuequ
P87RsDxM60zJ6/tow3fcVfJaixs6quFebw37Bfh+Fyox+LyzrCGLHrxPpZWyqSWIzSi+/CzQmFnd
8+aFlwylmOV7EgO6Ef6WSUuvkfnrL/z+mqZOtG9RqAI1WSShN3sfyVPWACpAPKi9NVt/l3Vp4+ki
Kpl5L8ySeaFt2OlU64/EqIitiWZSoga5kepWtsz9p5wHUzbLjZUdMdsUNSyF7G+42NAlGxpameBG
rms5cmgPx4v3J3el8Da0QxzB9HhN2Iy7idr8pVWEHg5usZ478lJrMTSGThhDOhsKRbkiWeMsMrLt
iheI87LxkFjUhGMnMdPZSsHby9KRnRT80yCK4T63Py5Y1dj9gI8JctA4oaBdfqsaBWPJCOiINi/8
yFnesmDzjUDV5nu5L+tGLfeeDgzcEVIa6Qlx3KBUbw0Bur0KypvN2m7p4x052wcvfhXIoI0HYvHE
dXOUjE4sbWc0DiDJ1dIcCWYM3D6vMjesAl86xDdmYKAvhCLLL1t88XE+ZJ1zoqQ4TuMB5GlX4phx
05YQ3lkB1D9HGOFhXoiR4m5FU6rCnPcgBj9Nsah7g9k2G5flAjRPsDU12ISSai4vnqjVvgLpW7Hc
JF6qOOwDJr/fBXWGwJWwOn1VrXTrdXCAnOl6SkPVubViSceHDe1Clrt1j3z9Z+TR4Maeet220Bft
Clia5SI2fRvNYJq0uBSnp7VKnSJOx6bs/2+mphcgAuBhwCpmHX1b2PBUcJftS3U8zHJXelHr7GbF
g7yPuSAtsAq1CsmWaWY37+gmxN9RM8sjiv42enCfvymWyWsez+X1jO31r3BDHdI5CQJR1gfdVJnF
OllKbdokHPyy8ZxXcy9LUmA09OSvP9gDCBT+Mnu6JAw0VUFY8r/f3tqevPzHdaR//fUKDRc0dWtj
F0Xgcojw1dPHMsYjPTN+UIsJeFTz1/xK5WcxI7nWvYBQ1c/ZBSLbHHxvRbhWbcbt37t5XrjzQD8y
+b5SubN/9NylBNq+A1VUixuu/nYmaSoJoICPPtiItFnIf4WnO3mZoKgBYe4szUmXUWrz4FGXv4pZ
g55bdBMzb8H7I9gC3rXUQAXJoBoiJH/tj+PS6VZCIFIiWfj0paKTG+5TwQDpHklwEUX11YTdhRqK
JAMTeNZYrDK6SVQYpQr6Q9oNfN9qIHhyEUI+ej+/cItLcYIbHIkfyEruB+qc2Z7VY01K3UgybEHc
OCC9/YkFzYmed4EJ856AwygXbIZzVqQvJkamfNysMwJgoTvlAyd66iH4cyeHHq/lYESQYY/SCtiB
UcRgdKbsIBUr0cHcWYP+4C8aJCRQFTIt47BtQOFL9gRgDN6L5dHpCNMwPmvlNL5fzPkrzUVd1abk
Td9a/se/2v/I08nZdQhBrl8oJUZFv25bOw6U0eWbJ1Epu+I0RCn6o52dYvitx1BDIhzw6hbaYDXS
OMK9MGkiZwC2UV1sj4ucrsMuSAjJSypSaT94L79i30QNQzIsMmABYZW/PpURtsVJcBNB1mRWRDf6
CAKxOQTrJoNiq6kLjHfApmhCqaxy/E8ll6hCtXwaYMLJXYXluB/e10ZySJ+7umfLGcL2KyaputBt
dci4S5Sd/CcLAFRYUX7nFmHSL0FxUYB0Mx2N9nhnlFiJZuBw5CVxAFisBvieWBBSopdnx1Dw6p+v
+6yyLgqhXqDUPj3vng+UdO/ORAyIOEUmYCVTsKBRuGoO2sAmVF7YkBZQRpUSCj4nFmjEoLCQsIiu
BBjhhbKAQlAxnVDNy4Ko1gt/0N+6uFkciGK1Teet3Q44hUiPZ621JLdr2WvlUIgt7kfpGR9nVk8r
Y/fLjBxiyDrdUzdsDawOw7jNHIJxkDfzLaLYmaPWRwOv6YH1S04xFYCtloFDddCmAfObgi+gAT+c
QMXQvV8CAP2wyYqmD+Rr7Yyr28NYNPE0mB+pWTm1fpJTERPHwpWBv4FtBBmufEhLSsKogwm9TaUn
w+SlXEygWVUXNmy/tfRocfxMUScjOYXWbiWDyhz7wsAhyNrqFUNLS6SVyr1Uh3wbSh2MxmtYRa7/
Fjaf3/zW+8Kud/ulCfQ2bNF1fZRIr/+tuI+MxMKT3uIzh1JD/bfSKB/dCJSUWPWhwgG82/tlu2Fh
58IhIbGBm4u8J+3H+PAm5XYm4gqEJJPboNTQu/XgvWP95gHL8BxbPCqdJVg8rzdpRkENJTaOVElD
l+eWo3+D8BakbI0xRpX2lfgWjMbROEdzD2R8xloWiKmcwMzoPbiXgfCilhi4qAOuibTAO9f/iI4Z
LIU/UEO+4L31BZv7kDTlO7XCbe0y42gNTiq0aNk2lMXmzkQG71Gh51r6EbzAcoa4yH2B2riE9yV8
qf78FswrVBX9mp27UW4MPxc5juey8PpWXgzW9wDJutMGiiUuNSuvH4Def7FUzMQksg/nunvXU9JZ
fdWkef4ZW6emlhb6SGUrOb7IA5gT5BV9yioOt6R9C2OxJ4kzn1zrYsbXorPlYc2duBiXp4tF859a
u0YbaTGuUHCaUpdWR9iY2XUae1JuC1jvo0AMRoNkjy5vg3APeLgjYdzxEQzZByhvb9S2njbNvobH
qGTKgiQctyiEvmEH8StDUtMei4Fmc1eWEZb/YYtT5qNdGeRXa82+SUlTH37sJLQZjMJnsj/06DnI
dxXU8NB9kZQij/BDNc0sW/VK3/nLV5/dkFvSfdu0vJgi62SYG05AlNa42dwEfag56J7K1AhYHWV7
lpZ5wvvWebgfXjsd9NL/Pf1KhotFAXxlHtKb3fLmXKUEy+VTzylluwxM7Lq5lEOMj5kwYvcvjOGT
GE3H0cmI9sJ+E4x9naVFx7cdAPSGO1t/m+8zfsKDDVX76cAXB8Kx8xTSUAlAEnwZL2wM2ozva9yc
V9m7fqfdvr6zxVqDx9vC1r03ozyvama8f4nCh2pva4t1OyVp2TbY+vjjadkHeprT6JLZ5Mm4ng38
PP2olzCvnO1goxqYXeaNYGWuIxg1tAKo9QJx9a+axZoCiBd5lRXlhN4QLZ/Vhl2x1loeU91j3SdL
sFOHfRZVPtNnXH+IBqEVoEcfDZ8hHE0//qaMz1SEZ+5ofVsHUsOBve3qRB061XvD6mKHlw34NAc2
kdAX0252oeawCOljelEGDAFQxDorMms/gzWwR0iNFnGm4/hldS62vWbvY3JxcZyFLqgnHgCv39Nf
l+2gKOi8IKeCesQ6rEwU0dAfP3kytqYnhKJ2mrm2cjSCM1OCsH1RkvgCZtzS+Jr2IDUc8BmYHnG8
OusLY00MRdBoyEObEtSbDB6IuMfwPGaUxg4d0QXCnqDfgCgjVpDGtZFHppdZtTvW+86pP3JLC77j
THqH24SG5ne15KXzXC1CJqAMcLh7HfKJTpSSRdwI7PpHC/dE7y4W1sF+/wLVDUKMlzCW6fEVCitE
o27uTuTblSqkMvq4VeviPLKAzO9RsNpOVHk/kXuwkR75sLmHXA/RehVl2G5cf+bnnqnpPDwLNMN0
2e2BndAlQ7qwE61Kwczd4KNQRrxaN2uUGe1nRc/x6fHD09wdO+/vd7C/rToI8EFF+wdXoDsGnAzQ
W+t08fi4PglKs1AmRCG9cebXWUmjQpg59s+9QbQEtLBmw24/+7F2SWC9O2h/wWoYcB7fuNGkEIvg
cbF93aAyrNYdUl6AWDQV9W4z+cgLACao3rz1BC9LrVgmy9ykwZGS+Lm2VeS0WPs18yGBhba2C1eq
cf3wzqdfJjVq9Zf4d312MR5QKIqAdyyc/pSnp5g86QQecEj07oWQodBCT57Umobu2RUs91hZIE2H
XqecucSudloQvPMhqU9vjqMjatxhlJ/4MYhuvSGgQWD3Vz6c7Wo2Rzg+7RV8S6Twiif5oFgM8r1B
r1Qz1HOeL9nLWCxIxsT7QPftxb4Rffi424iU+bdDBX8ax3gVbLuusJs2P4HnhK3Ucmj2ijKpCQev
opFi/dOI4Wp4IZU9T0/8PPsC0ZYDj8MoGIBtOiz4V+Ef+GpMMdfrjhAccb1H0kJgZPgu+RkyWGQg
CTkpQOCzNicBwzaO6RUkJDwC0Wz7Blkm1AXZNjIjBejv8rYYIxYHALyGKYwj9KH5eh8/aigsEHA8
oXPBn3YMViHwALHq3hdEe9sCCMd56TA1goy1o6OHVXEwIDbRxAO2z/kuXRdP3ZaXz34cQACXXTt0
noYBEwaAmLHfyNBsUd7S7h4ssEF36PNpdG8Op/lb5Rm9EjsnoPVNxecU3yciTBhvyXuz8XZs696L
5nZ+wquifFLAixuN6jnDPDvRhqw3kGMtKKma2fvHZP43pa/djIGm5mp2/tFKCy37gL0pxiQmhlfX
oXEZOK5T2wTdhh8FZhox0IbHa19dkkPgAYG/lXU2ApVJLLENI5XMJ2Lnq9yWP71Cloo52M6AbL1z
MM4Nl6WFIp7vv5DekDQgSE81saEzbeoB1I7UFUuzJAd6f/cJySY6QoBdFNqDbbqWcHDsayBLvK0G
k6e0YUV31BZmJUhAUHBoKQmTrUtNqsDbOqh2ztlfNgTDbbziIE3r8Vua/cvX1q3uaNkpCawgkCKJ
rpxJkGXKC5iTuhY3k+Hgj+5Y3C5pZ8j0d8r6d8cp2Z/qNYsKVSGpGMETNeG2P04614e9XC785XBy
7AZdSeCvmB6GobMTfdPenuTWyXLk0JgljVZzXVhUpRVC5VSr1qVVRKZHMzNlleIHiYzWR1NAoht/
vPe2OHW/QlG8pLWZ9HwHRAVf3YqX+5maZfNFnCzp5+KEPIJyTqH9u8u40IWFnHKgD4TBg4j7E7Ns
rfOCDvaBA7pUNaJkdDY0xVBTVJUEL/HqS06jqF+ln8oOy1DysBis0VEf0LQ9cs2L9hYgzm+sqxgu
QSLBInD/uAto2UUGxy/KeU4YuPP5BaC6JJ4OhdaB+gzx5jvEnKBFkIVqpNH/SAk7Xn9Ir1N4Cl7X
ArdMAN4r21dL8r9Zy6mkT8fQdP2cYIv5YZtcoursWrA7AZTuxOtLBmXyIs9qwPMzkXlrI9d8+LzH
bb9ltixt9RKYDdS5ifiIuq7VkYhdMAZmiSj97qNbzGRoENM5w3MxJEvtFlf57SChwJp2akk1AFvB
MwniHme+0zyFElFnFAk3DUWBpN2pFFPPyce/NxY0K2gq9GnPcRbXRznJPY9u4dYWcJQWRkZ1kfQT
73WwFk7bGs9yZ3TD9CKA0y9+Wem49Pz64f4H6Drzj0zWlJFSIprwEwQ2v1nybemZBXjxWTyIw4Mv
p5iuO4cmNSDjZKAKvb+E+HHo0YWCq7NHLKngE3OWAIrlFYM1+JYa+wQVU/toaR85wLX9sm7YteHf
PmXra8IXf7K0ME7TbF3CQ00Nyxl6hwkARpQ9rpx2ySLgPqA80CAQwdbnvWA+IFkXC1cu/hRtDaK0
RXNqOL0ztkxmE72HJ0rnXiRagG7rE+IrGz/dKHhdy0M509G0irOttbZlbjwcO4n63EUQ3cCOgcs6
DiLdL50n95Pgp/Ze5LOTAGJnPOP63f8c2InhH4junwUcPEgusbWJ0aRvgOVNT1NboOmXUrbYtHN1
GEFHP6GHvTxFLF3rkI5uMoxWUGjz4+apcNRLzgJbYf9IS/smlySq7803zf0ztEi0HnZYNP3gtGgW
VRer1KdMozPEboWcspBopkGLW8DtgQD3q6hGdkHhjYhbtWuyTMj27ovtANcYehl0zbfF8qVj0lmg
bRE+YIVyoPB4aTCcA+u3LKzJ2COLUjvyfNGGmxCHKy5gDYKvpikPaWkjcYIrbUU3Br55rjn1z3BR
Ds9/4FRbEXEe0cetFnIwtzR8XUct8wzxoP45NggH0QdMb1tFuIKW8bvjVsHzuD848b61rF+WSXsQ
lfSzwABumtLNc98WqTB9jZkWwAaTdJ2JoFpg1oUaMAYUjphJ713VIOJNed/l8WgeM+pe+m8oRaVt
grMTD07qDSWVbBj/4dbGooNogWZw7ZHQPW7iZPan6KG2gzrvXWk3kQ76cKY6sHQyYl1fm7wpsf8l
XU++hxXatcz2d+sh9GMPi3dXlUldy9MQWwWad9gdSB3YClTm0tj2usZh9uRC1CxwnXpV8zz0wFnJ
GGx8rs6T6Df+9cd8SOIGoua0bSZ6pGnSuxsejKebV4kr5mVpQpo0l2LXeaCLCYdar8VkYsLbaPF2
gVwrxy52JQpgLDuS039lCNidAofoCcj0yLXJ/x+8Tt6XiQaXT9Ylz+vu2sDmIR59T3QYAhCm84ia
ee/8AZu0Lo4GVu+Lc+YEt24jl3mBIvlssutnI62MEVtrla/qmV7sB+a3pZMBH3IqifD6j/jmgfKU
5z5jHdvHz+MUR4JiWfLklGMK+FbFZ+QrjXeOsjIXWLAEvEE95jWM3/fEAnRdgbZ4KAFXRYuuwN3g
0XPm5p7913zzYASBse8958nYmFvc27bRB8EsBVvPSf3YKwvzgjJ9bS2acvAFn7sEg5OEj4FJwiyk
qMXEsYXyKx7jKu0CrQN2UMjO5fxa2foG1vHMzZBcnTEsj6H0sT4gZVOVWdr3WZs64rQuARPjsQ/o
H+PEGJqPPDjRTgKgcMIK4jO4ZTPRqODz/ZCqqkmhjS8y14CXGHrPIIGoukye3dkNZO9kveTUSRBg
uJRaxEHnWjjwyXTiybcicqz2keTUI5Fykp8t4hF4QKRxniZJLtqfl046FG6PTN0yM/UPrsv0L8uO
cwrdZSTzMqG6ayPAIuaXvfLbVOTNAsOXt/Z75l6Nw2GRnW/qHyCk1QPFmJ3I1tN3JmSuWrf0dnjr
fu7VAW3sUbzu3ltVXri0MdqdZovxcSyzMd5XGgPmq9HwlWChV3gMvoZizvG6A0rK4ZHF1k0IziHC
tOHVhVgLmN3LqCWxWlGSN60VFaKd4e3Kl43ujd5zLDRNGPgwG9TJiVzt1G7c6uMZCX4gX3fzLtds
pto2H/ACwNcX1va/B8dgTKrIO0rmBEsYDhtBoO2TEYsjoMGIXMyFuu1780QDA+bquFqqw5cAGAgI
no+8xSLhaPGpAm2Z0bo4gZjSNI6cyyu1RfjaU5UjYyNVe3WZ9VsP45DBEQrzjmHFUKplokb0NV4K
Z6Xf3Q+BxR+04IDg5rzI5YAn/aH7ni1dfDXO+qhZZz1xw0LoADbq2BKpkWLQ5YLFany3Li6cDjnK
mSlRXkw3lMPAynsNAObltNAtnnVyH55gAaqSi19j1+csIjRIQf1eCV1K5kMlzS8SwlLzg3OnmIWO
sHVCUHdZv3oxgm0yeX+vBZect620CpWS/zHgaSGijueN1nhz5vML3on4qjWMw9hTEwJsalICYsK7
PvK1bd//D3gZcqFaAasxhCxQYJlJJZPfPAHcYU/kN71jEKLJ1Ab0BRrFCd8DQ3ARhBmDn3nOivjP
w1QH5VcKE14cPrvAdJ8HKY4jFTT11jRMQwy5D30EXAKRUgFPRywe6wy/ENJMP066g6SAAp3w+GcC
/eLLEiGWfMMernodb3EJyciEfqRPZeT48QCxYwAuCDn2DfPFzxaH15NEQQfzHrNr1O+/PxRc+BCy
iTtUYvVy64VA2xCERfIo7Fwz64qC7IVm6yPMw0I7tw96zGlEpfnd8sIscTH26jBpcc81QRnPKMX3
76T7vQ3cLmkl9tZVsnKxKdnP+cuTUvPf9t1fzg9kRP8h10XEe5woSZg0/1Vj/tMp45w9dj2MzjOx
AOEp/mQd/3Lkpb97Hp6pvTx7eJ1auvlYcdbKgCexXdpWi0943iYC1Y7U77ugANEkB/kq/vHrKf+2
na2oY+scaEIAwIGTTIu10RYK0KC49wukFysZnkaOQRTlKLcISW9/Wj4Xy0kw/194yx94MCxd25pa
ufYRMxhvJsZqIJNfCrKoe6mbJYAO77B+vGfFeCdoktMnmxJ7Ea4DpdTbr5O5Io4u6YZpg9tLvYL3
ERJX4GU9Krj/dmCqibrwyf9fDG9OAB4LHC6t+Y3H2DAomn8ALwBRhU7zIef+74JtfEq1FCuGJHXl
rR7YKtUGuKL3RFaXD9PvfEhb0byeVDWcabLiukOuQYeLzMBkFAAJul3+VNvfkOMVMPr9jL0erzeP
gd6EeX0jPilnkHl5cIPzNSCGfuX33WoYz4TWMpxcSCFfZqb52xR9o96RnYLXKnqD7fSFZEbSndFO
zTbVoMD8db63TknMchGmkVyj5OxokztBfkGA8I+tjjusAmqk+HpwRR65+Zw2ycTZAq/y4Itj/F7w
xn0t8gI5KOAtiSicaJuG5lrAUxC5YWD9Xd6NCTwCWo32VVCRlkQoj1nq4TFbdIytTU3mWLAxcK2f
maWDmeJBVYSpzYubcLlZWLews8+ROKVgWkchMEDXO+eTQtavLT6V3tlqlDRlA+9GvSZo/lB83FIC
E7icuJle1SecrZG0r1mG4hmJCauVCeyhRtdzakzKwbloQwBjtoS4NtIgL6SZvajee9u4oj7uR0UC
Kh5ws7CLaazy0ZmsjRn2l38tKDVwXU0thM8hbEOpE4gGxiHmEnbbx8MCDxwJ9ewf51l93tWpyjHo
bWQKlCg0lpLSOq4g+F0ZsvWgJMAdRhdzSfg/UTshQ0xouTwGvZyLXeDZydSF9+Ag6pOqef08SoTr
DaMhKWkmxribeSysqls192dWwPWR7IHT9tJHCaS21CIAQ6oM8Rq3xbwSMjV5+LFitFuf8wDBlF/v
t0kgqJhRg3F8k8nU9FYErsoiW8zeZ6AAm9Nr03sZVkZ/PNJxNV/aacLKqymjMGVhGxZ0TZDYglDW
qzeW+fa153zY3xeggmGQXlLZHr9I16bYfndfr9eMXAChW2qSkKRtXJu7O+xacklEzI7+ltfT3vkX
ydNI72Up4VdoHZbsg0lWR0pkMJhF+pFEb4VwgPM5HmAYs4o9VAZeTuFvvYmFJMZbaEy2Pkdm+an0
Dui33JcRyTMfCODwjFxm06ubGoU/MfovpBi9JJFf8le0RPMQHaABhaOY12NUPtyZOMfEAz1n8/Zc
TaDBZI2v3qEIRSVKf08lf6Rm/J0Y5JJWIKF14vvTj3fr9jj1fZwI5UqZw7gzr/rD6BaUsX/clX37
g2NUIx3Sdz4gOhVAEPUlKIf1LcqL64rDDR+B1/WXqCtdViC0NCvMDqmhoR1MfZB3Wu8/BXERZM9g
kzxS7HyIesFsRlPzXjSJ0WnOVspELXv6A9DmDCf1mNkBKDneaXg8nerFVzyg/3Dic+Zrav1wuC44
I8zGXGYLKSbRUcCDoS+34D9ZSJ10G8BIah8XJ+gQoGvlCfod6tttN3qFc/vPrQWV8aUTC2PIv0xV
1QBFSUooG62HtUYxbOd1jwqWv0q/KUPA6zjbtntwCQDvb/NklTKVLPNulPXKO80VZ2YGlYeaqQPR
FuFnXEE6aMHtd8LINxgfDESb6F70QrBsMVAuSRWNd5zQE5tvVt1iTCjD1RjKrMOTqRijgDGQe8/m
287I0VZ1R1+ik7X2jdNNhxqQHpMw4eWYq0dD1adI12EtEJ+3eyC5G8nq8RMmeiqG3eXFVmuzxxzg
OOcBCHevWvCQw6YJGxjFUsjdJj0c3367PcxFHE0KyTe4NrcH21zYrFPonhEN71tfFtvgOV6gpa4x
JFl7Ljm6OpOVX3scnb98Foa40BJ8CXZJIySgT7BTSsuGOeAmf4MWwQ0dwHw9dtF9MHJZwNjClRss
T5ppZSb7tY1m4jrCXZBnVozfDD68HRJq7uZGLKJQGLiR/u3gV6pGRz9RZzQAPUQOiPwNDR/b80BS
hcuI+tD1cz64D4lvLEYOA1eQr+2WIfrwd6p0jORnEHWtzKx61wIJ1JUmyeNjljVXHpZER4FodOep
6fdtAL52OeYJSvaHLAWMN2FmcmrxSyE+oJgHRGvRU4YLJ8rByTB4uunG23htO96g8d/YQHsRjUcR
vABDoiHl4bWaeF6zjd0bjCly6RN5/ExtCbTPiGECiPjNQXUZsdDSLG+rLRFAgY8d9OjeHCCgNycy
eoYVrCiergT3u1lqPbyPtwZwqu7ewPeJ298lCyMk5PsVbxJgyT776YHWKRQguWLS3ROPsl9oz5Ek
OKtSEsrA76gNo2jkhhaiTcWCeKtoZU8zGadyRUQtcDqCQoSuBSVDkkWF6TqKpE7gtqDdKTGo8rxz
xtyvNsuDtbYAg3CUOQDEf/IaKBiG0Ksf3oFxtq+WMz2tuR3Phb/DDNw+rQNsCC63O3uzAo8h3Jq7
uqS7Rrx5IVJb1+8g/U/ksPcozvgO3h2M4wPfNw6xd8HHak8pMIBjAl3jx2U/EiHitxHvAM+fqmqr
BoK1fdL+9X34QPfRldxS+H+el9dTUJbDfgQPTcmgpqqt5IsDJgVWzT8yUFAHqd7sikcKjZSiESbH
IH/Jp1b1M47xw6CFBi6IcGgi69nE2zHPWLEiImuoorJQd9p4I4EUx+wlc9LMUxHFJ0q63FRSD4yC
lsPeO/zlNhvsLzEcEgo6IAsQjdnIJqOe4eV+ad8l9S9mY7eGgHGPS/LsP64Bb7VVZsZpCRsqy4Yl
Cj2yCuOM35XQsQvvbc3gCcVCFTWg5AVsydzYsC3J+i9VoRzEHl/SYjI23S41SA7fKnjzvI9kyHlD
xoRnIyNpwlZI7PRK2LTMQ71zrextwzB4DpHuL4n9VJEkJRJIqlr6uvdFBACBG8HkIw1Gb28xZYmg
Fi3YjV+KnTNrdC5iehT0n/O7zm/xeCVVn96L6Ea6uc+Yl6Y1gjKbZv5YpjanrtbLEjlGmBaC00Ts
GVJDVJVs75tKxEvsv3VUNxXp54vIjqM4w8HusjSCRo5VVuk6cJo9byue67gW9OdrByj9UAB1c4Gb
l6/dVx7VKL8EyyV8dezsx1xWIsJn7LPxYeyaHT/dcopiaeDkI0qS9nYUvWMmMISsyAX4MHK51Lzm
majmk2FQ2FPE9GoUVFRYfOOicdM3D4kW8gFpvfOXhyGOywgbFfxtEUAhk+NbrYC+C+kLlbfNlK3S
In6jXnSTDWUAiUEzZED3hEocN53o7OFHlUyi4N2mtp1yFO/F9Q59aqYtSBox2IgxK/EBKREJ1AAu
JS8gwYhh2rzgN66MTyxv2oxIOiV3iJF1mzKlq6RQ84Z04vrr7TFgMXaMjE7mmpeOQPqPv4InRueL
WLlpHIANEs3de8eRnwA//8nZ1HO5XE/XoKVlgbOx3B93YmstuOZnk1YAKIUfnRVOOavGNaqeJDtv
sS+jGkXHT/eBVMh5T/qLfWaz/Ga8ipj/WEH0irOGBgl8sjANTg1ss33Pjg+xI626IlpMqBdxNe1k
W/yT4hmwaCNDOAcXjUy85EOLp4xWg6M/XRY6Gyz3G80Nazv/Xe1D/E9PNDPiPmDyIXOS3WWUeQCV
woqasIOrFYX0m3ywH9seIaGFzwf1jIsgqIgnpPLKJY7JD4ZewwZf5gcSw3A2HgC5PzHZYi3ieVx+
nL58oi98gmcOeFV0O70/JkW83tj7qFBwJptbp+C05w9SRD2Hn/ygtFDPDzHK0PdwtO9mR2GcCQMS
9lg6YLRswT764enA+h0d7xrtoNg1Xl5JSuJ6HSivdtCf8YoeaL1vltixxOnHON5MeTZmI/HvMB50
WwZwk8pXb/7brso+b1dXSf4GZrOp1kDplKl89pWQ9CdvCkfYfxeTIM900VFTJ419/fxBW44rK0XV
+vFYFRt91e4OcDTmZD8wh8yZ5RtCPwixrojmdyzLoilqOcM4AlxXDkzlK0r4tp+4labg2FVR0suX
r91Wg5jKXkQTmSclLyQf1wJthWX8FYDF4iDT+/0LsZPMqm67CmF4DyUsNzq1DEoOYa13gFSTDDHE
rfE3lH9K9mah3TAoEk05oCNW09QXeeiYKLPDTfbDwrDedWkiMoA87fZjWtJS1LRaUkUHAPsGZuiG
TGmKfVySFYQJqnQCf/wPfWOBG3loPV020mJRmRcwUjyox8IOlJzky8TdwUT5tQ/5UZx/M8C4L9k1
nP0zTPzzesaXzm/p/7RGo2OT/3Sbj2ujRVlzLQlihTWihQhfWXkir2v8KS070nuHkOQI9KuaEgGn
bBmQT5Uc+Ki8bLdkWd4qNE3NQnLwXuo/jA0GvX/ShDjVE7e2dtagcGK1JpNjv+6t/+u4pZgxK+MV
nvbTejvDKuC/gqHzc3i9dLtEqZ/ByXqPChooTjUuXYpXGYekPIfZ+5L+Uxf2oV7UY7PFKqM+LKaB
HDxly4X16i+3w8RCPFTghp0TLmJWFaUvbomQH3DmIPv/6XHXtRk9/+DzqllGoPdLRFIqGmUcNNmk
ouEYmBWvsBstokDyb6Zjk1Nrt68G3jRGwrVXPNikyhU44O5YWLofafCAl4Xbb797+HXk/pFQZJh/
40a6GZ6nlH/a7y+N/+pe2c46zSsNIj34dE0vsfvnAR2gVVX2ldJyg4h4KwDZusDTI2P256v7+l2X
w3orXZDlHyDhW6fo/3+Bqsi/rz9TjKRpchxOk3cZzNHPXnbv3OSvMwQT+3VEZZredyktN+w2pK09
ySqmMF3aaSNccWv1hIqWbvwLr0gBWdQfWdf/FmbB71ftclI2im6RRlMyNF4/a4ga12wfCOhiE8B0
yk74qtrK5pB2WJoOHdYORHBSXUWNfTUS3djc83zrAq5Qx0BWFZb2+dOSS2qqDLKgqHdOHrs2LNsi
Ji1OKjC0P3biaDoEsf6qs8/oESqaiHE05+ZWkzF1tcCxHtGP608AKllQi/osVE7Ej+2eAIO3opAS
Qg7KlISIC7/qdQFDPdnhG3C9zy8462Sq0wUTmRIJDJicXDcQJTvGgdtpKcOW6fLAOG/twcSfGSvm
5dPc3/Rbjfnj0s2EpRvbOqMSAlY5qI5PR40zR7J0bIy823UBEwFI8jWwLdYBPVHVtxmze4wxuwqk
2SLfsxFfMkGf203fX7MvFXWnk/4rCUD8REIzCzyGxtheEv0vUY+MeO116NrX1JT1E/b8E1WPh5pR
2AYeMAqKkTFPUE9r+ynQWf8aFUcA5VjlL4SnL/igpAQGppYPtVKPpaVNSpRYBuWwwjY+w6T69vDk
qEZHE/NympIIHrTv49+mvPRCM0IY2IJsp/TAMXgwOn5K5nbDGs/MzOJonpBr3IV5YnDeyXcdbdjT
/NCLcvAlo6HW0aQVi0P0avsyHuupUktWyRuupM/tTIyl85ak0CVNSAwRdAQI/8F191GbxhOOIbgu
9YOpkp9qZchun+33TyaPH0s2cmgKkiMJgv6sI5yz9PJ8V2kOx9Yowfq8Vl84Quv+qk8caLjlSI9b
kZJO3oFrHIthFFggEVq98KrvIsUz7hWYzvI/yUQUHWk47yfBXSDOWUx9dIU8/+uB5c6rmXwaR7JP
kj2Pyjy1NqVzE4KIaBC5wbU/1NkaAJWYxyupvIpEw+Hdyqoy53CP4XDjj4SdB0T4BxUSOOmJNx75
awbu+sa+wObqfoHVyigY/fuSmJhloMFn+zN+HEwV1DzMvJO+5Qzd3w6WqfXu4BV1eg17kFzXFu4M
X5UqD60we2/P8FZGarV4qJz2Y1O6hcCnL8f0N8NdhBvnk7LevTov/Ag0Xe0ihnQne89DX1gjSJvf
nVrrVBdPbpgp1vVlcIKwY1i4YdDE0rQ6dsek0BYReXO08PfLaOJnYrVe5FuyjxtXQUrIjYvtluMf
2obzKN0Si6QGqWcoE2CxtZdWFDskML9EIA7VLQ51Aki7Pwa9N2ss4uz3y1pFAz17AUa5mmOKeLfH
alE+q3DpVZVJdjhA8DTWtvHjmCDzrNlVEzZ1PxSariRbGnuQCUecOQRDnM1oclP4s6zumzGIONop
GQ9p7BWRIraeAc9rZehayZqOpGAp41jZq/ORp868v2qhnTJao3hHbnGfH3je756d9ApCreImkEfD
WkxFXVguKhHYe9VsAzmULk+b6oGo7J3uuG7R80CZt+l09hUW3m5lQZB4pjVX2BHAdXPb0PG1bwsM
B4Dk+6si0vhSUXJwVR+qbVFGTPKj4W8UuwlfcqEOwhFsFMnSl+On+oup56QJeKVBE+5ohWrf8ZO/
qjC/Xu4FFWIvaN5wsEcEEe75OBQ4uhCn1sIcGoEgCIKnmzxJJeOKUlhM6A76OdyicI1akR7IBY3U
bLfWes6x4NjveoLA5gfyEU0B7vZZoRMwj7fFsr549xQp6a97mn96HoD2mwUIdpfouOBQnTKCuU6c
ZAVLkabSJtfMcOLglmz2f6mIqsidr5Sf0JA9F0OmhluOihxr2XpgJz92bbZ0d3I6v++fpYpXwCKg
tCgX3ATX0v6f61kqEpViKhgm5bjNp91tMK9OSuEfFVCq6wEy+uUWVhnLAowO1vsC1II1dSWeMLIq
Pvl5rn/5TekhwGumOzC7KY4XkeEHoHURLlp4lY8IyPHskBXdXfVBR99KTnbM5aU3nYXPwsv14YE4
5XYyNcyy0VyO3Duc846r7sBn+53+Nud62B1SfGfBIVsK8XICk2Mdfz4Vfuob+Xumfh0AbIM7i/lz
85G/yyqfe9MOzWT7G23qgbpwXben5rnToCUA8scW2qd5g9ltx78MJ6vZK8bz8zj0I/jtBVC7U6GL
4RowA/Jv0CEWJtdIGyUqiJxZ1ovUCcrZgl8+pFmWZzBgS/iD/eOsSrbWWMBvVtXqXkLemd0gFb0+
3MrlkLWf6ZcxFTqSbG1uzA0t5EOsJ/+n5SIXXEbIMcOLSdPmP3ccfaHDrINjqS5eIyzW5jwJ5QU0
Ju0hhGdFZelT3KOvdLP8IENm33RwIaq3q6LnDJjl6QutcZc6VD7Tos5l6geC71UCpEs9/YgVibNl
3u1JiY7dZOgrsJB3/bOAfvWz98in6HBiZML9zY2S690JJ79E+e4zX9Jkq3gDQh6bArzA5dXDHstx
fdOFUXe4Gfp1TvfwpMO1U1Tvk+gh9U3M0RIWFiaW+5se0+mOC43CzooM/0bqABAoaZpbZ+7cOcFf
eVMJCqzi5hOmfQf6Fi2F7awF+25jzzsiOKjuLwD0itTVLCxJhBh6fmHFwUdmmeado8nbZ6eU9DAC
DCIBZ58N2TwQYdOi8QTSVkDnrYK2YUIH69h0VSJSLrlkPNs2xUucbcYSOxni66McunDyuB0Uag4o
hA0+nNU+Ih/AMVGXZb8OfsTy6Ss7f1lfpUiTeBnrShu+sJu/hSRCiXAr9qleXV6B2uOTo8ue0n/h
gYUMWfM4q+h2Kho+1MEHMvi6P0mUgNmloei/mws1emYpQ25Bs14MEnh4whtnS5W76PNIwCT62ajp
Ngz0Ot+L7SDpHxOp86B1Y7wXQv5u07he58hO6R6fWHAinpFHHikCEilGFs+IK69aDexa+SP6PGud
NPb9HLSAllBeO8zAZf8Y45LOVFsvxpZLeIqFOeZg4oxm3tm0VtphOS3oG3MKpMmRCovC/w5OZDlG
qTRBTh3bOWYfBihwmFkyRkgYbDUMFnWRSZA7l21iVQZPNcNZXpvq5IiGKgv/BiJ2aCQb3QiLa3x4
wXWKx8Z9esZJVO5K2DipySWELuXkbEkkahzlPdVZi/AuuBZokmsUmQ/XyjhWvxk4vPq2uvuVxEPn
jTC/PTTrsMiRbSfOqYRyUOgmuZM3Bkfg+LV/wwLUHfIDjtPZR5uMC0D3U3QQEKzzMz44txQ/qwaJ
jKwMsrSy98M5Ai57wk9iWopxyRYm03JjWe6Q7GKYV6BpLH7h/xFE/VFZaadcyCEM2qD4W8HKssvj
gf2MquDXv18uH/yI9NaGLajORHpRxyavScs7Qz0C/cZtXcckYjzYftP64hhsSJVDkhQ4Ydk2+Fi7
5PO2eScC+TATibuNlT6cNznJ3n9nSML6/jfJZOiuqWP+yfvsea2OaLCCwAopI3nHd3xEfUKWFd2y
P6cLfuCZBkP4IWJT2lT4Wb6+mUPYYuuej7VOh6THOYWpQ2dlAqRHRM2+ohAd8tc6MZkJRvt4My6i
rQqYQwm3QM/2zgj3W4tELxFdOX+0WTTO3Tvto6zzLSioaNfXiCe/ZuLyGpV1G4LNvaXLy8WaaC2J
w933kUV3ooX0F6669d6EoAQp59/C6OJYe3EycNYTd/5rjj/PCrtUxX/BxIbnM3xxh8/wm7bKl2iy
Dt4/Z9wIAsU1U8RMn2NHH4BVFaM8FYXrRLjaT/AxADi+RZiHkdFStc/GUbAYnIh/rCDjaXlJpcKL
vYac4tuwRW3kdNDh/ZvzJlReGHh8tYTiLQlc4iZArW61hPF8Ff5b50PHrnKntgkduOLwJWYoCORg
L0sHw3zhU7AtWKgSB+deUnv3JzeGHg+sStZqHoZ7tRyHdNgtlKM0dnYHU3QMIUvxuWIWPG6/q0QS
eg0Ydk+/1pqpNXWU1qN1vji2xMxvX+Bsy0MyC7YY6H7codRvgMJV/QxboGO0isYahV/n84N4c9Yj
1j3bj8fjVj73uG6KN6PBtCdYNXMFyIadJHYlePfLLn66YRvldJmMclVLr/qPl4DxOqLx3TUDQumy
TJTMxCIwJHPwJW0B0MciEAkbdhU7c+YydkF5HAATQqyqCWtTJYLOwLyC1nH//oUVz+Kwz1N+S0x3
zQDI5e3IHcRihomfm2ivs/gWxlNU38yLL7SP5yAVdNd/KEd9yF67R5r/fZA8L/LNMEv9twg3OuNO
Cq47DFiL009K6HVelRCvku5krqyldj3xAxFs0jD/xGjHJLOxLlttOlF9tsHTVM4xvsEFmwtt7O93
mGzwVLn7sTs11eDlKnbY5dnwf8LmxfDUHGVONqgFzfPl6yj1Go8v0ZSTciPlw7dGsexirY4xf0HR
FmhzXi98zkUFT/buK2+2OTQWrygi7XbzMX3xo3xkHMY821xsMJAB5ihByI2+oll8PeY7l/J3HIW8
mHeCBJzKY1z1BIwhVg5lZ7wKzHcpbwPVHsKgcVfXPG6uoVtqOvxy34aiRV7zRy6vakEd54qo73o+
ZyewTR2iuM8xdz4FImc6mDus8we57rBef6IjMLGPhZ/wuD3XCPl1hX1cNo4CsSFX9H10+wa+vqdF
YOu1ZlXAD4On3paHWVjpQSH38SmBJ5vu0aFEeuzujSLB5wRudEbzO2I8+8hDEPDWcbjY1FkbLCc+
z/2lyWv4bsoionl1JHf/fG69YqhDqZOpiayzBCV3vAK5LhoXPdhTQYJqyNd5PP3I+5sZxLNPZThQ
Pg5TToboce9/7cnXZENyCSUnoX2LyQNTJqB8r3kY9qMIGssB1k4UM8LuhiZxOJ6o42BgAz8YIHZ1
uzn3/eol6LhjjZZl5lUXh4RnzgFwRy5wlXK4X9iwiOH4diThTjwNqmJdW2ahOuRXblg71FQoYfQI
luN49nLRS2h1mfmnCATPbg9wgg+kaasVKGzD8ZHpjCSQhr3AqqESDXFa52DbiFuHouCtZ6iOGWgL
c7RUD0LLf8OjiSpA3EdbaLZNp5Z344E/EIs/Axk4HSdM/n3+HAce1ki97KsvBU10b+Epm1qWPFp/
VWAqDsJnklhGavoxoC6uTj9tzGE6UiEjc6WdmACRqzgyhE0/3SjiWV/3GHcHA9Pmp5Vg49PZqeg7
kx/vn7HjIPfukitqTWSxKzuW9lGL6fARUGs2yRHuklmiCm+xVjmhbpkMb8BHxDHj4KCjV6AuKlHZ
gRkUS3gmHK86HaTTURFw3VC78lOy/9S5JTPW/KqxFY3ecXFMZeU2y1iaQLWeA6v2cp21pusGMgQ8
3LAMznO5lZRX2vQWMA+UuZi3nM2iE16TDocjEyxT2QtexM6ELtm6RhhGgSfVshxSzkXQo4OK3Gk0
qrfo2LkHOi7XeOmVnKiJhAgzOSp02HtIfw1RqRRb5XIPXAIcdSHjDV/P/Q1Mc+EABUkQ5PwWVHPj
T7tIMv8KHEJ6zKRNa4tbEvVbZf0MGqVYZuBLJC00suehHdVftm+zuvUckXi/UChWyI1wNI5TpGJl
2HVfN6N0yterwKkW/BW9Dy5nKjlf3PcmcxvYSI0J3+a2J88hQEmOYfbD7A9XrNwvzGgts8u5BR7m
oZD5hsoqZAKq2qpiYyjntdtWvFC+SKKhV4mLyeckqAHX4emkly+AZKIfKPqnjA1XCM6Pl6ZWzPqL
iipeFBCxsMHFT6V3C14vojduyuvyKZvIqldJavTSw7po5O/fuxuCjggzJ3W3mNzdQVaIh9haDgQb
dbTHyAb8vzJLjF6JKo8G4t8NS6TyBcbDoYQT+7Bh9jonbhznSNVXYuQG7+xbelDnKT6YYWeinAsc
nTbHlyqugPxVTkiq1OBDQUwcNRHofWSxCddu0E81PPRZF444pMWVD6YGVNm0mAxqJ9bSG4lxiTDs
Pg75jFMSm30Y0xgV5TPcBOKc6qAsW0cDCgd63tw12Y5Zm4Elg/ZoWVBnA3WmIfT+nlf17akELxbn
WQ/m+p5YudiIC1J2oXdgqzuXLTFBOCovn7ub4/NDURhIyuk6q5WzhUQwuaI5Zn0GgOxlpJNwk3xU
eTF9HkcznsLixUs+va8frO83+BihK+POjoUKa6bNvJlxcBfOqGrdmHUO19eqrAHCk8Jd8Wa3BwMO
hnbLYjjNvwZ7/GaJUz4VrmcH8n4KS1cnGibTu7rF24JWKh/iCv7KKbjbt2O3SGPff+NupI3Q/I/w
aIs7JQJosp3f8p99Is+POvAkp+db9tZWDimDZok138gjDgJ087XFolSwVp3rLMSUaWf2LXoTm7n2
QE1nTKays54Yr2LE1yJRSbJG+/zZRfx4PVcwMqAACm7m6R3S7Hy0LugLvES6SSK8qV6te0liH2TW
5hVnnI0CHoDFutXs9j8cechZG4obvAIgKnEUmN/hIKu8S8rHnZQGt7ER0VqPPFo54KqTV38gBpwi
8cFSsVl0TZHA+Q8ArSYQlkTYnlN94Qny/03iqDFdfNxgYv2c5wh5/+GWkamUaXLI9+eIXMO/N9pr
JQuGDsqdq26z9eSyB2kD4MghFmLcrjjsb16rON4K1EFeleoPHtNX9EsGICh8+Cmws2e1r7VGNOhX
PaKWzsi3wA3AvuUBY9arPHmERV1AfHggAHJXZ4FVD/4c4PVSg0EWAaJ0yLsIYOnFllCFkSCEhUmH
14mFGLAa4/Q2ARj0z+ltoZgngBCzFHxuqM5DC8Dh+SiTLIsHQl2JxlxqcPf7sxJkEx2Od0rfProY
FKuY84+YcP+9Cu4TueMg4Cb6E86UxaTdFdok7v0MQ6eMZnjj1+gpd5lcJzGpzWPqgV9AN/bBeMB6
yduvL5rHNNnbmYfHOZu+6s8G4miB0QMongF2pCznVSwaLH3nRYA4uoqLhiF7sT8djkCS8OyVyKbA
+Lc8XhvofOE/0DfaNIAPhRx9pMrEIk/vJzneI9RsCyOQ/Kx5Ee6K3M5A/1EyjcKKS5RqaQ4TPabo
tVr0kA0V5qJ55WE0OsA3HZQAqz5uLAEOKPhOK0DGo8B+o6quoOtfdFIX6wllsoi2906g6mDTVXQ+
gE3eLTvf918GUfHFhEX4CqGUYkZMcAp+WlOknVs3qBkc04fwabUGWhO567y0DT2qwq3EWTbVbtgT
1X1QDnllYLhebvH353kuZdz2shBkpGfhboeulGUYAEYMk0/3N3dGPGgUi8Hi4hh9lEqBCQax4k4Q
l+IV7jl1Rgujz3qIg7RuDOX0CZORKOa6I/fMdh2VGygKjCBh7ZE8PcSGqXiRucB449aOkMorxwkB
DvpGv+rbhE/YNdk3A14M8dKyp2bvcpOkR0ObI1h36jitjyehde0wBIbNDMA3KXDEJ2a+AfWMl+p+
jygVBPRz131NcmItlCSncXIUI6g5j3Lr5goZ4aEU6iXlmQCm52ZtK5UK6S/Y1W+ymhRm7Qc34G15
CpN/icm8XvvuuBdPXmjpI3psA/Vmkr1LHnbn/KMiCdmZCSIWQSIkftclc6JJK7VM8jmo14cTzJDj
6hYVkHHCPuDqh5d9jqT7TrvLjmZR+e2kUhOGdOflHs3Y6eeneJEVMW4BoX9bPF+LhOGN2JkMWqa7
2jZQxUXhIwBAUIgSzsD4bDEo++fFLoozFqNO1vJo7dVPJW/7omxxD8kWyVhJo5eGrR1B8HS/nVYD
el6hSlNCVQBmybVBb+ArPSvbctaY5bjGq58mo91unoHqvKnz6OkqqnzpXC9pT6ClXWOS6Xkw0zd1
zwIyl4FTYXk3stjE5EMuxn/wSdTwCk+dRehyolvTC1aVeey3ustoq+IeJGygZdX9mcDw4JSWAa+t
4F0yDYtuH3YGuEqDnhrfCw7XSX22/Y8VxqH2AfkhEsRz4zqANUfvf8SUAz10R9vXxIMchuS8GWC+
yctq2sK858Vbfxp2nLWCAxYz8VLxbi7+Tx092dH0XbnzH5D5FTygOi5+8xHPhISaLcyeLqLoly7x
Rv1BV5gUy4noFWnkkXqmXwOcP7549YAztKCsac2zIGvyV8ifS58rvVkQpnYGfIM5uiGDi7JAcqYF
VNfzYrLnEOvXcn+DvQy7lEtmLjP6/ncsllLHd3MVYZhViSvrYsiVyj2eCK/sA10AGiNMv+/3Jtdu
S7zHcalZsKg3Qrm7c+HXTPenFAk74YIoVWidIZpba9RBugi7flPnbufvbczzZOHbe9o5iK9m1gcR
jQCegVw2oHtqyYJIgb4z2JPKpUpNOeZATS7HkS9mzHC2MMpI486RhiOprkSep7nGPWHifx5uuhFC
+OILUP0uRcEfFYyMg9MOcIHL4raX3nqI2c7YzJFfoH7wfimXLAZM9MfsCuKiqfBhQt5AVSGa4VbP
obobcNGNQxFXUUbWcEzu3L6t1UX/oNMnEgv7uYV0ibgweOF9WRctZeptUrAio2a09j/gWh3dg6gz
EmhzhGTYZEQ1S0p8KmUEbUuBqLNJHI3LqwJdXVdVXFrHVuW2jzjDPdhnIV/JBKmtlV8CHZgfjVMe
ePHTvTs/eTiKn4pSsV9bK/iJWH0vxMPZUiGnwsdR2Isn4nHIrwczM7bCNvSxaDiLeLA2MmEiOEDE
nsZCpz5h4rK//7ozk/wGDAGf3bQFiLfZGkv+pG8/lLR7ZM0ONr2wDNr63afrcog2dOrGKusYOp5u
AMF9sryJ/Wb+Q1anIoOOWqdDH/mgL0dvcxHZXX5CWYNOOzkaGkzZOyXIR6t/zhAKbnzJuQUXkKJp
wKACWmVDNw1Gd8rC4d14SgZDY1Yd+DuFNKhiO1xOgvBDHd3bvoh4FSsCP+p5XyS8gZKsuNfao1qo
klTCFXYn4q2uKYdK3ayunYQUcBaEz87jw+dSzaebzsPPOAKG5DdC0U6LE2cU2auibMhmTFKvAQUi
RnDcZbPZMnlzayZXlRSWeBrxTgXOtVI+TJGfU2Pbod2ey2H7PQKjp8/7n64M1hKc4ah0N6Ed6NZC
yVNn4C9kU4kH1tQ9+WtAsGNXTbvPqZr7czDPy1pEtt8Bk7aknXG2x2zE+3d0gt1zvJccfqRmFUoa
vLwH7gy1zmyq5jZj+lXetXoX+lDbUppdW6CfhpzLAt7nBFSCIVgby+/h9785kLQktgPsxc8yF9BW
Vy3f/QSOmQd/nVBClB1KBPz3nz3LdFMCFk5OL1h6HhF2lXq7L17Hl57E81o/frS0F+xpT8mqnNQF
2fGDO7vXYZf7RosNYeylKTj15bZ1cVZknvSQmIqOyDulgKy1+5FUF9jqAHKyPbGixw/+laB0hlTO
REnzvbhLs9oSVq0DSKolnJB3ZvpXOim33s2yzGqShP7jAtpmxQAfALFUjX0dF+orhYeFgtsBL5pp
0E10yQhwsMz9ysm2OZQIbhcW2mxT6f5GsS8QWe3atMWtZIny3kByiqmULABu+c1hkfoM4tx8ohYy
A95PDtX8kCxHg28A9nkrJsZK7yh4WNkjWvzqOAfrPGshjeQNMn14mLYpk88F3XVBY3HakiorUIX7
tqPySdVV00lHSLJlNpM22zVAtH0YBUcu6pfbj/m9gMWuVyVdXLwiNxfoo2hHnyzZxgIjT0vLMy6j
xc9quuyruQgZb8pFlJ6BVTDQNRXM06aRE1KUUabzTuShEv/5sFwfxk26rFRY4lNe7Mw2JdaQsviN
idtw/wyEkX6IxyjZIfFjqmCCKzUYUXBfXryuLalr9XR+msBOqkCbjmQ90SX0d5mRZOxaTf6eM1Ja
D071YRng6HD2C9rPiAIrSWpPTmYmixUtZVbP9HbqxPzXJ/BeXIuJZQlr6rihtkbvB+OttVFjw6fA
PRgzixwfGQfRnWycKmvsyar2WREkq+4IF38znEZl59xP9KDouMY4gB16kpTUL6wwrjkDuBxaVFvJ
Rfqu8RcEc9BY7zDhNbG1xB+AFedVRMdQPmiLQj7z0qlHYOmhLGBzHxATAqXmQKLOw9MlVpTtDbJF
kPXqUq3I8XTs41noDrdCCwDkbqyo54/wsaffXs9/DIvsom4HFR164KCTLHB1aLke0guS6XjfNKXz
Aeq8WuSLCVGCIEoKbEUpjEQfjbS7UOtmTpUvWRDPle9CT7N6v9G2Z2dIKH3iH19eAv95bB3CzF6I
LIV+jGiZA/0NVYZOPGCvJ5g2YAcStkJ4eIctGChHFajZgvQkQT1rR63n0357zJooJaBKWrB0LrWK
CSD1+MFx0qlfZW1VMgFo/M5euaWpD7cgC30bB5ZqNNdTHG2wmaIrVBeTNU4aexrQtqF++wVPx1fK
q54f5Esmo1HxKHa3tAfOm9KsI/bU8pLhkJyIkNBAQw5z9599NIaUiBu5lIjpcB4q0+Gw3N/woVE5
Onik1zXLhSqK8wbNqfMEVWExuEvdFy9CfCikgitdEyX7nhJqX/AjhyzbWZpiwTlFgwl1yNKTYDGm
gue9Rjrm6u+B7HYY8YyuqH05wVo45bw3Cyp2ZB1pNQxSCC14Z7f9EYJZz90nureCPryAUBCnx5OE
QEQrUHlFnHuyX+F2AxQfEvd17qjcJ2xh96doMvt5uNduVFFuaVxnEoLcE6StfdVfAa+6FjGgJbwk
2517hugWHGZjOYl0dLwbayXp07tVeRaJfTuCMkbACdNaGBr1Z8kWv8yg6BpCHa4/tYSEehX4CCfA
KXtHEgsT3zAvEX6bJPF59qmheJl+jH4aAK3PK0bvjravi9w1esUfX8wxYqLviWJ4pWxkpWIvpGur
rZb63oOgZkRzRr8miWoDep8FlKMdYUn+tddzArt7u8plSyC/iNx5WOjDNRvpVFpeESev3J9SxRQt
Y0tmsmhUvINQSzXGoSkV2LXw14cgoMWS+nDx5L8pwVTBHAssOh1Dez0iz5fkU+0RCKAycXl0B0nZ
9tn0miTR/W5VUn4skr70j8VDDnf9RFHKS62zKd8VCoSCZwOyEK1f0VPYjhvTyc96UIyYjDAb2kTQ
HTwkOAmmKEQqn9Lh/lJZugE5bTLjqHkGFWlg9RRzLOYFn1RoyOVbAzTSl7WQnSjLEcXtlYbFJmw8
zwcOGKYRchicLPnKSWG/NHy3EPQN0kN+m27wuYpg71GuMW38WWXSaaU6X3ae8b43c7sjnY4T6EPm
u8Ar5bYFxIj8MYMjR5XY8xEPSX5jcbVv+HKJMTS1llgxlfxf2PdGuwhgjav+XvkYvGi1z9Es2stJ
jT9dCnQBwRbYG8TODpiXlyDu5uI2fE/WKhNYG5FVjrPgnOe+JVGiSPXsFtt83DGxYo+k+qXqwHvV
Kxdrjb+KHX5cBcTvAzVDkSTZnkUln9/U10XqTJeE0hGt5pinN3D9j5vUjCbF+unESyuNLSK2Oqeh
bTUZXixcaOlMKcLsSLrNAXJhHnOwNgmru79zUN0CETCJ8BwVETSFF3SbB/kZjMfAB5zL+xxtgnDd
8PTE9f0CbjYc1ng/XlQXsQ+br+D1LmH2Dn2ENYT9ykcP7/LjjrVmJzImWfGXYVwbw1mkVESyaWP4
BAH7NC/mi8/o2ncjsMumdbD3jT7IEPsfxTrut/UoS6VbmJAK6Je07J88FkBcDGyPB5oT8FuTacrB
IigkLnIqtK3ybV101RvZ4qWYVjbuyjs5pFESjRc8dYa9WNk4uMyq+WYm5etZ8wP0cH/YLvI0cKxO
3Xh3nEVPNcGlAHsZValfWwJb8EvDhwfMgzg3bbHGy4VIk6PA5M04OTYEg7oUYcrA0i0B1bUVbrQA
SwCbmwvRdT9oDTe7umiObfsmBIoceNRpPpkUoBazb5GtwN1NQTqRTlMMkzx8BflVOZZ2NiiBEv89
0QtuAvbYCiF3tic+4XNlFWN1NQ3w8MEUjPn1k18JH8Hrfxf1fbBzFflAWSok/HtT9zIDqHj/rhkN
1II8TkJJsZ9Inm+9Ye6ddUvNP4I4AspeoObuM/qQdu4MoUmgFl+OA53qsNM8E1fXpeUQynbvtbxx
W0sZOJBIIZ9O82lEfX8TrLud0cAbG3DF2apoGBNK4DU+JaHtI7x7xIch76X7AmdgT1aNBJRGdolT
a/GtACPHGRI2PiKtLKySPiBkbMlIr69qt7Lb5qkj9eazpKeY9Ls+Vcd9hUbZf+0BR5KqDiThCMoy
ZtbCTJ9MKCxlQNw10mSneo8VepuUARdU661DYIdNpJLYCd5qeLNyBEHOOw7q2I1yDOsBQI0MROYP
f+XaOThmX27OSR4gdop0r3XoY/WVlAN4EskPqngRA0c5KOlW9f8Zkkfn8k2cE+5ypARLQ/wJk0i9
+xVmrnZlfAMZBhz05wh6fGACL9XARZzI391y+MEc750tDuh7vlV3JRoKCIIDm9eNCyKEk/X7axd5
yPuKr8gp5BlMd4+c+F4eYSRw9PQZ0SYwJohN9m0dCouSHeekOJihlSUFdre0FvF8HNxpjAi1+f1z
DbZ7Oxrp7VAIR+8h1aVebFGxMTIl6l//idRut2AeEcb9r7hAFLHkt2JYsH4ZvcIAeDiwKMcvarQL
6Evewm7hVjTwoOgeurU4AK/FIQYTZk5n0TEysbZjuyfOCLNTuXZkudM+KOpcveGU4Fz2Je3ziKAZ
3cfp+FMxW2m5O/IVON0DYvPFl2ztpzPV0odsuOo1DUA0jYHaSuf5xnA6p380NSRObJUm3ZCaxJZB
Ia8OXq7T8fJNN3YISED8KkQBrMi88HrQRctyhcz932qNp5k3Oz2cG96+7lRKy4+ihOlqlp+xsedL
2Kp7T1aHsd2dPTyC0GSvg26/0GftuZWcLJlyr67G3nofFhrMAuq2LBwkW1kqC6Op9l/X41JV7jyb
xWJijHT2amrYk3NslZ7G9OAC6XbgNobi47u/zNfROLR0RUpB//BgI5ws0q+OwN6YWvMENB69muPU
0mROS9A9wGrNotRlqFCzj+3pcWFcHb3H5sXhGsNs2q1U5wASZ6Xh3LnSvl6gVNYBiv/yWaA7bBwz
KDXgj6DiE7CIryj8n6unwlbEvUvF9jL3QWQh0D4gFBJbvMF4qdktQIymxNYPdppXt76Zql+INMZ2
z9RNohNFkmF/V06AI3ieExFyHfsglN3k3RaQlpmZszHXlJWh0WN29xK+YZfpRZ1JchW/erwtDV0x
1+6GtZrYWgHHZ5b3ft1tCxecUgGdZUuAJyrPbOlkjMMLO3l4SXcX0bdNtfSXZce18D4hGe30rpMp
OWFxsrQ6BxbtuQYDQaCyBpT9eYGk6pBmXxAjKFEjp6i+w38pQRqVZSURgH8aEUWE7omrUlN6KZJh
fLzbdkjIWKZgjTdeybGK2GZpot1NfU84AQLFsP67cKwrzCqMG09MHDdYCon1lYmpvA+I53q7wpmc
ZLjS8XgAFJi48eXbIX3YGqFrGN1uxdNhlFSH6K4Ul+72AEmyhIQ1uba5WteP02LKb3ArbG/zMibi
yBizY6OTm175DQcteAM2vQfm/JnJjLkr0KL9jAwhq09SRiQI1/pfFFhgXfjGO09SnqafCB2UR9r/
ape6JADO2vK/+gKo3x0Ts852uKK3yKKRHSZo+tmU5K/d4saqE1xTLzMHrYRLm8D2BUCAJCkylmQv
/VrVzl1/lRaUmlT8CYS5FM8jn2lCy3hIlX+8izNMruXj5wMsbUdUOfG8w+hVYOgdX9ptiBlg2RrS
gxlGvgBGzN7mjgPD7rB5unoEMWcGgumCr3vaF2KuOxXMdj9XRD+mqq1qlpDVED2qQ9e4OV3LIYtL
yXPaysFobaoT89vBQrCcXziBJ2QaAUW3e0KbP+KgTxYeFBkh12OwWCULLx8STd27TnPp97Z9dvcu
zTNKn+l2SvUxpMieaM01SUzU5Uh7tgmlhHfYC/2YgT6Czzxx1ZCmclGsyuhllsFWaiAW4ftld6cO
U0IBTghF07wEykoqCElGfwqwyKTof8A+cWFpw5qEs/dkTBsvoRRrGDJChybIZW1iFENGogQIj1s1
B7i+F605dpZE70XzWrOjbf/u+xojmi3iUqrI1qQUI3CcRi4WGgzk1pfdQBFNDM9wdWyB3pM4X+Pl
qyt+y06DEUz2WwvBWSL2NI9WRcpv4J7ZCeAuLpW2ZXI89oXMm8NRL2pp+HYgo9AJ2wnuKuv7pVwe
GgpASkxj6F2PBJlD/13XD/MzQaYVGoCIvECf/eWXP4cC6P1bypnRzCduXOF0qdof6+JE1fRb8Gj9
5Gq8p0JWfMDH6TF/+B1AJ+GiOmSUoe3NHlHS7Rx2nSXdwlZDsvnS5mFj2niCB8LXqbyJR2SkNqC8
mrKXwg4kKNM5HRphMKlCD17YKodCTJF5eF0OTus3l8b0VI7VsONMu/FmyNlQ1M8SDUqlsTidqR6L
ABkaFvnMo6l1i/G4pLm1WGpEW84Ad4xysLdLMbKXH7dCob5RlIOxW88R480n7xZee/7oofCNZo4C
TQfPMA4RIgtRGytefUtMQKcxzPUa+qDhXDKm2t4QJ+Gno+M5KQvAk/cwft0YGKcTaKXLFlCh/VOG
kKy6dJ1JTCM+e1cxssrvDc2OKVRaQ119bQ6yBnepAZqYUyv42Dxe6q5SHGeW/z2C9IQ5Z2fFnx1J
e5W3mmvICbHoSyMvtwZ+ptLC3m1PaP8Q/Oi1I4tmCulExRx4vE3z2w/GK2oJr4ZvLmYwF3n+5GWB
8YpeZkhsR1UcnzwWm1Tvm5li8Spg53dO/UDdErp2ygD1X5YVDbm4H/gqZdFEAUEciPm03+JytfF/
TUm/tMJUMCYVfQU3WISH53237Ky/w0xWwy9sgg2Os0zCUAIzGZUrFaw9tJaLEbW44Gnx6T2Wgker
lzJkLqYlR0u8j86RahTMoGiAD/fhANpsTu+XMXoxKkKOKtszEi1gdSJmbcrXHfdgjb/MgsKys5z6
ibnE3HikFK2pNva85HPf+b9UvM8G2VtiTF6NUxVjUdv9fDWusA6bSErPmY6ouyPJmKahWCVohKiT
M93qRr9ZBeyTIPxyLuP9/r3ZWisamCRsi3J7+UAhjgQ6adeeXKdVweA/zANDLSRhijMGbGhq87vp
jtIpbiPMsyLp/r3pilx/2xgYPrXo/UPK9lmE4uZiMQIk/Sz2+YItOm71jtWS/0jp5U9nMNTaZJiR
W9kDpX9aY+nZb+f9wyw8UKk9Z+izElkC+Y92oXg94oluLIRVmCO1c6nX2S5lR+iXshTlWFsdZQPF
AtauvZksa4KJg39fks0c04zUKfcED/WCRWVRJ7pCy6ql0H/DnMVtDPM3RG/zFCbxJXJdBgVkTav0
9TdKQHemNJ1XSYwi7uIeraqC5GqUQCdNm6HxOfwQTW8+R+Pb065zQpKU48nUQX1xO827zGw4k7pF
2wR6BMvHqu/j7Aa/XOnPiepJyUF8SuQB6SNRifCbLaTveIOLPL26fzkphTa+2uivoZMtcelxPKpU
sOpiF6r5GV33hVS+hzSpW6/rIacHohzlWIkGSY8QA0tI+nL4cxTAGi0V55rs4JH34DVzfnJ4DKxc
VPFftO+U6BRBpijyYRdteU70C1etCviWyXK1OGrfe3BLnSzoobYdcd4qa8DTYGCneRpmR9PG5H5s
Q9OYPgzY/XvBeoDenPQH6IKI3ML0MQVXFtbJ1YSUrdNx4+FHP7hvsMoVgFJToUwSbMhd0DqPExIF
TZsjGk2q8r71f/+H8TsifYo7i8o8/L4mSzlC0OsMWLGP7Y7zYh8TN0kzsFMyWfcMOgpz5HbblHwM
vJ9f67481YC0Nv/9qZEIo3dEABZe+DDF6oWEnBBZ7ZurR8/OG5Uo/gXdFgs/xkb14Wi0vglhOln7
n2055VGyfv4e0IlGlKnNpW+U6Pa0N7Nh3IFe+MgUvpJWzULHBrv1fHo909bJpnNmBcPuyqcUW4O8
K6oVvpAX2DU8l+cdZeA3fq45p7kvuGP56LGkn3DlVJM6QB2VtOtFrQZF62rQHKTPDlptHmTV7C+6
DrSmkOLx9XxD3kMbh62EXfeqaWnPYiWys8/7Ekbe0MreiNSVk7vA4tHUBdTrzauNrL37YpS0fuNu
cunNMrjbsA4Gs7elvvoQ4N6Exra/I5POKvl0i1lX02GZWlxoAq10zQ33tVFlLMyYvY5fEq+YuoJD
bwyoZC5CpKlhq5B+qy7WmAP91YdjYk94SGquWwa45NHuVs/YgEJuRaRjsjakdILzAz+Z4KouEy/3
h26MnS8Eg8yVJl2I//wLsKEgHho/EGkdctCNoGloMpO/FdJUorF6AaDFFVeDk8A2i0r4x8pmnrG4
kYV2ibBRvJJzl0D+6rzX2/W3WJVcR19qUZU85O1soznvGyOeDwiMoJQyHAT10oP07tUciT3WfUZ/
gy/lyAKNsxQVv3mV65TAyqNOccJ3vJXx5UrbtPsLNZEpU1+P25WSJowHnNDzize2muK/mGXx99yu
fi9o7vzJcbMvTtHNX11K9lD5OE76N9pLdrihnP4RSLcX9zUTCi0WVMj5c0+liQvekfx6AOc5lsQH
xGNfZmn26DUK98OWSJNEiLmd7jG8G7JzVk8I0vchqqpS98Axj8GUdtE5pz9W+I8y7gRFiYYH1aTd
Cui5fIY7exIQJ9P91GarLb7jL77l7YRR8OwzkmUTA/g0kk48n05ImeKixHaT0ugDvPj3aaDHbqxr
P8iIwJg6/95VPF0E/Wc+kVlWbhJKZ/7BzJYo6ervNPBW+GAcN/2hJkfTF6ZD4USKbo08EUFJJmLZ
UdS74zMtUnXgK+8e7Odme/MnHUE1M5iYRYC6oY+ydqzM7npuTbpQrtpZ/fBkpBJBLGOhMslXNCEA
U5Ff6Mg985HzLe4QtCjTfV0s8ENyfM/PabLDDlpSx7tdj+PCYYsRoBSMgDTiaJz6cX4gNUoefzoZ
eDLPM0fSvrLuQhUXpEg36mAJ/+K/EI9fTuAarcDhHItx/rhcA3FTais3DAGvn23kH7lzS+fTjbOA
x7cL3NG3sNLwmlTBvN1Dkq8pzj9sXHjcvyUQ8HitFbyFbXGw1QHQ5+dlllF/R/PZDIaEQ5a9hkIT
IGuwQ93y+EL3VIuE22LXvw7ifLXxOdBRF5+/ZgBCFlXomRk82aEb7ZxZrcYY4FLFTIfUu+KSQQIx
+d/dCNs7u9+Se38ICIGdWxLFktGdxJZHdC9wgdOjCZkXJvtF5k7VsMAV0lwPYiuh74bItb/mcom6
DOJpD992F6WLnsEkCu+hutDz5Sg9t0xrnglv7pvxIT1yLbsIzR5SxUQMxUzG/LcuKRmgv5mqtSas
R7KWFkTkAwN6QRFwTCS1KFWTQApR8ov9uVcsxV9dknUFwbKxdMzCyccZHaXwJOFw7lQZLJgYe3Sl
lgpHJzZfdOlSMXcU7kkETLjpnB55yG0aA9B37PXLTW4pfO28b4IqISzP4fXaFDq/WtKvpDvW0D1W
Pi2CBn+AqyAlPTZAgpqpaQ+YewOnjrj5sxs0VfH4Yqc7YeTHSavXgYD2vCOvjXgAZJyNLgu2NUWj
Dq5I760WH7b722yFBmuTNsr15CqfJmMWBkgtRenQbMl5DBUoG+iJ+sF4f5MKdZZ2tctoOKQa2UM2
G2kSY5dkmUXmgZvMcaIHI4v9vrM/jky5Y0Jcxes05RlU4Uyy021lbYAHi/rR9twSRLx6Lk52EDnC
Nxc0bCPxY4DFqyJWE4vlItKnhQr1wbNDseLH1KfG5gOEbv7URj10bb95nQme6SHNFZbKj25czk+V
tuxEhB8wUbSK2CEqu5V9Y2mrhmjgsjrg/IF+W6g9UL+7RGxmfQv2vcy6vyE+kZbl5unTXfxAAp1J
cEjH2Buo5xPROs6dJbtV7JamKu6Z2XOWjPWUihd+WZS2ZCwXnnGUD/ZV0VCvLl5OqEepABie83XR
/dCPOoyqdzgcCeHEcW57APe6Pm3xiJ7EJS2SYoRaXUzUEXb3Xhs+i8MLat2/5VBejLuuJWG6/Vxm
RJ5mpy58OOnNA68Gtr3yHaAwzEqlt/VmT6b97ju4a27eyLREjkoFf6hW/s6k9NbtZHfbB+Y/01AF
lMU4X+4nLSpFD07JA1W6bDyHLrILP+1FoVgbs01LQqHeafeyJjpLDeDXKJmQkeixsHK9NpHSoBLU
rr13RNa+FQw2EwVi7Y73aKOdbhHo29siyjNYGfZma3Xz0WwEw7jdbSiL9I8CmNybsYvp15evyvsi
88GdKAbOeqiEBgs/w7S3KLFXo5eYS6HoPBKxcCnNkTLzrSTYhHO61lFcB9jVPqy4Oq4JyoEVn7BA
asdMoaZiQA1NDPMZzA8f9skAYxJP3PgJAkHfTZiXB0uSVTDF/Xmfq6v3yKtX3trk5z6EXOVcZt3Z
Mcfh+PCB6uaDWuNMFYZR0shu+HB0DxQGVeEKrOKurDmyVl1ErRlrc2bLhNvRCCoVUXIK6RcxALOY
wwiStPBAecsSOp4457wOCVbGElvr+XFVe6G6mVLN5KNRiIy8e1twJA48R91PNB1e8vI6Y0/FYmgq
WRt4BXfj3mkZA8JQAW7SFNjdqPzXfRYKTFBl8+0+P4Xzd3LCFqHquMsfIOYuuEHuQbuJjm3uUuj7
+kzVD/BNyc8r1MwLW7OXdAMu4IWV1UJ/qp0yxKKroNMlXek8Vyi6GtrSehX8DomaMsdKtgSYPMP8
BcN12FMPeIRWW3WPN2vyMGpC1WVcIic6uHQUzw2SgCY1KmDDM4vrd5lgIwd0Y8f6twbmp9ZHvf2U
YFLYmNdfp+x5tXDfrQB74KsScE2YZYcUmQ34OgH3Z5RLcMwgTQkmaO90qmUxGkGKVu4OlbXxsjJy
DFrqW1CdIrmjmFBjx2g37JPHwnLeaW9PYTAp7MLwOvD5Al/vUiKcG/acE+kSFgumM5kItNRlsV1I
mz4UdHxZKhSR1ktJvkiNvu2r1OxNoG8jMjpP++x19RsJ+k6H+KI6ancPe2qtT74yXgsH6erzGqqA
oCE54bOSgWCzlWOTpegPdvERQ54QfzlIqea+ytcEd4sZTSgRda2qTrZhgz1ojRSvg2IPb6kJyeEU
xpupBnr6wf+UenWLW0tr9Mmn3D+OdGy8rIljp/68hpIiurhZ0LNsn5dDU6DVGVxYTaDlDN14lzCP
17gGBBWrPeJ7scpljzxyayBohqGYwAjvqfooPOLGF1FtlDVlzjkkIUd5cLrtIYvZcPodYW6PfiSB
MH+RVqqoupmrQyPMhOeSK/iXdj0B10Os83irnufv6TCYun9ojUXcbeQMtWGHk+wVRtAEtG2VkuIC
ffRFtMgP2rSgP0l58C7aFCfsjZW/nlGlOwX6DHAygNbC2twOz3Z/s47A+l86O2LMkJGQBfrL8oBY
RWFIYYWESu9Ilt+Btqp5B3iVQPryZnyftYdstzvqCTNauxh3FZucWSuAjzEn4ApRdfam4eZ+Fk/V
/JeRHtnzgCsjkla+rXYj6wTPLe6C1UkVe8tGBhLuMXFqrS3aVtY/Ogygf1/n6RTXwY8n3RnZrzDr
VHAFemRFqM1NoaZZwmCNJrXDABSRIwFtRHjjicPqQa8A2MDw1o2YZ08GjH5/mRZfoLsmCwFEMZ3h
keUx2e3s+TWDjnVmV6DVBwKPE1Zkmz/ey5nDq3q/w2sjo+XT8wLteYvw5bRUl8KF7gtswiqbAAY8
HRBd0DY/C0PHGDF7fvSZmBJzYK1hNk3B+s7OREWW67Ydy7jEACDBEDwWlYmqph2TkdEFf3vVA3t5
L37euSraYxSuAfE/sfITRr2bSTO7cw9dTrbkcm9KN3lKy9WPkqAZwyZOl3MVZ3hVUymA6x2Zkq60
SwrlN5CDotCptltQ/iOQeiKwEDwqCYWFkqJQCoIzyRW+YrLfqnopVqUZ9fpT1hlqvISeG2Y+E2ws
4i4KLo9vh0ig/+nsTu9WAnHZXNU1NMO2yeZ8Ow3psf2X+/DrFvkoKoC8HUU5OQUZM6YZOIe3pbaO
Xh3UhhFK5y3S28suEQEYBQZVDzBWE8gzdmp9Dc68Dcsb15iDnoFtzXuqd9iqJUncF5eNe5ePRP1W
MiONWRXPPsaaPqCq2FMyD5RSqPYqC85FFCjSrTTbb9K1xd7DyYf77dbNYsnn5ka96lNykG/Eh+1z
ovf0F3Be1rfHjz7KHBdqmpAvas2AlypaQP5It+jKg/0QjiiirEmSxIzYjJkxrzluCC5MAatCzGbx
wC8+yPhbrplnrcyNXYcWYiRGpwu3yBYx6Qqig8kngTBxOxjjL8UCr8rxhrJ/B8iuh6hunkGR+AFp
kvSXrWjkF72GeMbwNy7GfTZaoyGH+WEnPDx4+kzwENf56Y/jFkEgdlYu/ROscfHtPDLggjBf/Yf2
dCz7mDESoU5piznDgqArNXEMfhWaEyP4qUKqRKVYOqSCVyoMIi941GA/s+KKK16QbPh20a2Ai7M8
MhuTsLmB2uHm4nUuKPkpECRkGc0RkHWfcwOCeCI4cTbO1//yw6F6UGpt0j8FXp2P6f6OmKXSvSFk
gLXoGov0QQPfshE7/oXtJkl4G/vbQDoxGx1yXYjdHOCXtBRrFA8QLo/Q8Dr0kiWiD9srB2+3jisr
Gfwbm0XZTmZkAPbTn3VFFvuZPs+nLFyQIOoTLI0D6gPdDaGAGuJXMmL27hybBs3XWg3c+QblQsRt
sLbROA6DfnegYWR7+Gcr60NB5QGEKaQcef7TVeXiGmwnqCYNR3YLQxNl3SMbGsg0j8uhiPzMPEa5
XZ8yKcoN33DQd6GvHpQGFkI3rmVv/V1C2mkime19dz9BC+hAlj18PFTJ34fnVPmd5e6aDd3tTlYo
Ob1YUYpZG8DaawQ/ORFlNGxJ+Pf7Vts0vxuO4bgAdlyg2JoCH8bnsHBW4cl6Xkmn9oMgOraqngzG
ViLf+mZclA78GRJq8YNG6r8KHotH2clJLADeI0uXokFXvdEYiXP5ywFc66tbZKZnyrYzZ9cvw74n
zwxUcCRuy/VVQ1cXA3EX5CAJaGA5lkwiqKMls2DBVFeZJmd7cXiGiPzDKxSqrLHuhmUWMvijjMFw
ETMh6mlEegxVOP3bWCPE7oBSINBOkcDmXoVLCz+k6YjWZjr+f85a7SC9BbcJusAFk6pR9dz3FrAQ
tQepUDUoB2agfpHHHRnH4m1m75JJsnW3dutxhhQxiGZqPftZp+zo++0JDZzHfkkGULlROcQ33unC
TRA3Y8QlU+AQL2V4gbEF8ZrrBh8f+Yogc6Wf4/XWCSzF5YKfe/89XaovDL3PpSkWqY/QuA/8VEtI
hR+xg/CYOiVk0GjB0aWuKw7m4oryuQEq8q+SUPPKydBE9+Nb+dEohFASCZvJCfHu9cHihNEHzKzU
zmd8hHxUS0vHIESkn7FGTsxxMcNkzzfkSIWjYztMzy9QE7KcXvtbLe7U8PLfJwgP75TPv70o+UDp
PH9nTCByJb49rFMCZTjWAEkSdxOu3BnIoGDFsYMLtUZ7Hb8RO8SecppNtbkHkIbiiW5J6nuyWvd6
8ievTtU3ZaBXR0Ez8QUcKYiw3T+e6bLaSl+Q7D6F+JuWkYwndRNPk8paT73mTKtzhOMVLZXgkiDy
CnoEeEpQdjE6SlpSxP6CHTY+oqNZktVxvh3n7pEajt0stv646Sle9i5aGUqoW24mV/r2mO/I21Ho
dAZbZsKFXNcXpc1Ob7BCODRYwuVDs/fYuEpW0vZGgnj7luSiwtPzHZhnE6Sh8yGwULC3294h5V8U
R9qv+w1HQ/vE4q7q6IvLmNfbfauVqfPOj0PmN21sv1bwTk+BRlOgz9sJDKufXrnw1pKz+4qxWno2
trLmFrahy6tcj8citdwsdsSmFVRwABX0l+9Dc8ZWlTcfCfqxty1KPjE39/oM/zLGiXyot4Tq0+H7
HrZUtd49KWR3s9WdADuhyLR+khBFDWWRqOSFqAnuEJ/qiu0ELkhxSUYwF8lncqwssU1PRqVT/n2/
vKMk2/WECuYcJtKMcCcaUbP/sdAbO/EDULQOSpfr54Du9MT665pXZnLnC4+t/oSReqEoa8d90jJz
0Q+YOYS1jp3tr4/h3Qbn5BELwTb7kpYzBSCsOl7Naws8JNNLUxMi7G/NyPZ1vZZiu+dev4atwf18
NPfxQsyMDr1j289NbIBrK6ef/Rqq1PsOxxfJDb+7Ve+u2kUIJAsqdQRc94IWefpOi+KTqDbXJb3l
U1r9wr/YwyYUhkokQS3n0Z167IOUWCLfseN+dVKB/qsOdiwHAiIunSV4l+/41gRmFiyzrLTsuIgc
ver0+7YRTPdekZydAokj0jkeivaRYmIV9deNp/mvwK+vzZh+KlXx2cX8MlsCmV2blGDfel+hQ2KY
YDJXp22P15ChDCTUieP7XArvw12tsqlw+nrCvlLQLC2nV569AqqNJHPjFRkpzxNyqZTDs6DBmkrd
UNDqc0gSLbw0iqZ9jXsQwVoKXpM8QCPg4DTApDGTbiUGAiWhgKZ2Bw8Q5dmD8ce/Smh7YMNb+2LZ
lFclWnoq/LbqcO2kxRoYc18PhZEulDqxZVYwDAxXf56nYsHZ7Ia+joYyuusduogKXLO/p+KaSKrP
9HkguSxtcdwdrjAzdtQ1C5tM8HP9N1R9OUbeW4VFiccq6yyOZPeyl0VNGHVQR2xxbj4qpYXZjLQs
KpV7ESuaX4SZYSU8WM8O8BRsCK4Bf3d/TEjW7AVbPSjnY5QW3lbACQ51I2snan8QzIBSAj07zPCv
QucRehiTMHPCzEVlJgQ1cTCAtXUjsMk1B4joTZXsUmstxeZmfR6i0VQqwe5g5szFiA5bEsXCNstA
vw60FMqtr1kSUsK8KSrKVCno4VAATp9iSZSFtRZSZ0zYNaNDTIciCB4YB5dGLaKHOp/YuiBua2Q3
eFyZue0kL0PwfB+uj574HnoCZhQM/CDAUhpQgrKy+vXr2Y3ISmQYEWdAq2upcNFIFCidZHeyxgHB
B8xmO1xGIS+d6ejI2ScIx6tx+9uIPuY9XY5sOTaykNIvQWxbBIvq927sFxd6ENBSD49zZrc5Jy27
iwEUfTSJF8fzZ+0kdsWmbAlGnLJXNeDsW10t5K3S/gAXykDCkA3A40j2DGgjrBEbbfFwh0zzyLTq
6Zt2AOzPXSmv4so46tIHmx5r29b7gojMK5HfJ2riWrHeIO4PVEm01vYJ2ET6YKECuA2+oAAF4V4Q
jueyWYfm1sOcUUx4kwQ3g8OBBXoGPGrJ7Wp6EqJLbDKLkNf3GRpP+S1rO1ywP+bnkbhd1FVQyS7E
WTU3zmllWHAxzz5ESwoIzx5eANE+iEA6ObFhZCGpoz/zFhl7CVRFzOZ/ANyGa3J+mopiaBVqlhhE
yTnM64Bi9necgTIKN56VWWG4LCP8Ug1rUEt+/NcKg01ozXSX3EA1CV2u7EjjqKcYGaubUJo/GO6v
kf3nes/wxf/Q486ncTsCp+6ZI8Xi+NIAI/K+3ZUyO0nBp/g0sHrZxKgW8m8ivDDYaw6g1vSa0ute
nrU30xUE7EG5NdPki8SU4D2XpvJ4JZtdVrtm7bzn1BST8PZz+1gcWuy5w8CLk0MsqYbVdSH8dtj/
yc30n8yFa37GlGefixN/BT0pboBgvpPIv1ToyGABNnR45Urv80xWp1832bSzDtF7y6mAXPr42GfT
X+Oxl9b7xEE6AVbrOQLchFL6DtfttQqRXlfZ3a62Zw2OBLNSKdwvKkv/hKEflidOCoNR84BaK4NM
YsNM0lHgz3NsScMKy9g59qHF6B1mLa4bhGzh6XzQoFDzzKR2JeMm2wC8dDQF6vGkPfq9/jIq0P4y
Dr0gSoRyH3evW+SEcd5uzddVAbWyPEdxXH4n8SbVDA6HvwZKVBGg0fcJ0qV8MeX5JBlgNtzoZ7O/
f0BhHXBMchFyxvnNtUXWAWgcI72nxBNNBR+8KOVwoiFxeLcz8E0FOXuXsWjj7C3Vg/3NY3oiJMPC
clBEw3Lhz/LfpzmQ+j+2/zsCZnrLjdbziU8PFtvx/bAx0MSWjDx+1zPdJfWxhKW6RTRMeT53rxaQ
khahUSA/vLLPtk5OmDXdAgjCTzX81S2YHWsMtEoZgDUhR91Lp+7AU4SIsiYCEBuMIFOTSJv7/0KV
1FdQkwEKMRr0hY4JxctiLZD2hxV/OlKMzSZVqKBejBTh20bFMJoFZmIc4hxWTFERRuCtslsMnVlN
61+ZyuNxgaFL8EqnbqLlwGvgswYmJkAJmr85onf+dI/y16aIaEOL5cgm8xjxikLpjHdV6x1L5E2J
ubJINH+782CVlfPvpGALZe6mU/TfJB/RWNWSrrLyWwazxJKkJWbgNry+T2l93MarjO25MQcamAOh
BPk5CGudK2VW1pTLZ4Qy/fCwr3x1y/ZxLjXVIU8pXjF/CvujnqLhSMdTpgydVT23lHbbnvjoR2uy
Rxp5HN72kHuC1hgK3TbzLnGwiyaVbr0Y5tATN7KU0vICqnVH8EgiXwD2uLX05NlI9xkV9JD/Osfy
cXl6VAR4cjYokUVndzN9u2WSoX8HF+ZIRhyeEo6NLADhbm2NHMFYk6a6wj/98JYSCE4XKhynY42G
rPbb6IOF/YM0ElrUzJSvJfj/yE0SmCxaRseiDhz5GP3ZeznGLKdHuEmIF8MwoK3423lMell3k3JI
aduhjg8CFpp+b09c1GdJVAlR1yX3RvtzSKxfEboHu4efrI22ih9t3uxxVXLqIoavIbQNa+yjPh7C
mdLN7AlkBqM28v2sCo6Kql5PPk1BRP+5oNA2LZoo0B3FHpiItVndRRFpMRqnlTKO6TLWcZgLYhmv
Yz9Q/dIY0ExmTtwFV8DlDtubP2zu4PO45vf9Bl+IA2eN/mB4608fqXdfRVkU0UC/pk+I3q/SbXa5
/yu+C+mCe8i/iwwmLe0ep1nSCLJods9su8pq2AI0pvj7JDRJhuncSr+NGm8Pln3Dz41KzEZHsPy2
AhQHGqtVl33AkN5BsWzHJKg3gUDu0jMGwVTkZBLjf4Ins0+JMujqwL7MelIwNDWjjOE5Q0hJS7Yf
1Z+1Q5ilFo+NMa5kU6tbMncGvvKqFSGeRpugsnixenToq6GvpiPrySlCUIHFLg61YGFyYqjtq0HK
T22vn4xHuIFfe1RST8xQZtVWqEcJXjvuIiS5qhXYMWaXIQC7UGw8FJBO/2uDXn6OZcVqv4+8Bv75
GimYhpkqMajia/KqJW/v8ogSISMKFsedWAuP/3EHJKT04cKrqYyZX8qLNbQ/dpsIv3k32uqL/N0Q
aSoSwrGGLhMXCE27ph6G5EQaG9d/2xDjT23C6LfLYQlyn27jtdm7N769U81c6hX43P6Su4V3tf8H
/YFN08wEnk1vqQUDiEXSvggTkuU+TaI8aMspRHztMNwI1FLfHzdOrLr91Jkr84IigSwHzcLIwqhm
GAn1njdsZCDVEZT94L5o/1NN+c/p0lGoNrILvt4SwGh1VZhjErgnaij2gJIDJh82T+zjEdGLPYQd
9zBXx3MDymhif93EoMwUDWEsDNDOVE9qU6r3Dd0OJimaVU2iinhH11TF14rKQOg931uMsKM3HFyX
W7YBFvnh5Ol4oHnB/KNGV35VJWKvR1AJ/nopiq8n642pXXwUj5TfKM9v79kGWm/JoQ2tmvnQ6V6g
Ys4X773Md9SGy1JPixKdAMT//CVHvCVwbJAe7jK9Co/nB9W0AjVP3zj0gKB6LE34t4xOnw+0+ohf
BVB4ZdZprHKnev55cuMZArOH7Cn7YY+jaTw2M4HgZ9ipjrsWEx2e3EimEkXrNgdlfiIha20G6Jp2
UBTH7zq7CRWC3wAIZbf9LSDjU6tHASorF4NJ3230fkkdlGwOSPi9GDia3QvNuHCIA6sf0o6ldmra
kETqcvswfRfxwXBDkb6HsCQwiEzbzPJRhBKk4TqBZ9hJsCu8Imklfb83KSQNivd0ONHncY79ceh3
vJjzeYaorDwaP+ygCgDAcluMB2cu74Qm7CcMRRdvFcFTYg7c1xeao6kW7k8Q3XQqTq8aUn/KvXOL
HbyiuqJymawWVDoLnTXhNEFQQzfoLSVCLXPryB/v6nCMBdLLYC9wU4ycUrxoIVzoRcST99iyEJ0I
7gVwvh7eynIukCNrqXlu3lqDHKGOYRccTtww7g+UtGyCUHNxptiQElsImaRfr1c5cnHfE6MHgeac
msmJ74JHn3Q/b2MjsR55VuY5mB9KDuMddkhlPBT/fN2NAmoAOzy8CEbwDTu+Wcjci7R5Opy47GQT
lBmNwWdM9KqikvWAw9pDwNyoNPZ0GZFevDVz53Io4/oU1eB044d7E56o8PDE9QI/yTgSYQK+45Th
/nkZjyo1XDGPlG8nLmSz+b9Ypa9uAoG8Kxg486DykpKF+W/8rJR2zCnTH62zYPpUOyyf8E85+Y/g
66Iojrjb/CKSZtUAmhMqUa8bUHynGK7woIQE4j6d3VmMjur92MiU0pmQoiFP9JLRX4lekIc2sqJo
EX8uFEULfvLyCERCecbblZ2p5q+UY0YSKHXTOl9sS3oXWkIiYDiEyQ79AtcvUE+q2A3XGUnRLN1H
E7AiXYOcSL0zICG6GYX/Fe+EBOHXCxT0TxWZsQhmG36vG45b03xXRFcSD/j2YZ+tlh56yCwRN6ni
mSvAPQGabxrOv+zPHitC8g48txtGf7H/kLhFh8pgq/Vtv6qiPeuxurw9bjJ4rowrxCbwVer83WL/
ZZYwfrQn3m+zWXLNjZ3efZbwBGOrVVUsI/Zn5M2gxUb+2FssTQOM7utL1yhlOcNNwSvkVZz9CZEd
DApt/l+yAJ2IO/1ZuyNDCa0jXx9YpLyuc5FRlHfqN3qMNnkXzisMrHxmfaB68+nwDuJ92BIpGH5j
DqMqU7n1roJTnRyptcIhlyXQV6fECfIAx4NPOFQQz0ZIa7/QMoevUW/cS311lByVHAh3YVvVFjv7
O8LcYJNJXAYoazMYVm2gQm/0vW1s5hm9ugRqj5MK5cAbeZ5/+eP5NvT6HD1fSk2bDCrD8C1j2y+j
odXbWfZ40wKBfprtwcgM94/EaK7cuu3+qsW1lv5vaiz+Gtp3gKpPd0XTnIJZ1b4ALRrrrNoQw2a/
6R6KrWh0HvacW2BpQ2zawl1ldeNjyE/kxS4uzs/YDMFPkU5jIj371KtqNP3WUOBB7/fD/z5duDS6
iX8z2e3jfYoW/6VOXN5Mk7CQmxibVWJpOdPX8Lwv3vTHlmaqt1k5toHERNNOMwIKArbURKcOPKpz
myFToWNC2cF25Q+/ggCRV3MzcaRkUkwx2WnV1F9wkIsRMIO3fMhKX/VReFPpvhbsFWYV9LJ+8Gkv
crMAu1Xw9Fvn/tPPV5VvLd8WMnH6Qrnfo3DhR3KH9p+Ii/RdLDUuqXvTwSmiIJRwKbZHKdR6hAxb
Z0SmlTu3Ot6+udwmZoRhaO1GYbiWvp7gxL8dXLhyf4OlYJ6YR/RCz4Qp+i9VaWaPZL0cPN30yru9
MDnVdNW8aGZuQpNOuoLWA/XGEI5KqmLnyve1YFULlGGRhpKTQ/3sWZ8nprNEV4A/EQVEO0kuEMNs
gf2Z/6gUO0z4YInSUQO9TkuWZdMcE+nhRa3a4tEzR44uw+2RAGcwfFPE8LlYsEGqOExAjuiqrnbh
dDxBnaG5LrPvYk8yEa/q27A4u7Jucu65g41e8wtmhQd9AbpWREuHCMp1v6Kr7oC+IMF9LDx2/OjJ
+XHSAgIR2KsprWFauDcrAlDz4NtN+N5LEl2ijVfhUWHDlsCg23F4pbRpUa22x5t9sAofuKAIlC5X
cD4VIMjtMmDQzHl1SNiJE5SeFLQMOSgdb0aTk2N0IKIgtaP3DzMoKy+z7FVcBZXhIaywKPTJy2o/
VJ0Iy8FAQMtPqUoU/VQWysaDLfW/NfobZHua45tzLyu6xsP23+P5h6wmN3mEwH9yPrUeAAFW2qW7
5dO+msBfNsrr+SG1IjBbfHzL5qDgg+UVXx5pmB6tQGWMypuZQLM0WF3eppmg3qBWY1w7LJX1A6+n
9390YWEHDSkSTLDVk8pj50IC3c8ydPGUIAY33Q+tUeLUSE2FkFJPKqglAoLTFb6Fd1Qnai8kh9m8
PAww0o/Tr0pOfGajN7ms4vjXGFZv1bHV12kKB5npU+O9Aj4WPC2ykbc6w2iABo1hVyvcWHwMQ+kZ
6ilGBL2vDQNjyCsNn4w47TGbLMqUxMWR7FQwtX077OMtWDTaZTYGXKtwCou/ULE4QHscNscO8861
YPVGZhUFyjlZf9CT2efTVfoilzmZUY1rL5gD94GBolv80qdaqb6NcWzrtRzL9aiAU+eH4S74tAgh
2554+HennicxEybuPFNHqEH95dQvFu1hyOvNwsWZQs+61j0TbJMaEd/kGR412kDGQRWh3YO8zsog
SRg9B7LBjINpjEgNA74oLOqu+L2D/t27Kjusq2WDb8orh1oWtK9ol79X9G8FUi791dYZAPhG7jD3
LaKnf9gJfyVFxem7ZOFC8uyNCfYAI/PnZdNZHFKc9lXu1mnh4GYTlMXiX7ClsGWwoFZMFJGfTHFj
35CKELuVwgx84JnKd9PA6w2cdSfsEoD0WGxmKoHOpAsTjJPyVXvb3R5plkXgwogkx1pb0bcGHe+n
+yu8Y9RhOkcODfe0TSBNH9TtYreaUdlVJILFbRLsaSujB/AmkmVKXdi1gD+fPU544d6guJtEF1WH
N8dRPBDeZAcEWznjyUYeuZnJowMhNINh8JZOFqVp8YEOAb/GRuq//jDU3ZYaxvjHUSTccLHo6K++
m6aKLg+E0II0EIa8u8gnU5wwp1r1HIXcv3QGTg3G/rFg3OGTGtxV0lAe5gHQWVDnjVwd/yOg4orb
5oLA1RYheIJ/Qd3XzspxZpCkSBO6SBgpwnUUZFAcL9RO75tVkhTmJCvjImXnlZDIq+gaoQOlp5Eu
XB3PvLglerKYoXukVPXVbbAfmgo5W8OxzuhEyahzbT0DrmZJxgHxnw/tyVBnlPlyVvIjcsuyNoUF
5E1H8BteY6DImYOzYhyroDF0d5w8uyXtBuhD+E7v2P7FyfKEIz7nrJ3yAMWDU/4YcpBMGoFIwPXx
WEubYDc7vRcFEw76p9+9glBP3+aOe8StDy1m+63jkZ7RMP/WDUwzpV1Tf1uUh5NnCwxRQpfL3fNQ
EsXnb0lRdoqIFEYP71HKK7dBs3+0Kg6ceFn2KDEPmldjdOUl0l802hderUqF0wZpi/J7lbPqb3mT
7dTUD+mJOwk26X6OJxfGI2ZNzu5lJaOqFQJ1a5WsQn00V85afvl6/RS43FqKjoJU7uhwFSiK07qf
oACOnUK2XtWlU2Vz2nxer/TKWoCrzZnZN2p6NQidCSQnTLYC0x018js0WcyNJm842iTWIJ0NaytT
UmDXz3SHQb7hkx8U6sgT/TLVCqIoNNpVjNMR9keL4xlO5h7xDnuwB+lsXL2hPGKvzorFzgvP3YHg
pRSUrKWdO6ApSahmq+siEwQp2Cm7RdbW4FA3mcCT85ACX1YYiMFxj/HnMQv1/colhZ+Wy8s+KbaY
gAoGTevPAuiZx13f9IarqZ2HGLsHj34FfB05z0nH6ANVhMuJogL7Nia7QRDfsHvr+J7Knx+vANm5
vVTJLVkg1mFVroUsKin6xf7jWWd+jUYvvfeNiCex3iNpeAgGW1npUG19lVVzAzLYdlkL4rg7h0fu
3BgxWn2Tzbw7ueJTCgeYDu92L0Kcd+4Qj23czDd34pxXYnjMPzldc6vHdARe8+Hb02EkHGrxc39R
fdLoDq5sYCigR8N5w47eOuOBOiYDXJbpCMGYEYR+iZCMs33onNcQEmec357e1spGAhXSbIY3tsuC
hyocqKIpQsIfRrymP3mi01fWZuu6pbRlmmFGSggiRtFf/zsKkAt97Nej7T4eqyhFCbVieoZXkU8v
RSq/LfIgs36uxToUsxtc0Ou5w3GiD8ZHc/RUGTzASCcpmOWE2XUb4A5pMwS1aJLvWldb/8m7eoR2
IlrcwZuKZn77/nMrsu1ElmN9OjVeBMrme9n7FFgmmYQ+NONyWJT9gUHJzc5IabJePkuaMuwpkl5P
QFufW/aqNXk9JTPE+wqy6kaGt1KzOqG959E1knvwx+zeRrZqdx5eD2B3rqoplww++dJKh/A1XQXC
fTEYcpv9OK+P6eU52VmoZa6p2Moc2rYp5b+U2962kNVHPha6Ua0YsQ1Cqhc2SiQGpjgfmlqrpAS+
sFiUXWFdJG1KGtlaK3tjLlFr8prAQUYkqWz3zl6/L3JayQUAQKUgM/3Z/hOl0wUGsc1MA6gDMEWI
L2o2SJ2+wGM2CXd2syZSNCNGH2Th1Cqjce6f6UovTvX8ZzTB4VfB07MvweVsRGfA5t9qg1xmZrtZ
6/EepIe/6rhKsrHcbbOftqL57xP9obEJRD2etiOyCMkQrK80VdlnUfH2Ft5Y7lJdORBYdT0mjzqt
TavT1sBejB7qbP+mRw0q+JrIXGQtOaUsTFjRLZRwzlUr0ty6MfZZNPKqCS3ukNxNs1HXXAmZPK3z
qfoPXPk5heEAdC7lA5SoXdYTsCdTHUL6YzQZGGdFukMoM0tL5aZDXpQX8w8bqEP3NnxKcc/w/sce
6pEqKYrWwi+unSOjGTN3MuR27/yL82WVxicPTEYdE4/zsX8L3/1qPZUXbyIw1mVxYVJYKFgWuV1v
K//x/jlVaVTokLbF57hzqmj+MTmpjeWXq7bCqZV5mSu0EI7hhxEn6AKcGg2qqUgon+ZfuXgo7IDU
QDnfm2J8x4Vgrwt4roQNln55B/PBQksQxHbC2UYTtzgR6E6uBSimjHYdzQkwkTO+6irp0mZr89Wb
xjJApp8HF+kNkjqkaUCxhcetGnxqhxsWD0Zlca6VF+B63hMRn2Gp3CYviiJw+jsWKTcOeM2EuQK2
L+xT2SSwY6iFpHCgt7LAEkjmHh4nRf/T54vrRPQMcLAhyX+ash1UIfEcYbclTs8Ngx0HfKaMCyex
X25WpvblFewCxGvXmvZ+GEF/TGfqPMxwPXwIwhC1iSn6+NQgk3NtIFNxXwQ+/7OkMJklreTjwIUa
shzpXbHCbR80WX6eK5vcH0N3PlS+mw4Hl74k2jPiRvoqf5UQROxGKbTKubb7aQX/tkROZPokVh8k
v6Y8uXVgIdkaInqtfxBGOLYbnu/erC4pyg2FviRISpGL7R180o3C6VWaJuSeDugSmLXlB7DkEkNX
y4J9PSvzO9RdYPBNW6xiLKOFiN6ooFxCh1ElhH3CSIavNohVWXs0Bnuke6wKgdIopKbj24XQX5iQ
Jdhwf5YfGSyGK/2QLo2JegO2UfwPRmZp+YXJJU9ys32ARmpGvk7f9n36oIbzoQvQKySWX3xn2SKT
7hht28ZuTbuu/vbcHZrALxi9FL5/ZUa5DppJjOkrC/IQkYqHB0mALcegBgrxPrtp6Qid6nPcUjG9
U6JQFrMmS4mMJsdbB2X4DwxY6Hj35fzW4kxNTnY23j9PrHvdz8kfThRqWD8e21wGAVFHb3OwApst
xVSwvyhiJIF1HT6yWqR7V33+PWP2bV/lAZZF97lWvjr6TgY6BoUaAlPCol3v222Er5bdUXCagFDM
oFBE78WPz8mQjjOrTrvLLBrkPbarqcQb1R2MjsCQs7sggDEB9sAtJpjf9jL8skaE9ZdlBFEEmRJw
Zh245RByrzH390prcveVyX9Mq0nePmanPx5KbVSV+/NAc2GdBzJOfdNHG7nJWhAqibkroNSmG/3d
QMPt+C2gNIUjE3cmw71SdCNMja2mSByBW3cPJb7J+ZHkXW0SIIqADhof2RDr9Tp06+eJ6d1o6iGs
fINixW36bl1if7pVwiTTGwcOoeOFbo3V4yXYfR9Bjtc+vyTzurPv6LpFwcqH7v2XSCeFslc0OYBR
wSyggE6tljoKn/BUBAGDCpuDdOY6s9w4YUQHluIKllaby6s+8iHgSb/29XumBp8mHtgIXRliMc3f
TNctgT10SpkJBlXE6cZLMe/2YLgy5/iDXqmJUAOipGlgXXDzaTfyWY3d16Q+QP684r1ZAu2aMn8b
xv1zo9nnTAF38ZX8m5cM7umXziYERd8fIE2MNdCNnOBT/nsQ2aR4bL+lOxEma53MolomDwWwdzEy
1afDSmSGvw8pwqjIDGBJ+jSgBBkZhMzHi+nx3lqWDK0x3BIoqy6sPTCDIBZP23Xz56EYIaE/SAvM
WxyUBJhdSbHf4hAZEiK45Vue2mnsACSS0/BSBlihN5XdWrZTUzeaSF58iMdhvJOXuxC9gx74eTOv
xWKROeAuRGmh7uVlRuL4GPeu0sciUbIoyPt+KxB/9J+MCq2yz6HEHAH8AmsBgo0TZ0RUijIcn1js
ZnPBpxBhb7GPbRb8zxb6+byuYZoCVuOyuT+B4K7Ajl1PJrOoZQKIER+b2XoJsnKjPy53fuAMyrJ6
sXJwsiABgDK2Eh+5oNL2ioAalToYl2cJveYCK9NTGcJcwC4QW+0n7UjI1EY4YZ+cuON4K6gKhWmG
pVkDSCqK9MR3iubCGGFS4k7R4LhZsQDkG8jzyrVXRHepBTj5zKCVhHwiyuAGJsHhvpZ6GuOAc3AC
trqDBvv+GaRFjx4UGy7LdYFyJS2T8Y3RfTdwDZAqf4aMrzFfYS4ozajphPrbZAW6jxiDsEvf2vrT
4jsMHdNIGeSOeaVhmlpc9tiX9ZSq6vkTBQtoQDw9kE0bzduIvPJe4Ou61F31rkP5f4kbKdA6SeXr
1XvD1H4exf97apn/Dqh6u7Ag0w7fi0H7qgP+THEjvykJizIgMwXpjAwVQv2X8uvREoweqwwDEn8X
GiX0qwvDZuCWN+Me+t18W7jNX1dWKD2pw9yXjsNazJihL9ncobd9++A8uyf/Y78zrSQDUxMHUR7A
gYXe1JcCa0RuLVXtc7VVHbPkCHYJx9cp3e0mCOHBpezc5gGdW+HRcyequWQxb74oRB0N29mBL3if
8f0XDXEfCmrHnJPw3MU7LLKWzSKI0YQuYM0KYaEKc48Ye9oiJ6C4loy5OjTJ3wqAmgpl0CC40OLM
Lwv8UjB0CS1aveGZuLF2ob841muZmP7tN/3s5SJgDBAx2kp6G6da7AFVdcAYxNZYwA+vS8Qkp03q
FqfdNvkoSiQ2hSb8zTBMRyD+9djSWs05MHXBmqJgOjn3zznHTW/e+AHpq93R28VAjEsPLtJ8Eshi
0kJoafjXQvDJhB/fx9FHvtgtt+6BjLemkONa5nca9VXz1MAD59+8a3wPn10fxQYaxljcofigovx6
akccyDSa6r0+G/tGjUsa3yxbs6NFpLQpWL2RWweJlkAMmTxRarD9wDNPgP7thvDxkO9rh6VV0dEk
XewT0rvIiov/NQoItlqNYPmTc0jY4RxA5HraC+sv5AV19BE5OBxSnvdA9czJcZvhk9nhnj1X4UXj
UcY2TYR8WPvI2Yl+OF4bZiukj4qBJ1Yfit2nP7oBeKFdCSWzxf/uZ/E4KRyhIAVzZ37zyoVxOUEV
Amvum3xVoAuQBl+Q2Xpats4prXVQS15hLSe+dzo7vEEltHtZig/M8LAa7ic0MbzdfIH+uGmDcMNF
DNNBYeNvAD2ueZReEONZ5va1ehd7IeaJGFWCgQADGnCXi5ce0DYFBkQp+Swo1d7wwepaUKNl2zo+
8wxiRIC6Rz1DM/HQ2O6iRhbAwqEK8NpnLBe346gjU5W3i2N7lja807Yn6M/ZQfD4HRMeQuidqXTo
eTYV/WySuX8b2Mx7Jz1MtAjSQ4zWyFKEYqQRgU6ljzrKfVn7Kt8ALd/9gQb/NXOX51IqPVSxfUKH
Izdq5ZC1B/IwKaSG4VgtNpDQugE7DSAmslLE6I59e/DxdNI3ODO8oD/AAwPSjHlSZMgWfQaZUp0k
QAhvk0uScMtTX9Wj08Va7F9qFjNdF9xa+wySIzezjgy72hHfzUcJ2nRcIPn3Prx6tRzgOG2JeEdm
9NphY1HEUkO8CIWDsazxQCBYD2KdzuKDFe+IordWnJdCXUUA40Wo8Gss43rHbMh2feRRtKL+Atqz
xbcUAVHX+eqx3KNE2VDvEZFvI8XNvyC3D1caXu6P2uXPUH0k+L5QtLve0zwE6lyh++ublhe8bHFQ
MgH9y3aUDOwUUNlJSQ/pDaOyojJ03lh1d0unmliD74w9Qr+O9bfOWFZUfwODyzskejBGe2aGqF+x
M93lg4cVhlPmXIXmB5UmJ7bIfJPL0GUQDW4OeTP6ONTi+8sB4dgEzhdtPsEQA9OLhiKjhUZ0QfsJ
Twd3JWpNlYfDmbVv1axY+NtnSVdLu/UKNGZz6TEArCfTrhnvNFKrDUYLt4W8lMNhNsIR4FDEEB5K
D3Jm003GIEu8KInUcVGp8PzTS0H71Vtq5fW31XJktSzb5OV+k1JJHQEewsgatSG9t2vyoDlToit2
7V99m6XA5PPBm432bl+63aZ9ucJ14QnegK+BB+QR8lJj9F4kD2o+2QhMYTWmFNS790mALJ6riDRD
Mj+lhmKfKTkEQ8t/vG4lqYj+sEec63dhdnfmgPIv4h9Tw6H10IeeUjdgJW3K5GJjyDneHdjHRXmX
R8ce6OFx4xYDrDNeVMWvptkNnnPok4rCAQ/8N2T1s71fx1ylmWae6yyhBQD3cE9EpYUiwi68SXaZ
4Wo2ToN1khqZEMc9gmnxsKlpqz0MAd8T9MKUaQVSsjszSVcTXvqQWX5wRjf3bwh8bJ44zP8TfVVm
y5rURsSfeMRps6Mw2OPuGadzVy1wSrXmST/+0cHYwXTEx1OugdWRjumJ3VkszbQfujcuJHXxe8sW
dWU/8kcqKQMMfYsTbFmYaar1oFWaYoXDsfh7pEn4BVJWIa+2CeOaEEwC5iSny9qF/8pZuL3QHS5Q
YJXoTeapTHYvmdI+ARPxtPPGQ5EmYaewjLiqq9ObNG7lqfNn12StMo46R7v4GswfytUSPVrf0ONo
myLtTiaHY13oMyY8v9CGO3IYPSul15qX9rJNFzGIlc0+0U8AjraFKCpJdCtE32IcEA9Xc7hjuVSf
3S9+vnfK7YPFkWV6s+IoWtRLCVEPqr3KhL6m1kAa6XpOM7JyYgTBDGvg+29t/YUlBm33usnyR1me
p/61vgN+H/sloPHuQuNhY/6vbPu1qWwz/k/LhmUajI6Be++Fd0aNu1aNmX+NMiiyau9uq7KfLkfr
BiB7YLDc84KX52I4dwupJTNUjXrbpV2blfcGrv9d3mxA0sbJtZl4jIS9k4YPTiv7gNb2WwL8nW8k
TZ/guLyMREyuEafpyqqBQ+Txkra7uxTEF1m13f3hbUrp2QjCcxypi1K9YhY6SiyjsVsKfqluVuAA
hKwSeBqvo80HtfBzuxphFhzuUy+DA+0/vAHVwcmSzhoyiL8BPFbP1HNorfBKvKm8M2qE0fCmjgFo
vFRo8Sd/LPE/EYnwNNXHqUnA++eaSNp3Gsqz2Y5yGjDO6YcwDCfjA+6VTUkcmmcOBBCmew77jndt
EPWrJbG/tvcr6B4eiHtBblu98aKGZEVJCnyoq0ejmgCkNa2JJf9mgNH4eDetBYk2aTfKRZZGRtXt
z1Kj5JNCKwJFaZmsq0lgHCqLlRUvkeYirr1ZhBpdHYXy6Clk59AJjGhTjf/MZqBOEC/z4f/0xk5E
D8ZCQSARHX4+kdXW17b4PBdE1xwstfVJHj05Kk5FAKfC5KfbUxxnRuM7vwrp9XvlWW7ZAhXCUrJX
SRI+oqKAxMo6M9w1fkeo+ZukDAjANSiVhnV1C//hQP9CuH7BsrqhpW9nDDHVz5Uz2ZpWisZgVguS
w2DWRn2RbFzMRkZlVCcHdcKQWk9W1ikADFW2weB1/DxvS+khmcp27APQczAWjEn1Kd+ebhIny0GW
jtJivk5dctb6SRIh1j8rz6pjoKhV9hwhf69z8YIxPGTEXVJk2/Zhcep100pFNwojWbD3sGBkM4QX
leG7DnNfWXch0Eqko9x1jai2khcvKTuxR01oxvSlT2FqkdxXKkM1GgBySyzVwTNngut5cdX5GB+Q
dZRYD0jUPyUofvjqg4Z4tQijvJEyqgzThezQdCyl5dXFb2b2b0rR7H2pcKbj50mZpyOqQivi4Jqr
Y0UFV0RO0gTOKQA9leQTSIpjpTW5LK1QljqMhx7wqprV9m6OmgVxJGE+dr6Wz8HH8OH2Y+z0FJz7
OP0B3b6gbDeCAdsnkPciVXIlajsVd0lCT+Zugedkute2Zzazq34lfB3A+q8IFWB84Zub4TYT/8bW
N+vjWF3G303GN+MWbV/3ymwQPIp7/Q84/CqZoOKKXodA/GvPaDOKJkcd1hyw+kcusQr6S+aD78ot
S1/MmPAaZCx5qszmrFZ/fTkUEwqhtzQyw+fXVxih7ouT9FbouZarFlx1sSvmC4En/3QTt9PIxUJD
PpEsmQa2Ro8cFrwtxa5zJbPsdCJSNzu2q1o40fFamFyJNQNXFUw6iPZe3c1CtNV+xLka+3H7BxGR
+8hrRp6C5w7rlhCiVE34bvzC+ry6Bb50MMN5832RHZKDAghMozp8/ZeMBHG/KhYYStxKM0rtbLPf
s6c6AMKBbZ7UoWbNAvk3ym3UHboY2ixtOSMql22DYsbvIRtHHJ57ezUaPScFBnHrE2kR5hqoqm4r
j/ODxMoI+cJQMGBVedtXrdA+Ya0SwAc54MbBs/XvLXOTeUXZs8XEHNZTvMJI36YjK5eyG5BgPdq5
OH5npl0YWSVvUgLPD0kxgvXS6d9ysPfC08vAVWJqKp+CHht7nmsO2066gwZeG64XDE7gv2NtuJnP
XlRimb2RFaqKVc84oFTQYaYOZ3kl7jwQtfRccVKx3FsB3tAqiNFEfcmv8fWfsmFHJUC/3rzJWeD1
wD8BXzFm/F6svk/ydPRjoBLwvNwzOFxYGWYz/kf04Lvxsp8aem94QuQKzcUMqCYT89CKvrVouROX
MJKihyw10CGqmYGmmP0Wk+HWnqB2SflpWEEOBcvpgT6KXu8nZVx8Vu4I11NjMLEfR+Wf+bPe+teP
70dgTwE3rAvp8bVaI1oJjn6G/G/E9fg4io62/+IIFWmwQaPuKvc7lvNTR71zCuTPCyziSUjII4lS
ipHhQkvEQ1Yyrh8Ts0Wpv0nM2/6QqxF9WmvfR8i2BubUBpevx7XNpALDQypVkGsqCZF+nejt2rha
mE+VwrhLD2vZv3WixBMX4IIqjBFUAeJ8yQre2GnsA1AEMTKPUNiITlZNKw4RlQMEn1VCggxlVHuG
XV42BkALGBz5vZZQVol5ipOPHAmHr0LwfTWKaZ/oOjYTzF4rYUo9MatEyQtt6LsY4S06loEhXuos
FI9qvrdx2jXFDEzWFOMZyVAqgoIM4TkZREYjxUu6hPIPtyPMT8tLuIuGGweSj3eVAiip4Y7HUpfF
/h203m6edkeuIuGWnYiuntkbuI3/0VdKwnIgYvlcCxYv1gl+m6uPrGTZuhus7qpy9CeaXeY6/1oh
Bx2z30eBV5UYsY/4YIzEldA7YzH3LVJG+L8TViuAL976BA13fJRFcEfbp/UjGNFs5aAnk9Q01mLe
OVrEwbwbiT3T3DfItruo5abdsuY+r0thsV4vpZHfseKAj2pOoxZLR5LA8NgXPIEwlCtzqgMEkVWr
yskfMDT/Qg0jYceM2MICSWWbuFkJ82ddJGiUlNE84CcXtfEMwkacEs/ERwmdYvpfNG5mAOchlRNF
nqDmtGfdmR02xTLMFP6j55E1oCscsv3ieQd2sGc9OBcGtq+2hxbHJ/9LKK9qc72wHnPaEtPp6b0s
IVr6IakRwSavvDYYv7BmgVosEwuwk/WgdIdu1Rz7c6hWXkFPFChdH6QNR4INBdAczCPZGqEVmybD
ejHb0gkZmxXFHCvIFgogwTUFKfOkHfGWoA/tS6psR300qD5HLHVXmF2SBYLgl+AkpsnWBkE6zaDq
0+6SBmGlIrdm/VVQO+FtBNNDTf5ev5GTFxzMfUqUdVe5EWEmOPGwXdbOyt+IUWH4Tpt9zuLiEnIQ
5WcgEeoG+ee3NhK52G7OzQrr1BUtusobIDylb8866wN4XpnCTlAtOr+eG3KZzlLZJrAB9J+HdOKK
bv6sq7f0rvHyNMfdMm5HvNtGtaGN9TkKfWoSukt0iJ9OWqWPodqy6Gr2yeH07xPETmd/wMlNBSgv
MTk3p7V6a6fUqmUZ1c+guJBeAehtdkMfla8BOGxeS0EToHgnksoDx0s/a+O8aIlPrtujZvs6LABn
SEeZYeBO3SQkOzHbObDc/Z7+47mSlG0IQiiEwng0mk5o3MfLbiBhxS1igfHJwOcu0r2QwtdunFNs
x5pTuoiSADUQkQgU0NceRS2gWCDbFSwAgUkYF3XdseySXxH4DNSEhlrHjY2+AEtktQMUPD8FjcJ/
ERTt64++lEOItyFsj8DTQGci8Jw5mhH+F+JmcsXIUhjdmmca0fbUSehhmwnfocBpJrbVLssBy8i4
1jjuy1pOUYDFAyqy68HrxoWeu/sGDLlFPL3VQ17CyonTmzEyl+FSy+eHEcmYQiAWuRaaloUaiLlA
fsxNt8qeqoFwihVzU9Nuphej1QJYjCrFi8aVWSC+qbvOjFTdYe1O6A1vmbH7SqrluzepsPU8lrin
JApW9ay8lvb4Sxi92EFNmzVYZQ8j6G9pYTtlq4+8dHGjGxQE8M1VeZEKxlyn3+8ekm4KISXFYmeR
5jZ7IzYbPOleVbBz2jatYFBORnA/jVP77yBpsK3ylhzrzL5HnSjTi4hT2JYh7oL8vP/jsY4AnRkg
K/cEfbrEtBQy3VB4tc4lHsKdJPEfwuF3oWr+KOXC87vKaxRm/lLNeSZbnZiy+vtE+oU24wcyr5xF
EgBG3lACDU9aSj6YwubRZ4GLWDtkf68JEbXk+F76Fixzh/7RE78TCoOIBaz4X+LLjXr7a+EFlfqW
xVjMcFnUbBbaghq/fOh0Ju0fXcVzwrGHw3y+w3srEe6dKrxm/fFkINCANXRsM+Es6unO87FVniuo
RTA+4YBoFi3Goo/h67uOV8Mdi7oe6NeUx9xLNbF9nf0GDfrnE87qiSyzdSA61sOe7ZuAd+cLVpKj
3TRifB1PogSqONY5GjIcqQ2XlEzD8cNgEA5z33HT1ujaDjGXPv5wqZFTLVfuHp5b3Myv1ZT9Rd7m
IK5qzTNpt6fyTWu3kZKJN2XiTsmoaM4627v9384tSkod7nuShPq62A2Sq+DIGRcnC4ylzmHhgWJM
i75rYLnq9wlPvrfGN1JTITdf/+V74edxWlh0AqQ3YqdCv0uknc9Yo/9XbF+kfQpzBqq2ZJdtuwl4
FSesuf5MRRHoXlsxQR5ouydxKgjLJM6FFaxkTA0qpLDh3F+FEEavebRFyjd0W5Q9nR21qIxsfOZX
N1ez6miW1w3MIcZx8Tgxz/skwdz2M5nmfkXCtZD6fG/8/9+DANmf5gczxBbIdQxB2nAQqrCNL9Z6
uxQkZI05UOPoyqgoB5MdEiHoJiTrvnvQo8xKgWAd4LRI+Gw1ylqSb9ShMKYIDZ/9pgKvu3qzddzq
Tv3d1ZBKiBC61B/h+lLrYiWU29R5oWWHWXhyUjxWIipMnMQgLfSdN/bgf+70K/AChpwRM9eyTdkZ
c3iKMk7ygkM+JICLGtSA8dq2R0N6VKQb5Tjkeq8auyfSXaLs+0rRK2Mjl4kwZ9TqNqa80u9PWfnO
BSkk5c+I4ZBOY6mqQ38coEN2X3KfLgbrNUdODCopTdQxPZee++QlEgeqT0XLCBlo7jUNOHGBRkr/
Dcc6saJHSdaIIg0gSzwAM7qSngNUaYRZNfDEpChZqflPoCDoXYIWEBJvQFfkpKkOvhbKPE6AvhpD
3A7w0XmQ0/1QogiWDvwUp7s6+QOE4aQlJtsWfKBaQ1nv6SEB93cjiUPOpZlz1LWaS2J7wA1bPvLT
1BUNi+iINVTav4F3mq+jHegzRYWYRzvPB5xV0qENVj/Q1QFpzfklfF31rektgJ/H6bFPyT8L+10r
3/Ho+jA4eBy72uy6CSyin8cmn1/q28n0ViuCBjNNdztSyGFeGKTF9pd17pbCOBt0uHyUhJyy/jyO
TKApci56ef0N/eTAt7XZvW+ar4UVOfuIoxNhibVfenvijf4r45HiIH9fH8MectC8Eo62byrszbEE
NshxPvyf0anoplzqaKNnOvd23nmW/oKRw9OI4nOdk0V4wB81lY8pInxAU1DxdlY46Usn/KV/oF21
KzIA0e5OaOz9tFApfva4cbL27CYk1eJiSug3f/oA27RsyHCpe6OXPtqTrpzBlQ4HxJpbPF7zzsnU
wL+DiNoTEzWSmDYAQo2zxmJ+WhdZ4zL7jwNkxI5YEcmnbYiQOMwGXO6h4G6Dxc6hV9AN3hbTRDOy
QPIAXq6dQmc5V3quTZFvn/1/cOt1f6mpDWm+ELqhu/c0H/UIpFY3JF1on9IYdxUnNLH0oW8ZznrN
m2S9WJ3m3YTGEsXihKWQkNDc2jjrH+2z8KbcboKwcIIsjxC8dhMSuiXJj9p/UEQa/a3keXqOnOhy
OjTWlbRaJKn/1VOEfAcmnmKD8AuuRN/x02ZlNc80J375YqYIq7UfyvpIpU1D9Sy4qNsU1vM9XyIu
B7VcOrd/3WB0uATVFHBeJCrquWx+1vuTNm373HDmvoF/rd+YJifS1VYbjohnnz23JmgLZEDN8JIL
ZWoc7krYLP6aF/oKzYQQyoJy+WAI+Ey57mSfKDjj26WUHcNiKjBqiJAgt/KabHe1KM3phjkOWvdB
ignCC6PeoeCjOSyUxv25vjuMY5A/eZEZi1oEZBN4Yoc+Y2eQdC29RoOcxukiNkEFkeDB/sjXUf6Y
deJopidnH2TyhdUy/xHexQ/uAJJ5JrKry7yDIIqLYlyHIqNYeYhBIzxbWT7zS4LM12Pmt6J2bsuO
bSFFw3GnqdteLk6iq538Xyqng15L3hwdxS2XcxTu2GuecXns8AXaugdTB87wJzlPZeQbFERVT0I5
7PpIHuiLhwBbBMTiZ75efTtJiB+OF3ROdjsS8PdP+ReW+loMh7GVw47WR++1jNWSJsdhcRGfLD5m
/voPkM6CU6Uy6+qLfrWyVjo50EptxV38X1ab77OFBvRLEzBqU6ODw/qr4qJxFauwetnM3qsgPXW9
5pJMg/Z6w4Sc/WGjtMnAmGxuCgYqys+M9dhYFyRS32pe+rqE5m2t6GE4gIWp0tiSPFN5CrGycqCU
io+nNC+wkwJ2fib8MFZ0B0yYHW+NqBsEgzNhCb5qY/ej7EDqX4nL61hJE3dTP34hWHPtwTiORVfa
FCUmy1fEWeXfFCfZ9YKi6YoFOgnzkgEwtA8rmtpBDsv3rTw326DLEpzwrkx+xJ196o3c6bF4+fKN
CaQcpqRkV5/AX+8D2bHmanjdmRwLqCJ1JpVC3HiKxu+43aWC/aLgIvIN0okbZXBg6Pm/Iukd20Wq
9dovR+aw3KPGs+Awau5pNkeAArpCzAWjmMg3P+PjI+H8DiazrcR38toy2MaMC3hW6/zE9WMbbYNH
67CGwnnkbKNtcxXJO2xMA2T3vHzMdnKJTZVJFaRQLD3uDK7Y/fcef8jHWIQgLTZFGQKrmLrtQNat
sqFXnpE35z1p1QIET8aU9NyG/yN3tVovXV5WKMHPnsDEXncsBd8BA+QDdGVDlO67Gd0p9gpyHHgE
ezIw34nsSXvzztEwUb2dWpCksXzgGA7qA5O12N0flIQLY1HU4JIMekajF3gTq6n+qT9XpfcUrRxS
Q0SYHY9ZqriA7E4kg3TLSkbhNGnOouOwAwR5zMEIWvp52phpqGHaKv2Re+uZFRJcVO9PiQs5rfNg
S2kR7BkzTt8jEbTJi6CkTYpYM/rAgoZO0mZb+v+gOr01GW95/TPcIQ3ZvhuBawkK4WgHQR0GMBYw
lN6Bxf/ynKAsN+lzwpx3R7TyDDETWVQI7cXGW1tfjCMjvNJDdq9Q7rdan4av678d7KYLWM84fOAy
zkg0N2vDuJT0kdTNWzbD0lJpz03e3xCE3a6/8rIuKkPCFZaVuXZRqZYsgJ3+J0abD0pTMjgwx/JQ
mFD/X7S0fZ8y7dYKbqS6nYdSTcr1UqKDa432SSbwDCrOTdXSmAGhoi2Bd/iCkBPmQb7DQ3WVtUdg
jgAie4xL+exkEWodA8PAvlsz+49fKxS2ttRKc8hNc17RKbK8VnjQ4IVBbwOdH7upvmscl8ot+gpS
7ZpQOgN80q2ZG53biAm528AVCEAMDMK5mnQH5J4eBCniAj8gOy+tvCmIy9r0wIH62QEOonnqezqi
QpzQ73xWlFacGx34kTcvGGyFzK0PdF3ea6CybA6oodu86KYhCfj63IWrRFykvUm1XVDe38/2rzLp
eChBSCve8YwJP0VfgNrUrwOA3fKxi8dKomFxKtJhCa3rTVdbCBnogz+ACx+WR3eG6nbpHuADAgYW
hExQ3VuLEuNMuxhsjj0noUtxIqO5ygrQHeDc5Qzc+6S8D5hpq+Q9M6OKGM/y5BxaZpRk0T1MX/at
peiZRNZwSt3Ge4yt0TGNXT4HkZuHSXZBb4zs74MzsLAYXAIXSOpBMR5Lt8jtAw6abMHz4cf9WBVM
qapy6yH/n7S1vm22CxGGneWCfcbQH3fR0qf9LSw1ax2zC8shlbJpaFAFQulqVi+nZiPj9ZXB4w4b
MRECzZImQWVUaRogqNEP5lAnDgpgm8efHV4xiQwnzMxgoZw3Ncw3Amd4R/K261lELktIV9ut+QRp
xUfT4aH/JZ9Kkp2U38yn+Q+gm0C/J72lNXCN1tOG8V4XVjHSbXITkfO2bvWz6e+UcUJWSatQQBDO
mNrpc8feQfBnOIl1FZ9RkG7d5+Zku5mef0LOroth6qDwwgS5cEaygjxB3iCZt5iswz7w0EkZgYYZ
/0GB4iBgyMzMr3F4eWpJBTFcT2Xj0AqmoItQLw/HSvD6bDirY1N8/Y1+aos/huaQQ3AHitIufayV
VEgtBu1oKxWYKW4GPvqlI+sV7QAtu3WZKC9zMDA6eNYdE0XLgkRSVjn564CoKbqp9RCb/RzaDC5W
2YiS2MpFjBdvBWc7r8/SLzy1/R8UCox1KngVBFPVJm9Wof8F5WOlL04r6SJhMUeOYuWnjqnfLvYJ
5XXfNIaeHbu3DzImxxyCJamsjuNe/5pjqQxzbS0re1/cCzVH6+Kn+3ch8qeesEGaGgTCi+TXWb1d
KBBIDSEFQFbiqqGaUe+zVC4PKbUXyjbvlP+sGhZ7GYMsoX5D812wqgQL0M+nivnl2FrfJEgwzNcW
D94bXe8mUWldJcVGwykBycq/46uRryuXzRjpDtWqfyBz1UxMV4fkNh6oRzSaJMYwdqwrjPcBTY1J
mr5tEwQnlkdjocvBNLgaObG5YHJZbBaLzcQ47ZctKdir8jmyoZZPLs76cRIwHlN80FDZ2pM/Fqei
EOMtaiK0quvyLlr0r8FQTiNnPJ7hmM380HdKO8daULdahhG36hXT3qCXT1zORns/3KTH3BP+W5gM
dTwybKOhfyPW1hqoSoRIVA+PhlAfPiRSP604VaelLBxZFTqrd/wKdw5NK302pS9X3+2ZsOUUbvo9
eT7SYVFhZ8PL4XWVzGq0+NDDJEAGOkl2OTrhsT5CZ8TGQxrs9H5Y3w8oSgparMsgCyWqDjG7ohua
y0PPLHEwMlLmfnp3d4+TsBZj11pG/GbDy6SzeXWlyOgiOgPlTJY2JyaE9w4i2GX7rkUQNEJ7Fvj6
rLvH58UZn34eIGeGpZR8nTZCEWl6Ik1rE7hs8VGDZGSCJnO4BHZx00bpNVBwYx8sG6Nx9T6Y63WX
HGPzeA+tciqKkU1DGCEy9KdyS8O4Q4BPq0yGJH0odKdInJ2oY4wplRue/5nTN/D5HVo2q/0Cx7Vs
xl0H+ERMxbxgwTjNUOEGk7uu6oewMespa3t1huDsJ1iUwLorSXlKpfSz/RRebQB3mb7JbwPfj41g
wIVc7NR1JobJOj9f9IG3Frjp7i3NwQ6a5s8lmtxo/Rc1uxsYcvvA3Ot3GSUiq9T05JicK4LRqv76
plFDm15lXGCyIllx8Lt368DGoWQf4U+CofZzc6p7h9ICEI0AhB8KGI+fpxOdMZxHxsqCOIpjgEN+
wZsAzVCsDSYgiD5/p3dKcyQC+DSqPri7tgN5XUiZX2H25Yroj0OaIw9bd4Bo81+30sOsA9ivXihE
weJrU0zQVag460HoPsToJLK7Uh+NBwXBkQ5Tl9nM0n3W8qi6KQDtNKVFgnSE3VEZjyTsascOy7de
+xfc3sVfoguZnhinuxT09s4XxiagvqbKn05CTQffvjtsfpE2hkoh8YkxaxtVlYm5IzAWz6ITLjhm
GeofxKhiIIpgoSg5y57OIjz03mOq3Z0s1VvUySK9bNjDWmbeU41uys4J3m/qgTKoTd5nnLWhyPsN
gqfdmcu8eIA5XzTMiBZJXaV610INJJnFbeFJWO8vT+gvm8CfvgcS0Oj7tRxw1S6W1jUYlGbSGaiS
CkI3I281D+wlogA1RXhlSPTZQVm2lcgUxTUQ2qHKiS6zF+xI+PgsxCCRIiX5GIQ88bep/zJewkmy
NGvnFJB7o3JHJONQv5P3NOtfpC9U4tYiBATr5b0bSf46A4LMf4kYVRIBsF/7UVDMYBy5x8dEtRrG
bntdxKjO7fzYi2Aqn7xQTIkKijylsoRa++tEXvp+iL2qUb4+oOAV834sEIpjFBLVJ3ZhRL5E9YPG
yumke12UZRgz4RLeOeX7N51J/91u3cCF2DHX38bhr0C23fMfmripEHf4dCqpnaXk0pvLRAOHy+Tz
tz6FTCBJdFa/LELyMJw3zZ7C0Uwq4iaURRh7GeAOTBcx2T32kIj5r7owHsovN8b9HkCRxet74r5I
lb0IsyVUDE3ojx5r17+aJfO5kSCsonMOY/gYzN5dzwqzE3ThlqJPio62c9HZz6ryIHqcKpPzcgDr
rSyTK6QJn+6gyilASzXiMa3i/tH617jrPiOF4Cb4LcnfIWqIEuHsr066xaftgED1A+P2bec221OS
1fq2j6ClpJJB6el6JAJffHLmlkH2U+J/yKr3sHG5Tmc6jJ35+aI2d7eJWyrgUSy+PmfcCD1mA5/B
Z7+lGIIWy9JTgTiUpL0v/y5hqdtCbkWuFCZ7TdoDWAOJ/P5r3umNZMfxLYYi/u1J/EZ9U8v6fXsZ
eqnYouEF1iUnvhbRPZbDE0UrN6FSevCmeSjPAp90N6U9euQT2M/BUq/OlvWVrzGokBWsKz4++PJl
cWS7z5KiuF68lIAeiXSJjTzer1tC5ROoUVQhvxMiq4TKkBVMBK5fsjF8GXOmpjxK0RI2bf+ttmbG
sDSILAiBKjFErro92SWjh7yOOzPDO/SnrYa7yMmmIG1XYE5NPuZCxg8/1nKCxKugSihdC2zV7dvd
wtlsyq91esFNOYxf1kjBMnP0yE0ZJA2Rrdlx2W/MdLQIx2m2pVwaFPQjFGpnziiKqMP8oHpHpd5l
oMZhFumQ4cyy9glGrB0bDbBA/qRAVcQYx64Vp4s47zoBSAcEga2dcl0uvqRkVbgwn1a1eikRIWoV
tvtUUt4ZSHKW9ZPCuwNrDjOHI616qmCq7rXUqLsJCng4sSHweqVn9ykNCNf6+cgAuZsFYzmg0a1x
yatMJXUL7TeBlkFtSkf/aQS9S2XB5sNEfIcrwrQvM1xruyXsEL4NPu++40XnkbaBYAHBLLePJJcp
OotzSuMVItB8kfTORN4kgNc9rDKCaZp3ynvGAzPBmWyiJbGDh309XKlJeE0IdFpN8/j1I3Vnxh94
CwQltHDdMbDjF0B3Lf0pNKHjd2U1fAUVNVs8SvzLCCz1t4eewliFZk+cIhGp0Kf8qlo/7m3isHbr
WBMZVRmnI/OGOmtHllhIIU01TKzWRVxnu762K2RzPVxoi6tA7BapX0Farc8BIImvGcy8A5OQ6bB2
dRT3k4Hej5TWVYyYk/T4s0Y0f8eAdW0+JJPL3Dv2hRYhS2ARUMJfwIwmXmX4UzpjyAnchxS/uYne
d+eyaQHdn3YoG7kNFzeY1+pzZMyYz4Ew/uscCsR8KgQUSDeCHhTJYt17QWJp+Pz1RCppJJDMdM9G
Ue5p1Jl6om75EJKz9E5sTsHnDwGFWfW6IdZw9aNRcqYQFjieUgpgPmmK7vfN/9aucqtQCE4Xt2C1
P86GisCqDNAinneIPqQwLNE1cW2qCkT4p4cAFRSsF1FTw480gnTm2ZBgVRNsyQIaOJyomfl6pUyk
cY7Nw+z54EVyO01w9c3wn/dSeImOXCAZgf6MVjU6tI+htMO/GNqPD6jQJvDgpZ6FAL7NQMOYqxK5
1N4hAiPy0TiA9wf6Bixz0O+Kyyc7aGKx5FcIrYm/Vp7Cd/oeESeEWr2W11yaF5qyQSV7ebmy5dXv
lGCkjMyXAAJsGnnZE2pfpx6CKuRdOQ80pfQ02WGfyiYYQnbiHdIQc3EhRIuKsoQfT1qavarQY01T
63f+Wfbs2Rh11Muozk/byYEtQ2Z+kWNXrTGejcwovVarjLV4Xxmk7abPtpykbm7HY5fahAM9X+rx
az9xh91m7pcaCpQriusJQ7YOQEFa5kjTtmyiUr4AW5GzJ6729lbSW5t3MNqe+FDKHCoCR7cmrLT5
dD4Xr4UIrcHXw5ybWjrLMs+khqDfH7Siyqs+eq2Uz64nqXjuFkxoK3smkLvcnsvxJCiz3JtDofVR
bi62ug5oSYDq+Cqope8BbmsMXZ34bAIknnFNa384fra1nDFoYGsQmd1XZmiyS7vkToH/nAcj4ocO
0YMTdwaM6vPU5jKVkfMs2HkBl8QsTNedcBQ3nAd3j3rV2DCrlnyubwi0g37rxQrj3F0IG1pkuu08
x3LNspP6aWTqP3a7Sw/fRFKtbytJfU8Cgngue5mvT8mEFjOyl98iN5dS6NzAHA+c/AeDLGB75iZ6
MLPWqaD/Hyy1kaFQSodmpUW6DgHyNJXf7OJB18BVH4O2MBi5ZBERAD3l0Iyi8duJjc/7nEdJJP1D
M3dmIlUkwdPQo0zQAV52DgV8Pr51lwqAvfSRHukEoU3MVQ2UK54m3u/Rg+gtitBoHAKb45gjGXAX
9R2nVBuKeriR7Hgx0HS/YXm5udZXV6J9mnlVEsTVG93Ujen3FmtZYwvxbwjGKuezhgWE1NdwyN8o
LdoFF73jC9f3Tzdw8DAgyQrf/lXB1+bbfZPVZm0XOb82i4zdmfWxpOJvZAo/g00GfR6pLIBd/zG2
FDILMW00PxZMKQOU2XHH/rx7f9oY9he9mTXzk3YXF9N+U10St6MSbX7uyRGb3NB7maSjB/ghIhn3
lMm28Lv2RzOXysulLojyIK4+gPbLT20tdQtqvTgrdazWbUSsDEa1MrW4gqCoEnHyiVg8rFsjZAup
9aOtz5dMCpIbmnKio65KQIFyFnF3DXMgysx2Of3eMH3hpgwHLxa8yt/rvgZaeBJIe0j2Qx/ea8xR
1/i5jLgz0S0GaBgBdExs6bOpjnYl5w8450q04h9UGUXkb5LqcnYTVwYYKaaUZglVPx5ljSDoxGPB
0MjmP2dGKVa7kWpSiYS7TF/FeqAdBPFxMfCv3mzUzuT5+oXGZS3FjFo4eYAYCm2J+XKhFUGJ1RsU
ma6ekmZsxi5j7qRiC62Td5EW9JzNXVscWVKxZ0JN2y/nBgOgMzgzZ2UcbjwCYs6sdQsvm5RROZCA
SHUUrFenH0kYqBR7NC2Cz9XGJwqP1o8Dr1uKh98n3vEISpHwTu1XiDI1fMos/WbEXGjppxbEfuoB
raMuRruGn/CYbqcNhVbfy41v4ya4/Feg1etz1OiuNVs51/qt+4pmN8Y2a+KWG8JII5BwQENlL0jD
P68+nlTxbixsq93i2uCc/pRZdlGk7U0FVj75Yu8kKxG+8PlSPOHPpaVPaRcvT+WivtFf0KOxMbMA
v/U6AEpT3u+Abph6/Vg/mlINpxox4AeqPt59iqeiR9xpKDr1V2VB3qzjZoBKqm6+fh4aJArDwwnm
qYgLQbFOITDYnDcLOElJfsHIsKB3nEfvNruH+Kl97hJRwvgLds770whoJ4nVBRBoLJd+OWXKqAFc
sKVJcn4svs/OvJIjowBsj6dGSI0PuSKexPNzw2I7ssFox0z5Onoo27XlQqSApZZ72FpK50NaU96n
bb2UtQ+tvLHFgQDxmSyZvoXJ12WBYVFP4x1TR4ws7xjT8B2WldGuM6f6ISNxyKof70UOhndQNMCf
Our7swMw/Of1iK4gUD1mw9pPO2jaqre7GPJ3ct47sqqIBvN9ObDeOEXG/GHE7o4fozzsfPA+4Cov
/vK3LxigWTYNJLkvkbc69UzJAnV/do5SIeG544MU2Rlkd0J2vGYlVaQrCj/65H+aAhUW3U8VdEFQ
XIJXquPgJ5sJB+9UMNHO02r4XoJaxBD/O8a/y0RfikOf8dY6rrWYuN+H8fB/p7xLI+jup06yRpX4
32EQoG0qgRfa6JELEvSkYZLy
`protect end_protected
