`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
USWneqzJjEvvLVqdGUAaUajBJ2ImPLxg2/KLoEbPrk9eOwxHC2j9fTm9MA1RoJeG55pMYJ8+/D0O
7mLSBorfcg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F93gq8kzXTqGNouO5MnGLf8fO9j4iAZhWqIIgA0lnNb1UV/ene1hl7LfC+Ok65b5rNiCmCcrdko6
LASetg8CXTmlAEuthHv6DHwaI5CB2iGh4hgCW2dOtBuBKxaPnQuvKQMVJkpC+0yai1hPLkOwenfi
wQUQJkXdP8iH9tFN6Lg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08Zhzbs8Y5TSF1h3BiCDLmb0/WsGqS6qd8k96zr2RmmF1SkQe98zXvR/e6uUmifbJahpoo8BMNr
EsITo4M3/Xj3QpMHst+toF5NkVX2m61XEiPCQ0ZsWBDH7AsC+rBahkHGy16Iy3oVhBzAzo08//1j
zvld+n8KbbbCuHaThGVUo04ep4xfrvBIMoxDx9zWsug5OBEYoIUkcT8KSfRLVYMRtOVhWmKmjBWa
Re/zK6PhdRq/n1F9Tb6sB3Van0Ch1LqzntGVDPd6550ueapI5jaVjphuIjOySrkR/HdPzj2x4AGC
okBn1wQecGn3GWUKfQita5IikS4ZGtzBbuApBQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bhHPz918RFkXPT8bC5qOlslNfijRn3VAbXxJSpXPyYTz1oad6pxgJaO0OXuHU4tXB/PjGRzPWXOQ
ve4b8KJ6wnVE5rPfWn4z4EUL7alsh5HA9xBrL8lt+mljxTJ57UNo8Z6ajutyDQ7Tnu40BZPYcSCM
FQUj+3RlPVDkTLCH9+4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S6Tu1gelABFw6/flIL+WgFwGGJTENOQWgFks6OSNuZLemu4LJisJ4EgYWDLKHi4egK5J/RnYZmie
ZAXXCKgBWvsCA3v+ZeUWNuk75ITRReW/+NmslbIe861nkzL6CQhclPZbOuJDlp0USUBEiGGxVvmb
BmFjlUQG76mCVd4GiUxmE9ilmyp8zPr0TPo63Dqt/YIaEvCTfqvhryX14ycHobcS+qXweQ52Idzo
7wqpL3Gw2q9IeqGOFn+8TPYMSfWat67ia2zZYUorkmRKkNqwCdaPcMzqJpC93wxOXhGdaSP/su82
R7qA18LwZYZGBjzY5p1neLlT0AuD+6zW4DDRzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15376)
`protect data_block
u2PLW8zWWSqdWY+M07TSGLSxAOswiTeLyMI0W3sOTRysMYXFSFrYMLRexKC5SVS+j02Beox32aRX
EsZuyhQeNQwdvMwx557E9BmtlyyJLTQXNqKh1/wjv5MDOp0Bfb9Gzsl8br/xZHHmQtj8Pa1a+Hsa
kNVptll49SfiW43oWoxcwhPuAIFlu/xiQazmkfQsN612jSl8xXzZAvW6PYuO6qSQQBKvOz3pTNNp
bm3f0VU/dyEENaE7BmUY8Tz5D0SzMR1xA2WGm9n02e5ERNNmdDFVqFj7euk/AgqernRM4fJE+ue5
i3QdUwc6orie551ZEAE/VjrOCs8P51mgvJQlvdHh2UnK9dZyHMh/Ztm6CqW5yrRYxGDGoByHFrdG
6fCpmaaGUg7TQIFadnQuRA1BFK+/dauNPH1S8EL6mPaB47dG+cmHUcqYXK+7HEGwed3c0hNytgGS
XdLilVGOrI81KgDtiG6CwxYdYqvDulEErq0PT+mfw3DsZ3asQ/UsYhgodb4SpBUy9u0Epq41fN1B
lhBUvG2kQ+QfcpOJRElz64gwqYyE1gI0CeJcRk5yqruuTOLIa7uFpRuGLzUqIi040eymKyo09K2a
j5IO65TIyMwiTFdLSxVimUYXph48KDXlQ0mHguZsonOe+jCHV/cTpQxikjfib8U7AsZwTfcLi7iY
5iDIzYWdYkbVqrJ0/Et6owl9RBohuU8k1oCn9f1DMh81t8bxxVxezzhwQPoHZQDrGPPTUW7pzCgC
Z+ntO1W3g9J09qzCaRawBuS2a4zxBNrdSP73rNx3DZuQK+Sm7fqPL/jLxukgpDbhjE86AHk/wHZu
1GKbacT9xNHjUB7sjICturYbo5z/kJ8DOj3qEn7uFIhgiz9+aOkWz5YxbjTL11YYt+l0nAXPvi+u
1Ft6lXPmPuhbtOcl+/9hj6aYKZXYO2nSp1dex2cyy/wM04NeEyVFhbRjnkLdmfqqgKC/Pk8Lz5pe
6tl+LUK5HLIpcXcSAKsz1tsOd5/snUQzunoHzDYmh2c6nX4+vF96+ZXouwGlGivqjdqn3z4Zkr5v
2u8RRBUiB2K2iS+s8ztSETeVSh31BjSoEPchQdS1E2y0D4E9NOwWm8e9SPm1vHhvL315MqBRwygx
O4c18SApESC5LnHiiNOUpnyWa8TMtf9/uaxn0hCRI7v3pAQLrX6u1Pv4rcY8zM4Onbx+9LzOVoDt
a/OyP90gDfck0kmLgDmwpdDXw8l0djQy/uycJ4GTCKgz9jP0LvVzI8EsKgeoZrT3BqVctp4PMAfE
MwTU00tAXJQxw3vG363Bm/jTHLDv8hIKEuC0qKNDMk1VmVS2ZEDRqvd3maNYf+ZEOhccSosoDaqT
7xIvDL/aWNEbZcKlRra+GjTMkF6F2SDyeuTyu3Lye6pt7bspLyr1g9wElUggu93Sqal5KHnqVMrM
Jlzv/RESZTdoWRNdnwkyC25Y9+kdLUD1qknPouEi/vV9gyrbYEi/SQEt2wLJVKfJENsUgNqe7E5J
C/KfFIp9AxDuqnJ7DEwOVgAbn7P4w0MBpOfHPuoQgIrJidd+mUzBxB129x/LijvQLmi19Lozo9rW
MtMqFhl+ifCdEc1TOMWaHVL6/qF3xsOBHNrjnUdxrVFaM9Ka8F76NPhrpbqeN1ocYDF5nEY96owv
KlEpLgyjvWeBqxAIlA5IJEduiuhiGq+HnEgZJvhFgHtD0o6o2DqV69DjLIuHsCFFrqEBjQvTsZT0
4UUjmYNU5mxUmLELx8EFIzdvcDrdHrTRS1CWsZ7zfZZrsiKsI8tuZc/9yUpaXnQSAmG59PrWFK35
a0slnwMpGKUnqCdDk32jl8QizYI86LYqqs4NCYfNbgfufZHjHW2+TPkZJ3EMH/BAVJFE5aPBGOaQ
iQ47T12PHmsQ4eDN6OG4JkHtIuqrJxKKc0x45Mn+AII70vhRI3UWvd0sQ88hEbJAo9p+CL8dJUms
SofC+uNqSM+k8V5OB40Mvt5uQgRGw7Yz0yZ0dUzcii2uX9wsvE/DF1Em4+kLTkMstsanxa21ovhe
9eYz5tqVvCGB2WalW182dFXJmAGo7GbMI31hSb4lt6d1yjO1m1tb4U4vPezKVsvU3DEt4fT9ldC6
6oKZT+u8bpXYWS1QLZe58YvfxGJk1MJhT3EZNTPFs/LbJlxnYRo57X7adcpHl4nDl5i+KcoZHlsa
XVZbGKXiiKQU7qQz0VbckFjwJ2s7/wmYlAv4O1/l5MEzjrqJsXWTLkhPM4IVRrRO+pHb3kumwJNo
/Gfte+l9mRjqteGX380MWIn1MaHWQ2mcDFS+vnZGpx7ObKkkxmePvj8qnxt/fA4tDXFZE5vsl6fK
W9+mmA3dLUsh+xSxlgXX5SfQ3zhqN2JYKbD1MHfyjgXbK7qmtZYP28Td7uX3NuWwjmkpJRpEySqT
LtlvWnqEuuUbF8aluc8KJaihtJAcr7RuhbNWsAl2UGKuLDuPTxUEY2Ki06UMk1L+IAyVGxggi7K1
+Ila4WcGjpAUktl0/FdW4UuTPl807foKupBUEu6TDc+SXnkbDUahy7NSP9BTaS89UmWLHm+ndmyZ
RIKiSeTyxKTq4KcmECL5Wf1GsrfKS8KlvYxpZv7qT3xUoIlk4+ulh3qUVff7vVv8PqDOJ0ZPcKw7
rLeqCYvaFX1BMHtO8K2gSJ19MrfuwPH8dao07tzawkC1U/GecvtRofROZozJn5A+Mv29d7+gbUY9
1QfZno1u7X6bW/X79hbGotnB1pGE+VjRNiYO6q++sNGyzRCJ6FLgdB9L6CSnmInSkMeBxh1XaNix
fxKXv7rSY2jGRAV3eQbkxH5Pegu3eg0MSX5Pd/DB7ivCCKOF8xz7TVMvdt12LfObVyyB+G6VBWTm
meJq6CCc2sC55J5e8a8+iN9r2SvP0P5yIV1atWA04bhs0PFIKyi1ou40wZyg2KQ83t/S23hnpCSZ
Yb/Lw3U8a/TJyL3MVQR8bXWgadoZI5xXXLjhd9UK/LdLvqw9U7HVc+QttSdD6JF9MTWzCV5BzG+Y
SJcPIalp4PFUXcMjsKOUIEMui/G6NqxpofW/9n7CE9NiIVWUmAG1NybmTJMngjmC8Gl2zpTrFg9R
8ER7AcnmEQfIblxLpdjltrXfls6xeURLehp3OGAje+7wUzhw0T0gutkCy0jztj4i4fJy3lpbO0rV
hQbeWDnUKZRmZsaZcOanKPt9c4DNoYRES/x4/u5Xz7CITa5w+xxkkVezafombuz+d6P3Xg79HTfZ
MY2UL59V95MCU02VQ5utf0499GP4sslo2T59z6wqvniy/SSM1cm6Tq6BecT5iU8c0rupu5d/RCK/
kvwhDBWe54usIesJwCFx53KIrzBpU7ZXmE3fJuz9nP6453BWJ16HUb3QkFf/YhNUa76E3U27sSdv
2q+O2D3D+LBQ2GKydZuh6Rt5RzoSXJbcD6S3oG11cyriAGbLXCEUWx3iL7rS7OiMlP4vrRjwMEAX
Xyf6458VawmbBBs020zc4NTq5C83LST8S++6AtLsCrPTdbqUbfqzOv9ll9vfnFPa7M6TgEoym6n9
oDXC2ntvUbTlBkcgNTbd+XSbI2y+3NFqR5nE3nreGWb+mCqPJLJz+zaxlwrtIL4mP2oj8NllM/3M
Slw8mAFo28EHrf60yDNaYYZV9pcj6vQNcDcSmY66ISy/WBO3GviQenj1rQ+e17JGskMTcdTrphgG
XW3JIO67SjZuY9nIeO1h8hNY45KkaUcPrpRoc69/JB1gAodNQo9wZ6telNx0uGEOxyFV6/sueF4W
DpQIuTwI9tUfq9w+JWC9kIPXrqvyqIPiO6o1zO8q9xVzUhycPLo8+RmQbqCwHWP+N6wBbvLbwbaj
4/oVt4yS/e5rjStGA4elwhxa8nOqnc57QNEubLimUxMc1lgfLqczKcBPJZ8U+MyxXBqZJbqBD406
T0g+NdOWZVmilAZy19CVEerjjbtg2yUzfZ1fFBjyoSNa7XPGduGonSybMZz5n0ox49DUWEkcg3rj
bWW5+9KHlpidtNrxQOrNu4qh51Toa8V0vxEd0t6GfncTA/pN7HiqD9OF3orGGG0uoOKyhkdYDHWv
KKKZMNGhq5UYmvs7fam6sf1WC1QEBM3qKSWfZqEJSxjm+oC9z78aaczLLHEffhyU+iK1A+KL2nJh
EKY7nUmACHv9oGHW4fyfC6Vq7Ubo0uAvzfYu6f+lGfGBClNWk41GoJsFoDDYKuU88h6S8KnS13dh
bwpuAt0wSabRAn5OPVetHjZdWFtZVd2zFpXSoGTgI8oaFeG2AoPiSIRW1sxf1Hq2mzzQ96iTjSVY
U95ELXcqL0a/8CUVXUqGDQdZZrfdE9wRHsfvVBTg07zUr1zqMJIb6GWSkZ1pxfmMB2wuQwBZaNh7
WSag4zwEB8/Qff5KfDtU+psyOEItzTPwxohQcOpjC1gdUNRbhERstpntEgWUmhmOJ+59BYNLoHwp
Q2pHwxBJDmwAT5z9+ZkTgdhKjsq40wzNM4N0IwCLkVQpam0eQwLrKJEL7nYqSjp2pX1yMLAdKsqV
0el6Z6TQIcx19Lk4s/5nhmGHokCmZpdLNySo+iJ57jo1xjHO1zcllJ6rFWdEFGSWginADRl7eKTL
zXWv6sb6MliDEvoz5cV5ZKdPLwJsgXHyi2TAitSgKQfeZmxcC4IqG8rxxokHIc1Vln6vPKo7vfEI
LcsJvjAosGfdhCOSiJ22UhQY3oeLLpUW8o8c0xOCm4m7GJL8iQFh6YdfhS4IFiuazOyeZ6BIK753
n8nnRDZrf8PpktEFaBwbsU2X9jkvUmNuOqmcAjxaUBDAbmI+gAMH2nf2BKwcfdqa8Ds9wNEiMkH2
gXwsdwVDogYQ/l2BcNQB0g53dpNfqizBM7PjORp/7aIg4m05L1lbMlR5hm3ItV2IHVtFXlp9htPK
KG5cFi+TAOZUPTyz8ogZlU5HBuIwszaP4zYklj5rDK4VZkE8ajRJRTgZb5M/hCbQWk+1evz1I4+C
GgzmHoMK++0mtY+ON4jaudWy9eWpw+JEswWnwUDx4w3qJD1l/uu8oeERuRgTSRHOEI7DOc6XPqKW
/JXcr5n3sWvs+EoEjftA5pGXnVVXbWn7d1onQoxVkN9QZEED9XTIk8WczmuP1ogS56n41+Man0PT
swBvu60B+3l54FR/te5GcgvFyRHW5Pypd8/28oMoeipGmOBG5zweYjYT4VJVEQtkGWSbiApsaDEk
8nBN6+KQgQuTNTMLB4K3WVVP1BFimioLPZlXxzSWHyvkXx9OAAtbl5F4KqapZH84jI+kR1e3FJXf
uE2v/wOz06672kG8fO2dIxyHuNS9CUYBjj1xE++9LUZ8RLgAhxl1SbGxeTvobKcu0T6lRu2mNlVA
AczKz7mI3WvjbstfhUTi9v8Dg75llZTrT4sFGUbAyDskjq6uGpQO2botLIelLafd7WeodgoMNoo4
YZz50BgKuefPy3sN4T0xao4Nai5dCEjxNWQeCzONo0ISWi4fPqYn/f8nackO6L3MJeIcL3XQozqF
aCFLbtZ97EroqacrsX5ktEWQweMu8XD31JNzi6861Zs61w0/mjAGG26gldJNDU8YaUoBMLsBKNKc
95EmNHgTmdJJYF7LACM5ycXMHcCTYHMx2DsSkunvkoou9ELyyJlL8vQU9qUvRJtMyHBzaeJQdlvo
eNTnfSGs3ndv0HxbZH8rWpfEGhWvYGnH7kyGAYvgb5A7FZDMh4Yk+l5jjmF6OGPBiznICrk/p5W8
NEe/pfTNCYNAD3eAoz7tROdbfpNR9MN87nw7j8buSEugGgz40p/Wc54AJ8a1lHHOyKJRpifAFxWU
84FAs9nR5tbxmQ0YKNE9gZ7C4erLB8cll/Lu81hpdeJ7B7TOfxHJCmrSaJ5x9548e8EQeh33JQt4
NAe+nEe/nuHnmFuAx8v8nqzBmB4nZ75d5Z1aduoIHLG0r78V0Lk5PG8JkrlCShYyXhq3B5hRNbub
BFHdzHGo/3n9zQIM79MXvTbrdPOO+s0VUFoauEaN/EcE6W8cFjeoBoog/YG1iIJWXKFvfxfh+6wW
GGik+9UrTHB5ha8xUkWqGB78QBEvbQAiHafAjc3POT1m/bSpqXvJdgi1P02UlLQnLcym1Hyne1wS
d9wTfef31+1bFowg76zaIUs06RsSfQ3c4VISGgd13LM2HoJvNXWkbRKqAXeLOVpm5eF9F59UbVa0
rhywYgd4EMUyANV1cxIz+Ma1FQatd7LE2BWejW6iyIeJKBtPh7YG0EkyRGskSDiHL6ywx3RJaGTR
gtpfceDou5jUTgY+aUohGP9OFnrxnPc/stySEu32xAcAooWQrYUaqcOjS7fqxn6FDOH1KU/7vD92
Tu0CrnNPrU/vtO0NBemzMbw0ukZXe3rmpIUtzKvQnkjSnlu0VeRpzRFtX5Cvua8rR12xa8fPC/E5
OLiQ3dL282HJtH89uLtU5fsv3sO7qlbJ/Pqxi+n9pVYmaQZIpOSALAkS/TA3XJyVJEB+1o2r5VYK
hrN/VCqtI6kNKpXOpN8NCwszq6FmXJUj3kEsEGnU6tuIMet++N1vHe4HdCREjQUof04i/nSfI3xR
JoghNRLlNiNGDr4LdOGz6hlgG1JDoSzBQrASvFtegzN2lTag5J0YVNxAMY3E7bzKszvGUJuopZRM
0i7x27HoM+TvnEB8XbciJu5QzQ93SDuAtjWbaGpSBVspkMVp2rGynRvZmr+sMqpESLNHC6Z8dvLZ
K2W0qIpuM4/5rdsq5eGdtvIYw2l+OywXNJtPvUpRhwmfo5Hq4gsiJJ8fDFO1Vrr77SUCtNsgHSuZ
A3HYjknXA3kVRWReFENFMSwEftyJ/Zn8kPUemn2PlcmlMI7sHido/vPjg4iqWy8TqA5wUpMiG7Wl
l7LzPz4bT6NzkupYWhBq8LhfcLryHk/ahJzybarMRc/mpJvycA1t60hSdVRGQYMP5p0UJWBPDWLk
YQU/T3OrlmFHOQ6bS2zK8WWh3JjBghHqiV20/luT/FVR5t91akaJJ0PYIDNzWsctd+ngUCmIiN/E
fMr9w1KxRpTS1Ii7VJO2DBarAxRnXzBDQYy2H57ozKHVWVJ+NLGAc5FfLWTFoRV64Dti4eoFR35o
eLWe4ytmC75Sool/IoqUiKEQuFs064Q8WAGkCDcLyYHTVbcJnJJ8J8ULUBjfWVbuhrIi07SOKTnJ
1Unjw9lwKWH9ASPflvFHmktBcJJWZ0bBRLFTNQmlAgTmak/Vob+7N2Zas2z1/7z4VxZLXq3u3Onn
G35hlZOyD9QTrfIVXeH7PRRxjGuRnGyUb/qBD5j/Ka2EBTSrJN6BJX1WdisF+Y+RE4d3l6TR8Mvx
JvWMdccTeXZfS8HnosWIsJGbUsEz5xIn6TsMkfrXPSjnvgW5tfqpDs8f/+TcJV+Hn75d7LGz5CmX
R/DgBt2wUGf+JO9YIgsvkVG1BreSSt6omqnarnrQr1KZZzV+hN8UFdNCWIfU94n5xx+qtAyxLwoT
diQS5cWUj+pnhZ2B6Qg5KwkJNSHVtKw9anFyWH/iZlntH99wJ2a5RkvUlP35/VyiUnDFNCGlx0U5
ablhNjCXp8ZF3rdXHYaqQt6Do333xpIVl+WA05KUCJ+QUHIqdfkWi7MrPSFrQjimnChtrxLqOMhM
42V09p+kQM4GXlaHaD36i5ROvozbphwLt0zv56dNYZPOZqOiwUlfbV+LJPN647KCpMneRqjEJSli
bxuB6xIdbQ/VCijmcbzGdQfPu0Kd8mBwFispJ2puS9k1Z+C92fdylkwexF8fMWnO3rdZniaWxSn5
a+Nv2KMqTW4rC4xs8COrr/X8Nh2hsbkxBwowcFCGVSc0uu/ZyL/osYe1v7T3Obm3vVOyW7eh9l3A
KJn6SSQiZWAd1RWIuh5kf+emVgQeMEzAi8WesUis9isT9lEHcjxNyg4pcxa6KeCY4Xb/f0HuSJRt
Z9l/Moimcg55YQvuAx++tTt/XDLTUx6LNcmf06XGIioXiqPQFM/a+TE4ad0CKeebtPhl4me/7/CE
zKHWyMiHs6b9RzbxxhS9qy0gCLM5ucq0haqlLLV47gu2DgyGzRy+rP68YZTHmpTyBB2IaMm6THQK
pYwZa9myd9RFRjU4mrW6cqVKizaykzNkiEsQxjPwa8DbnvVP16EkrB7yqdXGWwPhqTNI8oD3vD/Z
MnYx28o+w9V+oYbY25OzzMPIp6n/YzCS2dPVIq843ZbEvTsDi6THrltAMmoQaibwHqGijuCNqWeE
VlTR7XKCVsgilSqaTPIH61Xce/8sXIA0bOCBPK+mUkkyL6RYZJMBNaiSz20k2NCkgaU7lSlx9yP4
xPpZQ5tLtUe4qPsRQeJHE6gvyGWd/944E82HTUaRUSM53Xli4xfq/ukQB66vOGNBT+2qlhxRFFG+
hkxfs5eHIljxj0ATE+0cIOH7DvV8qQe0cr9E0XwNtwL/pVWgxjEjQzsB1wLkYz+ORm4plocvqIQx
opdbdPFEogjxNaS7zXxmMHOKZkfYNQgYgHYUe2xoUPvVax55lovZxPNlKth3qXb4jEsEYfQbYotU
zgeU4TgG3UArRcAxsjEU+rnei8jUIojN69rixpx8zvHXNbc3oBPwJ6wY3W+Ugyjm4BOyfB0KStnN
Lgu+ygRViK2Rzj5O28SPNQjspkqSKdFEZ8fwfYxq1kg/7tC2XU33ZB1YIU/1d4fN4SH2P6hpzHTz
XUlovbkXEIowEekrFX+QHEjm7WJTLn5t5X4SoaZTHvqeu27g3l8IZkweUrN48LSc8SgJnC8eyPqr
n406QrFBj6xTQmY8J+0b75rAZkun2XYRegTeJc22e8+2gw+rr29IoMk1hcG8SwOx0Jx9WVO691Ra
uEmoeHOSppgV3Nyqn4e8m/AGSjLhhpuoO/KlZ54fhbCuBuRaf95Pp8bo5jynazOsYmjiqikQ5nvy
WZmPK+ILMxwiCPUYuhzR6iGvOoqR8Kg4nMsVryEKK9b21XPFqMFvV3I1vCMO8bgzxvGxm7rUayPG
VuxNeO6r0ucFW+tcsZMYE8GK0y25XOQMLH0kk5T6qwEO5vNNg8q6J76aFormT4EDDopfNbJN5qbg
kGY/cfWNzuO3yAnCl05FtIkYFUY8czhATa6nTo4nq6O6FUnrtV2XgMhv27tMry7cwXwz/Ra0zuCE
9c9u4ZkxdLupF8+fDd3U8UmMA3/hLsP+SUDG9AJ3JvDlwfvyV2i4QK13iaoPF6z8BggsW/EXI5hv
63rwaqvTmCwKu+UDHPNUzMkxh7nNKPDO3Q/RCizwceJrLeYUtwBYhwN74KubQJWVqAmVTAMF2TXN
bfdgpvN1dy9EWf/bvPo9akbrf5lBQCbBWTDieIblyxotRaYVGwtJ6ia3y0RP7PUyfMtRzikuYJjp
6xYoL0chkj2CqY4dQFVaSVnpIAQSEQZavDIDgl/ytKWGeURImaVLKEukVRclbJXro4cmnWWa5wxj
wsRMGSCNOuTgF3QR2EEzNYXI9eWS1m/FfJsT8Bcq0M3dYhKEymfURgpYflTo47BvlIZqLOSESKF6
SUukPxZYy7GmpOMPNED8KMraAxp5ZZ0ISWQenSjojB1kvpt4XelUr4gD9dc6LpXgCmg4Q8VdfovR
hd1KRL0KdVzMtQzghuh/EAcZd/CswwlZ7wcQRFUpKxcCnbqlcwxItaNQY/HXwg+ukQZ07Bk8asHl
raGNMKSveSTE0iZDKnarGKD+uvgF6k5iQS9cW87eREkfEvmmrJZmq03fmc3dpdQokTZSQ4Ax1oXb
AgrG4MISM2EG30epUvxAIo+wG79j92d0AOiqzBiqLUYqj8Yhn/Np/GhpGDG+YBi0AJxcUYeWi+PN
IF7ykXbUOYOYfIDZVCFyG3Bx7fVfWYPt1asoOmNodLBEilR5Vn4lfBSMssMNS9Cjw5hX/gvmbtba
sqK94Fh4tboFWAQ+Ekrhox82FW/IfEFOQi60+DsvE9ag5gwWcVyoiPoxuVskIaKgadjkbdSp/8XG
6BS1FErz6eO7ofaSlCMuUEWI0PVPhEfBXGgrAkiSUZCpF6nM9TYwlZQEMG1FVroDZtu6GyMkZqCL
Q/m/Fm5nz/oWMRHM277E0kaWh1272j4mikdigl79nqrSIKpT7BBl5nDWsUexv6wgsCvz7clekZII
OPA/99AZb7zXTPj0bnhytcUvUpSw+YdxcmyC6q/VrmUk35xsViZzg/xAcGlWTOJMmCTXt+mSFTxh
jfIhs+CEkETu/yWihQ1ONSnSJA8oSGrNKNNO8gucpW0MCKGyGBZd27xO+a2fewDSysrmbgK/muax
Dj5D34TdZmiV11Nuweoa2Lx4zTvtYbotSbV41qUvqIL53PXYpdJEh6w3/xkCVxkZhnYh+MLTS2su
dHjwgVjLHHagi5szVRTNWRRUaAWBN4A67q8WKMsjSm9ehNKgYWBuZaRX/RWfk6wURcywhXBpWzi9
Zh1lq4vKN5su0urA8JPZl6X8WlXLhy0SEuKrAo+q2SSirMTVpMM6wJHYNp0vyeWGAhVSf92L7r+h
IQoGlkONrFjr2CSeI4zYW8V4lHtc22slgI4gbc7i9rmeFS/QzXUKxE5hDw0fpCJliS+HOjkYWalS
/wXLnOA8JnVFM480f5uM+/TkvSgFiGGc0DBpB5JuQmwfwDfpSaFujDMrYqAMZa3f3FRA4h8iBBVn
AllrNoqLZ1GKB8tRsf+7JveXGVNYjSf5zDIJCp9SpwFznnhpTPD6OXmFjN+8R2Cdc760xjxHvJc1
QLwBJachccROML2chZwguKX/cIsNbIMyUIVsv/JrVr8GlyxXmNnGPUN7IZ9AFnxJCu+2KoZ6Iu5d
5HYt4l5E+F/XMbmnNnpJGngVTlNtDiVEKxvn8iN7adNkav9vIV6f4j71K7XPFb30CtjHK1Kl73ig
K2gbed0OhvI8dfv4DLzH3g/+UWtCdc6oQEnSXuZxUbe4tuDCna01wtGGS4Zb8h6Z5/KiHLEzLJeJ
PELT6yFLOUvCAPNqcFoXoiAMIDKUJGLEDj5l4cNtJx6jzLjWWg2SjaCQ0WKaNh8VIyczKp3+NCsr
r+JlKa1RTXbTV2rbVVTfbIBPSHfI3HCIXW7+OzD5D9sePpGRBxlbkqNFKyH8PmawadIQGI5786dN
x3knufTGK1iOYfnjHdPMY5/9Ofyz5ESm/KiZI4yh9SqGVv9Ky8bXgbPjrXfzDztBas3zvT2LOM4D
fixD+iI/RrTk0V0mBqsSf39igYoiGOyqQNklR2DuUHOdiTvUrdFc92034l2tjvGu/0Gs0wxjJron
bgsa27OIl+ACXEN5ehSu78Tcsu43LFv6pun11O0zwXbNIVlZEHVzYEL/eXSbVtIR7KwszK62ZYO4
4Cfz4CiRBRW84iST3eeFo2Z5W7+z9PY95qK4ZfE45y6MZFeSdQosaa2cEUBlEpEhS0DZPnft7xqT
FKkF+lyqJ96gpd6JzlLxIGa0rN6wBhH6MvfnP6yUjMDLwTWX3ArU2OJQ/2hhf1OOtJu0Bx3laNdx
uPCgTTTQmVJhPEERxoSNV5tvMHoerJ+bKQzOvr/MG23brY9OeyaXfmwnGh8NcXkBsBgvaCvT+Te6
KUeo9CPvgKrfAnNPr5poGkiZvctHw0ae401K4a80xw1IynQox1Nv7fRYHnHnNvbHK+FpUN6SWR4o
Y6WgdjYdmXBlk7Fro4LL/vKhEwOi986CMuiEolSLSUj9snI+/N70ms9P6mGYDItUi/vbGNU+Xa8M
a5X43tZd3q8fAKvmclMhQu3tBpLZ1NTuQnyOG9sLg0BC7IK71/wYbfJiKujU+6EaKYTV+wPAuiEF
UA4Rj9Awk+taL462g4/i30h6TIiKBCXcYkMrZ3pZmwE9HIEXbNPJjPHENbyqoQvrDn2/4/dy+1ha
pFLzRHqWQxNGxdR6dzZu4ZymndxsFYLQGbhh56W9zxvvBChv7+VGLjny49QmPwwUkJcIQd4jSCHN
IcWSUmgtG8ejmcy0eYF3atrxYdr3KJtUrtb89n+Rmj0meZO3dATEO1LQUfPrZ3CBbA7Q4A7FSLmy
nQQXAJUD8AxL+B6hBTEyQinZioi1Q/yqFul40VCbunqcL934/0j4bNmMqrUihPjSqscW83YMDUHz
21MwobouHsWWuFm4y27CoL2FqLyjimkUqG7NnQvOJ9xbAHf22KmG1n+wzzzRM0gaGnrKF5UuD7vp
tOyj7CVn+OfZWokxwmnbNPOqRxdheNZhBDXZPuOukY3Vt2ICtnw0RBmOEWmjWNUuZrCpzsD0qbN9
y1vO8iDGPPm8+bfZ6JYvFuCijgel4GfkqnBtBSXiRk0KbsrSjlVeSGmW73LJRicPdD00O/eQUO6U
TEGaBpBzfJ/7olIpr6jskB8aFrbpSwADDArp/6UiQKUzzdmHiX284e8Thwsp0Art+3TIoZVTB8lZ
LZgj9qrDbJ7CRpC1QiGM/59g9sZx7A/gBMsdo/SzRQN5LrIf9Abu5LJ9eQBlD/f5l9NdZNIOvC4/
25u34/UrasUVkwOdQ5VGbhJU0jQcdA2ezv7WYPJyw4o7mUEKCe77Cro+QGaCWoOPIpBFLaEoT+m6
+u1zvIqV5XIwnYD8stDELBp0JTgfKocgkZTdp1WnG8d80YTAPVHjt5eaBmr04v/5oKemXqFGqhOx
5HNKQUai9ASXm7+T4qj+OG5IXaOS7HFsvEgudsMdW9BcuSIhQaornuLacgQn7OuY8O2jmfuaRdRS
gpqWHAIq6OPwfbntTw8HjmaRVkX5JJN9SEEdWLdqYj05u5sdbIQxQhRjAj6vq7C4DCdqNpdarh1P
rote+OefvtxVQg1karqeMkyN5NaP0ovmYgQRdbm4qscSKEp2SWWLTQ7SUsu2kBwVBq2ll9MJDwtS
42aDzUZDhP+DK3wq2pAp4CKRkH/SpeHP7RmgYH3CIPVjNep5oJPO4JYt/SrvN3ZryAaG87uIHZ6+
FYPKQhSn9f54QNrW0KOAosNbgCuGtbjpCS6GYldZezec0NLSX9Pq1W56kU6DbmdiPLoXU1eC5avE
FmmlMTDGP5N7iN+eO8cak0Uqsa6UuJbBpY6j4J7abLTbuU1qid4pWHS5pBgGzH4hQ/p9ko2QHPwx
KQfrS2SSR7vOWf/coHqIcF93k5jhqvCCPtHCEN03IyEC6CCbGtcYJRntqwKqirNrA4dVcnZ4Ysxm
a25bzdDspL6n8xyXFrAX9Ph3dcEiY5bfHGHBhW5RClNXBZYBLQqfVi85GY+T4BibRuYoK9uYpuOe
8G9sYKmTheCF0MGV9EfZsIHOIz9mKyVZBRWT5cyaFSgciX2dT91NQH+0f1c7IV0bcwqyrrdvg5pe
4VOab/LAVmR+ggyK0AL0oF01ukZ08pJ3v5gzXzNGg3xqTQOzQJ8NlwJ3aJXPVftnuX0Q7FEnVpMw
KatpKGr6nbbITYxYqPCBeyKrJDefPP6QeXxiukGHK73ohJZ8zwbOu0WWOgdvl4A6fjXkHYghCGhE
xP78s60xzRceS/wzwhZO4SNmeEGB/ap4aus7ACjgzODxE4N/n4lFMBiJqGQ4oLMb6T2DSnLYDlfz
L/flLgSj3p47I5XZNNhfOcZygn25vAMnQgdo+80eN4OuphodGkgCB592ztfeHQTopRjvHTeW7guI
oqcOq+AEKC9iSOgl7DSQmlMfpfNGaFPm0OqxdQfC4y8rEIPM7TN1z5ESZYzzWtjByeJL+q7yl8n9
D+2XPYNdCT00psUPF80mF700MdDvhQIJFoH2AK63v8tcC6ByBHjXNzi3Bs82ivCiEwCpgVArbIoV
xGsGZAnKajVMF55RWJzM2jGXQ7590MJrprXCT9CnDIl25m62l3ccXYZPXhJno3a+33YvrMXCRrYy
xwxrad7FW/5G1bXZQwjp5vikUD+NPzJbvIYfT9tqO91KmWhZoZM1+t8JxP5qI57nf8s5cqlgD9Tf
1kbVuSif/zSWwfm/pqEKznT/lYoIFj9a7W+kdpGMtX/7fubhyRTet6oZ9GywZ+VfbSXsM9+PuHdA
54NcDfCRTdBdqw5u5Gu9EN/6IG2ABQlmbZnw3Ypc54qhZsRsIxg3uiHVTgYv43ueoq24/cs9hWOd
lAL6TfVzZgPmSxecPco53MWO2dy/Nn/+gmaxeIccdN/eQZyjW6jjMUEdHfFj0d8kKPqY/hsTFHiW
n99gY171iPWixtjtMGGqxbu4LKImBGAC5189u6zDd9W0MrAevGdwSHWv12L7+v9wqRw1sxp9TuhF
AUvIWDsNu1/Nj/qsL8Xf71dWR3WMOtGfsUO8A+0DDk8Gun64J5/MJJnFUwtAd0iuFddVac0Qeo46
9d0/BGH/jaaIHAmjXedVS0Vx6cdy4rov6UZ7VMBZRNNQ/+ZnimJImdtpV7UNQiEMitTGYl6euQgR
8BHN3ufgQ1NtQ+ejz/FG6jv8rGbJY9mydX1hQ01NDxPLhjKZVjhl0r87UoL8M8+a7Y0JxbZcI6k/
RApHYxjHGO21jJiYHOlN8A7fPBO4iQ+fX819wK1VVanGvffzf/h9XBOX66lxD+Kmd3K9fCkFVcNp
D97FO/dLPH1m0suKiSxjDpJG6wXTKzB/mjLEuxbLzfc+rGkL41I7zVh5z2Q09ojOXsG1P9MytHkC
2YLKCtJWRhR3z34gxboTKiuD9se8XfcJVJkuNyQ+/bqEnm3TopfsMGvSp2GCndPyn/BO+uo4Guuj
n781yLDt3/XHL23j7R2QGf1cYo+e0HN/ofNBIPXtDEF9ufpKXZ6vehB6bMTfP6i0mRGJi8d3fnuf
REcqHanQ748Qu1uujCdysW2O/+7uD2uzpxR71fjTJlJMrw/sx/zt5hp6SC/9R3gkCmNqgzziEVtN
Kn3AFjlGLG84YiObbkTKyzqaeM17HnvN6X4VS63WuOlPc5mM988s3BBAi6xRdmZglgJM+C3PNlLd
KS1wOT2sIECtOeLwRr2MlteRFVmMNeHGt8wfEBSCNlD7DgfPq+hizYdHhq8hAAIsotyceh9lgw2o
C95gHwg0UjncFa3x/2k4B50WwBCn1/vyCrinCrhvl9twt9JhRKqhL/xN4j1m8rf4qaJg4cGevXUp
OB7XNbGuSWLmcYfvjL3YuC0bYJuAwbIfqI+ELN9N6xNxBy7ZDhqr8r59y77Djt6RYm6eL2s/wdJL
1kE0v6puZKlpx44cTEo9LIuMlBsReim+AfFZHzEyY10uPp41ZaTJ+ClX1Dg+nCpibGRrDAnNAHH5
UCUQEwAodWpVGfgr0Wq181ZPo6CEoD7Inxp2+kHBHucAP+a/uOH6H09E9yppJ4lR3qUiElUoDBUl
HBIum6rBbFEhwm2Xc8KeXHiugZ7taO2WwWVJim0wbDzEhtd3dQi4V5z5ZR9xngpVxjQiWOMJh7xU
8ppjMKqKOiL0FXYnNOdNsAzWRWqb1kCL22MUHFsCUgVRBInPKoN7wHBDTx21SfZGaB4Ze9VwHYC3
JAp67sQNsJH4rFC3bg9qIMgt27EUWJuiAA6sd84rYFKReoz/DvHAINEc/bkrLol86VdFL2sBuWfn
KVyE1SrU/Ji6D7/HbkILzcWv/Vw0E4r92DKqh8kE28AZ4eNaeZJ3Ic9RxFmD96tijqBEubBSc8If
TlIaUxBqpNXAcpSDZZM88+96/nj1ZE1vMUKb6GMkS0bvWtBJmUq3c0px2tWFYaeYsQ3mRQKeY76C
Sl0HKIi2X5osSxW1XsHCtqWvzyhxKenGG5Dc1sHQKEj435J+95DNi0S2p1qSFfK477MJ/87+migh
Euag/hOraU+JrIP2de4LdalRXYzm1pz2V3CZfVKWsObTfOxqoBWG71eGy4FNdYqbB4AG4RRMy7mm
Zp+g7yCxjQq4DzRdqknxFNZTtPmfMgCwI8O62Qpa47lpe4RSHGrf3fzpbUpzIxIIJsoUQFsOGzgg
nfVeeBDf59v9Huff0bunAwfqdenZ3My2P6Pl4gsqa5tKBP63ypOepLuTIZtCDQTu5xSCZVok5BFj
XyP76gprSx5Ducdv9HVI/tQhUvewpRgJFY3m/imQoBISpWnURPxxiuz0io6mBVSYfxg7burKVCID
2A4W4pS0REvTiZjtfbH5ReXTDnNv0yGIwZg3nTGXhah8hsF/QVgM4eD5EfZe4T0n8HHwUKmNyMwX
gzwgE45zb6zCSYeKKCgmqnoYcUjInwPew/AK1L0vM5Vl1+O50Nmp6H/JRKiW6vmmnPi0xrnd1zfI
+kbnZZluW9mTI8VyTYCfrIzi3OfLdqbS7f6qA85/c4bl/GZTCP1m5obCxDqA2GetZAFamYGHfGZ0
9nx4NGnPehxLv07qIUsb5kXyLhBJS1Heot9r3tTt+Z1XrMO1UHhYrCiyc0gWs5Aw97o3UmqYV+BG
JrooJ0zOBfaP3EKjLYE0eABoufKIzbkr5BBddI4ZhKLEQ9J6evxamwDpiLE65lRTIPhGI6yoSuIB
EPGlrL8bYXwpLVhaOFNv5FoaK+oqScOQnL5ck/3ZRJsYAxdEeZ00cb2GRGCObh7M0sW6RXfJ7Pnb
Mr0brR7DBbUuKiiy4Ik7XomXl5mGdUFNT/uaNKM5lUk7sXSKA4pjzdijB6WTzlvyxY3o0joryrrU
esHHJQz/G/QuCYZ973api9MFLm1Ms3aOPy0uIlJz2sSc7ED09QMpXXs9/VjAPc5ad/tttrxdCbCI
myntoz5Gq+cNQHuB8zxigN7OnBqsotvU+rifuQlblgmry1TGSjOtONXn9UChIooLTChZd3rElemL
JS1Z5LijNBQFOdknYsPCWIQ9ou5MyZSikUJ5/qgdH2S+LVnHfSJIdX0iuNNnaeef4S4t10htTV5I
TieRGZZic5nAWEb1QtAPnsIZDLeJz5DvY25kZKCsHcLkqe573qFZZce1k1mozvWC4ScwGJk/Zmjh
h3k4UM6Jis8mI2jpSskBLkdfaDMo1NWPFnUQ3Ic6Y++ts0RlkoG4Uuf4JUejhWVFNBqWlmQRKltZ
KZX/S3eG5aVbZRPC638A/7oCFcauSWCesmb0QbEQhbdIt0r8Q0Iw5GsBFP0WNeILpmDYEWf30s5s
8FQDyal2hzNMuMlHhrhJo+l5ldHAO+LRuk9XrrnxE+/eCfW7qv9islMOVef/jNHmaw+JpSrfc0EW
JFReGuD1ArAGr6CbX3Y1ini3kzVYN7S6+qOPK7jbxS9h5nVUX95C6uViFFzFA40L6FpSiga2QjLU
7oF9M6hEW1Dw3jCoMahXCq2g2rVsoLwEWKLzr2xPpK6pDvIegg62TUWsIBK2fTnqjyKQPRZDOdVL
3i6G/UhCcwq0byUQg+gWTecXR2kyANwT/LcTws+9bVlph6JL18bRjwSH05KmleV/jaaogs83cS6v
gPVwICUMghtrAEbzst3juODnZSkQR5rCD55C/ZxNg3Tjrn09Oz59un0EJbjTS4K6/GDqaP0j4Z9O
b4yKqsBCaDsA6nmAOJkHfovAHn975fl5T8aP/9QroiISFY8PnBFFJ0eTbUrmwndcQ5lrWjDcCOBB
+xmJEXdqYnJvV127aFlrnl/Xr3Cf+1kUCL0jwZh/RHROH67u+H6SOjHGppVA3XQIumPfVSHaFSRO
mxj0MUxl2kltnnEZJI52rUNLRvu6LTM5e0IRh43Q5/mgRDPi1+XliH+GRwjUDXS2tsxkhwdIPrQp
fnjUY+yvy/rl5n/9wITo/xzXK6h/+YtubgEVEaPmm0zYZLXXd8lt3hN84NvchLMiv0Kxo3AdIyfb
Jx5zweLv5AfMH051iz1gE1CDHlupuYrlkjBMokZ4+EtLZymNwTC0DOu2pCWXja2+349OiuWUHQ/9
k5/cjqoygq7g072tpsGBd8kqUvj75sFOWhX+Izyno4uG57g5VGz5ro3Z6IoIhGHhe8BMCoB3Xw2y
l71Gydkc5AcNPcJtrkODZdOEgV5lzmxl7aK6YVDEN77AXLX7E0U6CadiV7iF1lMnsUuO92I6YY4O
OEcqvncE0gLsJPzV0HuJAV1Bb7+uGXlABXaCGvOJwKnk7dcACtWqqUNJgg1L2lQhYL9byHekl/5S
dn9h9fmfVGfkUiiht9tWIpwa3moll4EAKB1466dL+WAixLHeLLROAMBiqxhHDKKa8+LyVCo2T4Dk
VM601bvWVjM6bAs6YziFLfSeKosSdxFnnPo3GOhkjv6oBKv1YfW6gm3aYuhxtTHrDXMCRWc6J39s
IeE+S5CB5KE0xYdLDoQw/N80I/bs+UuTd01ydHxZxRdUSmVILAb1dqeofIC8VK5+OzGzh6GS01hu
KfBiB5KBwkRfFjYjHD/vgrHcujXraeTcH2vM/ifC8F73FSU0Ozjs8zY7z6gkfOvFzB6TInr+Z9ir
Q4nClJQVQPLSGmXFoSgPJRz9fFDGg81oNPGp1LEAOHGkka2AtL1u+yDiKB20mY8LoRrOefaXN//C
eV4HMiioeFiSu5uPTn/zfoHGMeij8s6TWhjw8ZavFwUwWzfaapDPMt45dEzKpPRZKD+49+l8xvPZ
weqoMr/MviaNeAX/2DV6wet47GYSA+A34e69s4Az1LFs8WgiHRAZJeQYzvfV8E1577CIQPiNKGX5
lo6Isn4+25iBT0urHFD1LlXiYmQ8CRNdI/p+WcmAVHaxIEbw22iVGZYmUyJ33zvWZ5rTPphqwB6k
trAkiRypzKi9D58DXPlaVSSLy7lOYuK6aZeeaVBvTrZhkt2MQ4JehjcsqdlDJL7OkbhTW52ZqSqC
Pn8kwrhjS6L0cURObbb4wRWUFvVD1X85t3OkGsCLUhY8tLUViCMFdLdNOxwmnvLh0/UNpHk+GCRr
1ixTYtp5GqUGl+dSD6zyJ9HFsfRkblHsZpjYqU2hvTz5zsRVevLAwLzUX+1as63O1i0GwitSZw++
PijSbMZqZDEn4aF2TGWVo2WIq21Y3fTA/eJWwBs/tnN7i+L2EPBjnYmtI/f8BvSQgPC6Rc9RvxfA
RClWzbgozdwpa1USKjm3VwnP/ZR43Xn7c+3U4MYd1MO2TM1ampEyZVUgFfNKUO+XtwIDfWKsxUgy
EPDLboLt15gvmrsrXg06ybotUIPKT/4Vic+zj7HP2UM9L/CJBwdsO2Fb+itU2ap7fpIO8I3oqCAj
HiImM0AHl+/hytZONY2NwX7F9AZdPp0NoYqn0sPc6b3bAt5LTohguxsgdeIEnIVHeNbOp2hXcoS8
rDnfGgaTIEmTOT0az0XoAEC3uocZtwEaz5o2Gol2eyfEjfYSleVv1QzF17KsD02KLIU0RiQmPtGH
bE5XWekUt/V9xusH9VKv6oX+UWgX+ShB2Eql1Cnq3zURgHtLVA7YQGjNPLe0vsSIlpKKN+oUuKWv
BAXLELL72VOFPV96AER3kBUseULnwNbJnPHY5D388mrs/7v+HH/RHuRwXIl9RijeenEnkEyLCqpT
UdO+a0dZcO0V181U+/p3jW3TY2kzpM3xp3GtO4luferCMy/bz/Q3RdcDHftBYEvKxOZoNWf+Md0E
keUxixt+ynymTC8h34cKlaUrobFePbMb/GUzsv7R0oUMbJSTuD5zle0UMWTZZv6UsrcBjiBYxM+c
24FVrC3bPfXsRRzBEx8ywW+JSYKiBKWIMk5AipZoDC8YuTLodGOzTFG1QI/YHI3QZnD49E3r8odC
q1I61kzUgZ/SPZL5miSP1KwsVwZ7zEPPIXAQgTUdOZKWMhcYe2kwuEWAwYOLhaqKFO/deQ6aggbb
4i7XioW34cK3Yihrg8ACD2y2hKjoSVgTZo8LxWE1CYTL74crIJttMAm9D9z5pyZE5bHU6XnIHLjs
s+DMkXEuLviuNnrd996xbuYaVf92L4pHwWCpXuk68Lf6/fG6XSoOX0Qj474118bpz1D5taDHVRFz
RK4P9TybtZtjKR98wLl6/CPDPD7/q1zOP+Ad9TdcZ3b93xxB5coQhV3KaxelY6PabZtz3Pl+PRuR
Kyk4qMxLc1xye9WkR1wXmR3MJrXyefMZwA2TSRqQKVMPgiYfTrJnz9/Y6y7CaufTK0gKa+77GqLb
kj1d4KEw/zalUVhWTZbD4kzdk0tm4DYlaAR5AR0NH6PXbxl3sSIhwSjiMrD87s8ObEnFVRFggYJC
3ppx9hOGml9SQmUVzZwJraIvFSQKHAHGKPzacjMb8fUVeu5nzWvxn47mmXYn1RI6maUh/mTDYYWP
hslgEEZFKeT7w9KKWQHuPC2Tt3/t9I0/D7V13Jrco6LrNne9Tj9/JxEBc6VCgPZOjjnEkmuv/LNI
pozimdTQSuA1zhCqyn6eX+2BctXBRnT4R6Yut07gN6EU/ugWl+4dUJ6CdEiQ3Gj3iz3fsLg/h2J4
VV/4+4M5P3LNCsBpeXTlIiC1esuMo7mDvC87GXnpiB7ebl9WO4VsI59ya5X6U/Yfl36VG4pSBK0x
89whtaLjwKCXUxv0XOsSLFBf3l8rqlDk69fFj4s5Bg9W/7e51tjg7JD42Q==
`protect end_protected
