`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CQirmkq/BKqR+F2Yg4UkWTIdFrTRgyk4k2iLzfwHOmDbkUM55Mewqizh4+Lf+dmwwhALeC71UJDA
8mCAPTmMHA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BYObDmDa8ddFsyZLooUzpHL8ns08oRugCcZI2k8wJ7bPNu9wkzUe6gLxEl5Rus5mNXhYLj63VAJ7
Iv4x/x3ytUfhu3Rr/6uxmrwyULLvv11XEvyVGCHx4t+Dw8cVgkM3usRkRQjUSA971GtmeHD/8MvS
cZY9jYskPE1Jpp2ln4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kh2guWzq3vblhcxdfJUid0wZnG6MC3o3a3YO1P6t3Zu5fbaVoJKIAXW4U451VmelQdzOKVHousSk
45IlwBxf/RYbtIg9YdXFrqworoOKKYA8Ps20E3y76/ejy57L44f0vm/NoFaa8+RGMVOrMaXWkAX/
5m2QReWMg9vAFlHZfrIsQnJM7q9vDbH/9XlzT7azdJd5gljApTrMFtiNcALEiKPoDWNj9DKTR/5M
z6fXEbBnQi7svJI++6ajKLfscdCdmkML0xv5aJaja/A6sBU3ZyweO65mSDcAEiF4/LGSrOI+kROs
k5jflROeFMl/1IvGNyU4OxK3jsBOPTmAsiyzeQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ybTxbKW8ZHek5yeUP9rGjX5z9pX54PPpKlEu/sk4QGiMGrMi9n6exyltQw3382l1i1u3uPUdj71P
S8JZfrL7/T6Wx0syH1SqEmm7l5ELtT4AmtRRmr7PjBfr1/vMkuv09pkrXQw9kL/r54fCF2RBbGri
s7+5RYH/ioAS6hXm/iY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lzavdu/+bN8Q3cXw7+sJQn/P0yOfwv/fFtLcbHiKvjYFgahsXpekRbm3lL0aoljDYfGXg0j67Y/J
CJh77b2zEDew+52ugEfOsJOLiiRpJwaOJF4CPdnGFr+y2s/iVHaTGQEUZijIRl8qTdOe32Iiq02f
mP6aA/zLN+yrK+T1T2VdR0v0N4rZ0JrKgq8LJ8s0nyhEoYbHdLwsd/ZM0u7jNcGRN3tz50VSRBLJ
ZurOPxU3vkWwEns7DOtGOqOqjnvGsm8xpTXRyN4dwUahlB3pl6We1goIcvF2Q5RgulgpDiLlxbfg
MhfQJZhd0vcYcyGscC4+SmhXhqUJfuRf0w9ZTw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 70192)
`protect data_block
qv8DX7tqszlAnrMMFQvAyjuEgPBHuTi1RS9pXGi1unSWEAcUzGPG/WVKdzHgqjKAr4iiVKlxHzJn
h8Uxlbrjn+yPwpUG1q4DV7dD+pBir0bwDUlYU4hNcnWZt1dZroU0hyvG2tTVvowG7er1i335kdAM
PjbFZs7EWvRnDRRHx10w+3OfT2mqX1VhIcqEuQlp1137UhpooiehRLpFMH7ZRgQkcKoYfaXEQqnQ
IUIXqzwshM8EyYFu7vhzl1dcgwuBz+zJe4xXjRIPP9p9zD97KGqUIWMtW/u06XQyn+DAXiIbYAdv
XPH/V+4cn/tM/L7n0Ruy5LdSgVYz3ETR+ap4RaoKiSQpBmJoz0pgsipPeX7eL9TvLzJgtPY5Niz+
8nt4dro50xmSfQMtGbi/bUVN+NWuzzkbmvFpQyxcU4pfVzKJBWQEQ4es9NxRaNZODhL7BApt+sUj
czkU7A2LmTxFvMiPFim5VCGFpYdUQJBlpII2ImAkiLermQhLeaHPwH1VBLHpVsxtxPvSBRj5Y9jO
vfOVbCifZHc3XQD3lc3bV/kEjZesUd4r3CH6oE+yNkwiudE3Z75ECvlQ2EGSJ4IvvgF2yw4hA53J
q6jNtwH0pfRSBcufz9ufnLkTLsY9qgu+l98leEH4Noovj8s04hWWzIPuvXsRdxh4UTh7nEfavqlY
QXRlge0hBwyvwDJEfzCVOn8dOP25B3XPE+0TNyIKLihcradJ8osDIWgzeL2oyjRHGfPnKw404eRS
fQbWGeZwuPbgfczaJzrf+v873pnVMpfXyG/z+TKaocSXUiEBcfrZuZyKkj0J7YihI33TZvqwzMUX
hXuqooGTfL7AQOzU4c01ykL+jWv3UsYIzz8xk9wXcSkFYg0SlTLdzexkb1Ypt9X29I1jRESw+M1J
KT9KIaCOkOF8pfXXRn4opxDfHzPGfULR52vhI8+zlzfz2SIfq13mb54DWslnpuZIe1wxuanmAOuw
fcmIaX6SusFhACmBKKFxr1PRBF2Ca5nUZ1wjxlSJFQAD+c3i4wa2MoHCP1pZ774TTJjBbXqJow5V
vreoe1Z1sgbxATUO1nQ7aTTBq51ls01rdfRy1hsLm6No8bLNmWbClpOf+gK0y6zR4nakbzHOLWru
q7Jv9X0B0ce1Zs8JqTlpOecN0wITXPAe/1/B5bRdGkGDRq/eVk4QrJI8Tn0W+L1uGvdnSHhekusI
n7CEo9hk4crKkMi53eVKWYCCdVdKNZHuCUXBokxxzOY9fgVeZKIYeHuMvOcQ0kviYtlLOzLUuxmR
cORyjkxsOhH2+3PFMh1VbFjOfMBdkE0j/67ExLxaeZ02t6L2lVR/nvLy40KN63zEAJ16PmE/BoTz
f6LbSRwbBKkBUypyPOABcN+42vvOfCVMtUv/FA0UqLOpHMPxG+iRl+BTRG+yiuLEI/hgTv7tmizV
UBLNa7VRY9rdJPIKHGhnFxxHN7L2CqGAuwFC2MPoycBgVbINDKlUZgWQyj9lwgYqfHygkDloWk3d
vKXE6IYI7Fnbz2m9gzzfGqnldHVsulU1KxW4EJJrhr4m+ZO3ci+6FePdx8fwgN8IBklvfk6Y1PT2
SYLrGF4jJhuW3AWmQqbvbtv8K/v5hE70yCl87GoudH2SIwz7tdnPmeiVYpfP1WEPEtUtb1/fZHbq
umg7we4eCW4YAmysVv9F7LqczqzwlR2nq6+PA4VbEPKoLaA9yXkMKigsoGJX92JYTzSGR35jML+K
wahZviu0eYtZgPsEW6fn9xVUjmvyeqmfMoHaD9C3hWdyaah5l+g4+HT30Rpr0c94NGaDvFZ1XQEo
8uuf+0Pi7EYgRC/XJ5a97O+Qv9g3udlHTFosjhaVhduZCsjeY9RUSkFRW7NZ77gptGZqnW2bCU4R
F6W08Rc01f5CyV6PXM+u8X/peNmhnqkN0JHsaTHJpu2tAD4PgcOzhI748SrJHqQqjd/uXZU9Rm+8
6YmaTDIok5CBVRHhh+fRVLR8igOUDbHytW6IaYhc6tc6CcyQu0r+JuVMvg4hTZ/AGcLAP1JR/DpI
OnWxPakZ1/dO6eF3kLz/+J7KOCn7HYzxvoW0uwDEvPgn726O17G8PQXYZm69kGtutGk99OXoqTnQ
uoshur4TIqz5CYrAyfe6ogV4pmw41x6hkyvEju1Y5B8EUTWnHZ5XmkHPFE0WOXVuCy2ZKAu/dn3J
Q6u6ZjW+RbLdpOA79PWVInmWHWgRK6LSsKzVCkBxcgjQOFAqrhhBbbHRddE6TCfFKRxq+vbDyy4P
iZ+dhhrIxL45Yhtxkzg7LcJRLWels0ALko/8S+HkVUkkVAlW/rVaeA8/H3TNyf9FVhjPxvThO97e
690xZJk44juOtiYybhm+rV+C1YYNCHRsGij9d8y3Zv7GPAuxou8oC98bt7zPOUeU5BvoBwaSVBOK
DhIvgr/6YoB1DaZ2VzsJGFL2yvcMPpXzjo3Y26v9xtIA2KS8Y1Mn5LXI0hNxO3dpKRIa3R6sTJrc
En4161UNxJzOvOyAHVRVA1RJEx5cXeFilNdj0VaIwprMZRsZDNS94lPrKzmiSu1QljIWMKWEk6DW
YsPcvGrmi0EKbMBfgPfYb5sARuMn8vFg0caLhz5kfpaZpcutCVOD6svxbkzPHoJ4iOg+HvpdUf+W
IRgJTmV36pNr6MX5OsLZRSjSIOCSSZToz+5aosRiQdN9FnkXRirVqnI3rwqMDuW6ra6InxSmdK6L
38uAocR9xHhHmHhmeb5+EqrYx0ClkYZumZb1A9thCjYCNKLEnSSmul6XwkEOu/8TjhvrMO+6Tkg1
U6mCxjbqdbXbtLhKnfpF8Wk1AFLLDBpPsZ9xHCzfsYGV0vq/C1keKbrNwULgUK2G9s5sf0KVqtzC
4OmkXK2+IZsalfXpGK70+uobN3HBM3Xb8FoF3ZLu3wwI1rIzJt/biYSd2nx0uLEMQRC1Y2hzz9kZ
Df6Z2bvh80IRUGTFrHGLLFwSGq5/iqWQbaxyyLoeLuuEPm3x2OdzTMTaH0f7fLjeSrdCIIAZzuP7
/YDza82g0+PA1fVvzs+Cod4YjIeXIOM0iIlvEwamWjf+Arnt0Ve4IfEm8rcp3r9+U2ldugZMayR+
CmBYLWV0VeZhORVSNr7gfgnJPWI3mEI3Gr0YqAGSUhBjhYxKflFWVRWxvwpCDXWPvEQ38BOU9q7b
feADo3ReahuGOKrHdyp11JoYl7BQdwSaq1is0SB6qNybvv58Cu+yFVDLMsI8T69WVG0yRics+2K7
f44nUZThSK2fbPqAHtLcwHlpooMygWo66fMMPXbjnvoO6FFpKlsZeBcG5BXkIAQGG9pOcNucko1C
qtun73E67yLuH3WqeBPyTZ65w/we7wxY2oRglWmnuMkxkOMx+dfPAB5rDBZarucamHmKRyicC/5r
fo6VX6MKPxxV5G7KVJApAGbpu313uEG0dzIgiJnKtd6yucun3mrNcvn+Kq4AhOoKqema9ux7Wl55
iDMQlm5EFJP/tIprau0QfaeSvGEMTLEiUFvzaM5eLy7j66QqTgmPyAfCyuRb9HFoF09JNIfH7nJN
j28EglvIwixYRjufkjSJ24MdbAKV3D54rQ2whcRQaZbrrrmyzYnnCfY+Z8Wt+vKeaL1glDGugAQX
CE+QbnEKrqbZRlrtIMn8iD7HnsDztHDAEJY1MZM9rXrjA+vlUWmsyMZ0ekZBVcRI+jgj+JCkF9FV
LfjOezdmdEyyzNsCq/YmerRPzRxNZht6zKBAKy/bJkToiqA1HWBMnMNYimquXZ49dMqWq7rn3oEK
AkfGwVDLEXYWb52umf1M82KFKqO1VG6e5CSiBmqYp/9lnTfZRuMQpqL5PUcsyIYZ+QsjystZOTQv
XMr+h0KVzMWPxUh+jizKjmTPAXgRNfywkvYP1ohkh+wOyTTRv15WBENWkarUHMTndS7waIo6trO6
Ud/KaBiGy2o06UvqFqIXmWhhNiDVdxSFiRoPhV/5wxLNNnEr7sufb+jpZRHFxmBcd5Bf2WSnAh9s
p4/z/GaDo+bHPl78nZDXQWEUp4qP4i9TPVW1qHMy7Q77VZB8meowo/LYGJtSbpcCd96NHhrWZh2F
rR5N5kGj35vAfQ8VObyO9ntKXme/RE+vvTrVn5ywVue+0jeplQ5YAR96RYBGFCbIy+pnh5RrWeCf
Q2yMOyw9HreV4eAEGK5KMNENKuSItNcYD5jbRIYy40PEZArNXedTtcXoqj/RliKD85rahr+KwH+3
Z8177wTleHXMhVkeD/uPHfgABdhsYtdeKewCQLzkupbozJ5US/BInf7r21H8pQ2X8YklS1sb5dDv
UiivCNwPdyfHLOw375Gs6VaKUNgDiRr8BI27CQhpJP6odfxn9DNTGyFfcKvsTvE0Kec67FAX0F1W
kpOiKXJgtK2d++1oJIr35VObu35/yFWyoLPbU7UvWZ8P2Uum6ZhujUZFTR1mK25XrwDZXviOrcfI
mMa40BHwoYC6gB1rPB636iB4dOvhDR8qtCFDEIodEDGLMzHFu2DZ/UIVG2AN5It8o6luXqrxv86T
bnN+F2oUq2+M75TIECsSfSloaASf0fz5HNvWww0mkYhEXwtqc2Nyr0NSCQ+cigSwcAfsElm/iIE8
YuTzLMGj36kaMKqvHNF73NIx2THSfKNGsY19BxZZYyW21SyLedKhmP11tqXz8Un21cIWOQ+wzoXS
a2fdJb9tNYUZ5g/febSs8L/8VYvpvREhaL6mNTxmSpQSki0Xr8JmeB6FTYSVzMIrawY5x+yWcT+A
djfCn/6yLqfogCq3jxvfMgauQKlqrEPGPPTpU9p5BSDCQOdl+GMbxF+FhQG6QiGVZWNZyefIOsO0
BtAz9h57dEl1kTXF2hDT7CzJdz7wcRDV/AZEae60HElg3ydM9KNJtLpg5YG0BdKRWOK49rMKcvm/
id8qvQa/jHv5Vvad1kbXT5uw1DS3U/dSyxNIjO92uXIf87VixJ3lbmDxn+vzHE2I/Q6o3XUQmB2v
me3L4tTzOJyPmakDA9JrO2dvN1VpUDvkVPiyivbWdblPbTgEg8X9a00wYseEj+ucKtt6F5xidprU
dlNTs9FKvrt3aMbjjSKVIV3SBauK3D6z6R+XO5u1fPjKgaAfZajsfdUoDr5V2oF5SC8AH+hJbVf4
WLjXE/oCRyhSKCiUfSa0BbWr02lPXD31OjqmXD06rf9QBj58i838xFyEMRNexaDEj4bYsS6o3w5P
Y/X1g/XqU9z2hqNS8OT2Cst9jiU7+wltDb7oxCNO3fyXkzV4cgtJplgSqCOVAgCqnHqTfhNhjxgL
gdjfOOKTBRWlxLesNmAnWPhgCADnG1wWQjUn3cWIIK4kROfEAsiOfb9M4v/++8OtIa2SPpMaP+B2
Y+tt3fVALgFC2LlkPOAMTHq8lgBdP2Sy0ZedigEWR0dooeMJTwHBgvaF0HydfwvxTYGyPXxugclI
oCKDljBWd0WMpIdcNZPhQ4lAJncet649qlFT5eIDVfRXL0x42A4bYgDUetRt44em1tiQNram+vot
UKu6OMM5WrauEtKj/JiB1QrGowreNyJgiBLpsPF17jB2zFyfa7rg7gnLSqZHPTTUmJUCCyGu8UMA
gQhALOFZ6BXuzTcon728E1uFQh0PwZX+v4oBy9iP87SYXDGEZXFfxoppEUSjTrDHwAZwwbF/JRMU
nC+Hv1LkKZPEcRIurV3nxS83WuOBkvQUhHWM27jSNfzGoRkgJGR9ATVJT0FRCQE+Ir2wp6saFEWy
FGn8vvEmPUz95zP35RRib0AiLN2QbgfWPQWXRBgNRRdgFIduR6ybL+axuR0tF1vnF0mk0zHzSjDF
TqrN8R3Xg4PSULdcqkvSRldOftiOReLNLkg7GjUE+ZTv3mvhTgKleotb5epgAv1w4fiWm4vwTiwA
kqDzA0leCha3fVsNZGjWmyRA10xng73QADPzLUS0wN/6UP/ONXIGKgmVOzmhFkaIY/KbkOk38l8r
pMPY2t9JO5vegVlWwpEYLHQDS09T6jNgpmPDRNLuyqRnOFOnZNaCP4GMN9N30Ipo4Z6+mqMEWEgk
ji7TNXrRyZcnwkYUW/IHFGcZ0LRIGI9QnHbZOS9Hgn6Km5EsksMkKfdlPnTC3WIOIuDA6vm4guza
upVrClGWFBT5TgrCZqggdHBd1T3xy0qa6cg38NHK6ddNBDKxvGubl0cBI+fMFwXkjHnNG4zUIrXe
bM8cd4VcLIA0aGiWN1Kf6UhiKkXR53+FfyFrN36kGUHbfHcL0sXT/DVccuNZZg5oBInjzdROKsrK
eldt7S8JFKUis1MRZG2oz1bL1Za9Im0YGP9Ysw3vp3k5/iJJ0TDy0NcrkbwuLf2TfG50NUKXb129
RFApJXDELmhrtO3TCO9gUcQ46pnEWn6hIEfL8g2rumy/CrdmDZvqHz7MrkvUYFVUJ7Ekxn9mxFLc
esPouePBQ5/2FlhLoG8o7R/URMIsAb8c9v2xYwzjhej9rrxQLhcKqOoKiOuhzpfG04WCW4JqS5/t
CG9aWSH0juyloYIrCJN63hIoivrpuDgMTBlqJHzmx1il0yqVJbDOSiwkC58MVAVdNT4VaAeHFHtW
4WRydsm6WLBaViJROzksFMhw7Cr/fSPVUmrCpZZETvf3XSkyyMi7g9InwCLFKPEd4DU218FLA1Hy
sOgedNUatDGceEPkd2CzLxAc86P5qTUxlJfLiitdxAtASYyppgbd+ODD93TfeHtVLf1elOr5qO3I
gbVYSZylGQqqD9QDDXEVzD8mHxBkfYJEmLOqkNvUMt5CvXt6CaSG8zhvM7YBjOESp2V2G7zpCzUV
bCc3Nw0b/0QyHvwPX5Og2FqLiMUddVkkR3ETDs9cW3BihkcDAwEOzY1hZRvNZeOWq86BK9Xodnrv
zAAYDiqXvXD9SlHxAb+rGQ9wIA+A2cy0e8HWk71SjX5PjM/8hJYacDhPrs7tZbiWXRTN6+lSYQvN
/97yXFf6/pqKP0fCNZdquL4SMgO1Q8paK0pRb/b/e5qX5WZcEq+5e5SFLX78oEcObd+FjuKBhQ+d
fRFrQ44/2hzpQ+aiLbEXhu8k3uZO3EL95bN2MLj7u2HyybdF+V0uZ3MnyJ4YybweovqCpW04R5bH
MGVs+7uyaHTbRnRhK97uxESR9Uyms7KDHkKBhKLDM7ibu9b6uFAuvGleCt8gFQAT8lBEk/6fkFYa
XN3vlz4DHRCF5agCLGvPVNskhBrYDK1bgaZgNtkEAqxMRwKvHvsescRiKkjDMRRoaxhQhRfZQoRu
R2jONlN50r8mu+1Mo6m+5yVOQnwD+ETWkHFRQiyJqj0cSqMHB9RRdhoN+KbFH7w+uiH7xRFGSsJj
voy0BZy4UlN+fuVjf0568erCsgua2rK8OwZVFFgZVbqqff0UynbVudfdl7RA+Y0AJPJGUH7GkiiZ
nsZF5rywEVAJr7aP/qpVkMnzdVNMzn0rIiokV9puU0Qn1OLamiCdVuQ189I+Bt9DyV/BgWTikoX8
3ztqk0Rm8d3Ia8g90E3jsdiz6qfWiiSRLjQLN2/IeNh9g//p683GfoI93Mu0I0GMJOVupRYgde3A
1lk3PZfX4q4JHvpXSEXfRuc97HHvZNwoL26g0384uZUJBP+s1PWCApOYqzx+8A3XLAZ4Lac0Ve2e
hICQGigqJnkLBbQywuc3dw/J9DIhgM+U6KKTTUxVRTmiNdjJ9MXsfRYO4jxHNgaM4m99D3hFl8Do
3ggQkryaOOOYuea9abt5DziS8OJUQdCvWmUk72B87qKcKaSGkAntLS/FOkoRsJIkvj2vwHW0HSaN
qCfOYKLugNOJroUkmEPPOAGraNyeiR88SKhs7KVNlqZTabZe2OHWZpHd/VkA9VD1TFj8U5ed2dX+
406mF2PHApW/sGi2ds5qMutBvxKBk+E9Xk4q0TbpLYoZ/TZYdoDPD6UwVIpE1xGWtUnLPxJBy1+T
8NTTqeZuoIc8kjjFmRoOWcDl5l+YpWR4TTg5kXfYmp5dNLg7nv+2uDmvyYhR142BHgVryMqX3ar8
VZecfaBgYOprfBI5L6Nv0OkkrWQYsgJagu5wOY6qpUyVrXdphJR7inLM63x7Co+bAEckz6kxnY5N
XyiIJkmDaRKatYu5yPIe383kVWmt2V2SQ3R34tQlKJk8SYiOLtLRZ0gd+ZDqOreu1gTU5f3CBH9A
jVJuyqeixzsh0qUT9kWqt587XyofYKBz5n/Y65GtsKL8RiuouHmxrAYmiGzxf2ulN3VckDwYxlTU
cmVYATye7WqBGgu81N3iJ7/S8VLMVIeHFngat6keWCLmQ4zEgsuF6CsUG65TILcLkkPDKH7trEUj
Or322UNBm4Ztfn0z3Ld+S9G4bt7FuvSYuCoLuweoaU9qwOp2tpkDqOC/38JCVtDombJT9DR4MY9i
T1o5X8i1U1zh6R29Y+U/2gykGyCf7rT4spHaV+ykejC7UTzPP2EXoW1lJsk1/wD4whAghB7xjYfn
xDihjonkVKOr6QiQhwHXFD6ZDGj7ZFAm5nvqCEQUO7PZ5taoAcMCJfiZJkXQVMqIJHjlcC7lbHbh
rvfGsd0WMjZFm+PKhSFEQOgqsJubsTDHWDdF0tC5yXTTchS9q0hboGuZjyVpNpkM6w1WakUPKK/M
GqBaF2U4jnd3t2glOS9PtGrLRqwq4fD/x2pxPxGFDuwbsjNXmIiJarlobFjLCiTNdlNkRJzXPNzo
ClrFmGggIvPJJoQtDZ950KM5YLJIR4+y7Eg7RCFEvQNig24/9szBdFWVhulC82LPQJoXdIVZg59R
wXTvn0yQ6sedmCMs4CcQ8Z3lcANS+mLo9XdRYoVmNrHc5GYtHUK6bt0vV4hN+bPDbvRTYV+yQCbS
PbwF0oG8oYje9qB7nWezSnNX+0bdNvtC5IBG3RDG9AdRqAIO4kKXMeSvQlR1ZFypnJzkOoWDbqVi
wTaZM6747cYG+wRA3CYp4u63tKbdO9fPkWuS6J+Me974gN5QUTxUsDKs4mBCoW0J6NjTh7JO57H8
6Guoj99uyo+k9BZg15c3AgurQLzIQVS83N1R3NnXkMKeVcxdP9epf6zTW9nE3xRbq0CJZRQwIwNE
ry5UGoYjQxWrAu7GDKPq+PXz7eCVgyxyxN7Recfh3DSDbmb7dSq5iKwBY5coPKnNIi73qiePT3Y1
5G2sTVobPdcU8xOGPhxR8ROzs5HHurcJkGrqaA6ftK1RZwuE95dSebK6GggIwuyN2RWewZifIS88
PUdTW4IKCZreYoManDhK28jXrfhxgdbCZ+HMc9bcKNynIYJTF2z15sFQh47kDFAxpLRUGGoZ4oVq
+2496oY4yOxhm0uL3E7/2OfoJ4pIityl9PSBjH/yna8efxqqBxs1fyp933AuSspo8IdmF2TnQnjS
kzaVLpBDBiLKiNP2GWgaKM8B8A2y26zvXTc9VN7sA6bGeGpi3U84enyIBiOHuawnUuqj//S3m68e
U07Pm6wvikeO7TMoHUrBzuUSOKH9cY1G+zuaFq5SEXsMKqV3O/KIRrIZlDG0uDyT4UQYyOIzHbUB
9u+ZPiVxxvB0nPZimP8mpmEZHINH+NTjezpdOjZraVsos2Lt/+eAabvfo57GewJf8nJ2yl2NcxDp
Tr6wOoreKpcS6QOzPad9b5il2ahpBHOaEY3t6S63gvDqnXlwbSbXWXLZ2mIFXxaMeyNMYCn+K9RN
/7aYc7WdlnLRUYV7zZAIq7sIOVVThlou/VoUx3lbH+PIT59SsFWLW6Z6lZL0i8uvGGDpibK9gra3
82bgPSA5VFnk/5Gg7gzHOvCiYswa9rGymgP8Fga8MBuM+CiTcwIhSLxLPGilXqiK5uo305eLXz1t
i8rSyF4lVX1sPTl+tds/aHJiaoyu5bXbTsxsFRCwV93m+iv7BSnXBh8UTiI1tvFSij3K7af2sjYX
4jYKHHlTk5aPqRYXHs2nAVTEP/oqvydbn3pyLN8NTfM0rmp3g44nTmdTI+uEjNCnbM5qkRNSNUqh
laNBChHkfyjNoq2uhAAp1iWrbkHsRigDWynW9tUsiYdpzNx/sKAIim+pPl1NjLHMAeDETQRL4B72
TrNDAZaFzDQXoCSGEpTAhFis3/ML8TN0ciZAQXrC/bpu1k+9fyxeroRzNRmQOMzy8zxZSwTJaRLg
DYXwIA8jozdImI48gl9n5S9JLugjvAXhEmPZkNLVFW+te58S0M6dzOqdcsqkPAnC+rHiqJTq2z3J
mCUiVdHwOWIRe/Ncv6QW8EAkkvcyJ416b9EuKRLN6nnbKP3sSOTSvYVRovDAnH4+IPAXj5/uYH1t
ZqQHAQkaCXdN3oAWxRH6hmJCBa7VDZn6mEz3ArzXY5BKavGQrs9s5d/9yGoNUzXkLadRgo2vh6y7
gaJ78TeSU5V1CkUvTTNO9z4VSpDCQV/USL70OTDkVR9EYTWY428KfuUGqGx5L1bVeScIixfwOTyi
WrkPsj6HpHN9bXGtKPWrkdkcjaI6txStalUvrJ7Fh0sxmbyaY8bfqphfbttblLmqfsZ2ABHtGALb
VWIN9RbVkzH7utRdocPvnE5JkAdhL2Giicgg5yWxg51Wz9J3sYZUyUd+gQYMRyM1EZS3cx6bbEhq
3rjI3Ku3fF4F0XQy8XLZyfc0RvN3dsp6FZnfRxOgnv2bm1mwwYlWxqSufQeVzNSmB2pX38z2vzKl
VEUhqEZdBMKYCgcDGDOwwOEceANsNyypxEEJaFlThFQR3b9GFNqYd9Qk1fCebYuG+zhQv3vG4skk
A4CsxCSnQ8IyLi+gEgHABocgP9zItptuZcVKlgfYtHcNC2D9j0ktnKpiLiScZGEHU/wyf2q6PtXm
FOnxoZgB9m7c/qeP8X0heHAg0zNFSl/nrBWC1K8hm1FdCEtBjT/BTY2hhOcR0yUqrxr7DFxvJfNY
DiZjiJ+tJAmSupaKOLfXMxhrf1ULhPMzEycZaA74hYSK55DjcF6wZeO7PpzF+a3IbkZPAVTrHVcQ
3JLWbgeW4TctGs185jtdT9mfM8hEDJfbuWyUWH0fwci5J9FxXVSe/4Bi022ia+x0A5xxguImiR+5
LcGE6f8rB+i0QIWP5JrbDVzyEVEWgHLjq4ij2WmGWCMbRpm6zSk1Mddx+xU3XBR9c03iBRMkTFMp
90fGJ55EeBu38wxyN8rvuRRgxZGOWZS8q+JddacoLTcE+W50gRGOTC6GuJAjVxL1HJ/a8MC5qY1D
7EURRkqj2BU3f4puCrVcNk39b9Y/dLekhU7gmp8LMLAUMsejiQVR30G8+se0kF7YRiafpAGCMBVG
wtn8iETqoyZ5/2Mlv6ZwO07BxG8ymCdaahN9b/Z6+QfNOYTtk5C3qdqLAsxCr7LYOxPEaNTsUS47
NBEHGaRyT/KF9yHuq7a7egKrC5KmCYgFhP4CwHwV5idda+Jgsn+Rngvh6DWmqvqr26FhQs6zL8Y3
WymBsR41EfnaINbSnH6KP47IWROGFs6Z9ibTCsnr0G6HW0ENCEjP1VzEU9FCR4GAqUgJ8M5ldOxL
UuL1oJuPS5ijHR+NpQXFNTykilHJ/OLkzQrIs7+vlv+gceDHj423xamKo/ZWpOTPEa0TUzj4Jy+a
R5P6NlwiIq0ZRdz9Nb70QABGFlw6Hmt0OJNYVuZhUuEb+5fVQb5yLlokRyJJpXfuDZOQ2A62sUUo
4hhGqBkxocw31mBtz6iZsQ9LJSUeHQkcE7UUs0rnKRao6Q40mBD12y4FD62N2DgEt4rvE/429fyh
5W2tQQzS0GB0OVBNOwxvc+cLCsMuJlE2Fw4hI7TJsC74VqoSCsfQmE+OZO8+Y0wEPPeYtvHjtu97
MO75CHOkYcihkPQ5amb2GC4ipdqsX3CWTyRUcIwibxF8nzWmUarQaHoFGLvEpT3ULPtq5U3JY9WE
R6Mqbs952RKkZLbbd4ybAH2JRYzU/GCCloX99SCSc5Rbou+XuyytSkTH3WVlZ1AiWDL/osrc2hV3
6VU6gb8H3MNwpkd/yX4rEv/3qtdKZCKnfzI0QKdVEmef1AyMP0we4+QMSJOC67zfIOdh2bvq8Z+S
TGfr+vYtoqbewy9gnD7+ECnsOjZiXCB61ZnFAdMoXzmhr31EWZb9ediiTC5Ff739vA/cB6nnRPqL
XPnVEbdhP73pxfPLG/BC6c2u8p6MY0EAW0QbM+eIYxjxtpbECrPCCBOoXBsbP/dNLBK9ryItabMb
NRT5tlLHcRa1iT/tnpEwtLyf1u72yVmHvjWAg7m8+H90fW4ZQM5SMKWZD/D+dVLur6kkUiuIDW0W
G7UUGYKO15ZmmVjLblVG2WrB0XW3tHu5iqPbUGRqutGJfbbHgyKKU74XsBPHvITOCWEN7aCH2VsC
Hhmeoo/GKTfwp4OGP4fZatyD0t0eBI8Imz81m1mYul/sNx8Kn6wpIhx9LEIydPOMS71xPXwolpVb
neHJzcqsqqR5U1XYltdnusnlM2CiSQMK1f8g26Zb3uaHzMEy2YOwL6Gko29zDFvGyUjyNyrAY5xZ
POAId9lO74PaA1+wQIFCtODa3D2YqZuKbyDGen+OBjriL74X1A7NqQhIJms9FW4SbgJnxpWOqNio
R5KkbR/kPZzYqiIi4JM6axgU8QqfyejvNbr5tZh/no0ZHXaLzJlL6YUMy9HUjfBylYbJILGPycGM
GSG0fJvzNQZYGCsyex5HE8iPUROvaD4Jp3nlcymTYN99tKgsm9jfZV2DOXiCCOCT2Ldc9wFqKwTh
nPvtYYwMvwyTApB0y/KVyje7mf5RxPHM73AePsW7GyV+3Gd7MQJFa2uDjWLL5RoRWYCgBNyr7+/x
7hSrVggrkO6vZ5/nLi3pY4JUsGviuHZPaJzfwBD8K0tFKFLPB9JGn+mLwKoP216KuRH5mcrPmkNA
GPc/A6l49MMJ4+nwTNY+K5r9A2t49BlNXWsghl395Rgd6WOk5Q8h5/wzIN2OruY3xUyLkIEog3dh
uMhoIGBCCl2N/meK/EvCvsKEeTqQ4Yfzbdt+vYpR06bMTi2E2+D5tRT6rTb85EKdMP2detihcymR
l1lCUBCJ4CInHQ7q7dElsU7u0uzZJXkxsoehCOwDFMpKkU+2B7Pg6bsU+ihqr+FAlMc793r7fqtm
hTQVr9YxATyqCfysAEvQlxXiyKUDgld6kzY7XOfYfqVUEVz640E4kKQdiEUtv+F595BPpq/oxCNt
ojeAPCvia0CmAhI5Xn9TwSxM8um6DbXXoorTUhScaT0nGPq9s+6FZN4mcRvJ8Owro3X49o2VtWb0
t3ipNCTldM/+eCm96IJQQsPmkyJexDixKfMWeBGJyGCUGUaZVB6v3yNi6UXSEoQKfUUeFAh4St/j
Br5lpBptjthb5iDGe1/K2rrcdSdKElyFpKJBOkwb2lbJ2Jp9t95pgwPZc4gsTdp4zdhlFD3E5bk2
fCV45n5tl074n0J880o1VtC5IQ4VBq07j6vUlyU0mTJxXoNVByWSyk7LAkwMI7Ac4fZGcV6qRY1C
1y/Z8nIIfT/NwCQIbJxkg0nkgx+oyXplhQtwDAqLtCxBcppp4XEJLh27C1SCHpFGH4V1SNrFbMu2
AJyVjaD4EIWbgrae6P81CDdoeteBg9npc7GVtAHVlrKIgN8WI5UmjbEl27tBo+m/FdmZGqZxVR8L
ZbA9Wa9sEYljd2/BTKpoTohfLWqvKaOnmRkZCuuq+jvrA9SvP3PKik1xhZYr1KgTz1P/kTROqZW9
ykWcVfr/xlJy49SPZG1XKYqomKY7CV2969E4BDXYEMeo5BTN69nvIzXHSv4RjsqnKgcKybIb/fXg
4RAy8Xf0qPWwZ9wfyPtAcxVJSTpk3GueBZRohYpyNXeE78Vz1uONaMIO5fnaeKXKjOhbMxs/a13V
5WndvrfyS4SK/gbCFcISvsrsyePz653zQA7HVl05dv6Paek5v3OFmEPfDdYLWaNGSJPz0lSBnH6A
nWtHZ08Eij+VNRxOwiUCX3mzxbMhDDgvNWSI6W/nBGLKplDitdjjGqllfDjOf9z0n4BRHbvR80n5
GNd3vtCct3FG5EZT+F6aohk7cTz2so33VFwHJUZIPITNlYfuTvn26RPQDkggqsZrEXaZQ9Ri/xOG
B6GP+e7XcPGLxLJKGYoL/X1eVdQxc5ztgSBd9SdjWq0Xp+MoeOtrPqEpwAiNfgnlJMGebskCG+CU
TMq5dRvlNIthMnPseAhGt59WMgdy+Vkd0dEQNA/kZxaX3xQOe8600z871+0QxPnPclVbqguDh27n
rCBjpJQTHNO4IoshYKKzuS6aO6OAt8+GEe4H1YG6bahnQUJAAGc5eCBEHG//NOcnv71/W7dW0w5o
r5umX15WEKafoKPecpeu+NoRPL0Vo8uUSNq3CGJRrLL9PltMlxcsGipMdI4uM1/k8phh7M0Nz5GF
1GcHe19PRJI6k0TBtFCMEuy2k8bR1IKWUOIdsNdtPKyVDoYx/JLfWrZnyUw0pGRf18iMyu0QTKVX
nbWYdlxfGnK26G2X3g3jY0NCL1RXKLQZdZZi6hf5mz8Pjfhpybrd48cBnSDv7R4AkP/wqTqj+4+l
X9jM9A/TJj1Hllfl1kC+ebwEjuqBsbqxGNovCblUpnHgSBB3PrBWjRxQyBjK0LXpCkoZNTE2WvXf
74brT+u2wcUG0f88ErRGYIAAVSIB4tL+XmCITUuMzV9qMte0qCua7JADmhA2Z8LMdfPQDl6yPvsx
lS0nfHU/rsCds1/yPwZvz31T5E9z3H5p6Jqo2ZWr7mUqqHwQrSHXtwRJedVDy1TgXUm4fkxWjLeg
M8/Ky+kWoT3HvWOsQGBVGYhxH+HtRzflEayIvfk5TCfBvzSoK/hg3PetFabUUWxvhgHp3Tgw0dyE
dqf9MaXwejy+/VrbVQhPxfcBP6ZLQ7E4QskGGmoH+c6e4ooWjxL4HCRM9w8Wqp4RNnVX+IJKdkJb
zBHbNCpa2CjGUnoiagQnzG51IXUsVPlxXnXVQYRFyhTwAwXpAIfR/cG+GHRSHDzohZunLc25kQVE
c9AszhFx015ZI3zIBejRiinQlFP9Vlw8+eOJA3sRLm8fBA7vHv1iq6sJzgfqVj/GY4+xGfg8168U
f72Yq36ssN2Hx17rt9yelArEeotihT1x3VIAG6OSMEaUsQ8VcjD0qFTCtCBYD8WGDAXYWgxQZ07J
k0hZAkr4LlVFW/sbp6BKdn9dZHPZXbv6tAb3wNld2SlE1ZJ6CHEgxsBt8a1nP0NdCnqx28Yf5aPm
3l4RkYHX6mG4ANbfqjBcFMLe1ZGxyPCZtxUd19bS5iffogaAvsdeSvYpMvcEjqRsM4XxXvrGMj2M
kt9PgVsXH2Bx93EamrVcjXJBXNcLmPeMU3+82mvSGsg20mIeZkJGps/n5XnwFHdFl4uRrsOkJfnP
esehPLEX7jzYA2KvANDRDF7c/Va/pl7wKiJkVJyMEK/O/6/TWIzLRpNkPb/ce848YheUxm/bzRAL
8o+eT+3ssPXvnCtQhwM4Yijrf+B9k53ZrpEPQ1rX5GVCkMNRoB0HfYx4Z8Mh9P/xAE9TPQhR5S6+
NDxRE8cmNM4UibioX/jDW+fLQnAr1xkBJr1T+LSod3IafxhrWX1s6fBvL6WkTn15CLlI5kCKhaaf
QckNw9m7ZoA2bStVgbO1b7WCKTg4PByJ/PHdIFLMxWHnt4M8IYP0N/XaspJmCcE+rAlyRa20BjbA
L2TvfCBL2+6HLBUl8HxfyYqhfOb6ERY/mxY5oFBe3QWVL8hjoBmWw/esSHV2hnTVPEgyR0Inhhvs
18NffxMmOC/GFRevAlOTFOiIoRuK5Na4AbEEqFpXnOD6HnIIbkp8vnCtJz6kJTwLxNV1AB0ZF35b
k2hEsad8U0uLMzts4W6HTUiYF2M8487klMa5VcONNLKgaSsaoY5fIp/5LEwlKeb6CxeIdJLnR6wo
IImwWLysSv7K9lomlrNEA23TQ3v0R2GDRBSzqAbH16COgIOCr2wUWrPcHfY7GzhJFJzY5/FuNrZN
etzbVVDAHOplpKib9eXwI3GJO3bT8QBS6/Ii/Ypsg92ul69FbUer7qC0wceEwcglKsbfwk/rj04J
mx/l/n4tTDC1yprEp4u+3V97yGzoLZ91E/UoGDm6ZWH+s3a6AIyyksV2oszpv+obOaTM0TqpMsQq
f0aVP+bmH4q2aBVazo2bldmQxOZkPAsRDdT1I0vEpnymofRIKXuNkav4DbkEl87anOWXAUs+BNPq
ZFgA3iDAV/lMEMJipPzqoKxQEwjAWbD1vhCNj8DM/ixvSPtWKjQW7jAPa9K7PcMTD0cVcL4GzFis
ouczRXZR6600UiruGIX48kasI7fMAPKi/S5MW8A2rsDIwAB9ikMR/4MxQkJjNSeWtRzjxSQphWJC
eij5aUruokAzalRo76Cfv36k5Fg2rs7VP4bPA22kUqSHH/t8ZqWQo9Wie2sdVgrRNxXfT6ME+3L2
vvWahefFa5vUyHcxH7nuoJ9i0uSoe0kA3qedfsYv7caYsdNvA35INQGyjM4UH44M7ullD33WCYT4
Spck6KkGWNkVCJIbjKQWVFdx3uhJCuQZgtHgLZKo0A38vEEnLEFwlAMhrghT1tETgrwjcxE2Bn16
Zk6peMRSokkWwEuznUtxKMtCYPQ4EOL5D/62Ii6KX8UPvYf6B8zr6x3sVJueQwUDGF64nvCGBPlu
cphLo73QGFR0JBhkfQ37BpiwLHBujP8Nm5RbRyO3BGCSzOJvgnL70Y1tOHwZrrryTHPAK9UrYfQh
nbOm7WOQWG5a0zrBkYuP6RSXS5X41tl0bY9I9utVq1R/xydn8vp4AyntsjhWG2oiWqtCs83rGIuW
7ErWYQOY85so0iDxvUElCEYxTPcFdj76mKjR2a5cw1fNPMCSKyQnpaPvgh/Dp6MfCRTKluETfEhP
hsVNTbiYpJgdwi+VaaIw//OkwqRMrY+bKI+edg5WJtE2Gm4WiKFFOye3QfS8V/nVNouLKtkLUtvh
lwYwcAKjr3Gg3Z1d4vsCkQni05gkDDx432bitTuzSZcpcT89ezufpg0bixPaOvaXRJ+1lcwpi5Pi
JojZYJyt6IHYq9UNja5VfaV6JQdVK4Jig/xiYJO7PcwECSz0PzXGKqbpg/K+3nouMpj575jXO26d
y+rSSL6AaZGKHWeVzogSXWpkC+qUHkaOvt8ygU5iJmhtuNSyUV6jhyOSEiMEj4D/lFXDcteibSZj
TgJLWkUQmjvcX9ikZA3Tb8svg6vnbxGt7Qvsz1Yfx9tBdwjDqkHSvQAEgKiC9GPq4SxmKw7LM0Rg
TBQYodMM58r6M0lJYeKgGwcTk9olff1qnd68Ffm3YhCw7at7jWMHq1z+wlE8/86f02giQ/PcTjxJ
no2612IgkpvbSeB0vzZCExiJjXKGA24j+nQxiGgyCBLIBHT0nGtdLeFCDwl+1m+1XvdwHxqdXjfw
3hy7leSVOevVqbn8YFdOTCdJj9r9XnmpRIqOyDjAM9lfoW9K04zs2TJnfQBZ/yg+IAKB/WB1gRmo
HcerJvNkIlgriiFKKOzobjvC9MOzCF4n6atvA2W4D5SPPnyx6e5mUBr5qLctvDHE498/pt7eNFNm
2Ot3K1Yurlgl+kW7/On04jsMYuok/nP4kkV3vJbhGCy1D05CJ00PVEHAg0WqHCaiD0OfzOtNyKWQ
r3P0TNdmc0u3bGaR4GweL1zRL54niymt10CGAWKMXuTGXHV2kWHQYXjRglRs8BjT8lO2NzxEJ2GV
3E0COVp07LDReJy9zYc3gc4by0oMKDnQ5x0OabuRRQI2BB9nh/Aj7++LSHsQ+m0V8j9sylKSXsh/
NEfDqRLW3nHwT6BQyV9yHPlIlbBq02OWkRlbtJShP+DxVYfWMcu+APd+Ojh8lA7Lc/AFo4dlz8J2
oCscXzkfwDp7U1z5U2jDrMVlvt6V+rKaNv6Mvjc8zVV2d4E8admWSNC5RPZdRH0VrPnQEA0WZ5Qa
YbUsLIofLqOuTp+5bIlVcdcRBFjkB3pU9rNEj+7wpjKwSxjbMY6dXSzGNlFlrevu+WiEmIwI6KaD
PcuKxdV0BXNJCYea91LPJm8vl+a7tl6pKFIHUaCn8Hf7gDmeJlovzeZB/Gb2icm8j+MU292QbEZa
ABL/LZBmyJzEi4xbCTvvvACy13HbCekHeeHg5TsKEe1a6F1108VqnV34G3z5/0LuCyEPJqMoArkB
Tk0fJteOy3R5N71Y/uU/O6KOJ7awpa7teTDWD/I5kosPACk0d9spk8w1cHAAlZCHHz3HF/WXF0OF
lSzG0YIFyG/EkoyVIMB+IXDpxkFfuTeqsGrSuA7Lj5dygNoNuwaEe9epg5ARFXURONFrMr8yUSHo
MgjFtWlYqnYL0gZK3G2iLvSW/2WDRvlTlCT2fh9zmw7mAlHw5sO2tJdM7baqHm3kyb3YTFwymSBO
D/QckjSSPDu+92BimJOoD9lMsnDICP13/xLuwFdvk6ksOwFlw3XyjXv8pz2ul7ZV7yFlkkQCUAyv
+jnHU32QZyc02ViXTAztFREusCt2pfaRYbV/cUehl7rbPd/DuQ7nnRxMk3mzigWdQ3piioSFYOan
CVHlTm7ynH17/CGvIYaDBncN0pJ4bIxuZC3naY5kYr+tAPXG8xNb1vCDLrlW4dKrTcZwi6bNNYUV
T4+NfJLDrXLpI2O/ZFceQfAUzaQxCYxNR752u5GwLELWB5xdx8xi/di2JY7fjpcXno7XUQG0xb1e
VfU6ELFdEdsBzctBw//+wOnB5BndfHPZmKtiKP7iUl5bWTA2lrhTeiOYqp3RXCKEr7ADI3yDjMNj
2Uu14j8OQ5K1Pik0ppVd/jDW+TkpqKGiECgMStgdABiMfPB3CPhzGdy/OBqFsDhRu6D9i+HiN73Z
uIwR/RzG3kwDSWM64hRE3y4wEH2dkNsOoLNwI14zKMlx5IbL1DfYL4mFpbBu3urWXchAL2y7/RxL
hVO39A8AOADhrN+DcXM8TGnSdo/JSkvEEO83ZuJ7nNWJakjj+nDHi16bt7754y4q53tRxfNK7PDL
TJzLsHjO9+UvlsDy1BnnqtmYB8cvWWHZXdQDK4zP+YGvZFOAz5T65zesDzNpJlZzRDc0SVBxXsAD
nMPZpkbQRiyUIY/vExVQmYf+3UemrEp9sEMjRRRDJjyML46HQBMYgJpmU8i4rkx2pNhO/vufxQL7
0zyS2PKn9UiLYyMN/tyKbwjQqgx103RuXo+26MtIboGcFQjzMOITMyQ/6e0VElyc72dehtTAqNsh
aRf2ICj4RM1aECyB+sbqBvfVRhzI9FXuT7Ihqy3Wqxy8CYWbSPtCox+q+MOS3OCB73W8bUUM0Wtw
CCMM0SmfHDcUWB0YpOwYBMpOT6nn25hiVNbWsOjrlddNoRNRDYdQEt5KIKvJg35RPKBu+ZHG6aGG
xmOwlg47QhskdQY3hyPW8B5zMx2hhL+zRkZGmET+LQCE0hlsbO2Y3WKm32ThrqOQw6jTbMSOATBK
GzYXYTy7rjc1lvgcbwKbFm7weTknAHo4DGBkG93euMDbiXIEXfo204895kTykJlXJTJP0qAiKtdE
5RpQvbbdvbYrzAr+aUD4AADq1OYImGlpk1lN+ZhBvf817qdHll95hLk33eeCnrM6ggmXOeZxW5hZ
QUW8/7YaLR0Rz9pugG0SS8MmI5pHk+KLBrZx9z7LujLc9qwwbQx1d4PBraVsmkPLXFOAAZFxdpHk
ANSE9mKA+NDNUlYbMnrQpqYfKOgG3w78Kz/7ZKL52YIsNWK0P379aBBs0eNkxLM94IFbe6vFdJJR
BbReQdBLBAJiT6STgkrQ2PHXRLyvvH4S6QV3Ykb9IOftaRiBsZCTScYvLv7SIpeCc4LlMQT8Ij1V
tPh8KxR7iZpW6F2kLI95ukEEpsSGvbZjTikig0xm1fHYILdMI0D+V9+0+JkH7yHlBjXbLc9PG9R8
wrRDoPOhlmIyV09jbeeyS2y9asuNmqzW6EzUPnRztzMqBEaTtRD1GVfrORNkTEbYWaQPpb4ab8Dm
ublzDy4F2I5SQAVd6TgPWRe66hNVXAzwoQGOGLx4XBPCF9RS1m1q7lWNcXDfnxeD9X5DFglIpdTM
27KmecfW+eHaSx/sx+j4o2Map/hpJyGsiwqL2FL1psqygLVBpfN5g5ZbmHjAtOmvx+Xz/TP4Au0k
oo9KhHkiUKGq5dsyWuc6mSQU1kMP/f0Pp8GrBpXHGYdsn9LwEovXLC59bgDTLcrEcij/weFyFEpJ
vVExP6h6qmTK22PrNs+jpT4ewzsKeM6jZMXRglJ1apqPNQjVtZ0M7yrp6RePl+aav9eWTRqNjmnX
Xnx44pkP1utqeQwnQfsw4pN0Ci+QXokWLwBOw+fx7/4zgAshiQkBHFvd408+0TwQaVXjrc4bn4Mb
SAbSYS0icPMYlSRQjMF2KERilc4xCcUaxnKvA2K663UkSD4RMEoSP7V98Q3ORr0zNrqoW9vLKJsg
aIA4aXRTgF+KtwxviSt1S84sKBS+UyNwvNBEXM6LrtXKmwpjrWcGX8lmC7fSrnHqTLe5gK2I4Vt7
rdKcROIP/7eDRsks0gQ5DDxn5OeBHofbKUnme7JZREYjhfo0EMcFrkjQySv477FbvqO+Bgp85fsB
x3FlWYhSBDTcFtFxo0vfC4veAj85SmGg1S2HiyAXpcPjdeWtRcDwo480b6HHsS51ljVs2MbOoIjR
FnSvVqF7XIvWMvV9hUH0JDfQvObxT7m/ryYxLvLGbIuU/1LuFYM6pUoOJQx6Q+woAUIjYn6HOojs
SWmgD3L+5zUaQA05hUkejTUqJUA8yDni7lbaa2jMdprC0Le7+5Lk9gcmTw0NY2Ru950Y67z+V0rX
N524PohJ9qEMM9z6ibQ3DLPxUia0Ftiee0bxJ5ek2s6fvkJgezbqFQenfhcW+7fztgN7yri14csa
Qc2gy0jZSHJPEU/eL6D4sTtQ1H9ItqGT7UpTK/aMFHTfI3MM1Vle7WtZ/TN+5Hzy3NnRw2nlGSOx
NY3D4cwCTAP6kbsNwS6mjMDGDeDh8E19yPN3TYN/XdIgUZ4LS2xY8vtBFbqlptw7TxJbNVAA+Wpo
q6+WOE2PLGlkZr2wuhJX0dX/aFZT736iWawrPA6J6J0Lh+V3piG1OAaLO3rAlsjPdhwAh9iMvsNl
i0SzGs+NQ8KGpxiA9x0r8Ejk5bccLFIXu7PfmGxacMwCPERDnx9vX9YwQj3yUNSLwFg2SmNO3AnS
I7cRNjbGcJ50j2pppUr+kpfdy62GjjO6EbrG3rH+6gJZNFntGZXPYYu6662PCcauQEvZAoZaD0nl
ASb5UvaIfqcMCXHOnqb96xQjbgL33Tep7Y7z1kUcA6+jPruuwOXgo34X9cIiDXLLxfge7tyjaG3j
6H+2ozqwmPzEs5bqJ7G4qGrbngGbA9FPt18Tvcs8UYmdaRGIW6HBvkhqqsGTQlQo4mEo8PzAqKse
mHO7e1PW8kxFw1JHmcebgsbL/qDT3xsa41SW9k6odnDc7NSTfM/ctX9ItnXbQnah/PO6JI8sb+fl
p738M1aILDmSL9n7CGeZDETqP8Mfz7U+04Z5k5OoamLLiCUKYAgDA9cmc0aT1jjpGRIrUiylW1K2
/0UkZ5Sv2SI9BDtGJtKn73EykvbYZ7cGK1bZPUNlECH0dNd7vnN/azqTeAadjrnvvszyoXIqU2vv
pVjOBH7y3sHgr9w8WhsfjbzMUtXDURhN2jUKrJ/yxCn/VfxJNeY8uu+SsuNQnVbjMhUmmC/Rbq5v
OcZR9/5d00nHd4C6l8ZpT4dnIDt1P6YRj0MSz93QdKa2HEOkobmaHtwtnisGdGKSBBf+KtLFT9v/
bnbWxEbAyJqBURLJnA82P7hId6OEzZ6fI5RMjvoNqJDu4zad7JeRGNSL5ihIz0JjAB8ZxgKq3Epn
Gk+q4WBVj1HH8pEg7eLC3iiAP2I6CtCMtBej2pWOyWAan9GEWURSHSD9PFrMbl2sN9h4FEjD1nIR
4T9ExpOAgOIsbAjyT+yO+d7eN2zFX/4tNoibWSAYXTMl9QybASpbuLBCtBb7/4c6Hhxd1COIBcQN
J6FGN1h+DtcIfz7IaAJRCHLA9s/q0UJitSr+2f6ao+pwmpdzZcHulIGc38vGUyrBkLKyC7UBw3Nc
Zr1q/mmXN9IU79asS+ESjvTjHKs32p8j92hbJr7BBAII13N+nJJ/JD7+tHIBzUlIEanqcwbJvGxE
6sItbytM/o5KnpnsmcHNEgQZEinl6GOmrBrswBB+zkreWd7Be9Q8M69tM0F4IqdGdTIii50J1FQZ
LP9kzOiM9bBNt+SmDabXezUV9bKzxhZC59gEVtXcI5hXCF8m46+hMwfO3i32oNEfy+Ql8VNVQz4P
/GLF6wbMqQBgtXsCaRTMJQGQ3wkBNnMceQiGe1/YklvtFGDB+Xwk+H4oqkH5KkMjma+FQYkCKL5E
9R80AAXWz3KQYj64AwoQetmqj7SgTiDlJKOS1x/FKQY8q5EWT1IM0RiKPNOWMA8Sxo95QNEPXNTw
AAscYHB0+Z5L9wNMT3gb5BRCw1XxrgiRUY+gAtmvxpChS7GQZYFcswvCO8W8R5e5xXbumPlso6Ey
mI3y/n/yeo6t0Wn9isfISi32ft/bh4S8gyRqaPL01EG2qvIcvmPnnNvQF1FUEVhne86Qkh3zGgBL
BgDBWWfTon32Qq4CyEDgQ6HO4n6mX8u4IkMgXt2KP7Eh033f15ApKrY4emw/meUJjx+6wBYRiRme
pqvJ66SrJ+kyFlbbw4Kr6fAuaWOxkH16zjR+WB27hPdpQHhA37ZAtIIM6gprmWqKHQrwK+Jog+fH
D+WqEtNrvYwfU+5xO/p1eZvS2SvvCDpvfM9PF+xUrTHK60KaWo+FP/Ok/2wBxIR49zmrWxCeEgA+
738vSbn8ZScTtKmYa4txHl6P0WC54/sy03X9AEt95IkK6qrVDSOtr8FPhAgqT5v5PneYIyilhXvJ
ryTYC/DJcOK4+S8njaZ1uJUGt7HYFshU3I5pee8BhIds+H1iGSTzbfUZgUCf/SC9uDTQx5U20wVA
HJ+eQYodQ7VMesQjpcmxCypz73x5oMTxCvsoIv6KtYCsmsZ2JuCadVP4GK9/OPfTuh2zDUMt4srh
P5CD02vNn8F8J4xMVKhnAACGCbSdiH+E3JZJEpszY9Hp985uyZI5tN/Tl0C5AQp91zz+jp3opPLo
FTjbuadzDJjWXlZG8t8h4eKztIxotzrJRDDtw8emMPgR+ByxbzCQ8yGznZbY9TZmV+YpSbgINngv
fRT5NpWW81KO5yirWIv3PqkU4/6VXug2Qv5i2wMSLPQPWzwDZS8kC1gvl/RCqRGi/J1qGflXdml/
AKysA4RBL4TFM5XcAtRmxJjpo5/PglYumXxXZMaRBaf3t3wWeBKE/p4kdxWNEEA34bDk/MsdSGyc
q8HOUMCxG8shUfWVzNVJYyUfe7LehOZ7T/157NFNEmyx2fGT7gnaYpiVBGg3XikYaHy/ixjkWMUW
lytJKTLWIgm4Hi0X8dOGyp2xojiF9MfcRb6kD5qfj4qCMKzN3xACNLFikUmEVTICLjM71icBH7oP
tNbeCYdp+7liqQrG+7M5TwMTkEKA2yY1bVZ/5LfXoBSVR0juTrKotLX/d++FUiESndBVzQ6vBCau
auS5zAO6j6T1Z8d0KadNFgblrabZegXHI4w/Z13dfyjbuMYP3VoninhK95KGsgaE3uWOl+jx3x//
vP91+8MbXZGnn3pU87DmwcdFWJNNLyLgdSd0wT8vZgQsUAoBt4s3xbucenjfa/F52NUc1I7i3WxB
LVw2sLjzitLjBDKJN+xtZr/83sWt/+R+xY9EIxDcQN5qwa+RqjJDpVESWrlW/PMbtdkB7Pd13nvG
VdZJGXTtcKluO2sNz6c6AXTmYJ8DYREMoHDtDzEiOgILebUNUOMFHhLR7rtJ5jqarKyZ8fih+64j
K3+4g62Rl4N3TlodRx9smByuOK2Or4Zh2iGkx0+AhyobYrmtOgsA2i/ZG8d4kALKL/TwYT9X5YsY
wf3oeKvT+DMohVUkC/psPScGCMx5310cD7KXtwsfe0w37mik/iJeQZ3lYqITIt251LJe+8KWYl/U
OQ9Uu2df3lDlFt6J893RL4vr5td+x1Imt3Hf8lKTdapjaLEDycxP2tumWRAn599XRLouvTCFijUw
hK0nPSy/hKIrKLuMJlL/SLa8jW4OV+ma0+DEJqfHzYioAQXnOpkmDfOJ1cVLt8GupjqzNlexECOs
V8yDDo6uJo3P9SzdZR6G0zHNUEVmx1CKS0MVoVCZpIt1OU9k+MYIsATPOqqTJ0qoWuvOt7aHCAkp
ic92PLLGwes2NA8xdTDjBOCJpJMzl9EH1eKOHJ7fyi8wl1tT6qSMA9U/JEzcUpK08nuV8hS+6Hnr
cKs6DV85IAWBtrARX/48kwDp//hEMd1jmTVt5eBC4W2flOqeVq1REOcQOUG7yLd6EQ11nesLtKgP
sei2CW0ts72DKdUWNzvaPbT2iFVy5QpUFufRcoxGNT/ogGoEVv1BNExmo0ypD/+YyYrCT31A2Wnd
unjXbJhWz8AD8UwfpbCNjps+7t/dnA4gmndZBRcY56Hy7qg8ceKX7BElkvqqoNdQfU5i0rMIZGqE
FjChWD7W6PblOMHTCv3CTOROROH2p61tOHpCTmkK44wCAtmtpc4VoOQ45xCWLcf3YK1YRNsAbChF
rm8nCK67ho23qfVAJ/LYC/I7ud1cVCBqstAJQGfKEW4z+QtIy/YWMfZkEUre95QZ0XulWwHsC9k2
eaN+3BxG1LrbpDbs3gb9NPvFEf5538JbdjqKwbVbML3Sd6iJ37los/zqCj8TEwmg7wbWcQfRftvi
f1DWOlc+W6xDRAXO+IqYZuiD7SQ7LFxY6Nf3eispJVtTfWVKbJLVLn3zDa/qZB/C9OfxkQw0v9br
7Pq21HnEq83haAELJg01pX6gNANBHtEaY+xnhPlnY229tLfDwTV0XMNPMHhLsrTc1LUr0Rfb9VOc
1YPREuntV+Tz3odnFne8A7pXEVOO6fverletZ1D2bJMnHf6jtZGcrDRXWYQcrwWZ64+ZWtAJjUef
XBOtLAKZCFJICdMKXaH1Zh0Qh1jpmK9MdRWI5WHlQ/AaVYBVDdmgBkCyTf8BpnBnWm7wpNb5GdvS
WvxnMKUjS1v2s37Cg2rGvx94jXbfhfeleHxkYt+eKUQOslqb2jdZScU+DWzHtL3zJXuC7eaYF0gS
h1i/hhq29tFw6+80R25K9JUD7rHl1XGFQET67u2sZ5EYwziYs/t5Ugf/BiAle0gwMlIQyyju3wjB
5detMl+kLqcO/zPWdiE4fgFERsmx7jgjvyb2VCFDvlz7FzoXasutccQ5BUPtN5JpZ/ySpJjIEGz5
ecTNeWrgJZmBNCl3JFRDA/4e9EQkBg5Bs+issN+pgKnjd7r9rjd0+OjDOnfKYcFF6AvRwLl3XUl4
CNK6dhdyknMiOjZI7XDuD15kcZD5xojiWbauU5+bCETmMrl3xPXEWbbOj3dpWzPlvdT1Oi6Wl60T
HbpUiapF+NXEoZKQHLHNNsuxa5xvTZ/PgKOIVIkOG55gySviaHlOrdfw4ciH/+Wb0JzSrUtAr452
HT3WHApFHvzz75QIi4E8Cg2eOY3788jEKL7+WV8xXowqsySetd65yvHE/dyyqBeooWTVaSIPc/qW
MTc4SsLRU9c3XfnIXoKZUhM1whqjhpRhTO3gExKs4N1EoK8bB9bB9r3xpKEgdUk7EBf9u3TEK89S
SE0wmyhO5nivJeqAi6nXPnA+MfBlu7cN6ELbhlJrx9Mj7ZX4vL4InXeH05GpSRTBgqvKBPJk4UFa
GmwxdRYNXqgF5YUcvmrZ113BkdfMebfoGdmNxLqGTgPv9Yn1mPheGsfe4MBf/Shh8f+2anleGl19
DMqlKP122AMTyxg89sM2Hgi14C8anIC/oHs52zrL2JKK5rOE7WxawMJ3TTTgkCsHlenD8WxZ51bI
X2OZy9LVrYQINJMCs0Rajze+2RrjKYhXwEm4Ibm2QStxI2XY8JzQeNZcAMM5B+jaOECb49ry6geW
oJzxA8kge9B6xEG88pdzXHyph29X6xginxniyKHJPRIUS6N0U4UO8LGBvs6PKDOGg4j67Dp2pasz
iBZ7AHk8FhFOb1LicTlzO2ioYgh4SlwiYjCW6P1tRNNK/G65tzWK/eIo0zMlWaVQJziM+wouleTz
pu1QwIns7UpmCegG0UtEi18mvBf84qMG7uGfeAxDjpz9NodDGUg2UUCTfDtchJ+OP9NKC9G8H2wf
IosRu1s4rVu5GcHvpTIX8lD7cwkY2DRGm8MchQZS5zPYF95D16whDYcN4ZSOIBQtB5cxtCrorEx/
Ge7xQrGBFxHpCcsBYatHeFpqkjSrMALpXhuIneFFQ8V2M6nWQwySwm21EsD6AJS8F/B4RPs0X1Sb
eGblKs/Kzujb0Hmq5crejGrydmoxg/M+PqpkmRzUF1zjlmvsomLSxwaxnJ5pxqUgGgUDwMj1SsR2
yszVl7blqkp/wWCRngJb2ovnqSsa2sKNSnuB+69nL3idIrRmahMz98lI1n6fOKpst5pomgBaCR4G
CwnmIJiTVcdDmnxE8Bcvtw7x4v0mYV+n4n1/UmpFLdEKVlfaRNipRh0Aeve5eroQiKgxFhi0WMjb
Tk/aKoCS5F1AKPkUWCFBkx2FuWbuj//sTS/wEkwPIiNUiiYUGBOiatoZRo9f0m3NT7OJrez8KH8R
QRzQiGptsGTwv31jEbrt8oaomQSTY+/8+8nf4D7Q4T7xNLzDN3fnCVLFmH6R1LrZ60jZOaUmXa/I
1NtYQ65guHPlyuV8N/d3XrtUpD7ILWu5N4JG+pjy4GIk2RByjAPQN96NAgVY8Xi03bPO+gh+Yfns
klOR8hnPRMIegyzxP3x641hS7kJMOjCknf76pr3K/2uUveOzh/2w7fxcYDYxVHzn/Q4KfQRZGIEp
fN7HZJMZ/CPWJOYECLj3czOfam/5NpqQe4XeXQWYYYq9elPlZD5mYVLqXtYt58MIiR8mSES0RrQc
SW4bP02ehr69mywfpqBg9NXqll0Aa2tzPSbmiU4qjSjcsPCGM7Hd/s4kBCOJJOtglEHwmmCh+c84
eZuQ430/oSoG9KohK0cMTf57R2kZF264XKU2tkSaW9hBfFTMUBhfS8BkKP6ewmDJKjMPWXse8PzX
fxMFyMXAYrPi2U8aHcd4BNFHlmsJCDvGqD+YodiwWesyv+1ApgP5/ngjOueAhOgBzMnsYZdHT4wP
477uiJKBYJIpig4Je+mdU/cboJJyB7C2zCVr6+mAUwz8aysEF7LU8IDCWt45Irh86CtRIPep5/T6
qjoPze0Nj1xhtrWi8s4ExsR6hfcxA+VVVXxAPAc22/IhVjmVYMEIc39fPb8RY9L0RxXKWFLlgbhS
smhseL6mdmuUuO4FUhNrTVkrnPrZtyyU6QQ32/126Tn1RYiGvKCaGJ6wkDnxDINVwQkB4Y6v41jV
1yIYAuX0Iup4FKyfziCpj1X9YXM2T+gQoseUxRfE3ZmryomQW9zTvsJjpwiv+AInZpuplrtWrj3K
Zw4GlgJHcBY3eRJ/tlultKGncC8VW3dvl72VWTSHIqJzzY3+phwlXA6iVJK6ifGITFYtsNAlflx0
bGc9R7nkcIJNWgY+nY0QsIz2382Axkfe8quB5F8WN0Dmri4rNZ6BrGWL4BFrjr1r1okYNH11vgJ6
o5RpJkfnMta1e7AAwmDLwnPZMe/puAVKAPMZNL5wkF5Dy3l2BsLIftB9xAg3efdsZoSKfHoAiIK6
PkepKLTOiA7XL+XGSGw74TNvmt3TpSeaqQm++DSd9Li6NVA6CT3PbgK1fhUewA47Smlwo73AwW2t
+k8ddVZG/gP9ZelXVPMSfQqHSdjV2qG+FkClqCYi/d0pVtjCazXES+uu8yEwH9529F+uIF0E1o3X
zwX1+YaA5yQZQXowftJhEiRrWABXvIkH7VFUzdyN0/gJjxH4iWw90gSiMZ46J+dQSv7bfSkm9Lqo
G6dKYF3sz5Wm0WpJeXAI2tXWndmFWRa+FTTGo/6fLZXd76237InF44RJFDTQTO/90B7S8pJyD7+E
1pxRZpS+9Z39U1hg0nfpCiCtV+TX2lUh6AYv58OyotHQhlWqEVB2wm2w8GN8IykH+3DxJ653T2wa
2kO2noTWgoL19t4pFSGKHrScLaBa2DbysrbJocExr6vdh/oHlJ/1oTkBLNQjZe1fKnvcliXUemBa
ULKqetqtRqptPLB2r6VUzI/P7js5POJUXzNYvUSMIhS0aP3/GH2ZVFLKUPGJLij3rHnpXHfidhVC
US5AXSNoeqHGNyQ1inP7KCtnc3Z7Exrjy/hxJrytb/F+Qw3urS0oBGOv1uZYi9CmgmNGFKWT5VVC
lYgaorn3WkWL1XwHmEs26cEDzDu1E7SJ/sW11ke/gE+2eOx6lj2PpOz3mWXGUXozXGcjeo9bFOBT
Ho5/8tO5BRjFRyKpXlyCgGDteeGpU0ZWQO+AhIk6cD6UFv9aVYmblwOWLTwT7Ue3ZmZJyo1TIR4s
nD5MiE0hGEsgvzuzPuUF12mc33tCF9jupg8H5OhpzlWWJdzsciZcVdB8qLQ3QFgTYfe2yiK7Qr0Q
bSOx2c5JlE4JggS6P6aX/RnADKeafcI8RoxbEzl3aUO2GlxYs1BWq0o5w/vDGUhrnZF4aBQ4p4xt
DkZBmV9XjX1I2WLmXsBfeK4qzJKSgbe4vUBLogCaTJYC2568e+lD2AjEvaFsGWr2h2nu7yJ5DSGR
K4JGFWcwu5tcHVnd5nCU9rBFc9LqJ5+wcfhfz8IaR88ksxeGfP6W0PO9+QJVxszMCudbgdBfkm78
8Bb5zhJRgyQmA4kQc9ySHmDi+exDbX3nNm27HaIoFdxckikH8I0TEQ6MNrcQsjlMQ5q8PrKtwPqK
lf6RLiUye3zkbDgrmgsqOuCgdVsrtky1kFcMFl+gR675XWpjyFBiQlBbFSEgdjNtc3EHf3eyjHxo
bdsZSTp4LMvE+PraWjMX+/hT94Pj3LiqjJcVIk2zbVQ6m+QyirZGcc66z2f7NeH+aiq3z9zjhK7A
DVsWDtlql4OESatPXLkEzA6nTraftE4hLPxjORwKmDKzPc3U/aHg39viorYrVf7Y4gKBWMQ2vd1K
yIHp4Qj6wzuZoDhBeNGZxr4rlAUu1vvwPspC+2pE09fmtS2ayY3dMEL91/WT7Bu3/Lw7gbciojmr
eCM+S3vO07xa4KkPZVdds9LahT/OX5VwCeFbNxHGy0N2n5wAM0FKrxqtb49B+G5+rG86unzw+Oud
T9P0KKGGz83EB8YVId6V8HyIvjcNvVM67aLwTLnlrcBt2Ieu2NWLnDdTnfPqn7aG0JeUYYvWVWqm
4omnU5o4Xk+00WgR5EEqSrGxRBOx37E9Dsfx/tb49bo1oT2R5WTbNhMOKikAXqvxj+HxfZ1DCGLC
PhsGyBBczBh2kI8rLs073iQvc/9OEwhucGQGr4GC+xUvV25oujqxnlZvCKpflJRQYTn9QsXElPrL
ZYAXzkcc4PP8rWZxxH1M2IB2OQ2AF7k5DESm7GObOuA+Emq4VUab6WINBb5WNqDsubYr0CjgRVra
KOEt6IbDNXqIYv6hvcIrCkPvUhb/K4WLNxr04RsEC7e54ZXVJ8Rckb0YCHq9yjbbT5GeHXamCXYP
lCmiMjsCbRFFd6RqTqqaUbuy7Mqefjo6ZRK/Xz9E05F1PveBkcnDB9EzeLQriTAGPy7zzzYk4x68
RUp7dwEC3jOjPGLBmwU4c98sc/67RYcT4SZu1TecJ6RL6gRneqbcTXbrkcnK8nplSm+iTr7yWkFf
SsP47yyYwo2SsXiCzdCteCl0TS53CFrLyAS2fq8IZ4oAEeKU6/HsZmfFwzffyIvWKzZ9MS5q4aiW
MOrjf6BOvzHmhhCvWvTigiwMqsYUVtHrF2MAaHYmSudc5+EQG6qaKG41bLfZIG/c1V37OMZBqOi7
ebUmDNXhsUOtbihLMXpb7JpifNQRkKzMuHGab2SHHId9vc+UyocDFq43xQDkP1Occ5wZbmbCzazh
s/4aDJ/AATZSssUEmp+N84vtyYk6ZETLSG8f/xikGj/VBt7eClVdooEv8//q4RPUQwLo2bxsGu4c
3YOpQ73ZvJi73HycKE4vOdSLt1rMxkyYLws9FrndUQzLQK977lArASWR1yjkwyCvdLTaYZd2VWMB
5OAo1p8VumhSJlHqN97Zc7JXEcYWmQJOsO2wJXtjJnaFLBjcmAOzorF+f70e6QRNAfR4QHGZZb67
Mv9h5ElNzRKUWrxjtPgCNUfo6ZTqLGicvQLaOS8zcpxUYlfrlWUQZOFlxtGnVnuL+GmVru/cmGh0
dZXEE00J2AJdp2+2pXvNwbfIYxputeKhE87aU+MKwoXPkF/c3nz45gMvb19G+QxlW9+qWltGM8x0
JQYCyYriVom5sGWohnrhYbFtnZKGkZaYX582NjQZEveueNEs41op2j0kdgvMFgzWSLVvLhJoDDrR
EKx+xP97cU6bMBe3ae065OOs9xlDe6Xs94v/NTieWD2DTmcZBgkLL/I6ObybI5Hvmt1L5iAixzcv
1UVykrzgT2Qtu8OT3Q0FgNwi7SavsebQ0PacCDeyZhY73hJJ2hdf7qYgr6fyvB3UpZ8OaP6P7nXF
e4rxVWOXX7q+gt2yIu1tvzi1LXgEaY2jEnl8OGfhUIJJLJ4io9a46OtH+azOk2pU5gzD5ZWCw8Qe
Y2oONIEe1Ah8qjzPVsnRr8hjZG7us8Ve4O6WfU/PLl+nHRKOP4HwgnctePiGPyQrt2f8Kks+kZ2L
5UpNHzJ6yw0R8iu/PWhepgZPsAjPiImPPpO71SlLeLhaNE0I2iE2BbyNjVPJlAEFDMcIZbZuI0wC
cVH/JpnmLK/dnAlj4jsKz61GQdj85Oh4E3j/ymEg/WqrQ+igC5EW17ZaMFEXL2CoK8ducWEZ5YF5
cjGWv9aO0p6Yx3Ycs2XUTX9H/mNcNs/koa12vDTg2hDIaez26E/SaBw7vWeQDCffwLH27j82OjUs
xVvzP4nq7idXdfINazS7Rz3ajdTP37TVLCql5AU3dcqLr+IR+kaCPDuMUktYShoalJL8M1daruVT
nne2Y0zZWI3nVGjufI+tAqBVmO0aL/y/Y+yaoBhKkDctTKGj9xixtkBw7B2yEVb7OSD0VlgHREva
qb0yQC2Y3uEHyAMvbCVx6Ye4lE723ivSBsaBVesnqePyeOYFiDDzyX/07U7lFJttQKjeGxtB85ZC
+fjjgu81k+Fn+SUth3rCUouduXleSOg93//dpwmBSoMxFmzbW0jvc/8K/znju6DRZGbT9ovyeZIU
69hNGZ2UQEDv7Ocq5n9LfkY0nbLbt8OqOZZlsgcTr/RgQXWW3uoA/iZ8lGoa3MU3S52mEMrvb18/
3n1wYjJV8yKnY5miIy9/hDI3s/pieCAAJL0Cj1iwewqhTOfAuihlD/dCSjePyC3QnAtbyp9yowRR
z/ujB/iQy8tDYWnLvAj1dVp7c2kLq9vHLeZ9pAItbP/W6HeC5TqqgqZatnBRc2YyrENDYwZk17GW
PGAGU9IC+aVRRknzQL1hmuVxPHbDRv/z0Lavcr7bijhUVMTmU87fj9Ozg0ADdDhxlJQ6iKEkVLna
qQILnu+wnksOEBvQySgygyrJ4apMz9BPwL5BBcraLBipXl+CiKwpQz364kfmtB+iaVuiM44BqVKP
I/9vsNchBKl/DHmc6oRvMycY++djPeVMRVf3B/YCP4G9lOBW4I0BvniRaMwNjcHcxdkpX/2tLYJH
drXVA5bnus/ZsM9aPjGbDQ0FGFRNSIx0HkXdYkN0RNCMAvJKlgd6giqkv5ffG/Pp11YOfIjlDg2g
RJZqKdGMuNDd982enDkgNCx9cDGjrGXvgfHcNHFEaFFSuoUgrHksy4KRED1r5Otiw1GtVnucjbyC
IBFL6ynYV7FxknZyl1ecMGFCkUokN30qwr1p1u2cjm4iIGrIa5xk/gRn3zM2IftRC0y1oR0uV+QD
1TR8+w2L/ySYnOwVEsn22OQiU1PvOfaf8iqDKq1qSC6eLIKRSIfrTMSeHXAmvKN5FWXUfUlRLQbx
yl7DqV9YaZCxM2T9pEJhBoGnD35zW9OV0K4WvaVhXQT9sLKiJWuPT5EscI7n2O7WWlLBcAyMQBGO
LrfofOSZF0etNab+iCJ58vX1/VAEGAuGhLpC7C6dCruZIN6ariK2ajV5OTZhD1uGOQpFVBMH5k7P
rBRZ3YlH6HCHinshKDZIiwx6Kgq+kqfdxI4SZdaq19Ss7MWcJmWmEZDxUNJluoZP5+9niGPmjrHK
2Pc9G2WIXK2YmRyMGJd3EWLJxPh/U3dMxgvSj5HskgvpSQx6w2FYH7LWDJrt4Z6aLjyx4iPVhQAQ
KgDDIzu695p9xUghQuR85ivraqiI/sALM+qvBSw3fYYsUjdeojSPzXtYMK9wMxXD0q+YL8xPVzPy
KALEnU3VL5YhfKg8XWSZZ8JqM8PdxPRCfEqP+BVhwFnO+Hpcp0Yt9m7dFbKcdpn/KiE978+G2Vu6
/nLrynWRasEyYQz9F3COCdzTmnjxzMfRhO97bmNYerEoiTvqbYgL6pko/wG5QmCJauU/9nlsKiy+
tWWtx/WmNC+CInVd22lQgkuM0ftlwVGwG0zRjlAVD2wNpCLyGe4B+NNKHEHx2vVtBo409d/f556Q
PCmjuguG1kNZZb45GUxOTc05/eIh/pw/O4zI0PK3iuOIA4DuTo++sPIC47UB284UvU5AbawvX7m+
0hvreQtnCf0D2wt489q8ddDl6U9TCozDxzY6bVMfDb1gU9yJOYIPBB/Ww4uTtiEvA6SXfUcLJInG
dIQZBut3WDuwiDR7D7lUoyzRjAwe5JrHr2wNCjb8FBkcXlVwKGJNy3f/jryXnjmOluuVNfzBkAws
MgwyrQwIdi9lMrhUDJqiC4rMThnLIwh8qdQnH08/tAmT+B9SGPnsjyoUA5Zg379QeI4GlHSRKJbH
N4knToFZqvwhgYMy4L+l59Gu5Jc745zEyriSosaxyym/q8gMNP059pf2nbHtH/15tqNWV71HOyxg
VUPYhU3w1N3ZvFJlwepeA7i/6AegqqSlsgU96NzMQ/eRtfFp5tn3CUsE/igCZ7pGeBkX4abvjoI1
71xvZk4AocQIu4Ygl7PjpVloM/mDxHRfS14Y0rtgdsP+QLTzVMtCUa3nMoX7jw8RGully5A5K/Ft
ILNDpJXscUw4ELSfbPIxRQQxoQspe4ui2GwdJ51RYId4kcYI3A9nkWOQ2sG6XgHLbFrkLTRM5gnR
5mgvREki0OO0LmNbzEXlts6Yx0sa7KvlBwxQeoAE5ADTuHHXnVV8lfM7sVl5v3RzguMAfC6p4LVp
ulWLj6Hi1EbhUglHhot7KY0QPK0uby2nQrXI3p0LnOpNmoonYWxLpv8kOKLYOSEtMwKIa1ajwRPV
iXUEAWBg2N6UytSkV7/uCkRDI/ZSi7ScUqakATUJpVaAJePUiQmx78fjehL2QwcZtO2UlGteqawp
iHcNEPn4gUDCOgnbXNSDKhFWkeatf+k0iyaHer2NmfFBjRWFeaqG8bITdHaJlJe/Ky+6smaKgOT/
tRuTZa8nEo/uhrpB8fA7y6VeCVnE4dzISedQYjzT4ZDwO1hF/hKwJCkdU0DuvKHwJq8DHarZZkfw
vXUu+xkX4RsVbVVt7aoeNLRhfHmsTiFJG+AaU/vrmUz0R1kPSj5u0zHwRABDGgE4XYKa+FTJ0lhC
Nr7jeIRc+t1keh9G9e32ThQ9f1vDHJ5w1zK+5A8frxkeNTjHV4aWlaAh56iDxv1QLo1vEe22d64w
Ca6AlbjLui1yM27MC/WQQlPipoNHBHQ4oqUWLL1rq/m3HrQEnGjEDapHs0V68vO7Mknn7JgPow6q
kxXDETrOd6nztMbJrXBkLgnoBWAeQORrkr2DMPX2VhageZdomTqZNyq+ADqbeC+MRDn+mvF1aoFS
vFEhyg8EOeLRIQNASUzyVWegVlijYSBFnZTcl3ijhIdoOxHFqmqeA/rtmNCey+ITDOOmsJPCgj+R
ZNLYKsvL8uy7R3AHS07eQdJUAxHLU0F22tRUoSoib6RcStbWpH4NdY7ThQqfJ8JHTDSknFspI9CX
nuM+WZFAYu5GMHAfFMyzDnYKApF2CSoBGwyfHVTX2wYrnAHE+31fGL8toxAwcWQFq9MAwLgoB6og
S3xfy+63k5Ab3jWKoKQf4YUBqHbnZLtvxCLYO5CbFWjbp7ze2MZH1ZnKpbfdCAvZ4Hx9xgwnEU4u
zgnMYZMcg/hKCYFanEC93Ls4u6EhqNuGEbjChwr9NeEvAJk+3NlfUeso3JkF1DNWwec0pbOxcjUk
5s8yDL/vlvSlMAvGYy2FxKpMUd85FzAf6D9lTDjlJgqlrV0X8E98dvYFWD6iyHVonnsgUNKfYlQu
91wRa37jXPt9gUI4k5PrqMBqFxeaSlQWOLfn+t6g/+r8LLjddfsgLA8ieerTip8KMmX7CnA8tkEv
nL531icj/hAm/fS35OCEUmIJaXrh6L3eeutMJhWF8xPWL+8ml4/27z9hyr7AN7LJL+sT7YW9jVwS
1cOhToM3YaPQmtoBVz0TA1IeGRW7z/gdtntmV0qnCh0awKp51QwfeBcb7+8JHbXlB0xp0iMgtIao
yBaZ5az+5hOhZ9JRSyGOJdk4sLj1hgTbj5E9b4U6lqnqkBv3J3+dw17xho7XaGAbFn308et9zkOC
Ji0dFGbYLatfJZnQUlYKE/rR5abKM7jC8s00Rr/xIgC+FLi8CwwFgOYU2HVBiS3NJOlxuy89vY8X
0pFWh3//SvhLGD/4wkpo3e5zwnNqiqWmvly0josS1JzZmMefBEr+oJSMjSmqStlHbkpCNPLJWFFI
fKUQYY9b18xZbQXOr1earHTABfQIC6dTuIoXG4qPYzyA0xuvPl/5jf6HN327jNEZyGLupFwJoe92
vUS6ZKVOwEmf+jpkKVK7PmC9y9OyWEYl+YFxvdFdnbkG0N6HyFi8YRvrYeKGg4t7EZPQBpxLlWV4
6IzLT7h0teDVu8seiiprNsn7R6/IcS0/oiswkiEYX+3Hf0Qifq56hKCjyTDmonpyj5fVxtvTcBgB
CkDmhB5rTORFEFxT22fIodPeXWPYd90Zn815wtp2q9xyP1MmmJX0TQNW+vcMLaTPTTi3SXztiBgu
d6giqw8vVywVrIKf9HpvDPrx/lCFXhhaAG9ZKUPvW+6dpNHZrvc5ssfNY6HEr7ISRtXEPhYxlzSH
RM+5E5NyfjtwFx3SYleseOkKgpq1M10vdUqF/ICHReQDPljduLrMiqRKgQXEh3sfY8A1EiLSERFJ
P7H9pvVneEVmLcHSRGGaHnsHUsZ4M1qdFT+P27Ijx9su41BmkTZzY3wZYdbcFYhYXcmVAN5hICA4
yKWUs3T80ztI47G5+QipJq9AZ80FcyJ4P7Yz0zVH74PRa78V7BjnpFxfyX79KPmkZcOhX/jW4shI
JwRXQ27wzGCmwGL6VykJ4logqnzWdKtAByivEn0dw/AtUNJG3C6/o8mx/4mBdi5zJWWRvNO8IWb4
TCiAGJcLwq+bQXvrydv43kQxgkH/73mGyFwGayJJVtIO6bbf4zL0mVdQZxXwItxS6HeG9/m1uYHj
5mz8/W1zng92xG9ruTegVyebAYc4sSEiFP5AGuckcctQAqRhOWul+WVmtDseIAZ8RAZoxR9o87yI
/v+X0VNB+C/kM8bDIT4NU7ShATSGtFypC5Wz0f2QEfKWFF4xkQkN96hdDDXbd/A3N/MLhG3TKubz
3sXEGD01MmgQ5DUSjiKOFZc3pi8aEJb0sAiYc7oWPoyZUiTADR7UhYYnNmyrvd3UsladlvwjD9r3
kTpWuPDNpOsdmcLj68DsNqO0bHbRgT8YbRaGypbNWSEiYLCkrnbkIeFP5f3vjvAmXKm0tW6doa71
zQcj/oq1EAp50srLyX70TgOOyx7gYlkK6PdLDO2WN4IA74y7yKoc7uPdP/aeWQ+6eqOL3RXUA8C7
ThKvL5qD6dLhdSOU9NCDqpFTxz2ur9hk9fyRbvtFw4ls8Twj5mVUScyRbUSq6qJRkE6IocA3XqmM
zT+ie/Rl3xS2DzrChWQo423C8Lry4mARmrTIKe77fJ8hCaZP56wR4hbghjsXkgo3r5jHYwV4XKdB
hEZ2x6QSy/VqBVNP+VqF7z8SyOTDejSO3W9IKveUeiPrXUoDEEuMThAhYoEJxMoBaAkhG7nCCv9a
O2eMLnQKrmslDbG8rP3M+3DnVUaPkQ17eN8AGa2wHh/e99IiAqGSaqfR+7LGxREhJpjWYBlgU8b5
MNSHlTKi8CEAmk9kR4Ah4ZX5qxoQftPozvRHQ2TuYzpnewyj57KfVwFzfeOLv6KWxJvFwHitw0sN
tGJzCQo29nmzrwtdPliQ3sc7mD0cffhRn7LO7DyGlYwERU51Vc2YecKEs9Z9x64s8dC7Jnq2AC8o
lVZA7L+J2yJKVu5kdIe3ut5Lk2DYJM9ZtKWFnUgvmnBZ3b+K/A1WPYDp5SoWKcaF6Cq8MHRNNxUZ
gvY/IYS1Kr9xW9TcD6rl/dZsw4iWHEvZp98oXGy+tSyor9ukv/NtGWeaT/BIaaXWj4m5ll8Upssr
jR1vbJMvO5Gb/reK2rHftripfXKyze1ic8gYBo/ZkSLHi+tYfCPnoDD/WsYzbncJaQjyMDuVhvHS
KAxi9XfmHmflSomrMR0UH34IJoqWiYRj56YpuMqKNTUnpiHS9IP/zTS8h//C9SKmvh0xcnzlbWmZ
/bQWJp/dBIiA6F3pF8v0F34uQJKGhQeGKBxp3SS/g4ezbRxssBpRSeVgEFs3bh66ZevYqKk/V0cw
GRsQ05V3UTw+OFkSJFtazWif71vwI0N1aFbWss5B/L9YQzYIWooVf33gyzHS1v1GnEtuEp9Lox84
CWfVehvh07gtVrEL/ITkUqDE8PinUskm7Fagg3yyYj5VUSMyYknTn9SyyoKNTShua3f9MGDOaA5l
xgkhJLtKTRznoQ41ObmhKT2GjiWexgCEGJ9cE8IXqEEQkl/K5P24oesPcvaH8TWh+bD19EVsKabU
hTRUIq0+s++/XZn9+X8gbm0Sh4956RsWdfWYxW5yuE2Mdq+YLgPWxAdjmjk6D1nC6MOR8kvDYous
1/VLLVLtJfvuucSZHwfT7UylgXFQHW8H55+aRMkpp/z4bLFugfzRRej8g1fsVqzweSHhJGXqqBix
Kly3NGeDFcVvVHxzXOa/S+YrRcFibq5lyLgMEwD7dwhssaUPQ5gUnJlG4C9bWfJzt69PQmMDFExa
VXu1QwageBoD32cNvqVxhXu7V0QImaSuYZ1EHOL9WEnW+F72kSGpVeHWH6/4X7keAgS/IjKNDN0z
SCv74kVvOfbF79jlupMKWZhZ9ACtfa3UvoFnXKtNPPJ4uuX6+CQpAtS5tUxDinfU8jiYDu+zwnnF
fgzl2MprTwqxOzcrhrQsiQ53OFapzOgy9BPCP4bfnEmv1Uh7PQWA2vhbcR1IoMImwXB0zxUVx9xT
P2lElS8JpYw/6vrWgzOkIYBYBNbaGcI0BTw6t8Um1BPinphvy6l+x0c17tqaEk22Z9Ft2/ORxr6q
Z7Kq7il5iRzjpXakl2PLchoNDEJhL/GuUGjjdzAng+KDpeGK8cAZfNYFIc6x/sFJWKw/cT8oyrQd
pIRkTPWEc078xaGpbB8gzQZPkP7t6lepkK8PFL3twdAJ3dvul5WNmmGU0gUtS03C8vmIjFDMFVJw
CqKBmwYzEN8+77mpcUn8JC9GIzMv0olNqeMbveOIyxp874KX+NUSkT+2+Z+eXI/3lJcJ/eBPueGD
2GLVFT6RnaZny1tkS6kgw+H9g7EzEAVS3wAGSeIHF6dIYwldWU6vly7i2Flqox/FrKLU9ElopfGx
hdvpM6QyhJBy/jlYahnibM23615bhHcdlgt0GqTAsJd3yNsGqXCFzS1slKwo8edtAY48VhOdYaH5
FTUhPbA4DbbKHQ8mnFCz8tBWwuoqf/ztxOy54T63Ib8JVnbwmIPOntyBqahNk4CJ4MwVypO7g8ld
qatggGPQHGdNo4B9+7RMhJRAC2Fdk9Qdz9sNCQIvCoxOqxdN4tNaBX9dNpPvWVF0bM7eXAXDlFv8
P2dY2CLeuOlHRCvc8YpXaN0wB174ZsHQ5cU94Xz4DXPIF7Lcnj1MBLiqDU4L85dG1ATldBmSBq0G
dNRnBsVYZmNdbua8hp/c1yvgTE6G7tS6BHm6duXnopPdjfffdedzDjNvuHHFyL3xeOkFL/xT51St
JXWCeFEPwMjjR5BRrfzwWIdjORferj644DyO41SiBHRqdViVMDB6c5Cuzp8w9EpwQKLrGl8zFdgQ
VyXPgNacusWKNluRDbDx5vM0XXKheXJNMYD2uuuRVIu4llN75ZYu5+d0eajQOIwjBpC9JPmUtmtg
TAJAKroOd4JQ7+9ECmZ/8aery2IqPqrM3RdF/YJG5c05NADDUzvG1z94NumKrmuJYfcnEzs/ARDp
YrgvGGwAfj7EL+jSCtP2GU4uB2RTCcRe8HMShxy/IYmQ6M+JZCOqw036X8WXtiLkRzg7n1nQbq4Z
gMCwQ40hgRMkpZ4YGjRKGQqHOXb8fK7OUj7gR97wAmgE5B9l9yKXlryWD+JiILJVcikIANIZcX6E
Iaouxucnzjwod/B9rq2l0RiDe0FhAa+ctQQ039BzzaXj83edu+Iy5Nct2dzobK5YRLOpRbJ4890Z
kf0wti3hYwHY1/XTvRuaWZzL0DeO1/KboavDaBXTC3caQRTbkDz+zF0DY5JSmWqjfi/iI8AeOEao
FRe/wjdhKEcAUe3rdwKVC37KR/bRuL8uwflmJtsK//GiSe1i+j4T/ztz+Hh4RUdxXN5zuiP5q1IB
/Lw29nlE0AvwtvzP+9df6TmHM+3bPonEBryEWqiC7Ugm8geQ/hrJVYLBU63yKUh+8E3IX0vkh+t+
ZmuZTMYxLkFiti4dmj4JmwIQdxmHouNbNLJKnIq8jwuRovir5y92v/b9TAU2ywqKEaBA9w1xKkhk
ITgogkOTszjvDFbnvgvCROmG6FwbjUPH1ci6VPyInaMgaA6+g7U7SJTNRSn/d/+Y18sji6uhj9k6
bn5yIkAxyXSE4dKyfkE8S+DXjm+7Fsk9BSkIZF2ULmnyS4qi28BGOThdnrAj48tO+ReMe9ucWMQ1
RMBwlgvlI2+FN2lww/vyNeXPoAqQiBYDJowzcFZmxBBIwUlHxeEIjg+hoWbAQcpYSI9n/8j5kTHL
Zb+EuEaaq8u3EKoMaWZjF2Qbp0l0nROvBxa2foOfoAWOeZH9SGp9/DRvo4k7BlR0rCOXMhHH/Ku7
npLunkHUXul+QZBrIgqcbUt6iUpPQUZLTkdMiAY+FoxKyG5YhjMFrMsyjBb1EanfzYA4bD1Owp4v
O88fgO11yv5bsWC4H8fkhsKZApfRotIBQOsCglKv99/Uw9lORdhXwXsLE9yOM22zYuWZFMczvJMv
1PPebobrg89LKsoMG5Ad+SgUNv+Q1oinUxwc882JLaM55tTt04STRvUZdLO0B3M3h9avy87XEJwM
h1+9E9QOZ95nv7/BBnSLCLPArDVooVFKa3DRA1bsadelj5Tx4CblRxXuq9+V0kVwn+r6N/xWFy/4
XEHNpHJakek2izyGasMKhe1fNIQCbno2IDT3sDs6vhiOyi4UUQG0IJfIAFkeErz+azyNLMgNq/sB
BGlMe85vvvs4PDeUq4GbEirKSeCnU6YnIfrEDJZAxOrjMImZiiyoTknMH3Kd5A24eELJ/ZXI9kki
MIOxpNoIPJqGMt/VYsYVPxtbOWt5ggXff/YnDkfVqH3WJtSzhZM/B3HZ/zCdl8NLiX17P1xrGz5B
7HNWhelDLc1xYB04ESlB8JG373/5W1bUJ7PINJZjpmXC81PTL9U0MbxPNJogOFkcuvAtZMf3fhPH
hcYMe/dIsEhWDpcg2w1XJHHMZJpFHnuT/lSu8ySll4jAbz4T7+zh8xTVqC1MYXZzyHZkN7ytxmKz
M4DagK+Lz8meDRGLI0oGcb4fQxqYwaLDNkZcHhAelgj2uCAoAyHjijIOrJBfg5HhSwYvjG13fqhu
AlImi2hZhIsFZBC8kdlnH1f14K8NqCXM/vOEFQBy5PnVTmcMlG4/zawLXDR6KD+HdRxiU+5MVNk5
Lpu46Ax1pOwbK4SiCWFj4LaZDTVplRZDTfpbQyV9Wr1sW7HxWLp0q+YXHm7sdIt/ZdpQWYFNZ2x7
vcWlhKH/lg/KBenQBidbkvdlRyifckkHgmF3uex0dqTQaczEgC7wxvTZAlzRSiUNtM/+/nvyQNZH
EoszYSIXu/WjnPrgRF4nN5+4Ed+bu++3kmv0CaRiZcLiGfOSX2wKhvYmntzETtQy63YNPuWeZxPP
nj/YLuibc51bBBnyDBg/C6Sk+gHDdfuhe2Fbx/Ys8vYRaLJjZVEus2PtNfyRWnyqkY5zCX0I8Wd6
XED2kHqS/5EupF3rGOTA/tNd3fhAvBJMmBnc6mai7OmnlhilIsXTIyVa1jLN4iG1SupWAUlIchvj
4WIfH2YSUK2pUbjNM5Ya5hECmwvVjk0tijmHOnZszcadrvXcJv1zV6xKEroDKn7HyUfmyULObT4X
yc44CNqX4UpEuOPEnqpQ7Nz55E6x28gIXvbBIs19LRSXjagiKj468Hke0VSjVbRYdLqSpW7kcqeE
S3u749AQWllonsH4LvNpYipGjfW4TeLblH8qcSYIjO0qVeU50iW+170bwuxQ6nyaQfHmoYvxa2av
5EZdYajYZPjjLJkFWdqV7iJontMhx1CQYjp5pdfUhTp9t+hlFddufRTQGi6tBLkDxpmDljJZA/oS
aIADv0leGgwWY6kkYTJB6w+NE20Wm6NnYCLEnBmCoXJmNptCMmdZaR/VAoVip8B3I1GvfzBnT/FE
FJHziodbYr+YABA6QqvAG+QR3gsQMESEgkoGy/qS61WCKwpVsevNdTw4rkhsd3UvTbHUTxo/0GUx
VxitobnNV/aVOVwY7Y+0L70Gc7/MTieBqx2uNgPQ1Wq3qbDdy0iw5ho8kwZj+tHkjiacV6E5zh9y
S8ls2/td2LieKRzNMfpt8eh1GPg5XjYTUhfdLGDVXKMlSRAOk732/1o2FNwdFw7yl9By1Uv6elkv
x0DD+Xxf9c+543WBAuV/U8WqK0kGoSTfQZUkEZfwPIpASQdfFjBzu7LLhOoZSWrKCjOlzOp9YEIY
Z5/dwFN+egG4Ib/3ay5OfBdsVZgBx0+oPsigMpxGHIRMSnHYJdyKr//pL1JXoKk68MShBrLfie99
JBTOWWu+uHJH5EUe20YHXm/mhnu5HFiubyKcEKUK+DEKVtgcdHVNkItLbrewRDEhBsTIOWqSpcfe
vwUrWhvzDnSM8eIfBexlJuqPpdk+dAmIudjTlJ5Lb1SXj3Q3MmOKuL2k7g3gMrwRC5Iw+XL1sXjx
0azNDBbIbEnFxkEtPvao77rcZUGCLF2Ocbu66P390H65qsVdjtqQRDFdxLURuHC6yIgZccGIxl+5
z7k1uS/b5qLzN2c8aN5j0vaDXIHWZbMCq95/Bl5tmumK4IXpVdPatLHJyRSyHYqa5NWXKDobkHXj
WVM0zjzxwjkB9EGEqEgDGtsOGoJTBKZDiZt27MhtdJNhCpVQAtnjgoWmp7I2Bz1cToJuf8hRdy9t
BFlRCjWfbazh4Vf4j8AnaVGkmAFkAbKhfZplzynq+SuYwdpQDFFJ4mPpSQd3kjVktoQlUDtTvwMa
lt9mxJHID5MIhgAuTecxvx2uFDbQYTS4LekmFfxauuCWQULrGrGToHy/QYTIjS4XyqjtYScAZsyn
gZZeipxdsDtNnpDARGWmXvbLbpiSuBSixJ8pGV1sQX803CW42q8yROCCdjuZDCa1V8HrOeyaJ45U
NV9mgZr/5ow6ICiobBjAblAE35pr9b9V7COK5OBIwVgixilzQoI9K4jseTuYGOoLxmUDPA6R/xtR
DCz1tgM7ZrXMmZUfC7JZXrwR7ML9XsbvIGuwVmH4SNVI7RiD1fkkYtLfNLMIO8slx6gvIIQIBCM5
DpIRR/1HeKHPMLxn2MYwIT9Dgltine83kZhcdTDKl/DzrnYLw1AVfiMTVj5ePEhEIMUdTxkPvmHa
mdy6P4MiBD9R11g8HZNmvUMwepQKajuiuZsquABJm80u87Wa8yrjtqiEZh8I34NqZkCAmDakGUFN
2nv+/8Vez9uiZSViZwvcK0o0Cd+qrKUDWX0sJ5yRsVOVUuJ0P8EDS4vSnZMuJVyQ9nCy51i/u0li
QHxXYqL/mMe3+CDjYZQl5hqDHPVqL8HIr9EfhbwVG6zDiUninLs4OSsawTBFtbUZlg0ih1hh0C4f
4Tk2rEZy6w0+vPNU1gkFVZj7mgnU6pK/NFgOvZhmRr5/aGGkLDvc7NXK8mmC8eZ/MOwoQ1EQS8v2
z+qefmT0BWoz3vZHGAtm3qz7fUIXQrH2yzA1cQqSRINNrpAK1UiD4yC2Z/rzVeIH4BzSsGWZQs8X
6gaFnBmOYcJxrIsBl9EKNtrSC2rRlxStjsqJ84S/5iTXCSMnT5fQroe090DXcZIjtv+w7ssmbTvg
TSWMRWutWATioJuCHtMmO3CmTqELUJovLpwG3pZO1p18caDYFX+l3GbA3spK8MXT9jNW6fxqdQlo
zoOa8z3iKRxaC4ytfIq7HmWhoPT1JkZalu6q7wJn5h10gi0VxG+aiJbd2c+JSzn3rbd9n1nAn1uk
wg9MtSguuqOvBVUdBWK3HeUYE5SR2NV0iEsiXPpMHF+tQf3vkUeqTn98/eWTxFwC0JplZmSOWhJv
/yHPXjmuhkhlwKgWC4WYucWh/+i3Ye3wjTHhwU3ChN9PIu4LSXHR01VbgtrVn5R29vs9DCn+YJ/M
6vYcUPcKmgnT5+X/A15YiXqXhJkFzjAmC6gHRzfEMrc9ZNSTMkElFxdg5nQ41jfMr5OWK3Ds9Xxt
6h/IJCXw0EW5WfyUoBqW4Zypa2dWitVIUvo2SwppU1uWBi2GY7n5w8WJpzyeK/k6MQOIxGj+4xt7
ry8EHHobN/Wq6wLacy/eZWDQnC3bVPygdeGRCFBynWde59ctwAYWJ72dXV6w/LsfbuHveQ/FbUEf
Nm7izXTOcKnOfFrD1I5aIEqadmLvEsH3vduLFVxf2BHz0loD1ArTSHzl1ZaYt+4OuGvv88VR9LzZ
ikH13UVQUblQOjbUPke4V5zvDhT0JQDcxTxs6+deKXYmDYAEOzuKNCQgLKC2Z9BDUlE6yxYzjP7A
tDFQje0gWSXNsMuv4zi2XYuReMGDT8HFQqScTXmgbCSGoWQUi6isH/V4Wk/NysiLnetHoZHBJSIH
Gu84odQ1QQZSL0dmv3dPqauoTLVi0ELhdaJjiTVFKqvljs06nB9btrcXByDTpu+3LcskPLXr0ym1
IWA38ezSh8eg6O199uUacVPVY6l/lDO9WSbYXLs7xnIw3MF4xo/fSSjz9e2Mmvi4xv8guHkUAlRQ
xYuzYyFIB8bSk5Rn6Wdx9O3248nxkkv4+FudUyzPVwlXEKXHnZa0v7Y4YG2ToYRefJnJUtYkBoD7
bsVUaI44FOG9bwsiBPxepTEweTlyrvdstPEa9e7MxkyLAT7HXuM1TimbS0SS9gfZ3FRGOiDk2sGv
GF5UlpdD+EduWkGaTJvewDkoPR6bfxp5PPakXDhyCUOKJwGMNCnnzI6xWXzmWeX1OxLhmyExO9eH
PI85ugXLBz/GTa/xIxJldo4nyU/+lYAqcXQ1r4X7LrvkXpqyjeIuIXrJIXrp9sriR8a/AqDXqMy0
RGM2Y+zj9hNKtl3rCcARFeM/94UNDgvgR8JxPGgeBJdda6Ak6KwOlWizawXN1YlWVF9Dv0mTZH/N
4bsGMctO631W0WD74iz3vwg7IP5jG7xjre50ZhrJ71b2z3gR+ZuBK0D6f3q3JH8TXlhbEUqvUdx9
Tg7+beM+pWNsGu+rJcooyQt9mSNdXv3CUT/i+We50dtv+G3AeJndpsj5MV9582ivP2SOc7qRXU0I
JI/FuzU1bvEW4wRXEn12CWg+aL4xOkD9jkmx8j/RYKeHpYnQndETteyLBE3htmLCwd25LW3IQ62x
/ZXBROOGHBdunTNt8/BF656v3M8f+jdvr3nYgsp4sCceMOugoU/lDlhol8GGMmUsIYdrwdc8X0iY
EAhFXoKWqGlZ5ZgKnpcm2J4MCsjK8e8YbiiYqeZcIwJzzgNUg/WsOVzLxq4qH8i1DLvrp9qwiNzB
x4X/oy2ojHtboSLkRghNgEedWzDaxfNOgW7uDoeWySKxt/YTFLiKtHWEtGxiQ3oQk/P3LDeH7uyn
GwVGbV7y9V+Ox7P5y8fxt3GcVFRWRuSw3Cn4VwKCx1sEFldlzEPJUZcK9CCHPlSGdgH8jpdgP7eg
od2VHJj37ZYk3DEXeeoh8pxscGCFlLcGp4lACLmxXa8RuibktOBjn8l3nV2C3FsK/0/49pGIiX6s
oNj+MhmmS7KsZXcQgeJKbFq4Bgo9F2nvCqkAjA1A/YZlUv2mVTS2U5neaGK8bT4R1S8zurcoWapf
Dfw1NoKfSFrr5257hP3LDnqNETriiXW9GussYhwAx4DXXXM3SKO4aIBQXkCavtIr2wRHTfMaLYg3
1p5r6Xssa2Z3kc791Zh7wsTYYdjTwZYofur4YKEPS8lLOH0S0Sl6BisIHS9JrYFu1zNTKBsXOP/d
y1nFAstaiYd7wkW7nqYuyJTfzmQ/ove7nWpzp8m8j9XmDp7zoeDxTzlg/LhYmp5xd5B/MFdngPeF
5I6bIBBMwnewxgTPj9MRcDJ3Eoj9HKRcbTP13Z5lRH/zG6wQpv7EGJ5Xd0atzxywphQexmigmDbJ
4vZPugx987tksHq0bHxzeKsV4Ewd+fdciLrUjSvZi3AIYqrvDRMdDxGgPt6j0x5VZgS1n+ud6bG9
Y/ULUQ5SUuSHYOdW/a/peqUx+0qblWJDNfu5ALpLu+Y8XdFQ4+3cyU2sv0+HEkmOuf6PIG9mQwvS
PG7kYnNpWb2CUcgbxjBeSxLrhWbu8Vx1jYHlKDRDYnRRpZrhTIO7Bur/I+XayUfBH8mrVaSZal8l
ctMLsNR2H4VqCI+83u3aFabtWKuz0yiFdxq0IYxPcTjsNsrx5rgK1PaR6CgqQyKGfbZPlWKnjZyk
3ePShnzPC0qRnNHpvs+Q81VUSOLQuRJS1x4DmZ1R0SfaYGdGTzLfMewEH5a2bexbxDnQ/LSORpPz
FWJHhnORFd0NttwOlBPWJ6mnIK9VA8lrvurlx/pv+ipwrfWVe/q1adaHq9cJ+xVy4DWXcry3rx9V
WO9/FcuVjDIqBuKO++ViVr1fJQf6SLzR04GXQNp74LAoo/XZ0wwXBwYGZu8jwhNsJMYx9krLFet+
P5KQ5jnubRxeortQnUm+8Z3E4CmrnlKIewG91PAcKgYWD5us1rCdgcFfUGU04SwE45mJfxLG8CZ6
3HdEsPuY8x+Tn/nZwL7aJ0Bp78N0zVEzHfs7Fbe2QiYVEhVZ/CxUduGhvfc1IhgrB1zMIqbo1J0C
P0S3XriZcKknNQZp6QV+xA9WKBsdl4/5/UlXbSYYbsXqBLBO+p70pnZuyNrWOqZpB5b2SC2Dn+14
H/KVYPRD/yvrNhmm15k7mh6RsdPnAp0Cjc1YLDLvtBepRdzU5xl8OvZudGECjkvHDj7scwC1zk0B
zwTQIqxxF+UyYvSM+e3eJlGl2u+yN9iDKFUjqkpo6OdGBSUwcATL8CY7kizyUCqXfyAIWqDlcs0i
Y9arHBsbQ1uf13CcPRvRmP6ETFt85/5I6gWH5aDKfe1NZrAkhp6R8P8RRD1zt9dNRItPpwvgm0k3
vlvV5uTXWUG8tSN9CBoeE+lRARkOooAWru2R8dTESF0j/rvI72tmjE6WaNxin7OOio2jWNtQsdFx
ZQdyd0balQ6UL9Zkn782CufXO1pzsrjAl4Fdn8ipzVYjSLmyoqp82fVxhkb444Me3jo9iI3Fqrar
XsJAOvx+ql5srCUrNnobWBTChraGophgkpaTYzlVoOKS2viwM/bDQldUUj+nlREl30D08VtPhW/H
QKdVQ106ufFcnSXYbnLxmG4KpAFW6fvcyhHe2G6dr7+h7SUPRct2eYBwLfDfT+vuPYH7aaaADrh+
VzfPWoG35NcQmbnhLLuXb1Io7fm6aYN/UN2+0F0DZWeNRkcBY+o/AxZZwRmFBmalCGIkZf0j4Dv1
mHrtdn76S7mfyuJLnvA6wQZOc6NwlqZDgSPJ+3Xz+RjY8u4BJEPUKRDCugVh335/ZBYiaZvmR86p
EalsqrWEUJeIKUBv1kotEIiWFR8F9WQ4OdVgRcMs+4ljmHb8hOvKsXu0wsg5PaoMaNyMNf4pHa4N
a49pnaWLWAxwrlNw1qnFl6YGL5/Y889i4/Mlp2bfEd1xi9W+dtKpKIKc5gJYUy+f+lWkqWsHMdiu
5S7dXdCxwQhZyVMvoN8rtfVBrKqiJl2DeRqqZ7urj1QVOI3IS6SVy7E5rSnYohzsMSmUkzttECdA
LNLeSB0TNf9ieRsommbMXD81FSFdUmCdmWlu4m+J1o02uKLGNvZq9EF386bHPR3c4e1vQCm9iVTu
emo632Cjf1njKZQCSYsJQOokrrfpsVWHMHGB60EZKANsqjHXqMmYFcAJ9WmWttji2C57+ncY1HGu
EQhV0e+PajmiVEiAoq7yLxGVaG9FLddB0YA+dWRbCtF8GZ0IMACrXveIUnlaVF9QAisCchfrxVhm
D1RSsdwkGH14Q2uNTNIIRA3pR88Qpumk2Z2/PddEy3Al2Mk9Lm76t9Oyb7R/zvR67BURZxe+mnlb
pvrNrHFqATKBqrqraoAyF5JHC5U+UIntSAtx4mkT3cEL85ZXn1ImT0T8tnwwUiAeoueiuOwmYoQf
lzxtq1yiRdlmg326L7dG5gT/KktV56B7VqQtn2YDYbbyqDMJNYXVF+UZaE1Dh4eGsC0i5FGhKJJx
YvjGonMeBJwtTNnXx0e4w8iXQ8y3I4ICMz1k64eijz3fhGhyzV2PZx0BbKd+B/pLtmYbeSMQ/uMb
ZSjER03hoKr9uKGhFqR0Qdv+HTD2QJ2CxYTHOqQVz0fM2itwugMU1xqBM9sOxqIJs9DHhDo6Cnqv
N0cFCPkc0bntHxBU3roFYP/JrU+cUSbFDBpK0jRB6L2uc56olZYj4gV2rD2Y+jssMMryJJGd8z6Y
qWeRcWmWw0U0lp08dF3FZ3ZRPyeI/7REX5fhzX6KlQBxywd+W+rPV8mjsE6yHUyVOGGqf4h91bzA
vTcuNtJKfaCd0fIn1MnbYFWgDFia75KkxHsQw8r363KtOaXeO6rlcnrrnFza13cubmbEmCo9K56p
DtOAC0grFW3WR3m3xVx2KGEY+zF8PDuPV5zrkvvlx+Qq/wtswFUzteeXb/C9QgYmDL8jHEZRDBOq
s6s7dFt/2VF2/WckeVjXCmXjPf9jI9f7HO0PfCbSzDJ9LaBHHDJvQL5mX/n2ojlLJp2GKCVRG6hs
C6/Sy1l3bYirVDM9XOqUu+x7dSdwJ/IZ+oADK86BLoOsNVYl2u6REJGZeGr1gb70o+X6sp5rnyU6
xqO5iqGC1FDyrJ4v9aTpVx4XXfB+IXx4fGRESiodfzXOAyA2leQ4uq9DS2N3tSr4GxY7c19EcPNF
gb+zF2XdvW37gnasZaEbc751XTebPIYKLrYdAV77EF+vW0V2qYMLoalrgTOIYhzDJW73VNcm+wxL
+x9VNK0Ai/8uawOdc6e8VV6w+laIvs7ui4Reg+WzC0D2QAaeClPJBtw2k8ZRNj5ssn4lAbnbTf3K
D94k2yt/1MxtSRfYCwqVxDnK1nqRSDqxwUE75jBKOepcUkFa3u4NJrQi3m2nLhQp1bRgsaoG/UFW
F7OoKyKH9Ux6zUi5GokcTgO30n+pRclpk3OSLuqpp8V9LDzl98o4wkvD9aOwOhDCzsIfqE0SSUai
5AO8eYkWHmwxEDilMtpxNdHyz3AGx1Wb6/97DY/6DJjc2Qu9ir1zYuypzdPcfx8U7OGbzDbqVMXd
6e9bvaWdpiydxEG4nreyDknXpzE5plgH1OZ8MobmWo/PKwr95DgYX+wx9Vi2PchhqXoOeMY9pxHi
K23t6D4rwXkBYHUvsAxNDx8ngjHJXLh7UKNlMBv7PNipy+9nwz/Ol5rzfMN3TfUDwCcekAXKSFeJ
lWJPjtdVPhqoqA3yC5N3ZBdcJ9GNQi5MQFxHfS7mMrS4xCopgeICIFJHqw/7rMq2ueRLomcoh7ji
z/6VbG4S6fshAytN0A6bYD4AZeu+E6uvrpO9FiodchfTmXfLf0IlUmv2gpFFRRh/idY56gjRq8vA
QuLx8WprTlu9/CLX9/a/nPYM4hnGHI8ID/E1MFeTL7b3wZU2F/J91wzdUEtzkX1NhDED15wYurk9
uKIOgRJKern77UOMs1KtcKRyueK4Woh6FyAAed4uHhvwL2J8LhfJ1UCiwAQjQee3Ghvy7hHCZmKb
IXGxgy43PoWvRdy/BPjVc5mGw1BDHubXVP2Cns7i0PBAZbrjQlvfE4UlFIxpoch48gVdr/MNnUDV
6RgXIwoyAIRdjN7hEvWIWZsFNBB8eeXyzvJ3jZIuz6KegRcgowPdHXLlBUm7mhPIbhYzdiDy6SmS
8dL4Hf7lShXfiN+nAehZDeM7aULnx/4cQ0LxQXfiaIBiv3wD3R0yGJubkVqGKgNj5kKzMH+qFJ17
t+r97fxLKL3BmmEu13SyUhAhcWxBmAb1/5AIWqtLQ6sYF5Pji9vHiB6249D8gy1C86QLO7KmhBFk
WwNT5Lge8UXl574j6uSld/G31maxHhNqerak7H8m6ZnWFddvetQp5akvlFnRktBZ9hFDOFuHYRQQ
18Pv85NOmV0Jk+aJ6LLvdy+yN0jNUlYcmQTGWT2rYhM+dM6K8tTHptxRu4BKl9hWk8GJlLU3aJ6x
wh+qQvf3iQtH5SzihDVUUu4RaK/M9wa/3QVK+SOewBvazR0u19kQULEFQjY5GSEdqOZDo7uJt/HV
qw2sHquGk3XZiyPOem8ttwj8UQq/GS8noxzg43qiDJzRknfB3++ygryAj1Hq8cGzihB4ZDrLfTIH
dzG4LYQCCO10FzM/MFolzgu/lP4NZV9osalJoKj+ia+GE4lF2VXFfGU8Qmue8Er/F4pFBGtR7sgE
WYIQRckgZfdXkZMKjsIkCuy+4mWmc6lCI5q6xm3QmioGftJQu/xyzA1+zILr/fUfJvcqwbKjiIXO
Jx1mZE46+Zf4xdzzMGE5tT+u0KJK2zWNkS91WDoxvKnxoCqfPI0P+D+Di+hE9KA1bilI96nj7K6R
ZiNYxKKekDmDxDO2a10jISU+zewsBLrE2yp1mg6ry9GeZn2vJIs4xsJ+QV8JZhTCxOF+37O7aXtq
Br2r+1CN72CLWKB2LnQ9z2fDlo5XoANUX8oG6wvBiVoYwhP90dOYCP8Eo6MeILnRUfi261Z5mRBj
v17wgqmehrWX5eUCU/RaC7PJXqXZ17I3UD69PcWyVBKeoju2fb+/l+WvUlwDba5KDIrFgfbqEXdC
nlM7VYeAHnW2fZYFtp19WpvjLz1fIJZcZf4JaMLgGmaspRl3U2/yH63gVTsGzTKX6UXFKrot6FBL
I0xWpBMwfrfx+WkgUDGnht5B8lQQL7Elq7/s6KjatvxRofwrjt1E9xULuAVbxsCX99IPajC6kh3F
CSk2kME3a21nXChcfjLMxIVuKzRgv5QlTRfEdhAv6bOWRj8/yFgE/5MLo4UuE1KJm0/jIUcE9eIb
FJ/fm50CKtYJuu+tNAqwzSYh82/1LKjRjCl200x+v/tXfu/ZmxDNm2o2Ju2MVUWC8dY/P+QY8YBl
I+lS55BY5AnRZjeH70kgWiTVkknWGW/Gl9JRUxCQWx2pR/r75/WLoVbGhsBKIpU+I1xjItyxx+At
tqR1Uo+xceCGafjLpQY4TXQVkwQZPKjm+GUV6z76sOZ7unqIF16ZjeAOqRXW/1Kl6R+PW32hU2ai
OotpOE1c4hSDKvV0qwtzU364cEGsJ4iWkWqb4Z0TixNU/EKJiETfXjNshgOasKyPGiWtToBgjwOs
/eON0F4TNHNWrGihBeqlkHoERJ7l9zSsgTMGrGQtcBsSkPUQnzOFoMUsy5UkY0Ojlx7jAZc71OM1
LJyNBfEXwIt3M/37+PRr7JjABphNO+9KKp/+1tdmsGlK9pgSNM2hjVEIzThhQ2X3cZlCP7h8NnxK
xi7bQLqULSa44r1YdNyjbBrXYQpz1DRvxiTR0IR4yiQN/HwZu1P/uFC/dLCdkLhMASWCM1v/Dge+
rd1E5voz6W0CtK0eT1ekno8tTG67/1AAICTFqwWefhHy81v1sv6jOg863BabevSlwv+XtFlS186A
f594hff5ZbtLSZvkm7EmdGlXaIjNi/S0teSshlFk5zHzR2p6Refa+UQhG4WOuCDEQZeXGm4umaW8
lKZ1UJglajjo4O9J1q++aIArIwspDQlXpr+7d+sp+LQdWUrVR2GusO2HFJ1icdIOa/ObE2W5TSiy
j8PwDRKhXCJf36kBEV1cedm+EJDzjFsxjMziVAB4ULWcZE69blUWn6I1TBxo1RGYeIq+BJMyVvTk
6+9jUFT0XbwgXf8VS6AWcxOL5VI7hRjPnO76i080MpMx1G2LTymSLZLgIEAFmI23F4f2Mu2icAuP
il9FLM0y5iRY/i1mfusYjsZZvFcErOXktkWJX+EbnwE0KxxLKxYdWtdz6rjJly5oKkpqiulrLJBt
78NlBT+jZY21ivNonGbGspJcvWnA7jTERi+zUeniReXtEcD+I2uT6Ciuzx1eciCMzL0JEE1OtiyU
4+O1+IW76chnZ//VHncEmPnbnfkd0FgqyaulYYIcLEeh+IPuyM0EJ2N8Ff4de+TY7M2XpEaa/1jn
eOQ23oRlKW5A0kQWjUx9SUfn0AZ7CKIahJ7a61Y/v+UOjsxH3ckazgxjQ3kUcb+XA7DBZqcxnntz
y8p48CzlTcrTV4WEgm1oqOyEOC+QOyruZrasPEnbu+MJ7/lvirXmpz54k1X7zF3XZvSrIBinANK9
CQsjZm5IBMfnTndNSmGLmjUXj0gWRZPDntM4/qQf4jN8VnD9FTx0i7n5jk9M1xUIUIhAFEXrtMGk
IYXo3k6y8v8ayh8Lr6JADp44bxzgHIwOm6fmiazopuoXxIXWBdT6UoACLKt22zf55aAHhzNX9DfB
WttkgTAWf8htIhKxgtUycwg+X1wLKbGXBtDsYYF4DE4xpOHeD2tLLe3m16+rQt4HOQ5NUR7S9Ooy
4x2iTnuVWt1kLNjTqfJg5fR/B4gOZhHTX8++YnuX+Ih/lGBX18U/kvBiUX2ce5X615utKsWvx3+X
sRDVwd4B6YTIksNgJs7BsQiUWO04d/Brudg6bzD2Tr7UF4lmKA92wcw6z4VmaaC5F8WYFH/0YOhz
3Qox5ji07zGr9/2TSSIgrat6UmHnbhOFv8Q+Glp4Se3VYE2eHbBdhSCkB2h5G1Vav3fsOQPSOddp
+tTTZyYvYx43suw/I7nsv15sOMm8jlJO/JePqRfwzbWuxSFubhwF1RFRukpmHFg4lUKU21w+2EVS
KskueBYibT0YrgmHcCTFDxwUVzMQ5TOUFnEpxnG8PcZJn7LI9rJi25vCSJve7lMm4q3NVY/hgeYA
MmeE8pr5JAE9XqbLbQIsjoUJqIRlffnE2wWDQ09JL/FgiQG261+KtdSYhI1aY6XCTYTTxeCmQyEq
/3OfAgg2WzU34X2UISiXATxTvyX6VW2+tiG0BhIHqtc+KgL9kKrNV0oSZqL0jPMawtLth6ilET7W
JdjFZYMOE6v7jJ8G/41V+Z9oo+wy3c8kyYrv+5REL/1IQYXB3MVjLdAs/vrl1DTk3gE1cClubTx2
0yETYYNoAXMX/kixg7WnEd+MlofBbar4Lc+AUuggbBaTd8mcqLMEBkRuPMWboO7ftnDCl5xpnRwt
5AzalHfixaGad5iCoaLcI99vSBzMs40Lqlag6n85xR8dzIM7fTKqUPAYmC5GhsP7z8dDY1F0rEp5
YkRwUOZNvAxAvr/uOR8DRzhOhZSq+XnK0wSlz9X8MH9A3nrRIzVZCcyEUk7nMCgxM2/1s5HoSfLw
akvVhGRV0HJZ31dcR/47Go2BaCqoaY2HvrPVXbMIarkqmuxbNkUfxEpe8h7J7vQgFrT3oKmK5y7k
EP0C1Sfd28/Yb/vL2YOBhgc2qekCq6EAsy8UjRuJzF/ps9iJUXhWeE7zZpctn+GRdnkt4Dlt8eug
jNcIjAH4oDHAOAK4AkQ+cY5Oqy09zcyHFh7NBrJjIjHF6mqukV19BO+rDv9OmPz5JH8JHFXzqItu
60kQnXlHe7ig6dS/Fv5txyMXJZ5sDw+AlkIfSl9EdjpTIGZaFXUxq4HQnBbFei6lTa6V+lID2Yh7
YBKJ6xKhkqlUhzmbb2u7MVf+aoPfhSI59ATigs12DLUIXMqwhvgqHQybZJfYilEuLgCfzFsUKW7C
j8vuWp243g3JIiFdyPt09+F0W1Dqh9Zh8KnJ6DbltD7nsyd6g50+wnrzQhaRnzFsgKOLpkivYpP5
AsTydZnbj0jPp7yxKWN9QEB66whkAZBmu6AOCtB3Ta1PqaukZzXsID4JHzlYDar29Zq9+vPgA6bp
O8QcIdSVy0RGL8H+UHJ2pE9RlxA0T9BtWczryDxc6XwPhGsGCzBqPKNARkvK5eVnK5F6Y0oe3/k3
h62k2euHDTVLT7fAlf/P7oZgE4WwkiMKp6Yje5HdlQaR4K9MAbV4UslZPHWkrQ0NrbUFj60VMLbL
2zqJunP71fMJGO28R/MSJP+FsJnNeobbEnTvvIrqKSsEjSQy2oTr5EKc1tAn5caodpr9BqYdqOJs
wIxorI4sMjDSYnIJ0+WakvVpPx8UVY+hNXAmmbThpcAvxo/f1lcJWuTokC5pR8S6U6oOfc9iPJti
xC9HYAQoMgQK3JXHgTcVP9dxsdUwvnLaRTu3RkwJzgWZQVWpYgL7bGnDoGVVKQJpeQRFy7LjTLGM
ZPovqmm1Llzy1dAU9WpZY+JkycpzWHIBu89BH7gmDTZrIxrhv8cho3hvDsHzcnGJUV8Ii5O6lU/7
PoIKXnqZU8NIv5Hvr299CsrxCjhgHQXvgLzucU0+Hf4dYJVL5qPH4AxxCg2bF9eu5Z1AZ8lrENPx
vxuB8pmabI4x/LwQpYTPo1UKRtZgpRns9NSzb33UaTGj6J4paXtZIHzT2KkGq/8A5TBPVnvq5t1S
+ko5+66pz6ma+pOXIfi4mN02QZhyXCFBlbuW2t3Ta5rLl7SWu8O945YH21KoQIQGksrCzLyNJutP
nqGv1OVDqnGqgHE1cwrUNHznmQEvDFn8YVN+6f6KlXpbQ0UgGxjH0HvkFGAr6oxV3k/q4dUsDerT
Apy3DyH8TNMuS6rJmK6182gdi7WyFsD2nOi1bDcDdSmXmMGzcaOkVVYzcsQjUBxVmRIuJfOnNHNM
8KQbmDey5/B20s6Dk80Bm+C4HglplcP0/KUppzuWQjNAUjPk1VFALwe2nyQsCjZpBFh5hy1zePfx
QN6DLQrYJUMOyX2b7ZEjZLu9l1LjfGfMIfzDmTQNaVjk8OtLtw2iHMR1JO1N/+dGd1vnCSj9ueCG
ppLYQm2fEKMaM5kgSVMvjw3ygJIxnsAl69VvvbndiOko5Q34o00ZGRMkxP5r+y9R0l29Jm8DyJIw
d3Rfh1BmCHltIFXeKa+2xFDTQV43x21js20+8uEB8ez2wdyuqTknOvo4xxx8+x7eGVm+XG+Osz+m
j5GmihNXLf3dn6eANroERj7LTBA1cDgpxOHXcx4tTwWcpw9VeHzmMiRmfDQTzMjJdejQDYKtEUOQ
7KTPsn5h6y79XSfwjfg8VsbIYT0TzGP2rKbX3horMh5kB1tvbO8Gg4rt4QCL0uoulEDSeT+LycyF
8wsJ8ulJz7xAPpUM/1xwqxDBOismTjJ3nFyODW9bKQ3RmD8Gpx5uo8XtuH8mzpVmhzM0opY1ml3u
1uYH+6wsTJwXDbZd8Mqugzj4Op6MqALoWdkQV5xXA0Rki+zLIelp2b7B/4FcMyG5Wqs15Kof9Usg
yR3oodK5drTPBcp/h+t6lA+0U4vNQuTbb0+sBsgz90Mui900cS4cN5k/5jUn+Ls1ygCsf4mWa8fk
IEIOFoPVtTQb//gHiK2KYkpYghs/VN0gw8wNYvgFZzJNiupr8qti/dwW029cy4cKuUdrwiJWuvHY
5y/IN4pHUSYI/Ypfl0fgORS7Ab0g1oI8zjmXObzhrwG29Uth90ocyj88w3UdRqDTvSBKdQnjyAR+
8c4FUov6OlJiyjg0us/pcIz5OzcA2Sd85l53Ble/z0g6b2dKMviXCP8FqAMWkVfM+S4YPU5Vys1H
tuswuJEuPmM9ip0VjJd0xijSNbQeAemxbUBL0kfQHZX117oHIp+obRybHQU7o0h0Jls7Agoj4C4B
nuKMv/gryPIlTWyu2HWobl89EylkIrI0+z7cx7XXs1uWXINo9l0CX0BEnZx4iuYEYaSA44LI6pwy
blMu2v7Aw2I7IkeoO7RnD2j6dpXPpF9V4C37/ccotxofBfAOxvD2k0ztMtDxtXA5GJG57fmhCxa3
4TN3E965D6uq+U5deOjXB1jkC6lXvGEgjcyUy6KaA8AvmHc85xCTM9u4TcOTcz8cnlSHQ8AL+75j
x0r7yAyjkAaVRG6R/MTkeHzm0bSVzwmo8GOx75C9i6kIZLbLRoAAtM7aZ+qNDaDZNy3u2wSCDnvD
xtVi9iJmZgmR8f0Nw7kT3FjZEBxs7ZEM2b1lBjj94T8c/UIIemNSUaXCYKhqA5SGW32AxwArK+yL
FcVNr473r5jdyc0bAPblR0rRV3BbqWwn/SaH+qujObMcxY1qevCkINUKP8nwjVzZEvrzCRRTnIIt
2SwULMQewoLxUUuudKEkD+dOpk4Wr9iTHeGqJoe5ban/60InL45gpNU2wcH9m3ShYp0S/X8ngrT7
sbtFDK1j73mva+s6hNmcX/Wn02abby+w1DSvHJyEr32lNA8eqT22LlnNa6eLTxBVbxQNOaqRNQXc
e1KcADUgaMqyr/G5+UF5rfH6A1oe2Hf8iCmNFWv5ZtYR6l5mV6pNn5hPB8vfkVNIGMF1mPe0/VOl
9Tq9Pc12qwRQuurfCS3XYjZInfiKnO0ZdO//VmGfVuIg/+HMz+qtRc/ZcXx4BjwSkWVSIks1rl7A
jATZZmBE5Cn9ZuZC4tSW8gKVzCCn6qQ+5ycfJ8JUt20pzH5PXJqk9qD1vOp+8qoeDt4pkk6/il+f
qqYGBrBdAJluV0+o5YeYfJdmTxqWnUOX8jcoYO2Tnb5a5Pp+FO4I/zYnfu3sddJjLyPXQQUJyoRE
B/tLh2lLdccXqWKCI3vaItW77cyvNRj7mUO71XpuZNIBhLU0wnKQ8fVvA+3H8jm2ki3iWlUEuKRO
IijjFSjtiJuxYrrEXKKzl6f1SNmFw1sQUTcCN6Y+LWp0/XututUJLSlMYrp7s99jUEUjS1Zqz9mE
2VT7+Zdj0rXZdZ+/cnKLBSYqG2+EIGaq/hZBoWhB42Rx3QzJtkCSQqv6Bqg8OiICdruWoJSwsorc
vJbfWT5+xBezdrDrxJiMTTwEEeAMTIUK3w6PAW09o+3IayZPFeT+6+bwloCktXNIe+7G8+DCf3zx
lHuKVCe2YAqcHgL12lLI6J1cx8xi/j+B/Ynw7X0CQqgeHKwnS/qjf94npePwfocJ7dWXmbX/s6pa
02B6k3p6yN1hMWjnodyEtK7QphhaBG/gxocJ+VCl0OwoFtRCPZ4AzTxcX+CBmwgqnXvMucRAmPD+
95UbWOjHC9kXUjbPKnPuhh0MbuIwPX8cVd/dC66DOmqwmPv+/n4Yd2T76D1B4CpNHYi15PztOCKh
5S16EBcDnfjA0jX/aqNW284vyPrHy7NdF2OY9Kc5veJvIOFW4oNMRsi+5pweRfcrVo025k9QoNEB
yDQcDX1MpCSi6g0Y7j7ZeSwo/kU+/0JFq4XgjVg1juqnml22uMv+04EWJ7bPFY05FuManTwe7GRf
uHjOLgGpzrVIhLKUULK5KyuZVlA7NzCgZrp6BbdzZEUO/BCeSbq4zU1n0FOTorSurAETARoki3F2
qV0m26xcKqA7QHrPExFNsSuSxR/VH6QcuXr7dpoMrVXNvY77QuC8r7X4hzysPF5KjgW28YE3DUjb
NFfdZVMzp7QX6Zrc+HwguYuznSu7Y+xbdDdxmoHVqmnO34lwRHkqiXYrkjLd69OgzWenlkQk6a0F
Rti5mzLU2IW16OA8OpRtCLhmQRzRlufLwUDbAzXgkVispXCcyXQBXtFu4paGFUyMPBh+Hz6hH0nj
sL8A0Xj2A9Kp0ndpZNY8KqQtPws6FE86+YanEEu1MHpEPQREyNQSfcxtqnGC27xBUzU9YOKyDIRl
EHWL6ITvk5EF7BZRRWMgb2TFhkUMGgAKx3C24r/iMXh8xCwJhANMyGZh/7hb0uIH7L0+6Ddumdrx
EdEq4WOU30exoS28UvmCDvh31yDgZnvAsCkp/vwuyo5ccmhM1qDD/nTwue82pqa6+SxHVcOXjJql
/MXTXCMJ0mX9dGTtWZSPmAFTvhyBpaU19TNWh2HimH/7veP6FG5+8YVBHrjJihZvEmIwZqLuWqef
YadRjFR598NUsXVXzIgKb6dWbOQoiMmI9R7wCCVP7GDPeNZX+cH7eYUeUqEzMOJrE1Sv/074DbGV
NaVTlEDXwLLLzpds43flW7yEYznx/ofN8WkHfTWT/8bOwDdLA5F21LQgXK2Rpf8s7Z0dwOwzqpMO
5nbznQXaOEXvL1P8hrlgEzvANsN9mqN5IPry69G4MRec9NOqr00/bn0c6hCCDgMhRv1khVQEaSY5
pe6BYfyh4EOTDlsj/w5xCJstvZxsRfibKhr7TMoyO/aAPWqbHeIEpMqSLNTMavlZQvWkXLE+1Hi8
dIN9r3oMlyZXkDLUco7D+jO6f+ou5tBMvDFRTcHn5e0nWK5HubxyVFfAZOgz42ZgnFnDyUZVnvhA
sT+X7d7Xjz1ZxWeoPIzS5c86ZXC/C+CybdVw1D6qN7ROcwJf55tXbDoTL9Hh5PTLNBcbAngEEKVo
pD7+vC80lprp/cxny5Wxd2gczkJQk+KuN7aop+aPghf7R4j0CipNCdMlmeT5V9WomfD7/x1kvtAy
EWtZc52skZ/g7cTZgTty4wOw0fr4k/Sr3ilGswi5islgLUMmEZmW9MmIJsGAB7gw6mRxUNwyyEtR
0HYmnfdvTrJ9VRdE8HOM+x/coTPKH8d9h5tcrUOpDmyceZ3ho20L0B9bFGxMFYUQFf97binafNd4
lRvkYlau38ldK/Uuwe2P9HuJI+ZLO75iNR27YcWu/dqLCk554NvgsyAo0YdzCZI1H3TtseaGANBP
cDbQ31FL3IT8PNuR6vYfkUKVzRDST1NIhN2GZlnX50YuhS86+Sx3Ynmaq9OaHWfwiWjlbF61AnKe
eesK5MObDHsaM0Q4rVjK4ROmXSX12RywkmSy9CTg0GYCJk02pltAC6eNCARbeLozvDO0zS8l1/GN
nWEQO5mQnziU8aeu7VeQYYxizasZMmxpmjBlHiOLtEVMzrr1+Hz5Vtd+bsViBwYPumIcdLa9eUGv
oVSnu9KoKAGayANrJ1iCm/riLhptRLQxKZLNjgr4JLxPolRfUGXMxzQmYCSTulSBFquXY39MWwNz
a6HqAp9K13Lb9GqdlKabdw7UjxQKWY1XoL68oYvxPQLNqX/2716YAsKnX+a7kZkduocWGGYiOZ1L
dbDEhlURJg/gTjHvHf3WlpIfldtUxDNgo8z0lSIiUXnzh6UMRnIfsLbjvujKspLwH3eQFiyo0LoF
HX0NZg6/AWTnGx0QdZqvfmQeJZxRqpZgrHS1ovPDivlhyLap8Bf/eGRLlD/TH2une7DVmrwnzu+S
mGWp8PGZ5V3jRNdzMBNrWnl4hwZ18mHAM5bWkpNMBpg8O9uXz4gUkNmNfmFFFGWcHjvu1TlGKvvU
XoiRcLi/HnE3usK9g5WuoziwwXplpsgMU584ZrNj+CmFtPDt9g3K4bu2JxUoFKQT76nAJt66VtAS
d+0e6cZfgoonfEwqzZ7EBSf4XV8mWkcQKxOuncDURRe3f+0hmThuVLagepJtse/K36JkHefPBR18
Ves3SKTaM6imF63/iULeogz4hECeVgYPWJIkxxiapd4dVxUltqvLoQ2zWcGEqfzI1jR0RdF3xcJj
wbFV/QnW9xG5ikvOGVEzPYOejrYKhdaBLJv7vPL+XkATD1+Iny3B7M6ufXPKyHkLYftCO+AQE10c
2IynCxRdih+52Gdz/+vF26gkCl/Tqcblt8USMf9kzAyWhxMDjsCA2J7zJEg7y8hCs25cozqUSz3t
Z+mVb+OauTGqQvOX46AMLQR3TlnDC4YujQJ4c5kEpfr0MlN9bNw//rU1pQzjaoUGgGoPoTpnFG4R
xzpK93KTwO4RGlkCT1o5zDjW0APgRFtV8RVI8Jz+35Tpa4QIu/jlCNzXAQ0pDTmI7nR1F0nqUvRk
YiyRc4gAYjQ9S3oehCNgwjjI9ALxOJYHEi0d93zbZ4NG8iFLrCLI7EQqA5Gnsx4JSQ+UCZ0lCtNt
0jK+qjPRP3NdfsJnMzMlzXuMDhH7sWEo5fOxZYTMreQmr+Z+wGzWOmRqAAbVM5uYyGepVul8I0OD
TE9tvR/djQiEnRp3JeG1a8Md4rbL5euLbLigItgWDI7CXUO+3okVoWmDzDDmoIlAuC0LUELTKqN8
iMf/tjuaagg3sU3nA5j3XMtesxcXFaXozz806tDR12+9/Azc/B8cfQPQoSXoZH81zhqoCv7+R4sZ
K5rGU+QYlkR0E9vomSJdnSXsZa9tO9RV/paSIVUus85cbQ5rZaiyFdJu43Or2BWgLb2TfwW1pvBW
cGCfB16rDb0f3u3G0Ai6Gq3lzA4/CnQVwAmA47oGgTYE/1yYY8cePWwrTaULh8NsnUR7n3NuRmvw
bmf4WupwuTmtToMXZdCXpkJrAwiYnR4yrR0zZro5e5q+hGN4I7B6nYnAeuQ080N8gLEt4ZiHk3K/
cUymvsYYA9XVxwW5uVsa9tAPCA4wcRR395Q6Ijtmmj9qNnt4pCpR1CtNaNwcGsB/mg366LZATAv0
DQv4FFSc7iEZ2bagCbob1U8ic7LzPR7KakUgnnGqPHm5i9emQSZDn4H23iUMcsWnwhZTwwBpuxrg
AFLl2WfZYj5UPKepmq7/AfeAP1h/o8iWSy3kjYUjFA8dvJ4LCo/Hc+ULa5o8l/PLoiXRjERh9rzJ
jXEHRv6wPEmqbXXcCW7UcY61H29e5RdKpU+wQ+yeyNAgekKes7Q7a7s7Upl/efd5p8dBk0pXSYOY
XZNkSczXQxj/l3ga32gnlN/RX9FCvl69dP82Rdd3LrrmUu4NVJii7nZpacmMwheVAGCEMIaqpLSX
AmmnvRgu+hHnxwWxrXdh1cwKkbSni7ojZUYMnB7HurzgjUxsSqGFW/170As9oy/UxtK+F3Ftle4z
z/ifOWDaNhbJf9pi/NIyKS4jHwukq9ZwMjUmptnC3zMjEOUsrdif7cTBYnz9WwuNVdwwsawc0Bl0
5OeYG+yp3HRxeN5jiiryKLy45C+bh4ER+RcHBk6rUA2uq2bkApWfi7AaS6P4Rambt5poJbQKPl2K
j9mLUiWaFEfGoVj3OAvWGwc5JxDsTPiM9OLYrEzqrK4dISL7pl6QJt07BGC/lLTh/FcoWjsyNiHj
9Xd8SP+bDywXNxaYd2c2sLbLds/OezWVmgD1QNsDKvc5v2tzIq2uNoSVZCHZ4oW+PQ6IH8t2NkUs
vVJOVvPYN0zTkuNWK5KbjyK+PtezbjCbwN909Wy4ygSckmS9TXlTagLe+rOjbZ+COf4841kCGMeA
l31hnQ6fPPvqwymem8H66fKSSA7MHADXLkrld4QpzdLjEAhbsh8r/cIOQ9Sg1VgHfILkcSXNPFw8
F9mTXtpti/9Xx7TtqtHZoLpOrHSJ2SNSct9LvUuy3nPTKEUkpD9CmhkDtylChUHVPAavRhUCKOwr
bbF32S2BHV6cvH7rV/HP++oBXPwcnxcYKAlEOAc8+6Gzx93wHIqMU5LSGPnQnoeObNnAVSQcdEPL
wYyY2FwUw8RqMexW47pjhaV9xnqI8N4yt17+d6oIie/lBP9yh6XNfS6H8KEAVcJaLXaOaz+kcicN
b9YHQOI4pJ7QJTV2NgkAbmuASWQuTfHB8/R5xfG22giz+eTXvxGiDt+VOKklk+mVBcGLkwcbQ3/5
HxzqwYVCI6tmvQfbAbU42Obl+vlOyG7y7Sp0XMt8BoJ+HN6OnMwF9/0A3qO4PuQ/EtIQ64C7lBIg
NMQtlERbplvzgShFPWw/qkXqscbNBfaLYQJVJFtvmJrVatF7X1GNhKo2yzKg4bkyx+itxViYUX0k
nGZlBdlfe871xKAoKksjqHsz1cnLSo4UhyeOaFJgbIP6eQJY/VqUV4lfS7V5x9rEDDxhDxO8p6OF
DamOlEIRLJdkYztNX5zKzvgM+xDt+jpeIIlgPr5+ePCJ1bRjLdUewYoPlqYV6dlwCd2eoNu1gWe9
q3FI/LRmvbRVKHssz/OQRt4yb58/fHoPdJKaac2ptL0XX28e4qsPB3TlBNhkLCaCb4w2O5P8pKAK
V7dCoTyGpbpSQerZLaiE6Q0t/3YW0Jhq0qDwvYkhr5KJCaKhSKB4CJnw49whuMiFMGz7zfStZQC4
QrqyAGHDBMvYIKTnGncBQ8+8zmSUNI/p08nR6Uk3cgeqCVjpkMmwx3sBIavJqpCZAVDPWx5/QXnM
/rnn8cbjieYI+OuVq6Ix+SvNQqUf12lLY953PYIulgRZicvhAV0XvE7g/Ig4qPdnTbE0YoEAW6+y
LLCEiwjdiHpD+t0diu9sH0nsWs68rIP8agN1ndUreFLcvYdTm4KiN0a6+5pM7+Ll3elrIh6AKJyr
heTcr9EiMZm5tCBVr/0yz1edkWSluqGZpS0QK5sMbHWEq2JaCr1nwwyAqBIFywkr7uiGdGCt672X
xOv282v1kA8xQA+I8dHeYDxSNZLGA1lMUDWoQOaXWncK8YM4U8EKJw6TyVx8egQ6v5nq+llulldj
wofbtOBnzH9xluPPeu3QnvY8cxhEAn/hMec88xLt/fyePwHUUJNj1SkmKaEwP/DmVUGlIJ4wolH+
/sYXE7kbw8vkPZn24cAlow79npjT75pjl8LfZHAEE7+IY42/9NYLlgNljvZYaVSGws00ukpqq/gD
kHq1yMb6Msy/RIyTwzxRmbsDNjegEIwlZYghN1o6Tt3bwkqKDHByb8CVfKvfTtxFZ2v/x7ng4799
pRfP+2FtJIqEFn7K03b0tJg7Dv2T+tacvm0VqicaG44/iPkcFpwz4rM6SPX/6kUQd7k2UW0VFopx
y+rs+eaHx48hSEP30mB6tzejBZ/yGG88s4FXsvmSNzYezK9NisBUISHKMFqmgojMGBrjRpSqUsjZ
Fyyl1wUojHLumPdPj/1YDQz5E0WwTS9/hZpDaNWY/yvs3RUEbq3cOqMdPtEY1Ff17+b4M5rSOlPf
4SdPX9laDVDZf3BNUwzklXc+HKW6kQevqNwNjbqzs/6XQ7gslZoKLzH5zjmCwpGZYcTE1lye+6tI
YbPmncUbKvntQS8yYG9xYtHjZI9yd15PvFtp+c7lYcsRuMVnWhFPwyV7hquqI0kkEu8vjNuDEOVC
2Vt9DCU1dhmWthaUsxypGR4Wef+eRtaPpcw3WPzO1kFyw9accr8dQgJ6JB0Pa+C29bUevYlbhyqV
2WuCmDRNkSrYhKrH/KKwInBeNlt/mnaalkTLP8MmiV6Db/hG8vmW60o83lGS0LvMqrgOPogtzdcQ
qCoFKWLl48A3lLHGi2lfZvlxavYwAxHuCQYKWUT0/dF/R6Ziz+mg5TsaTJihX80L4A1kHliiZ5sQ
rxl52wtLTevi1lrJ6z0tcc3oNo2hfbZT6BC6w6bfBBU4OIClJwlB/Qs98r1jxdCoeIM1BhcScM8E
i+KwFUn4Vn7K2Td5STyA05EUAz4KQBYcQChmChgB9gNsFezIVtJSuRTtx5MXic7cQVt5r5/XTQNh
LvFPGU7pMblbvIEttVThQTtXTKMq86CKLHmXCXO3Z8KwEus64+pXTj3b4do/0XIDxVOuKn68hDYs
3jv0DJwghwIC/GfBqVe9zfdKKo7KRmGFaiiP606asT1bsyKn3mL1mGUQwIVIa3jlRTFA+12sUgDz
Lb8PljFLNnOGGtDqjeJewniw3BnPdbi23c7GVzvh5Zlhy+rzaK5DUWjr10EI/CNkYqgPb8aMyNEh
DMJnguT70XqWStZrKbVR9UfpMIRgCqsKKAbsYaozEeHr3vMXnu/T3U7KvrRN9pyV3RYjoHeKJlwu
LQHJ39AWiDNlmxQoej07EOARnZ82QuST5yxPy7UqK9R8NYht8aD5GKWlxmynyT26gPGSnqx4l2GS
dVKxp1tTxMhxaFD9d90Wjsso/rYYdU/9ZzSe1pYxXPfb3JnJXiNR2jIuoLtOEVbZ6v1pSyY4Zv9S
LsxVicSzcGa/Uit57IDbEixEqb3CJlGgCTcUybt53Pdl3a96rkBO9beyrpa5eJlBWrfnZzLwaN1+
kGfsCgGEyARF3mBV9CbUhEueKcsPO0A2kOkuFBOCzHWqnSUeJQp99mLLmk7Mo2FpPw8YdLKUggZY
HpDcN1hVhrDNbnKwKaxLwtu/9dJNwm8+PnX0TYd0pbDGlyDSmYAnL8N0ndkTi6y9v78DpNmeIq8r
FwuD82THefdBjEntmTYkATalcJJlHcV6j2neJwB51SeHpQGSexYBHDkWT3wvzK60NJ8Nbp+MOHjR
kLRLC2RGotByRm9oW5xzr7t39h2evxo3KeF0p5OmFv+z3NIrq7Pm9ahvMu/OC7PWkl8Lkjapi+PD
ALgbcITJoIGJQ1KRBd/HFLYFgTOyyZzP7j2kabRgyJrylIeQG9CvfDEB7x2CkG4l4nhg1DVIbnDp
qoxaxcQq3Dl7rS3vDdhkWypHvLEykODquDcF2Je3J72gCClJBo5jroFQ3sTJj6WyjOzWUZkgdlL2
FQ+gx5wliFK/7PNtP5xGGC4f5Vg2hRFrSiyf2JFQcl4ysM2+uURzdv957SaHh2cdE1m5r0K3x+tI
RguXxe0343k3PKDXc0vJzjwjSTbkta4hrarpvT9UasoTmmnTmnJAktCBY+RWw1ivk5jzK8hCc7tA
4am6P1D7bwBg93vO2vBLruJx2LaXTBOsXe5flgGEVPOpo6S/VeTBrrD3aE+Ov/mZW5d00sHgFCMt
19U8fW/lfCwo8hJIBHrNWUsPpiOgfbIWDYqp0uNUkj9gEwx2Y08VGcBkmp5f/Q0Jk/9ueVNgxoCj
QKTX3JKqGe2VNfwdScqxwSSH6haW9g6vfKtXT46dzPGKTkxPLPM/1akBja8RZIZRAlrWZJ8OSBbF
lrIcvKCokzSR4kSUvF0Iec4w4DM56emm2779VTccrcwMMPCf77KboCF3MQgU96NdpWRMvVzhWxXV
a+jCUGRFsvS71sCMiy556MFOc+7hc0g519xQisSzVQ/Wr7DZAQIHQ8w1be65jXenk0QKwx28G+oV
YR07BGURA6szG4YdvY3q6weEWkW8e/XiWzsQnsWPBNUkn25AWipnnHRYts/VcdsKXU9u3wDTaDLp
Hb4kaopuR+2FcmadTjc0XpqEOT3IY/YbfPw4wshVIkmbQIu5tzcqn6UpPZo1JGCtTFRg5VD3un1T
jZPieZ4wp7cExo0HCNjhQ2V+5OGDwsGYR4szG9ojSEMyTTL/LJ4AEYQDX1bgjEgkDgipR2h81lVc
evC+n36k4PQOI4XwyLc95Ea2W5LHWmCggKBlV96KctJws6g4wwcKwR19Diy0tjXzD+dK0kRWCWQ2
mORaiBIv0V6ccpFGqUB3HqvhBE7vOkPkLVf/NTjSCoqPhKNROANEKImqylUJqrNgm73dvTuhH7pd
p4F+OvPRRAtoxHHXkvOvFVA3T6BBtcQxGLf1+gdGJo8ndtKmXNBnfCnFaEiOnmoTp+zGkaph8VMJ
fwF7/+K7zmtygxl5PTthNLkjIaI8k1VKKcVokUZF9sRB5JUMlNz4WmsdJ0ONMFwEl++ZH+p2sgLg
qEpSa2NSCHCUevvyZW0wnSXsbMROZ+qNtBo42byZEMIzKCEYGpiJnvve+B0og4o+tWgvyjNjyFWT
rDTx6rVsWTQR/bJ3V5e9i7TuUqcve2uZICU3w+fX1jiCGINQttXAvDF8vBnSdYHIhAvGJ5u5swnq
BjTLYHNSBkXSqERW+86uTGokZkAvKP/n1QZcOXb4KqrmgEyaHn0lFt3psDpsy6z4L7WSpcYz7wcN
8sHR6ORdRouOSEySuyxFDlMU2ye0MqTMue6H2+lFDPWacW4XHADzYaK+PlMSYZNf4OuUWv9Glqq0
T5I93p4BuMJ/5qF/FZag+jeWxNy20CTU3UagIT9xUrv/EjSe2SbtgFMhwfl55fQcJzif6mhZR68P
7WjoQ5Do8fK7z81v31BHdxPjKZIFMECH1wbJap0qyjIrSobf7TvXkzDPbzRtfJ3slca00msmEvbE
Fx7Ni7ijGHF/+VoTx7G2OxePluhP6TFhcwgE1zSdVYVIPWlcAkToXzntXGGg0C9Cx0v7K6VaT7Le
le6xadeokbzHvNXusvK13vzDo7bNGxWhql42PDHsdhA1Rvk+GAkwT+vmsah4uPQXwLMFMG9gMwbT
h8DZZ4eJfWyJxSjhL3lSJUZ2xFqa2pDtoUV5JoMeoGvDaVI+LVrSdUvVi2FZKsbqp2SX8OVHK9vk
KJpS0q2MInWdOf5fG1AkzAjM9BVs7GSTG/cfAbiywLfHoVb2Xt0B7G9JQ6pQXZURrQGXHDXzPxjQ
4FIivPvGn3xndOd21S0rXtFMjX9QOlDY3Xj+77doMHTDh8PQWF/FoGLyyGFE5p7Nzrro+fw/han7
Qe2AEwMxy6Iq+f6WM9LS0YBrc1/8axB8Q4gRi5+AOuiW8TWC495gY41TarMj+Crpf9RtyG1C8elb
765Ukwy6Hj+Z7ROUat5cvYTfshS1+K7+MhzIUX3+06284TwgdzkFKfP3qP3UakMglAP47c2w3bb7
2E9dp/KcEg91AzLqNtZEhT46RFZR7O9KIW5RYPNz80YWnXZtMzNPFxRNnpw/6xqFtdKqKc2ObVeI
jZlSth1ktqLaaTKQBZPd4qmSIipBZak89U2mwmaufv12KdIUzIp/1BC2OdiPHPRqZMJRYoA4WcIE
z85pi1fQB+OkLmtUmYmb1WfHIReGLH9XnBQjQ1BvE511gMMogCuMdtEqNFX8O/1myMZyENOv7fZf
oNek1CJ1u4JpDhrzd43yTDDliA2/4nnbbTU9QLECU/WMDwKWUmAZCXPSeVq7ZIBPW5D30CRGO6WM
e1/CMhsRMDJGyBEoEQ90labNaAAvGsLyPqS6b9rwyvLmOnkZjkIAqPOFaIY4C1pgJsjhYpcSfBBd
aMZmx+vttVa6G6Efs8avAfDhtyOebPs5Jx6vPetJ/L31nQ57xAaso5HL9/sR5W6Sn+gOAAYErR+G
ekjafHBFE6L7/3/n0YwxuFydvIxFYgCjCCiXLzYBbXbIGXq4t9CvoTBpUBfaSF3WvTOniyifxveO
s7WMrcmoXgXSewD8jSj7eZqrWGk/0SIxnhAYgoyQO9RA7yHWmYl4lf04/CV+c8YXgnJqqHbJFMsr
h6L155a5XWniU3wiwpdWBgcfYygU8OZhs9FAGZO8Y3AaAZau5KnhFvLM56sCdUkcqyjCIGppND6X
ni/jY8uUTL8BpTq9fiwfXUOvs38frIzl4+aoud8WvAGJZwpEzjfve6C+1migB2WyHgOgfjbpqFZi
cKFimGnkbuQROtpojaCcxpW2n2cS0REpKhxLir7X4kWOteVYYymQrNNgC83/miAuY8qsN7WKcndp
AW0uXoTZovWQxKY2AtYVJ4Zh4QQyw/RWCsVFf8io0KXeUjJuSxJe16wQMz4JiJOn4IwmVC1J/oet
TSfZ11U9BA52Vl7n1dMgbZdtEFi0gy+K2W/pnpmLOu3iQV2NDSSslTtuvAGv3OlexqEj0jfXmY0w
/WkMY2vKmEWW0f/abCTJ2g79RJplr8nhGuhMJEWaXbizZPslEKD2t2dGYxI0C3fxTasjtcvLfV4N
Z6KWBe2awVP5mq3DyE3kGd/BDnXCXZ6WmbpfFEUCwtfHixGsPfYtJupT5NXQwN9wVSY+kzCey1Po
INF1580Pqmq/HxLcK31Z9uT7L6T7JtNAFEgfXb8edABwruqML1H216cFO0/pKFvY2SyjR4NdRNJo
x+z5TCNeIMh8gpt2+bKg57fztOzX+l4mPj8cqxWF2P8jQMnGV54ou2vw+7RkmhQ1iRznB5xb7viP
9NnqBRif6D4tBa0lj9YoPCkshEebJBQgJ/RF4vwQCvlsKyC/K9mQ31bBFaEAKIbSGcRSdQyF6zgg
aHWmv9GVG30K1LSVnY/w8k0eTX7YKukyfFXEswqh6Vyrpey3AYswfs4zFZTILZ+BqjNNy603eo7v
USPOFO4gN7qMIuCKd2Ip+O0KhqYblo+RLO5qApIhXgQ7AOR9auv97pFKPmctrjfB4ormf0vxFLl5
qSSJj/lZMFYuJB+wKMLqdMGcrBzPTIU746l89gmNiVP0U65oR9TBBmoaZhqORIeUNf3Pj9nyWZOk
8cdY/NGUu02MLQIQJqwScmVTa3BzJrx2Nd+Qua4tbdsq8GOIhuedApEgB4s3G1j+JISwKAY5jgxW
aUo99UdtMADXhKpi5aRSxFQEMKTzpPDx8u+hizOD7gK5qQq+DleatlkkR1/T1r9LXT2OPi9AikL0
ieFjBTUJQ3svzLAdeBJmzYq8TO6UvCGrb60/6rc7neNzNLG8K7izKeBg6gq6fqYzx/hO+K9oImln
Lqu++NAWVNhAmKVlM1rcvuzXAvnrCxCJq4u9vYrovRuTMGIMx9+2lbveIbfZqyE4FwYJeCtgnKqC
8GyZ6wprHO4rISgi1coFW/gn1Jo40UAMR++grQZAagzcjL3s3FLCW5gkQjKxQEqq7uArBPrDcfO4
90jBhCUho1uikjEv1/cG+8LscszkVyKkGCPMvieENwagYKHoH3y5SlqgbEUCIB6nhRqPH8DsSdfX
4QWhRlss2tribUEJ7dO3EeS6oCNvOjx7FRWsxShIYohhGJ4XXL7iDm/ebtoTNFdx6SvrtwC4GCae
A0PBd5t9+7h0f+yxiATWZvSLkW+laOwhKf5eiKQRD2RfBOFLQFXnJQDys1ezDaLDUex1cGcq24SJ
F0Kqy42xKwPySjVb0+MQSc9Hyycr9nsNwihpVtNhMV6TyMwt9u+ENs4kf1PdSq/vZ0Md3TWoeMuV
h8Z1ox8ljPqlJxfuLxbHkl0sDj57hW5ogV7/RQtoWSFP3KrpEyvSavFoFhJpc93XmR/h95S2eqV0
ihjjRiDd93lc3v5HhdcA78Qk8s8B+zZuIa6L+xxIjIXcENFbkp1ADVbKl6Me75TWCSYjfqjoVocI
o1UWPcvGZZmOMjquVqMowDoL362XbLhDDcv+oxF/AsutYqvwvV3hDXuyMGvEQ84iqzbnLxjrQzKZ
4m8J8Nw1KQDoCFdGfKr6WK1cva+rAEY3820pwaSi2L5To01UoQAwCRFyS/jPoYJH2vNw3+/paA3+
6VFI/SmX06zXz63P3iyJZ7jEHl3Vu6hFnyO63TzVy1UWPb9FBggDucyqMEG58sVtkCud3lkyt1LN
6cuSwo9CTK8b+FxEHb3S/fEZ7fk7G6KwIFBAp1+gTOdwMGPX1N+PI1sUhqqp03RRRwfQcQABQsMU
H6StgdlPoOnJr9AIzITCy0UYfug7C0ruEFidCSILbpGiXi2A4aw0d5QY3iW9bnkv/mz2CUlLhpkx
btg+7IYdUjh78/rJy/nT9dGnCSwF3LNOnfnHnrOvOKIY27gA9bE0p8iQN2iOj987yZJl7ea2mpue
WkhKeU8Pgm1j97Enn0Mqr+2SbpCMnHT3faef1YxyA6XDkKY/q7p+Tc998K+OGtOrgyf4lffncthy
1FbH27bp7zDP6f75EuzUyBYUWSbqPX8wZWG2/GIvMZS6Wfy7mWF9pyLz5B3P5bjKQEoKtD8C5bRS
fkq7hIHVLOWxJN1RBqsiTt1hhVnPXRKqOvj+p4wbf6E692J6C178fJgsKtwsaXIvjUO3y7faWKmZ
xKyMIVzyEov87noK7ZGGCzGlkLXTGYaAqdamNop8aIJGKCrJ9Q1jxAYMGXKb+FUYSfuUO9Fys/Tv
9jBMteUMrEA8A3Dy7VjVSpqzP/6O+02LF2y6lhw7jp/5I3Xl3vw9uWIe30V/If1sj0h7Z1AiWP77
lehutFMyFFoR56fyApbEDWIirk9Tn22JmxeD5veDFZ3ywCW+jz8ErZ+jskunGMocENd3T0HTnrtN
4aBHH8Irk2zBV1ygdOTLtUW4xycVxfQg7C8CarJYkk5k4DYmp2zBP6DIL3ZTfi4E/886YEgXDJJA
gy8GyJYUaq+IMdk5hgtgQ+qNEC9yKrKhpG7EjwX0Q5ji3w67L8/1GPBe2DVpb1rWch46bB2o/a46
1sJLdhgCBAa79bfnt4Rv+K5i1Fmgo6M+h6D4V00EKSI/DNA+WHSyPCnpyszcblPRC5IDeECzc6Y6
qanutUymp7XAcmgE7XSW0jB5e++AMXBFlBOxfeD5gzSRlzVnQKoretPFfxIauSPILtx3w86ZOpsj
iEGTSu9vwy911V+WMS+wdxWe152yBSiaHMoSIsK8TpReHhFeHN1KFGLGtgBQEBMuE1IL7eetm2rU
RZMo83enmGGbAhJc28wwrdNxiwW6iuFQOHOCUeXZzMGWfCC8gdwCUX8AzlsBJGk0Md5ukLeNvnlL
9YO16vhXhLrMNcCv84MRAgAK2XxMhfItyhYUFYIQbL/SjYOTSZv73Qs9br2o31jL8QFdk0ux7EVT
lDBev8LNVocHzMTxcKJER/bMDQnNvBUe9wquI68ld4ZWXE9i5eW0DAurGNwoIp3omKzIvTnhm6TM
00rYZr0cc/cwRUBW6Fw3Pjwmyq2Fbshxoi4rlkTM9abQBMDQxW+qYOBKwhh93oGrq9pkkOtrF87c
jYUk6UNC5/L6KC8bK5hfnFKhVmJV9pbxBa1+M7HHiPOHz4LabbClusfW8bTWzeX4SbTq53bbEozd
fJhIYLt3r9dIYTPMVdFNVLTpDoJMJRQkSjnEhjWX1bzMOsphO3U976TswB0g29XvKjjvhZnTxdDa
oL/dFD6Lgy6KXr1yGNo4yjQG1Yx92M5dloe3PxXBEQa4rJNqLG1rO+y2gNoLGdg8QwlE+cihgZ0h
3AtbOMSYxdK7l5erNeYUmWWYr5OgAW4IC8zOVJbAAvT0boOPddymf4xNzQ8BZfCvklqCF6Q/bsBG
EZNQbeZ22Db1p1tQRmQN5HXJwLYpoGEzXOhsjh+HbVAWQTVf/flPHX9/5W0SjPItAkwkaaIdgWj6
QfvbG5zlViCc9cbSdAlE3ulOWFu8/oH4yI+B2RLb3+TmypP4YdZVg3JWmQINmQ9/IpIy1iKPQt2m
nvGngvFJUWl+Z0fW1WCUalJ0q60ruNXjFm4mHqY/T5QO02SkFZ5dBJE6mqC54i3xyTCXeNRFTlWy
DDFdzAfPV/8t2cm2nfh0CvXdN5Y8ayfp0Vy+FFuK3kUSwT62MNB+bcT0fyResCYT7l3IVu1yvKBc
/C+HDUxLQpR/YMl4h2sp12VG0a1Ei+QL7CBgy1chKKm6UAN7K6dA6/1xZ5O+l/ku9qJFPXrKeX5y
PwqxFRSEIhV62HTdM5R1dclTRlvlw8tuvJetKg58DVTPKobMJQ9SlS1DCoKhNjGj2tSkpHEVbIis
Qzohd5Cecgd3EzTo8gqZ0ol5R5GShHKhid3nkwSvBegV1wmMTALqyEVVS8a4baUE3s2cwfjU0FRD
1JQZoK0+5YGI/KotSYKp+YHlIabGTF2mpT5icDfXXRVJmav7bQNH1Xp/fscvefqc+sD4aRl0DPL0
yl4kQKtETN9RtGaMkOgvtMVXfV/E/0cB99DQJooN2RpkKFiFkczoZspOvlHji3KvhfNjezaN4mIa
q7AnPbA4nEmxYWR68k63Xk8dXaHF09I951DVdMpj/kfdm/QJYivXKShDfDfcCnx25dfU9vbs8sFl
bgQ/Si/zqQ1P79yHQ7cxA90WzJpjF8vwdjKExrd71B/lvwb6xam0Q3aYNsppw9GfzYcFzWR7IGNn
Ps/kjmUKU0L+9Jeip2Vyi3boX6JYaL3dXpUnIH3i0D5NtGz0KHkhZCMtbDJI9UiicnGj6hvUw8Ux
X4lENRjs1WWgtpQEjiNoJqSJScK490BXZqBOtfZn8oC3X0dLLFiOmo/htfbATiAhBta3+hsQTZei
osKOWV3MtE/Ov03yFyqqVAfhceX5j9w89Y+3KGYGfCjI7oSrRsuF05EUa9QsdSPrbjK1QifqZe/0
dtX4rB88r+Lcm2GRCLV/QnU7zbyzvZOtPIodFae9DqNtmJoS5Xi2URTmCU7Z9VyismqiO1iWHeS8
KTXgDQplah+MzXFNt8vbot4x6zsDXeGEQJ86FJGD+f8cEpQ/A4E8y8/GZLwjrTIyVRQR8FWLS3oe
v2mVRqQuiK/Cz3nKkaM6b78FYfLZHyDlYppJfketwQNB5zoV7JrWjLV2iH/Jc8X5efIh/wFoLtYl
SRrVX8OWbr4GbpAbCdBBBPNzxhUL5zNyVKBtVz/1j37XiX6AFmzumLHyL4GCXXndQhKeT0nzUNrd
dt+8Egmpeebtb+oWubRPAF+DDkHaY8yWKpLXtfTb/JcbXZvkx+eMuRIk5KpobmAdieqez/8ScQOb
v4wzigqxrHgKjKjmij52e9P7fSmDAdI3Y86NgQ8/ZVibLbt55gwzq2hIMT5E8YVNs1KJlP7Am5Gc
1kAsl+HPZtF5w3uj7uerGohgYR6ZUgpZ2tzEViPU8/xoklWcBNvojGwCY/2w/QknAkgvmR0VHhU/
1ieKNsBJYpToRbhq+LUwEIOp2aVZMK+BqhTDyl9TEi3OszTQG3zwWgwVoUxTGn7SRQ9fOcEa81ng
ZEMrNw6d/HHOwhepouS523j/R7y1mAQHALPCoOATDYFps5bLnHWzXqP37lPLyyKbsJTUF+GsOHd4
nI/Zocl618b2lWPjDlYFgcV3QOqhAFs0mhUYvOOoTEjiMATWErqk8AU2BXbYe4DNADJWPhiXHor2
oCnTEv27zOs7i27Wbk8K5DquhqAu7RQkn0QIpKVNUPXFDcGGmBbIOTUcXaXdaCtrTmw3f8uAsZ0x
MtUJDhNh9XEebJGk8sGL7Y4I8We4Mx7B8jazLpJQW/Joe0DMvT90vP28N3TWmKVNWEBjU9Lybort
WvGNMFPOnOoHJA/1Spu1zBh9pkXQRriEmjzyvuHFqd1E2KNRyRC2JsZD07nRFg+Md2Z9eA9ZMVsP
/wSXEcgg1UODBlqtZt0PO3DPWNm+r7PUu0cnwyG9GFlP5xGwvSahpQhBUk1KOR+Z4ZDCj5s0uwDw
B8Ap2EM/V9CwYK5gkRK+F3R90HxuoLZ9OuCht5i+zLQYw9GuYKXhmp4naIX80jNdNhpSudFv5GXA
gE4avAdxPBX9uCzzN6Okh8mAHN1GufTy1jvPOtAPPvvNaHyP4649nLvRX/85QQVrbEVQxZapuYIX
GxF5vlD5/IdSSrR6kns6iX/Xl2Y6/PsSTU3oBRjw8L+A8Zwrx3xGrmb5pWNHgkqQLNbE1nWMVPd6
hHIPHg8UVrmw0EkWs6tMLajZ+p+96Dt2fgYWglTqlgJfWyxOFVd0X54LUWtWENYrNNPcS5K+Egie
UrZCHkxnj5Sjt/EXHR2HO+NeNjcoSW8Z9L427rQoXi9zx6Ynqmkfb7U3w+jYuxm91vcoLDY3+v6o
jZCGk8j7BdDXIrtMcGnKDtsqQ135Nx8r3rNmt1rNeR/zov2x4+XUkC456X+lBllzO8gf6ASgnAuy
uCPsnZCq/V3x6A/YU7lbqBY9VwjiSsJRxbbjUkFmhEzdELI5QkYoVfLeUxlNN3l1Cx8Ex6vvZ7Pe
C7RANQZBfX/bRel609x9JtX5QoDn14aDwu0seQwb7Jo9eeylSeFfvT7nUgGQPg1dRInTXVVvNjjp
QCvkc1wpLuQl3Sm1fdNqvZXmCwqS7JayutoLSn7rj4Vf7i5Somr9F0xvgtVXc11BBAG7F3ZCJZTZ
DAUiIPxWDzzPIJEn/R9p0pUFZhghdPEaW0jKPRn5rrRUHBxseRv8h3+ZM1EVsciw6yASx4emGgoM
/fOl5b8Wga8Aqxm0qNx/y0dDoa6+kUeqAvpEUkK4Gn0vPWS6qaVZfcurclK8nIo/Do+9XkB68iCI
nvJIsEd+VHpW6sllKyJlZpcItYOkVhfxqJecFLWQlYeUqZqpw49zttcQkjEUn5gODhaI2RsrhD6x
SW+STH06dq0g0apXzGuM7rtb3aGZgjXkiWDd9ER5jZsKE+fCz9+QbB6aJ0/W5Tt1x72pQmBTexJU
2GoeYbwzNbEH/FiVbxyr0ajb9mPdB8UGr0t1o/GytkUsQS8khCrx7Vej0ZcLqqqpw5YRpyRrbUWV
/v4BVHi07DjMLRKnYW0ERSZXGA1ijhgeL23b6VuzCdSQMmOkN5oXhRT57K+0+NT7iCNcZlz4uAJH
mJqlOKCOt4Q+58LFPuXgOiJZWmgUGUpN0WVEhplhQ0+W3FLtwRghkGFH9sLTjHGh4ts8GflPR/sI
qVv1tAvHHLyxfF8JB0/Jkosg6xyapVTtau9lBiLeNXfSak3tAKWLowlsCYxSlHGQjF5mkJTqhQvu
4rXYcDxztAwWjulW2q0Tk0yyp6h09Cq5k01H1k4+2szlglye6wy5oOhj5Q2XXMS5VgHrFkZLJxDb
+dzJtc491GWcm1Z+MXj9l6onfwOOHSckrSTQcuHrFmo2RNcad/sG7VkZ0gzZIUP76twSxljD0mdf
Q+p5ADTqWG+TwyT9jcf016ZcejI/GNzzfGyX9zi0Gy+adBIn+G6ntlSh5PCujeo72S/6mxR/IhXm
l+SuT32o8VCpuYBFWumCUCnFUSfgz9JDoFL0dnjbdwGnXHZS3oM5E3EfkQrAQ58tEPVDa+wunT+R
kNMecJJYK/zRHI1mo4GMeGbmZxw1M6QV4dx5PgvEyByLMJOg0VUxi0PqtvjGPe0s7+ONqHs6CzrL
dSP1TMAXBvS5ePbPRvoHrUZbTYUJ/sIxN34l7Kuzm7YD4TmSvYBD42TtFFdOglZrirvjFuYyFOQl
fVepSNmJKAGMIJDhlYnoSvROwFnU+jJuwF07nbvhvOBifYQaUjBm7SHMpzLsBsdpIcVB0NrsGIIX
+HD2DJUCAHDmTR/nmC7dAWQ4ubcbHtSJNxEYGrYAHiDFMXRCYvp0GPos8CuceTSdzF0yqWeGdt6t
EhR1o2crfvLPwsl97fOb6VEphUGMsKcdyTq+HlDQ6Fjx0zkf3sUQFi88W4bXhd5AsK8N6LT1a1rn
rTaIEgETSRBEuLjMLgn0aGnPca45BuA8g7+hOJrSi/YwPvypIXh0ese6AKgWNxhocUCix4llwRiq
yBD/uJDuKeaqHLf58rmRxrXQ6jIadvUxeyXM70hWMJvLhubEFbv6u5NyhjhXmQdYRUVRktks2HIt
Sq7/vWpDbGKRtYOH0OrWpc3Dcv6Oe4gu7ofWER9SrCFYe7Im7YnLWeCzTPfdV2ppFSVgAdydpJsA
AuxSJfF1Dzcj+paQNveMyZfKeYmipOrr8UWmcuIWZzpTH9S8Kiewmm5TLSw5NjLQAebNoCM7sGYs
iLoNICxo+4KW8DpL9m+gEYH97D6NfIzRrdOyB00BaLRHL6c6VBJTLWEOi+R0oUV39w8O/FBD598t
n/pTIlBa8e76A1CuVKFTKYIIPbFJJoL2cuLzJAVuaX+DjU8OTvpJ68K91t409/Hy3lMiL0pF2hTl
plhJLJ5V2ZeEk7ByJlSwEghddY2Sn8BMyEwPoLNlvvr74p08ZXXWKScGVWGd2tO8C9PkzFmjssfv
NheDxAMuV+OyABc/zCNQE8isubk6KWZOoRD20FFzhUZ5/rud7t0QrScdD69d0S2tgFkX117UA/gY
3mlo/Xp0k0w/vIuj5ZmM13wKgPInQ5Gj2g6j5UZoamfiTbzXqPmpMCTtlxyE99YvCip+FbE5Gzs0
qigSCnquheAECtHpVXNlGpRaCUoIHZQpEPw/yqBqiEWC7B8pZpJl7uBEBA/MwTRaiqxFg6U1sj2b
r3DhaigVnc9313vojTDv0cMAtCDHyYNJ0ck+3OVkFl2umiFLAUo0L5MANokrVn7gNaFZAbyKIs2I
MBolJWLjvkJ6HXEccgmhUXqpIoXagZH8B3k/TMOIXsu8t6s095+WQL8/cdxIPYMw/g4oiUUQngLP
jYyx9g+eQO+FVd9KtlALHVbVKPhhWUlriAmUF82HZ93ygRSzT4ImSAL1WMq/HwEinc3XUz7NTC+e
+2DjbONKeoqglJjQ7yzy4KwHUJD6pKU2zcEmvIr47wNZNzIXbR81OW6SiegCfIFkc8AmXd/pKl4v
8c3WzLgpllVMKR70q4KOwPm22UeqlehhwPYmYVj5xjQmxdeHirzoGcMOWKQ2Up2y4BfOBlKu+YUS
v90LMMNNCQl2IJLYxdD5x96mfu8ZXOrQWvEciBLORXc+iingzdYbkInAoR/7vPAd9HTfPpdpOOsp
kG9m2X/6WHUcGLwWZB40o1lBFkfteMwVr2960VTyeS7Hhn9cW1vWQ+KksetEAu88ahbY5lT9aOVu
UNbUuyOOCmi1bFEW9baIDu78UNip+8nQZDWTwChko9GQbl65mKvZ7GyorjXN1zJz+tRwS/vRVY0/
xdrcG2wimvd0yc/6KBpHviof+A04iqCENpY8uchSa8lC0uaflSeNE2YTQEVt7c/jADJd0AviozU9
Ysi1LIZnq1/oBtCVK3qWm+lW7jbF+id+6EfjDTYWvJGZ528Ijj6NdUQ1UCNEf9kEWOTfsCTmgNKd
FFF2h/4lyiPUZZET+GPspjJQkWQmwLp63hRVCAbGbmPS8zr7opACAwx32UENJoMzD7A55hbll/Xi
Js7HVM4vVJq3XCDraX/7gTEb4+j3fZRMn0XiaVFDyy53RDDXs9L79BcNUU2wl65ztBiTu8dGLS+7
ooEG490RAOIzDFScCvZh1hP5n+3wwW1fBDy2kdpWrmNmOSp1ZuOzZk7TRaZCKFpvLBFO+E1JCHEU
c+bdHhb96JIvdm7qzankqdqBwd4gX7fwNRN2wjx8M8ujFrbElYLbfrhO3J6n/K6mQ0yHb2CDBwkR
gGPclutaePf1F1jOyZMZK4/M9P1+k2X3rIa52XbM+Bi3PyW/Hy1VoRlPSyx3OhBAklQiXGQPCTaR
/RtTOO9/aykP8qExWjewhHD6m+yosMwThc0PoWTehcZ14baMa/FX2be5fis0OucBtI9eZvEycXfy
qKk4PCuUOq0ySQ9+OEX1xV7piskaOtCKAF+I6dcSq/ayWw5FD7sVXBE6u6zeNSzPzZMdZt6tgLmA
gFM4JGix8PP0jO43WT2nQKq28o54J0zT52R3t2ueVFFRBmkPAk61zkmsuCrQMhmx8mtf0zLG/76c
znWhEXKCeciPR3T5lB1lXe9rfwTxgDxpOwDUGhUCxGatYilnqQhooLkZFREskVp2o+07/Rm+nAMS
EG6ejTgPNzAhtm0oZqYy1Qiuif3ZL9FWU5OqB6SR/hl0NqMaWkKZLtkc3OIiHUNK/lTscvw98Ni3
ztgMNlNrbX98uqZwdccZNssIep/UT22qpNObxLwiN4WuWBdYghyE3rpqmRp2hxqiYXMr6+68lnN+
vV8055nliBtiHCKfcmMH6e4pRXYWuk1m1rSpK/8/LDQ8eh97MBrCGGe4UhQaw10rgrHw+csHe8rJ
YkR2UXxLQHR90VUo7b6kiMrEldRYQ6JzeAhF1NnA+72f9Y5/tUQBdCi46dXLFlJ3pfe4/l/pIzVg
ilCUQjqGnWiRbfSB8C6gJBGF8Y+hsUDaLxA46aGUGhFFhj0/4WGkgZWCE7RUQ984HZVS9TfEMK2T
RFBJ+0hRqhDGkO41pBCZG3HJUKnfl/fnE8t5XFnRcJFMYElLv++g6RdgVfE7UHJOkV2aelYbRYIQ
eULttSN1rTZpwiNMXT1X+x2W+MyOM7ndD/o0ka7eS/9bK4awrkhHYnjoM23673Az4d4CntjeJxcG
j9rcwl5onovO6w59iIxS2itU2DCChQjokX5dREqsUpUDrdlc/TwYj61slP16Wolp5AdgoScX1eaf
OKIX7gD9/hdTDv3eslg+z1GxHwsqJsk17TZk9BepA7TRJ4UrxX4zHfQm61MENENvCtcmX+iOVlNJ
PqmHw8qdO/wNXkkKyiJqpc45VaNEtDgG0EJOhGZ/3FoYvZb3gYG4VkPPqrwU7OTORT29OW+sBFr2
KiNq+w9Skhznwh/uby4ZD/6lvCVwJQ17q9pDzKQYozXvBAh+IFRCv/5Y3/l6HA26X9PMxB2s8UIg
CO+Z/hf4s05WmA9s3CyuN5Hel8y1qeQsqYaU4lAe5OHLPDHftXXbli9Qd+0uJzRigUbb2n33gG2a
2UVjgfA25YaIS7GZpoWSn3kgWMyaF022XBBSYqEnS77YnZl2VryjHgLdb7hcx7SyeCayHRK+ggLg
w8rukVwPds38rvhAK0cWd3Cde4GWF8mD/KnyJXL4qA7J5rJvu3IqLbvP6TTQ3vETDsKAlP6/ZraK
pZqVuMDQjWC9IxjlBQBteN07jK2s4I1SGwJ5B/DxXeEHcPXoP7LUr4nad8xt2m3p8hUY40Q7JnJa
EUfrXxKIMsZLn630nNe1vhs4UiTYF+t64UOyVq/dBFOKZiwtVI0Ef8cykM2PTP8A1nJRK7rD4Nvi
+ME6q8xulopUYOQz+fR4RCvvli9nBzXjRhI1aZIFLmz6vVFJuq6jyje611MhTaG9cbbLK6Pa+c92
8DPEOmYJcIToJ/NI3jKBdJm6nj5mVx4ErhNkxQOlLkrZv7xr4TDGuz0Dw71genl23IMHtPjyec2J
UbwT+7EGD7U1RM0FQgVjutWA2jyOvMi0amsgo+HE5ygzm8jVPpRCs7y3Y83ug7fpV9bi2eZQI9Lj
52PCGRnk9z+oPVdxRznSL2/nEUCpetntioeC6ugESz9Hknrp1h4Zf/RdeKyXiYwQZQ2OSDB5dCQj
070yZwu07VaXJwBUAFgKX8F+mM03jGMlXZY6zTS4YSKJVXTKVO+/71QmvgjLnfFEzcMojpAZMjxM
l0zKQ6u37OudEhRwRdQEZZB1O0i9Htb37Ibnbsclq0sW22NUSMz+haP3nAkgx6BIuO2B73BAdibF
V0dMNauCNYP8yAj/GkIRHTFM9fm3zqBNZDjHkzKR2hanfAJ2e/NMnWWBTCmBCyweblP/3CHtiqHZ
TJkFjVqX3+R4CzbLYuf8/YIprzmumhoJVl46OaFg+GXo+Gc+bEx+B75BsFU+FNag5L1eKUnM+C2S
ujQa52o2bfNMX49sYIOQxEr2KijmWwpacM0mGp77OyBvekB760sG7uw2SZ1/intpy0CBpQroNkUa
JU5ydeFtHqzA74kYGINyREm1S0C+UPTcrbiSkcxTP4cviJq4ylefjOqwDXbRWJSxom36FtYE/qHv
TMSM8e0tNJS3vm6yAwa8VhA8FDVfhAwK1yrzwHf58WT9x13F9G+aPjCS/O893gQ0MTFtdrR3LcI0
cjzIMn5C2cBB+vmKGPMRqQehOif6dUxJH9dPrpaT7+KIQ9p9OTPapiuampV9+NdjPRQolhV6IwBA
gSQ65sWpMuX46ry/r9xMkcNqZbxjTUKUX7Xg72Kn96BD9F5E+1+B268cWyIJ5kx9BUxamJqP7fWR
BRhH2gnX4HS1pCSIHjHV8R3ncwrVicel9dSiL8k7We/I+pTCORmB39LCkHohoRqmkJGMKCgcYbCx
l+MIezEaQDy9WwYPAN/y/LGyH/jGEl3B3KZI0YuTZm0WzTrBZ30/AgGkbUKMXjpG0oWlyK5Ojy5p
njesLz+7sV8oOJ2+rT1KYJTFKyd38NpS9OMq8Wh2llAZGn/Ekr5KRBoYQxY5aXeriTle7xJ+bOQN
vsZkqaCzUSqlW39/5d3FSuJbjDaB2Adve7Cq0E17XJ2O4xtHoq2RZoJ7A/UbCgFn5ju8SwbAeAAm
css6/f9lFFy9b9hs2kGhUl7TQP4z5jKxAI2MBd3nPKsdzP+8aGqkQfk+PYwEIDC+a+EjFNFYkkSm
jzfyxOSG+ZlP7LHXWeWhdmGw5A0ubkUHLB+ZCzARJLuslMQ2HE87rnPqgBRSYYSLgLumjuVLHIW4
/lKb6/Yp9mfLFEVJ8ZeIfmZ0dOO1GrY85QCf/seDAwU6P2HteUR2XHD83+6CtoG48ORbUXDe5c5s
Qg7Fp5OGfAJWaGFzYdabp73VQv1LvlJxRfvv3ZmEuVsdVPczzbE0L9EOXBWfb3qOLb0AV6Gmr7g+
XZo7m2U8fIAZHSiBB4VCkLTNt7uVPvVWtwsAOpTDWxk+G+8K6jNv1QSriZrJwDo3e6OUJxRwnXmB
qdh7S8n5xDsFzBHt9KUHMm4ChZAGd2aQRCvkSBBw6I2Iem/h1ukAeOEVsqwaEmyDDYbQ7DWp1uyb
3MA0JZvmRUXnbYLJqosZ1tf/uCRQFxjOXrPBPe7pG8rwbrsNL/f3ZwP9N+dZ7+acQIsBc+PENCjh
demA9n6FjAh2nTvOqudg19/ikXEhVXU6K3iark38JFl+ESY+UTwvfhaKlBYs4onsAxiBYjEvT9lB
m8N/wy1cPdiAXUZBInFtp1OI4+v7EETs32iv1nMcF9B0eJsng6sToyPPdLkyh1X+Kk0giNc1P6aO
RCJ4MI5VDD5c8RV3e00WK1Jzqzepex0PGDFjmRhDbmu4+p4q9l0aBbFnlMIpRwah0XxlvIlFdGET
F4IcfaBNe1qHXqnZiatu+eHplMrvzT1DMWaeNRMRFj3WPu8cR59BIolVKzCFyim3ujqU+xHz7go0
M2KbPH8DFZaBM1LE9xAOj3mHJnYS1EoUKfDz82+S5wY8we+IaBUh0UWXqUATb42E9XsvBPZ9vCx3
/aIZsZjZKIQwJ0cef7/YFdcWNHvAGn7HfXDVFEieQydhf2tapEhiOduEx4LkPNEx4GrYffKHsaD6
K4kKewr4kmrKHJwsJawBkkTPZJ6+nIttgDloEhSnex5/1+nM998igFpZweZoiYlqKtA3CUdg2hg3
gdPgMWEqvE/pb/FvMo/AhSBdA5Gv/PP2kcZQX/GfbVNFKKA+p+etD84pm5p0jxrAnQDh5sa7NPie
q1Ds/JR1S9fxO9iiyY8FQq1OXYK9gnUGtK8GDBErlIhyXRjHz6Ys6PCGig3pFKBhfgdOJXaxZ7Vh
ArrIr+F1MQxOBwsW2lXRPSTqf9N+LWA21YGzXXiaf1CWueDW2203SHWftBFKzaVpor4nKRmHv0st
Mriwk43rn7cEkeCYUZ2ZUVhnZlyFoEC8AlfXcfW0gR3APNlM9ETmp9Iljl8N0QkH/E+gw2fC3L7R
75CBc4ZgoBOvj1ApFPuAgdGr9qfF3lSnOg3exoYTkqW3UacU/GGT7XPHqcWyDwdVAn+voPflbUjQ
UMjv/RsIqjXDLDfU2P7j7Ez9EoYD5MZaiiWa6tItP453/c6SMtYng9WPPY4l53FpEWwiAr7hWFCE
lfUqjV0DpKMWAFj9WoK1GKHwIGsSKtNIgjk9r62XMC+Yty3pYhg3ztq7axaTanEHt0akKR9UU5x7
H+YgQA6RuQiRW8uT2to91oFO/xowEbuI92PvyFP+RT6KtisrcP/w+AYx9OeQ0cvG//VkkhHOkOKp
mFd8Q2GKXvIY9ikmQnA6nUETF03G1ifZ4FY20+PHVfaooqDcNP623q74AFUCYv+4lw+H6BoFHB2P
sp/TQ/LXiB+NjMzYKGatSPzdmp6UNEsVCPV3SC8sXlGTcvjVodCUd/y6suLhvR8ZA3d34fCmy8sQ
a8Iis9Dx24twaigseV+42zTSi1U8hmeLNknq6uiZiU2oOP1qjy+3mqNTnhtfZKi/zIwS1xUfVsAR
a+mI8cXfxrSdYqJhgzDcPEgKVJAaxN1fle3mAC1DLT1kY58Vtdac/yvziC2TMYd0hZa53ph4NCCw
c9MGPnaDgBjoumprZqYwYdgRcSmCFMnWFInuoyFDf2mEfzjI/BjQTI+YULoRqjHNajNmXbxhAPmt
Ji+vS95qC1bKZ5Crv/7uAq59Tsj4oWCm6PnrTHJhHkvJVqE1Bb/qinzgiueuGUtbL505tY4jUphC
h8DDTPn2F+7aCEME8O/GYCz5HwPZ/9IeE//w7U2brMTq6eSH4yA0XzorOiZ44FBFnDehn+8e66ln
sWkXx/+uREue+DdTMXpx3NbwcEKzpdcAgWKRpD1Ip3j2mK+oK+p0dcs3HotsyBYoiQ5ctKakxhDz
eMwehVy0G97cTFcxlKx16WgSkliYudSbLdueAgHsa87o4zIvWJUHyYY4gBgRmQgkwJUmgPN3QAVA
Cutf2zk26H4TgiUXtEkcZXeLwreaPGHiY7kfCl0j1McOkXvr9KBxtPrVxSAY1GFMc/VgWPTeDXv7
COUmIZb0PpkossjsnMIQnATaxtdgq1vjEFizYHkl5XvxXfHCL3CyrDq65pDu/2tqVaqUiFC/t1tz
deynnAi1/AjHIPOsohi4oEZ526HDLeqeQ3QHYGFW4eWdYG8zo6iD1mBEmDmI5fnRizkQV0lH7+cI
kQ2smeyMmOHtzewz67f9S9j5fgrHtu6D70+EkNoZ5FYMe6sx31NwBbdbhQzIs9rlWKUnUhk5iSm6
+7yuEjvre+++o+5jN/gKHtS3YEJU0Xsb3kd8zDraxDDJBcUKPr/cC741SertOg3EZRwufFygBQ/b
kD3dLbdjWaeNRC+4mdLCbDFf00rcXI+MlFg3Xb6hrWE0tmjjxu3QK06zruI3O/j5NMD0kVbRA30P
kdgflReqG0iA5mYHNF+XM6Ksvrzlq0P+n0SYJjNH66JlStT3mYAlApJU1uuX2luyZQT3k2zXpdAH
EgwYH6nynQSHCdpqsOUfGjvq7TXN3Ms/Bi01FZzxySeia8kPD9rasPnNCGDT7BVWw+9MlFPbwhoY
M2HHzRvmO9maSf4Oz6py1T7ZyzTIy4VfdhZXybEutGnp6mzJZR0gu3dv/HSf6+tAzipe+1MuEOxV
HEQU8jtiSjgCoWWskVLx7rEaICPHyzsD57nDsLTKV/vDMIxOrqD3lAeTG6e+4+whShRPCIn2Own4
1J8VrlrNyqVh9Y/u6MmQMxxpca1m5KI9RkOy3wy6wUWcbxCoP6++yWZ+FOGPvIPKb609bso8v/qH
nx7JwKox5SIVNflcoGU4ygi5/p1N+0MOuEpOLvjaxzTZpwcsfMosMIpbicPcjNpaqTyzG5qSfxcG
AuyTKD9AkC4nZSSvt6GIOPe3fnNVEfJZbZUqEXuM6GDk6gZbzlH5w+/hcyKq+toKyLk/ppMsmb2O
slGnOTxVWYzRMjch2SuZrxN7XEhV//FkEGVFG94JxYYEkJMYSnt0PTObHq85GTy1XAUpebAdANBG
YDume2tsDssmOJqH9M0b01XMK/Wc7Lsx16KhONYThd5P6N/4noTR6/Jz4trTst8GMVuhMT9sO3B/
DIxqtAa+6TKdKEi0gHfmG41BA+Hp9gTBxAYE7geZkowRnRCOQejFMqL5eNVsCdyNGbg8R3G+DzN6
vEIF2ABVeCWXWLwTflyjvG9E2nsRBnf4i8a4tVsIVj4Ph9/kg+0uCFgkl2XrrxOodyqmaoW4csQJ
pseGBKPpc2V+QdRKKQSAVIqZKXQkZVUk4/fZUHavhrJlBrzX/mEDhE6x7cyWL/pwWfRekeC0Hx8I
MhjEQ7QZuXVlhV16DdsZmke3KUxGuVJYxJZ3Ht21TAGqGdMmj0vcue4WU+oxV36BSvTYRTQl5Cdg
J87Ovtvq7x+G72pJUMdD6Ym9qdWHwb0jtA+JzyP1JfiJ4vIsAZf9seCikvCvMiKZ4ixsarWUDO7S
HLUSSxAKh7BGpewPZGVim1mE1/qeBzuFqUcZNWMI3b0xxXgtsPuToLytKhabQ15icbQuAM7sW+QH
yBdW7IFadHkTPNES2j3upQ/zomzcKwRBd6PbSGnmJfSDTJFryl/AlQqpuQIkp1qMOrInlP25bQlr
JSOobsN3sOauBHzCy2TZkUDGYcHoMe7+lw5JE9VyXww4XvDLx4IYW336pejDjrpIu/SZoz2I7BWB
Cs6kDqvPJNbi5xkdQW7M2R+P2eMhDu/DuBB6Mwa8PsrAt5oTQ5NuNJs0oU4feZKcbRxBzykBUyXz
8pVJdD/kr09rKWMnxxwzRD6BFgZqb7Dl9bzr/SEixXUzPJ9K3fnsQJYTdr7ZN2az1QrvWAkFNrHk
SdfnuJv/h30qKpPQdtfTWAJXkdaYMI0WuX9IVfuFSbe5MASHa8DHLDUh8jTeLkCxzZ40vU4gUNco
z1YWfE2RspQo3VUmfddicfs2yBkzPUDOF9AsX6XypTcDQrNzrh2i8tEdabTazJkA0WidXpV5cmhA
Sts2UysxKhujwmeZOH5+yvZJ8Ja77f2o+BjElJlTVgAKv0QI3J4vnM0FadpzadgyeqsVDZPHGErM
ebbE7OrqE7pD8qlhBaEZlPs9yvk/zQlDNn9FSdHe7wqy/UCJmrU3CeX8GRqgUWdtZklHTuXgCCFX
85BYuG1sdj3Xwuv0XLSmMZYepZ0TdU/CdNGktzT3x+xgnioNReUaScv0l3Nd/7iKctaxPCZSDyIq
qVYq+zTf/LTnSheqpcgfqTx0GGWXE50LPUxrAOJDC3uHAXw0B/ybEJ3lwt5Mrotoi0VfZxSSUNuE
OOMBOFHM0y3Hynxi+ZgPI80n/9X16kidsyTJh9sn+sGBRPNL+Li/nlyJzKSP6bt82z3FjJDZJmC2
aF5jsiLKQ6iGuRxVEdUG9L9/UiUgoEdzpNGkXg+Wlui7RcdoykOWU2F3zTh+sd0qqvJaKpDCX7wW
f9rg6R31vNWh9JeFOroprNna50rHud9x57gqF9UicHmj/w/XhEoiyy+kOKHP3vh8V6ElnxoNOXAx
xNhx12aOgguo60zax8pAMBWtRQ7Hvab4ov79hjzm5Fr9ofWRaY/0KBeqkbxO07X/jLLdAUg3sdE9
PltPXw7sFJdX22ZMX2gjCMWjewn5xMdxdDIG3UhwV1iLfRJQkGKXe3USfULIr7E0FtQyI/oQK7BK
Dokei3karhEPUBWWwZ/PEzWrFkLcSsEStf4A0HqAxz+M/yuSzJeh7AtLCHo3hCiLqoZ/UyURjF3b
xTNrIcdlHyXx+vzUhT7RW/7/5zPeWD2W5pK02iVOC/Z0lH2jT9pgxhnPiyxfJg3LWZNHySleXtQ5
h9Q/aVoTchL7MwjGTO3OvloSd1npvz5PWdtT+CVqRAkvOWhTSnFS4VIUmnHzp4lgraW4S3kDkX0T
pcqxF1CKTApOSugOngzcV/8JrZ28pMaqiM9Npnt5zxXNkM6+zZQ1jw+e+PDqMZQa0XcQkviFT/e7
pmlruQgeT872jVLgkZNj1M+tx1Nspy769IxC+49aRc1gf/QeP6IAUcmo1izwG4DJPKFpINunaatF
HZxBhN2ev7L4uaGOVPReAPiTmzR/0k3OK6gyspHFfWbhULqVB7ehwkGBQLK2ctI6GfwWpegfRrJD
w/aKaHAfm7uMhFKcu/0gf/lQqpG7IpWoBQBB3W1ysN3ek/TDhmVT/ezdI4gcnRMhLizVhJVK6syB
lnjmZXpRMAtyX5++jLphUsdm2bVkWVUql4vM+2zQdg4DLDz1FdKI0H4RW3leTA5SIbiyk+DWYVRR
arrxJXb3p72fgh9AmH7Ggfe442LwSzjOnmwGUXpXBqbHL13LRttmQCKK5PTSyfsEmfJPaS8FCSND
SdC9Wms8DUqjbz0wE5fHth0sde3EpIgj2j/duI57XlpDxyBmZuc/VAi5LJXDxNJsx7Fq7Cch54N3
sQyXxNNci49DbZrMu4MjQiiYjfU73zNqoEVtzanvi1D1esUy3i/9SMoH9S3+v73Q8rcM4W6kLKSR
7ZdcxWxpsrzQ0YHjMbrI3h1Wgu3LAES/BfJTK16H3SXlBKJpGzih9RiylPhyN8cFwGzX9JObyCXw
ufAW6ndnsG+lPfxxO5TaN7gELNZAAbN2cMmUPwIzG+l2asThH2kpcgnlUWMjYmUaa0qvIGHddqQS
5h84Le6aHntp5wB/2z97kFcLIGjUkvvhhI8mgKTaYUu04lyCulW5EA02muzDDZAEuXaJvb3+h6pk
uAYlsg5LZBbw3BK/ND1qDzrz3ngY1z8cz/1DBVbnx8DW2dbeM0FUmM38fP2wd5Kh2tFF2oreblBr
y5AbXtBh9NcyHudOMk+ymSf3e11gw3jONENknRlLCXdTikcg4pv82ikeSUyTAI3RafIFWeSTxrOQ
vIZrdXEVqZonKkB+rKCmkAt5EFpe2mFsuuiDmEb0bAHaQGYjLHuUhx3A8aJVS9+Lub5GG4P2x6Yr
YVquKh+SCx8UOczrbDch4jxgFg0AO4AF8iunolgWjz6pRBkGGFA03ktNuQM+CSgydP7Cw6jFGSYy
5PUwtvNs0aK3iESJZ+1NoQMGCr42XbKlvcl7aTL80gKNcfJPYgG9AGeEf9OnZkR+FxgWAC1s2tez
vwc2GpMfH6rVjEbAKSd6yftPXx43SvVF9CbtzB2TqaOa5pBMg1K+j+bRwyrZmN7zQjWbPg7vuCXR
Is5kRBA2TOt5DSZNKTwy2yBC/fZGr1Ps2UXdLwNVQqcOSbDE5hOJ53ZKgzk0H4RILC3GfUrA1YMH
WKYOyRczSSrQ41ArzqWGywOLJunIOa8Cvc++MwvWiwnf7SLG+ZVYwDK7v5rWU6mNPFPkpchNknL7
qbP6a+8xvgyLtS/X5ivWW2mmK2X/51QUcBYuwjlZCwnhei5cm+hIN87/JHVwBqKA+TEZJKFTgFMf
yifNa8EoePhaTBbVENM3qrcWBnmXAJw6h5O4CJ05LFkGpnEumQazVjy61DyFK2/c9yYdJg8x7swO
XTPWQmiHkiAAepIQwnn8TSr+DrFq0wr9wljtXe9BUR7yrKvlkg25901yvouX0bNSmnkIMmx8ClM8
nrp+buERaHGjqMgyTmgiq1SSz3kPaIw7xn2NwhacVrWGOY1iY6+/7D8dMSnq7asx86RWApyYD7Mi
jcfvqIJmEiRmgNQKLjd1azM8ibgYPKjvru5K8gE+h2C4HU0e2YXB6MyhPO7l+RU07YSe8J/2Hggm
oeZvj+Y1AGBVsndQIrTMn1GVLk5f9otkLluDWud28Wfd6OkX6ruVbvzpMCURWlmE/yINDvoJuRLS
qtgqK7tK26zyOIUvpcxEEY6kwhWdOksZi/tc22Q+AdNyRBpuxThzNpP5KhS4Dv8qx0HhwEd5JOVF
SRMPjbfI2ZpVm1SuOaVBBCvXJaThZf/kE1wjp9tuXzNd9JJid+9+4GJWFnrvspkbq5ob+U/VXodm
DJVE5DyGPy+hsFzJixspMLcDGx4W4UZ4WKKQMgWB5XrL/e1MZP7nM2n2TrgTMZod6Py93iC5KowO
hdxcg59eDoqEJym6r7g0SvhRU1xq8Bg7yaq/lgQmu76VGnnhT1iIaH5WtzXoleuRJmnpV/sE2BOA
ush9BJlCsbEJTMqGvaM7O0QFi9vEmZFWNCMfo2Ez062iz2mJ8oFact7tcKxQPle4TlfdL6PsTfEf
bBFBvTYtANAksmFR/NOWQGaigezCfnv3mlzobyRiUVx0TMz4NkTbGkWtdVdmjJtL3NdGC/buQ7Rv
LKycMddm9u8LiXpvGAguS8QhByf9Oiz987UKIAOiaJ2g8trqsSC6K9ORA2xgMnxFbkVHdjnY5QR4
samHMcgqFPKODKVSW41hFHLVDfqugW7qVMmPq5yMY5htq3POKW/UN2C7d7Im/13bV1V0gUfHrsxw
MQerQbT16Z64EE4jJZfxAxsy89HxZoeqjBS9sT9bHpSD+0p39dxKnKvn8BEDYzzv0ySOYCMUv1ma
PSZ9XdmlzmHrxqdscQiG9E2I/J4FQDKyhU4wUP2CMlMg6NomqhT8kdaI58u71TxQpWBRNdWkysgi
hpzUEmCJQ97mjq6lIBmLAkOjmgCI8EamBrVAT0yms8+FBNBVI9QXFJOe8vLG9SE12qFp2O6st5Ib
qFiTedCGBnxPtQVaE3eTsHLJ82NvI9n0yVtoyPDucM+pAn2pPaPl5qvRfaVahLbPxvIIcnAZ08Jy
Z5YUe0FoeWHHhlJ/PTgR+BFxAI4zO1mCAltgjtabPROxxZTN010/n/nyAzEhu0su4oRWIFF6uvHx
iIdaktm/FsPHcdT4W05SHAMoceiPb863otwHWF3Ns/u0VbFC6+o8WEI4A6/oyMm6wQquIWUExwa/
j9OGumTzF2C3nNMpSTNligcfyku59YKxs4EhwHnKdhHxKHGS2xEnXx8TdWgigy/3K0fhRhJvq6ra
iF8gSWFA0kLTB+7OhB2wWxG7byIhdcqqd1y2n6blo4LGfME+4gYKOKEyRBGBDv8sGu6IZMDJZb1w
LNRLTjzoFAJzqqBYSkomBc9qF1QjLbagLrosqN+S6M637Num9wIwrSDwh8f5wK+2u6fmMjkRk92Q
yt3z6yDiUY7RtrHClXwPek8mOdx+Yml0k8QqENKUfGLSav9NfjAkSV45IQG1N60be/FVdqZWD2sw
+NeCws4eTVFnA1V3ZFtKexJ8nzcsZjaFQCyEaROYiDkqrrTWnq8N1mqbS3iLJlwJ5nyuJjZ6lo57
5ev9CCy923N5i2D1O3S1HPIHjitcKAi90awZMfEad91KD9Lm0Q+LXsrIE1tecX5VcdwTitV/BEgw
aa6u8Zd3BZu+pXD49JQvt3bhYabFqkjpBHPuUmyAd89bmHK7oXNhPtasJRHW+GtHHzBlYKy75u/R
W+P5v/ynH5Dm59sJTq5N6bVzmtQ9t/GqfOsnlOWObf12DrtwOO8RliKYlyFWyRtYe3Bae+udLFsv
UGN6GlMsI9/wVsNbFSm9dl+qR+rkW6R8IGCN98RDgPBQhCQJunjU7SEFen0meo24qaYfu7ZLCjUC
QzfPjZb8JoP5WbXUK7jgbSu79ig935WOEpRGW1ixtiwXHpKfRPrkPgRxOMUvLs3nEPzon95hS1HH
vc+b2ugSuzHH0ZpCrpxzRPOllls/x4tqCBP+Gm5vap/lovx0XjXPpigfFohKqUfbuNTaMysBuL0v
kAa91W+9/F7+bU42ZHRMtwsjI+M7AMLyu/L3jptVHDd2oQnDxRn7npOmuYPxFclqRnZBV1B+z5pZ
awdB247/QMOYsMmdaVKnuppeGNDtxnACl2aZzcidxzM3JUIT5d+S9K/FeBrk8HzYNUrhAs+Pl49Y
LvGC6fwTYnvDrX0f2pIIhFRTiYSKrENVnkVaeRbeVVeKIHExdJpxa61mWWoHjdaHwgjNAhs+GUtI
5vgHe+zUiYTNluMd5Echim5IG8wz1gDfRkOe7h0c21UYE1xkLz3dFLLcjoT/CIVFdabriQBAbibd
Ay65gg0EPc4bE4qENOHx7SMFVtzAepakyp3pwjT6zHpyEADE07fqcfs864dk5OcVL123P9jGSaEi
mvq+XP1ErL0eJt3IS2Y0oEaJBz7xQcPv/sdA1UbBUu9PUBJxFtrVAAtcWe8H06BPTZW6f1Ry2fAV
9V0CTVTnxszwV4pvioYNa3Zolm12/j/7ZMgDxbmxy1rCWn67izwl3DKSLzmg3kzCBx7G86M4EICt
5O09EhYM2f6k5+kqRUfZGYzQDLIw09IvdyJXnwzCPVaAPv60/owrnV+3w8THVkniy6nSPggX6vSO
7ONPkfuu0p62t71unniM4JM0ORDfBp+jtQo3rLG2Dv/XMp8Sm2aBOnuKIem3qpg+bHZ3+/Om6d3m
GNyZQTPzvbb9HpByE/FqyMy+2fzDP8Zp7gb2t93t/SziUHO7Wkt0Ut82scioTnjx3ikTe9FVNEYB
3L+78g2CElJstwrFfQCsJUjjQd22yjTUEKmDOSxK/AsqJSd2weEsRBePsaN3q7khnbFHeFD3sMI3
/heZlCbVYBHnLdQKtOee0PWCxk1hQl0L2zEZQdfY3d2h+wwTJ06Kco4c6rMYJfJS+0lfPGttdV0/
JXYewr3xdEBS9gyWdR+7UboMCV+St+wMysE642DK7WNsx+5nMfu5fAb/WoB0kdosFchDfenEJgdN
eeJ8tswHTlLntiuWv3NpIYDFnIi8vIQ9z/eEmNk74Ewf+Ohlk6iBWhYyeUiwR7uDJ0o2FoBvMbzV
D9TFaSg8shqhZYOjrwkbqN/OGFgbA7w5NvSscMoXmZrn08ANWisfAHPau2R7CAlPFjIrF2CWJcjW
WpjrX0wuhM9R2ZsBBoGbeuetQjWh4D+asNTt2ygRtUonlFeNCUE2xh84/bzcpX6Ma1M2eLimUN1Z
px7BDLATo1jdoQsZtJFkF0ysf8POfL/XTlUfuh9MFdjuob2XzSLr1dCIrSLehHqjQeyvCNy/YiKY
3HLB6VyOAnyll7LjRUj29aflhLTuLpWrKsy2aiz2xX08uqdxTXyXjgtii+m0IbvW5kiieS/1FDJv
cDXLmmULpPEn92gpPLuFJOKDboQvCtoZ9wq/Zh/rW1eKFMtTCeOVLB3/tC9OLMyO/t36vYPG7iH6
nuicIUsf/IXuBkcqdhw19537Jy2MIY+cIj+ZcF6gqtiJ05sld/74Xa52VzyTdPkCvA/tqPyPFccE
zEF0IbtZ3OnFjWXf9NZDk34SRZLaVQun2zLrAoPd0GnUUlwiqKa4J71uHO4pNDcpNQpjW2Z1KlJV
ZQNKhpaFvb+J2de0sb59EPbjuxg7Ao+FOJi+F5uLkl05ZVpumUL0bIDB7ewdBe7C6ZeHsmaPBS9W
ybOZGrbMuaJ5fTtoKI48VVZBU58t00bXF7lSQugP3Vjco1Z7kdy5FJx59w/AE553opHjrROaSmtR
mauxs9FjzbGlKgqnDcr1fbhWfhihYrHPh3tJHsaCJQVGn5aag4kO9T4PlSlqsKGHCAxm81yquf06
h87dEZqBA67rF1EuX0zoNbSsqE2dsTZok6SmI3NSGnV4QfQY+hCk78UDoos9clm1YSXOJILCQAl1
JUa0HyTJTUWT7WQ07OZtXeRzQbtnycE84iIlYyWeIP/u2e1v5aFnDw50+owjc6JvxFbNBalxnb4q
VQ/7Hdahzs6iukYN2UxfRPF5Pjer4OQwbP5PxnTK8ODpn3Eqqyw3UksMH8l1BlD93LU8ZfilWvmw
OKGpo05/hpsm674vJcfqYRqCh3hTmqUy6kX2+gKRDe78m1yWQJ+ro+k+983RMpVkVGWVLwbqdj1T
v6oJ0JOaxOpJJ33NAJRSvXfyAFbOKz9LWXXha0iO89qVKuh4IrzFR/5qUKwnKHNHNpqUTa+nn7m+
wO9S5yI8JNTD8laT+m7Dvhg5AIwvfNufjSvs63gg93XAjcBdF7KDvIZhqVGLptxKua4hSRq1ztwR
Qe/dAjFB7PDtYgpMB1+Pa1cV7FUme8r2Dk9QmkWgz6XnSbkzIFXpH2DuA3X+NtKj73PJm05rTsrR
FpRNJOg7L4ZeQNm9+7xLCE/GtKpxkbk2AVAV5upfwPt9z7aaNRmNigv12KwSpu5wcx1P1hGiL8KD
6SnBFmxR2ZU/Lpd6exUretHO1UHllsFA9DjZGeT5QtBSIckssIV+Q0Fq6mQEACb10zTv48TqWTrF
N/DWB55Th6tp/zjdaiGzWhrqfshf+wL6vxsWTy/v015Gg6okStRUpc3U+J2gzCnPtzxZLnC2z1XS
UP1D9DyDj7BPimOd3Hqn3GYYFUw3Wm+mfgzMd4XhBLTcVadHdXp4Svc5UIci0XOR3f6K3wo07L28
uDTFzwJ34hawXqMlkAaI2LSYwRwa0MPmRknmh+9E+vP/NlS4kl5JSbYNYTm41SwHKkNiZBDQL6ff
uSXiW9DyysdhmdbckrnSAUJszBuZ2Icuq/m29v/DQ9f75yRpvSbgmw2/S7TZoC58QAfVWWGp51Kb
VOTP+g49I+6/n3r7MgrF1YU1i1VwZUPZ1ODcoWFTRdolidbcD8SkpXP5WVOen8oYqG2UWwHH0co0
SJm6ACsyMskdVI2syLZ+m+puWbKcrhKdZISmnd/U9++ml5nNeQFN/YW3bqE+rMGhPzVMz16GOHB0
Kj4Jyf+pKfuGPKq5HQlwTvDqSmfQ9+P9371GI5ZQqWJR1fgnWuLzD6yGgdHXnXhlFSaev6UBYdTG
F7P0WnfoJ9dqHGoEnyLTfeoodCgt1b+4fS2ZQlolmFn77z/9qR9F5oa8zEkBdoZV6ryrXEiK3DdQ
i+zqjcnuWbk0Nm+q8zLOXEsOVh7FWruAfZeKHvd82HJDSaJnFKDwAUJrlzScFW3tAVapWNu1gHqZ
EKfXIUNxGcLI+CNdZCKVq/1CqEW493k9H7Rk5/HN5a1niTPgz/9zTomltPNObFbiGDDmLZDJBiON
nqevMipSf1ZhoDwgDpyYYW63hyr7f0bWOcHIFTyeIvZhW0MnHMmSYANVC/pfO+0yxhkV+BNAJTAw
7E7WJBhDGKrlxwOO2cqr473hf6CAJ/O0CmMKhFVm5jkd/bJCBtPetiKNoXP9fI7gsmMgwzty/zQG
GC0jQ/odA/sXb9UPCsAoCyv9v079/7Lm/f+tv+TIvNfYmHE88dOg6aMtXum9455Wc+9X1AcHUQdl
lnQLLZjHAct/8NL1lU94RpkQHAi/lAO08m1lrxRjsaTLSLezNB1JANdNVtk5wg6k/z0EjjDfrIWL
fDdK0/4ItbZFnCA4GmJr2bmEMujMwE/5EqVxyY27kct5QL5O/MwpMJcCfclPrmBxh6ByiM37s0xa
Cax/3wCluOAGP3I4SyqGtvK4E1HusvqTXmeTB4CVdnlVYs2BIA53sxRuf/UX9V+SpNRpacQZoDX1
bQH8i9xtSE4rqmZZD5OKS6qmi4pLX8EX+UftlBFiFPtZx4b+70qD/omDcPKAHitG8JNxNP/WKr3g
vJuqRVi8wecLKWSBBaoptRVkU1m083c74NT+0pEdwuU85nr1PhRpCvJu5134iP9g99l7bX574M7p
4JLDK8gzYDrZnv9dyKzdWZ4LpyWnT40li5Z/uQuzhAmCLKV4GrZf7vxDjrkwez01XvBsaghQDuah
bZwVdWdix60Y376M/csUCH9woSRtRRD8yUwGQ0ib0QV8r8nwAFymG0ihf8TDkEIyjgYN2ypWUJ2p
ryA8EnmT2IAehiuB1wPD0+xxqgZf9JqqsPvRDpo6X3DIcNwqGzlzpj9dIYnB0SnAoNjeYo95mZjd
lTvSyEgiTL0ulKorsmSqLB89Yj1c8F19TIWHByEzhTw5ow9aAAYFsb4hu2aH/57oko+L64tvGxJR
tbR7dmrB9Eawd59lG9ijNhEqTJH4lrCImkmpvlm0Q3TAl6TAYuOAMNW9Yu7cFuqx3p3HIIvEnhLp
yUWyC1e3EN6AaC/U0b94K70mOGOd0J1qm5hHu+P0anc4BiB7HwfiwG2H7tWEue9QfmpPlJLR1ycE
AiEsk9X8WqUFhHmbEzIJi/J7RPJSUMAw7XqlxPWDMfn1MbHVWSs/cw4KiJxp+RDAz1toLyWpiPDY
fqkUodE5Bv9fvL10YpRqlyag9p9xFJBPdEE0B0Y0lNkKXZ5EjFkt5yNHVP4RGGmoMy5xjZmKHo2z
flUGQxFSPxprEvsG4MsY1ti64h/ZSBGo9EU90tmSHyz9zUXviNbJLeUydTcr2w+mnzZYMyfr+QlO
lXZSlGL4rClaOIH+PlYPjJThQGA3YneTtIt84GTrTFhbtvSsFgUhJ9mnzHteJnFi0uVNyg57K5ut
U9oT4vpUJ65awrtBTQLS/ptGboVzOtODqt5HjCrXPL8Y3EJQCagzdReOl/BFfORdO+psRk1vWbNJ
ThTckRrcyUJLtzy3OzbE0W56c3aRwaEt67VBEOjnQq731XkuCS2uhgoTgorL5X2G2jYpiPHV3z33
uypeQzAX5Nd76MPolHG02BM1Ue9zqX07il/IxrjXZa4I4E1zAPChYz9DHxKNAnpOEY1ZQ+lfN+0F
g2bC4sAb5St6ZTtKBuhL50BOQeIBmxsFQYH196E9N6R2q4fq8Sxizz+fvegPyFqrwHMsK0DFKOZn
BAq4tB+Shj7wm+RTnzyawR6JE5IewbXUmPFFJUXJUxYBT3JRkiCJQSl2ywpdk4u+Mp8n9Ret2y2q
M5EJAfFg5WJG2tBm8sex6Y7YQs4doJb6xpcl0ojcT+EuDct/w1yCzAMoe9fORmfw73erCW4DAbvM
IigWwTyD8JHRIfLUGYpHWKAwU8ZOwdq0SV+NQFZrjzY6q9Lhog89hnPcXDpMKs10FiiqP7jy9tLh
pJir4VPdoBx6zcMSjAp38f4SpooA5bfRPiciaagPPGfMh+H27dCPtNkUOG1tymylDwjQqLSl1AHV
opEW4kNXdteiNqCpYjXa81Ph1COZ6VTRuuXT6T/6sIf1gtMkKj3bGWCORHbSl/cbtB5IuL2Q1U7A
/RQSsq+M5ksBJr+sCoI8tglRNbwfV2KJm3c4vGCze2KOcidkfEmBFXEssk6l4sJb8eq3wvbslwNS
eAyL5uGp2wp6bVwoZBz9ZAxymbGrEdigvM3oWnB4Th36YMwFnfNac2D8enNJoGtC0q1vBleJCkkr
wd5xuVJ8MiupIkCvTcpQYqOYAABSu5OfL3yoH5HHpAnGAqNwS6MLzCteX3AfsX3nnsYiTpjkxPJe
vwiYfL246axjWdic4bsTVNAvEvacIFxpZvAXFHq4x4rWTnTXFIz3L1fez/gY6PfUqcEt3Nyk+2Yw
LzwxPbTpNrAhV/5c5/kQDDFk1g7ZPLInW8UxmmUdbHy4dL/kR27jMtpM8Jpx0oH2WJzz2DhVMkCc
fZj1b4P1r84ziHBKsn4zFUOTj53ApMlYrf3FhJ7Z0Wz0hoV4bPIXpyG7fT1drAv5kMjeITd5QfXo
E0IY8hlU19wD4tCAhW1tlCPX93NmjTlucnglSUC7ui/OysZfO/rUxcOFqhWLYRmVYhaeBqCSAFlK
y9iTYZCBnpKdpXsNOw0r6AZTmb93YRahdw==
`protect end_protected
