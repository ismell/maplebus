`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
V5Lt5UpXNvrXV7kDzX+VYpDXf2swykHFmwaZqN+kD2WHF5WXsIR3Q9RlbZVmP74+5YWxrjKhuZRV
YD/H6Qp0Kg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ES4/7IHq/EFi4IOvDvJ4Ggnt4WXBTfOvbdPp2TTReVgfAv/Z8d+q2v61xgWNlqy9ecmpXdqzGzUZ
PAnTh0Ecj4qb+HzLhJVstKi+RA7LtxEPJiEF64MyU3ePbL9G2EHFjgLJyBvb4YuCU622CjY+s4Wv
LWClu1L5Xe66ZBIsMpc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yqv1SQzT6DcD1EkGaCCOo5uts6yn/a+kzOK8KMRIumOJXsu+Kdkv8Bed8kvngCA0p/gpZ/qL1PYM
6GXJdr8CBRRrMNznfyvUuqgsJXr9YWw3Th89Sr6hTrSnzZ4YK2EJLG+efz33B2i0VM2UAUiqq2ix
XTcC7PFudgXIl1XNkIAqXHtq4YRAQm5MDCvBzqc4KGGzdwrXsHxHnsyv3h+Rcn/jR76R7lafeJCd
PAPme7qBNlxzM+3lHLXoTAJ8gaUpmLTXBss0TWigFXwxWJR9P+ht7pbtUGecqrkTYEZQaddW8Ww1
CbruPvD+0+7U/6hIodujE1fI5w7hSelFnIN2gQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e21NYxfh+NL5f7nviA2qFEpDfLAqnKhmtD0XpL/LG4LHuEMNoOzx+BVU2T4Sub4UZsbJUsHyTePd
nVzHXRty+nDCN/FwlIOTc9jUAElkAVh1cfof+fYz/7c9gf+S/wFzp3HFmliv4F+83v/ZOY4kkqlJ
sqVxjSlwkxoLPvRdscI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pCExxKLZ3hQgr1beezULVuF2Xgv84x36KC/vGXB1I8PK5r0u32ztmp3q9HO+uAdvd0alZXtkq5NZ
Lcxw9+lStxduLn77rhvNuskhj0BBl8jpIKTcx6nhRAq13Eg+iVk+RYJxqKDDfOMYF8RJrEMNdP8q
DzW3MFKshGtIHNIkNnsI5mnOpFTipaWgVm4F4fV9Bk7A8B/T84lLgpvCjM1X6Y1b+mQKPsygiN+i
Pxjd608fZbo/qhlOUXAcPzGbfIzyRI41Y4LN1716JmKIWSwdwLOAFVW6wfO6qqvV9d8qAgsMobxK
XUpW95V7rw1zc8tWxWlOsGv91I0vp/MR3kO4Hw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18544)
`protect data_block
ScdAPD4RjHQZF8x+HWKPeVFbgXVznLdeb3O7WoxXOcq188XAv2FOdgU1Y2091+nuOVAShPSxsC5n
Q4Ev23A0IqYkiQXhBiREFGnH7JYnqmMb4Zw1t04KlZmS9YghJSyqGY2oeO5wa7j5YHnl9dHm+Uxp
cRK5Hkm0jhp2h9E04K9N51fw6p/TV0FeqF1phV7ecX9E/JzTnLxFAriSyA9NWug429L/W4E4K/9g
qLg0zc3H738NTWMZs9h4ehlWwnkIhhqsl5cOQnjOMQN9ogMZlDrdPOPzhPvFc4AVJL5h8gGAagER
GnlmkGDA3azcytBdPDJ1jWGW6ivb8/sa2I9O1P2WUK4Xfomf+opd6AP7Ywxtx+AHuGFXwQj2as1c
O9DaEzQYSUZtNpsuSDC32L2WqUdJUuGgNGFyZ3Zsp8EublT/UNVX6GkyWRy4UPjsUSuS/EmgnCjR
iF+BFbpFze/JdxfsCW97a7DMiP/XTnIG/4v2+GddJ8HaHQfRzZcv6DSBApgTyW18NqzoTDs824Dz
MtSmlnF44SVAJ2tosBFTqA1xHUIOhY+E2FBmRH1iZ3NHgq7KjNnB99bB/wBzlW2h/O3R2m9gp++x
sTd48cZbnReP7xKCZQTO5eLhIrCoEZi+DXt1w+4Y2kM+oMfOHeLdHyImrTH7qcY1Qkm+WfJjrO5l
u8mAAM7CeX+CICyfcVSASNl4nzElg+lNFyM71SRBx2oMT6OQlv0eeMAiOwAnm+OxYFTODTfQGp0I
cTIlvuxz5CQ5NPgp1SUSxVzUVSJa9kNeEFcslGv090/N98gjR3zUoN5gfYhKjimh+1T5i4mHoXIx
OB/AlAadViOm+nJ8Xt6SO87F7veS7v37+Ubn1DnQVJhybCXwQbJaWtpIe1RJlr16iPQ1lnlruqDf
r/D891ZkVZRUv3wDu7apZnMEkMg9LMGNVBKdfjLSEp60T6/IgrkqqcNc+07wYx1niIHjGV+zg/+N
gDnKl6F2HozITPAGgGhHd78ijMq6uADASqVAVNsffWNnqtTNUkavAvZBNDlWrY6JckvpcLywq8xd
KW6hFIWJPmnq7Ldz0eAgQgxi9662PUNra+4DwryU6/GinFZSOK/GMcqo7qlV8MPVYny8WtJV7S+U
wWFb9nJtYm+xvn4PcbRoJDvsnk4hYSp1SOmgX2EHw465UQuPom6IUxMA57ZLqCNVsBPzaphqtZVz
GSwJTq26vptBauKgvCqY2auF9S7K8OJ5UIodvrwJ0cYAtg9ERgbbv546By8T6yXx0lDJoc6e0Gv9
kO7BQhUN3kPL67DX1lyP6bgRvx8z50cuvc7ni08cde81Z/Xl9bUetfP6KWRLiJZ0A4aIRhnv2QRG
f/rnyCCW8kbhUZ9YhkCSBoC93mOp5OKqItt8QDunO03JPg46nIRqQbglpLcAuyAgdLVFPJatcHS6
+IXKOs4K32VMdi+bxee6xKUMTozmoZGN8OOk3gBW/7KIdewWZyxszyOYxjLkcmqGEwoY1lq2H0Yd
vvkmUTn4cfKdTjijDjXwVKk0hDCtZ7PhvNKr44nKnsADtRcun7nII30SNB3bxOcNyeWV7vpaaK/t
DPguJY0Icj1PAy4Q5XWYtI0NzXTZcMAH70Z1jzQWGTtAuce7I0qkJoQAq+bAJKSvVZpJn8A0BRt/
Ai9jxAk8XZmixnJTDDDEpzCPzaZqspcLycbNev/bu7OOaul5kYGR6NLP8hqBUCZolDWMfGGSFy7Q
quDLu2CmWJg9mtzDiMo22lDG3a2Y6HTqOvhanGbgDfpogchpMAMtOh6P9cszcCjfZMSJVz3ZxuFp
ZZ/sOn4lGA3oV+s+flP+uqe4fxma+D6uh4Ah5N+LXTr5xQrtwjqH2dCLM6sdfmcUe4/SeVss1RWU
ND2iPTuWyombz68slSKOXcTJLHLDmMoptOCOflz9Wh64IOhHbFrV+G0IxB6cYKHK/mSKzWK2n0xh
5gUsvzJhmPOxMk/DTmb/YR7GnEAdfoYB1alWE8rvsGOIf7DL+NKurZM+9BgAJuaufhwI68dQKoeS
qGtbFeJv/7y7TcAV0LvkTgkkrqGCruaiHHbEz0Ns8cL0VRlbLrAdadQ5BbYqW4y9CZ0PKtbMIYMA
w3DNJkXHvQUcOSOCDTNWxszSWonXPsFfv4Tmj4buO+3RAPCmL99Ur9t2meWkuz9wwlbeRcKIMrQR
mhkiasNTZR10M8vd2N7LEyc73F6bJ4BT2gegsGbz582wd8WIbYb/dApIC9hcAg5Dxa8js1vYIsPz
tpJQ0eUolGmn3VT7KH2FoYWii/MzLN/cLmzAi+WNeM3b2O2eGIV9mmtUppWnMrqnzgFHTg28C91y
pn3Hg3I7gzwV+aj25hm5nufgC0JacGmCtL9x+3MM+TUaHOFEY2WyOcx8HZqsXw72pPDcxQKKMzeo
9hDZlTZ9nXnLiWuJnVSmwvzrKlnJNz1TWZxBxvs8flPmcXnw+wscXiIBMQH92IXfIe+/+lPzm4QZ
O0YyG6ZThPCh/aYEPNzRpQgaNy1uivTm/782AET+jWagsJSpDmtwJBrUB/0FUxBYoErwveA00opG
1JoIc/L2EL7aEaaUROzC/289na3jxps0DqGIqLpCD6ZmQbK92m+3u/vSLzf+J8/5GTWc74OT+Q0I
eEo16mMTlosFETpWTwD+XM3GDlvF4A1pVStNd4miF0Gsio+KtnbAoxGti30o5iauUw30Nn7EkLTc
L8iNCZiCjT0U8XrKIu5BoF0Q+vlP5fBgRtpKUpbHIPWcJlTWmOdzBHrxEh49FlVMqfFTM1g6+dRA
4Sz8sefKOFKBZxHbMXr/H+bB8DF+UPQSGkeQxVZWXdBpQxNoq2Kdi7gWMsBI2JDwNG3daAf2Q+X1
czWx9cdT2o+3Q9y/gdXcS6MtPU0SktL//L6o4JFdu0WcgG5HYIQ0Ca2ug2r/dsEyoabSQckaKP7z
aYMODGQuLF4V+jTBgE9mAY6LceNdIRkwGQo7DqadaNcSO7eH1Zjqm9+uVvZ5u0s0esA4ummB7Ivs
RZ17E0U7UA/cMWgfOn2rBglkGxSzkXRittu647xkYrU5xdL+dlJRfceEqgIoeIkyLBbRML6leHwV
llv4if7b62gg2qaSui6YQsqsOGBUUU7y7v4QfasZGHjL/QJzxD/snYYDFRNK5p0CyyOt5uOfXHD4
1GO0O0G+Dxlv6ZakNHrdz1VOkcSLo0NTTboh1goCihy1R6JIqlge7eQt2pFVyJDmvdUDtHqz7RJA
iS4RW+CY/q3kZsQ1C56JCgzkDxye9YRTgrhPMcZ2JWUkrSf0fTk5S/6LOLv2ZI7Osu36k+g/WLJJ
D3OxW8luxtxEcpFqFF1Jlyux6oRduO8DXmdeGKf82P+mqDCTiTBMKbYoUr+k0iSabU/q20pWnqKk
YH5EX5VK7bd6z/9VlQBKmhAeJ2wwFZxyNfBdPjwjPTpcG3RBQL9wpZZOvBtVeUeJPTvFedMsXXb5
Tu93/0IDfiyPKrs6s9+cTR29iGgPD0Q/dPBPaS0xzGRJOnlV8WfFMHhTfwqriBf/s4hKJ7gTYPNJ
VN7OcAmN1AidKJ6L1zMY1a9HSbjBhIi41HfG2iDdQ/mqYxPfbry3YT6lCwJbLqzhojAYt6+UzFyl
Dbhy+L5GgVVif1JQPr9i8iMq967veUICGMq6xjCVy2czWQDEl7tZxzRT+33B8Abs/EbqRP5iExoO
CFjvKB54TQo66E0C+cM9UH08CHoMLE7y3SHeAMY91U54UvBHNaU8cHQgdAmkHdOaX8HxCDbMqJFy
aWiMNO2tSDr5Kp9//mD+20dSSuPYsKRL+CDdvUz26lv/Ju2cTt5c5QV0yK8nJ+h6tP/eR/5Knqpm
JkShZAf/rDCD//5LDPLlS54cfWBmzLbiKWzbyCsrUOGU8xGu/b8qAoK18DvTR3Ilzr4vddi3pHHW
Hujou9/4ZGwpZZjyfkj2zIwkSmG7lIflmYW6aYcoZC36HeA1SDNEdgQaP8O4in6YU/bFQJkmxcuM
kEJQSHTgZAK4ycuas9XgnpH5Y9bYqE3RDHYrCG0Z5qWqCd7xq4KhBd1rbWZeQXU5KWzaUu1f50EB
RIJIP+TT1c507ntPMDzChG7V0BDviYJZVGA9oMtfXeIhRqq3esHLk3wmu56f4Ry9dSE+rqd3CkBJ
9lxstKl190bWdLMlmdrMhulM/1M+AfRlw68SulgrZbojyPkf6HirLfB6utRZFcbQ4QmpzMsR4LJ1
zzfuh9aAMwiD9JoucBRQGSVBPsFNCSt2HLPF9jT88Efw65wDe8vKPNQy26jYTAxb0MYb7TDpEBGv
ZHK1nFP7lWjisockwCZjG0HKLMLw3Yh6nV74Q+aP4bHwsHmtSp6F4wkOo6PwTtMo9Hf8aihI7Ms5
WYDkLIa18yulDxKhgz80Gm+IDr2P+sxAkDSCdUhguS3Tx+GzHV0srhJRAy4kGnJKWlhTUKcP6um5
2FnM1JnnW8Yh8ZPMBeVklsbCgBIZ2d8y0YKTXRlx8fSFPmV+G+y+vSdsL+cN4qTb2+52YhKZ/EeO
3PG8ztbglcvAqVjsMMqI2xLQJlVqhlIeApfAd55U86WHSUerhKXf4L9cx5f9wh/AyHbW87WXo5/+
UpoH1ZuawWjZUAm28dNe1FFUupdvnO7x2T3o5rfSpTk18LzYqpuA0uEykfC7OdIehfBIvhF7UU5a
VxuAZ+nIOjqzB+isJqVlwjY+IQGPEuFw49jb66PWSvSXip6paCCLeqUxdFZbTQqnKK9bi8JfgSBJ
q/xDKoT1XJk8mAGWA3WyJiNJri6ytQmXLLnkuugNJNRdlbw8ZB3tFO5IVgs/XSlRz39nvy3gyIOd
l/GMybJlwslCgDhIn6RwZysBpKmanK8xBoxxh9rU7dWbZ9Eg6d225K5e5x1nN2e4ZLaB9udUPQ6m
TxbGExhWHCdg6RGEjEJlsRiWZg8xDcXHDHVg+i0Z9qZDKdpXanrZ2+wH+YgaIgZj5Hk07NCYHhCk
kWe1lfeqIAcVGpeP3eLcMu/2zil5OcBK1an3oHA+uTMYc6ytIyF2D84D6BtJJ94LroTlJZIzoCyj
25YWfYEpv4qAoP6zj3foaqYw3NckkClzJ5yN5Xf0HIOH1lUIQ10xNlk+cS0ech7HooGl1KrS+64/
g4OXfHfqrv0tj0x5pFvCTSiVKv09JiQurOCjsgsZWNNXZHznFfUqUcAbMPLQxxhFxcXIbhrXAQzc
mqP3Z/ynBT0eS3DXKlb6R1Pv96EGCK0Pk2OT/2cFco8SHydzD6h8xf45n42CUcu3YqzG2doP2C01
rXPqG1GicEDuZV75lrq2rNHAHkCqkZm28vgV3RpF1FO5C3Zwt0V2Uo5Zjt+eV11HY04hHeKQrQ+k
fuCkIFc0x1oTBhCRLVnC2BIBhAIrjUqxcwZhgz08AU4iZjs7BDnuiU7ReP+otgShBy2wi95/sZuG
Sn2lpWK/0oxaeP2XW8hylgZyRfVccYjAVZCiiQM1yDgpNfzu4mZMlE0jLT4vEi8w46INSo0vL4z9
XLqRrjKFlnWjG5+kIZF1abKnciJTGkjaKMIWvtMEKzW/oXQ1TrsZ/1hH4kRuvCCqNgQvuI2LPgbn
bOGMPssL4NJzBnIwnavmR8Q6IFEpeTJpn/6/NypvgvkzMsbQuQwQuXYXLWKyA+GaV8bSUGxlgfz5
LvsV/ULIdac0Ncd4ps/Johf4B7O+SE8PD6t/HGj221AX5bo4B8+DqgTcDELsxgqJqFSR7Cy2tF2h
QKc4cLKSIITa2xkOIA0tJF2NeZQKwNEfiuvVbr0/ofO3A9xqBt8UWYesMLaHtzq2SwxrnOV/NHno
VgHBCZKrqP6mXTCLNCnxPHIa/7t6HcR1hJEph8hgV8okjKsQgyaJyqFmhDU85ponlVKfCYVCrI8/
TDCsm6DiBMMTlMkzbeXf8KIGG1phtpQlSJ0LRbG7zZakFJOhWx6XxJyG1Xbwtcq0qcOYgp3inPme
kOYDJvEShKyrxjoVy9u+RvCXXNm4yA6G+4EtJV7G7DjPhsGGSKc/gheUWXALvr87D8/Da0bmMYzi
esKwvYGdjHOJhArFbOoyr4MFLL+zKlbQGhGtXvg1X/tlK54yXxMfdhcbWTsCvQ8GhowyYSQ1BKIv
f1k9MKOGrZd9bSszd/MLPDTMxVdlCifnQDnM0vKpEAvKibpCXVns6kHMv3zGx22R8U2N+TyXJ5Wy
OXorDRTsFAmZ2WMvgWilXQ/TX4WncMU9KERM8LLASnf4GBrsWLAINYnjvB8xYXnapOlx8gTKsOYj
/UNs6UaZs3BeDQt4TbiatVVQO5DZAeRXiIxhpXLyWU2weMvh48Xxsy6oRmI7tIXE8VX2/3mM3CoH
+PxJd6VTtHLxR+wobSnj9S1P1+sNYFzRpzJbFOUr40Q6Bh1H+JZO4ynXZ3CzeQJaKGw5ggAQKDtD
3qhqGQKoSepH3cIcCqazDxoSsa5hAfTtTf4sFZ7DmB2+l2HF4D4tSCamaEgmtlH+jDI5nhs8RpqY
2GN5C2kd5YaRQ+uURxHvF9L76IcLhRzpztEm5MBIXx9H0vYJs9ixWDU9nMXcs3jp6+IV9VZ5xNSR
NzR09wL3tGkSn06r30Dse0nrEwoXkBeFxX43x2gW6gPyBn9RJKJFFFV0qd3twwI95hpeavOL62oH
hUV4V8Z1urInE+iAOB8/UqNsE92c52KJyppy0SBNOiRnppQTY6uvTq3m9xUnkWC5OVCfnCty5BB4
b7etukxrAB+7FJbVu6KQLfNA+0WhJJC4sfr9E3HL00T11Gf6Zl21fHlDrrmT3emd211/93ZOoYra
ztkqi2Pizdmr7SVVXzFx0OTvWrvvquJxcUW7YhW9eZSsbS42i3rQB4h2wV2uBijyKa+9nd5X/lGl
mJrAb8NtPzYQpn1dWMOPaTCDohk3D936g4hm1ffpRJtNUwvuvr7MtG+8Sf3VAgGdpL+x0hxvGSh9
6cWWYC+PW4hP2iBm7JzC554dOY3/wtJ2RmsQqPkfHJnw3j/wAbLDHR2lsWKxxNySBDzz3FF3Pjgj
KFI8O90fLQeAziRmuvCKRMvhR/CwXjbSGoOn+vODG8+JEeRNQlUAcr0XNUVzf/zmbUB2V9n0KVxO
7kD/O4VW/hqNKPrIfoK7NyJ7d7mozYKZWoYBHSn5XC3nt1iNnHgQoVJAJaxe6VW5BT2JCOs/mtiy
8iwfDr7AYn+QxJbXacI09/2bqXr2hqZtGw5Z8esLg9ixhrMlUQY23W4soXVHdOjX75hys+YnYcs+
iueu3kFN+hOyHJNuDsfI0fq+xDhgKA2J9VE9Yici9OYMhvCfYAeeuqGY/CM3TGX+1SjRUNjoLRrV
Pg9723/uHiQXplE5zEqSX2XV7y21gg5JT/qoKs2GkfZWkZwASE1dGefyY5nMxgz1ALjHVXBPgi8Y
ixIySM5xjqMVWIdKURPledDHyl2Bd5KATtSjzGcH8QfhXW7lVn1KtKMXUY3M9qSIryhP0VNjYEuY
QFh5SEXeNzpMXVsU1NWiHGue/akajxz5co39LBFu3r8OIllwo2QxcQxSOSsSv3e+dUShXouPDmZh
jmxPLy3bzwp0voJ/7PONM2mddpZCC/x2+Fz4aZq0giA0zvI3TYzs9jLpJkelCZSy+yAlYCXpjSLi
W90VUFVXTXEmb68inOwHxDQ6het8NycagjoTATzavMrJ4E9dd5EspsyWAEN1prApXbVWnZGO3d+k
KCjGwUXIcRPVFd5BUUsMiC5yE32VAE4cqYqUtPrv9ba20BZCtGzd1PbvaCSyJq7TWROKIeOvlVSL
aRjjJ5zioe+95BuzTy6xL8nZ21o0Ge3GeENk1xWM8q8Be6xcl8kam2BH0tAz9Z4YZEzrk1rNR/LZ
WIzl/1Yqs7gsL3qUXd3BGo4UjAR0S0rSXN9rJs44tgM3u7FoClpZJ9MsE18tGc9rn7WxQ99QEj15
s8uBqXfQIQhcTrOSk661aFSgthzSg4w+KIo7LP2XTTQ3M3cgGsvuCjNKg3A6wgqw8OO8tg5cUXxS
wPL8hm0zkCopgbYdDf694j0nBS3dhIPjIf6PlsbCfLRXsaQoLeL9rujNLTEcvSrQMKpqGPf6Sw0h
xFvBjUoiYfHnq/ig9YS+1fA7515fg63WbC2C1qxFHhrRy06CRVhP8l6L5Mqv3BJIJPqEY22H52sj
6iQaCPnLKgrI6YOw2sptqByMdblWcYoB5Etev8pb2Z6+5+aBKGB0YgAURMHaMwjLho1tmFvYDZZe
nwZwPr87brkC1zdY6J/lLqthIpeQ036/7x/r5MoGk5ZCKE9p+C14gpy3dosEuLBx8brnBDaVVvuS
yDFXM+6ID3Ik7pMBSExTe9Fc5E+OVtsyVYpyplua0d3+eqPLaEEg7OWEshY7qiPRrywowBXFpgYr
LDHaBEDasd4XbMaOJbEKFF3YzgptmqB+A0veG27t55YRls4MOBV80kHXdq4zj0gmc6OhylchWrzS
w81QF9zuoaf/IYSysz2NK6tpXln7K64uLb6EyiqLdZwdQn+RszXpwj8JKpR6BWRapsVxNwLPhY6F
exyZDVQCY5sJXlZumqNLuo2j+Dzb7YE+mXu0bvxn9oEudxspOl2P15fnGhVp6pw90K2m1aNtJT4y
UhUy6K8QbOhHXt8uq1HyOlg+rvOQh8o28yFpWLgQZkAtTC44oQQ6ODE+Va0vQmAd2TmdZfLdAkMp
1opXKf6oePS9cRmHs5Hu9B+0b3uKutwe3wNlVfvyGPneEdmdABQHywG1//wQ/TpE7b3HYgfjo6oV
20PJlXDOQ6z1uI9Yyi4GPPY86bFDei0YqmP0kSrEgJAjlSDF8g8LLFaUTe2vkSC6Ow1L7mcQBtEH
OATO4BcDlqNHjgH3c4cR9xXzggzi/YPfVGvASxPxIXlCz8wYwvUnoOIfyBaYHglW8h27rfrhu/pv
IktX40092wiFXDJmRyNA1W3u00c9tNxkqxBbSrhzhcjWwjwJ4ALkPjmbf4awjORuwZnu18vA3ulv
9VW/8gWtNp3ZdYH0gvbFuzl9fzufST19o5rVOYza0vsusNm7OmBMHSvD06lnwBJ4doTgeUl3AqQn
xUHQnRJ+8H7uD9CU60AICObwgeprroPp6YeNBWQFhP5Pf2BfAzNbnIqrpaj/11MAZAc11+fqetb4
pHRGWziaRdnBFgXSpXjJj8lvsOJDbhndhe4NUPcN4yqASRJSH/POsJWAclaX8HBBY55oaHPRtjwA
NjVwkT4OvvrL2t4yuminPEoUWZ7AKJCHZHVip/Nh+lqd6/XaLISu5UHWxJfnhHQm0IFkT6Y3UH00
YAalJVwo8kQupmYtf7/+uGkJmbqTGY4Z3lXoXCWhiP4f7MPHHtV+dGeyAJIlg4GbAYMdJTH81G3W
Jlu2GcYyv/8WtFxFUijbNuc9X+7GbM/yYAp4Nigsdqa8DxQV7t+A2iw89+OqY3KuX/Cf98fA1Irg
BVKc7PO+eyFoEROe7gfQpmVCAPXHJsifJOgUNn+J+bffSj4whLIA1fEP4FASlSltdvIVBIGMKGgQ
c+XF4ZZklzUU+6NMDKnUBq8BrNVCd0tLVhv4pYx4O+2g+Yr3k9/CE9ZyPc4es47vy0VHfuqPqj+P
c5M4We7Ls0O7S6A5Xxt1McQ2yoEK9ru6xmW7PNWl0WpIa04WYBB4XR/aHR6ScI3I4xZ20t8sb7ij
uIMneuYsHHRDHfRLLajHPPhLdmOpfS6nQyEcRu1PrAdqC7EaKIzidk2e/zJusBdPUTyj0KbJHo42
hHWmpwij12rc55FqsUNKJWnXPdF2EusE84pwAv5KJ+n630CIhMld+hMs279wncq+MMjduGjDFLCd
imcphTPs0Ms1y2nD5ia/1mGh25k7P5NAQjyQPg2UKtJEfnI1YMW5rP06pq5lleYKDB5G8d6eGQXM
1xfvc4Qbe047YnGNUWaOCjlr4yXe+xMWNYPxg7qd3yDCpqvXoeizpbXT3B6BnTThlsDfnH6F2BjQ
XWaAuICahBD15a+OKxK+Lb3gu5n0KG3f4qQ5jks3hfrbzP/a5CURv3zk/lEhbXF5TlyFkwwD9UV3
MDlhoc25Go2dXGfB/myymSheyMBUUI3IMGwYJMW7Puuqr0b8Z1IN6GwPsgo7mExp2vHZ0M3G1Z96
zuCDVhg/NPlPITVCXwwOlW/64qfTQizszyezAomCUlVosZJKN+M7CD/m46XNxLtdYYVJnnZbl22Z
mD5ekX2x/xhWpR1zPXyRxhSLDM/E+JyL+TwJLPanydzAZnf+lr1BpNS4YwtCmsMfHbV9c7iI3gxb
Lutl/BX5gKRgnLv+LeQuwZV+SOxVe7tGfrmm17qqQaZO5Sf1rfKorRwzZXDgjWzMnRb6ujdH6nPP
6ZkmxDlW2dZEoU8bShxJjEIe3u9nDJdl/aMroc+CPJap7C1q8KFUFMdc5qajPwm9arVkLoNfzpF1
zdjHh1hHY+VDP0tBh884+fguNPClqGWp7+gmtzGNB1zDIQ1yNdI7wFLrDaZ1SOPq9aSs9LBx8n9S
11473e+b2VpqXApr2Ox4ImQ923mdkOef6f0XorLbd88j6j1BWfXZIVJRSqvXAE9LG0Grp0b4LV1d
P/HgdU8L7fQeu7qFEvfA4of1AeIIKtOSriWhxSMkMj5wqloa7JYQI2HkDAkZpxQIWy5zuvvfpb6d
SDd6bjccKxoR/FFprzQudOk0m6HnikSl3BEkI39WablHw70wLZwhX49KI9NDUypv5wm9JzTYL7oo
ZmQ84aZ2REyPlnYne4iUGBJZqq7KdiB7R/whU1Qqgo3loX6sM3UAXfD8IKHUrE6OrlqcAEFa6YMt
Rv0isBMZN4OgHONHwAWTIUAlyn0177m49QwrmE9nSu28U6fGFPhMyKb6+ZXUmlCzlk91doEdr0Lw
HpovhnLj3ZC/FLXh6F604FhSEGwgscpKMhNmDdI4f9VfW6+XmC/1tcVSGAguq3u+fwnI2hpAP7f5
q9iykGhL5c6iNv7Zk3dH8enKNA9JsAMemNjCmndQX6V7VFHLGOOe9wkbYN3W75FPFNb82k5M8TNg
SVQwbSSKktQehr2+9RrPLKKiTkwr5Sn56FR++TOvPVODs01bIfsdEBbhUicv+E2pjRttuqB0MS6+
HBXzIEORdMiHRvaJfgTvYqMLoSnJfdOInglPI4nY4xxsvUS5zZi5QaShWZfhmYbdNI6Ru5cDxVp+
ZrppwmOXL7iiJ3bNOsCduDiydJpMvuwfK5ZNZGTJxN1dh7jNtX4/EAhm17sYKVWeHe8id4l+nbnw
yFIpkcYs3w7xXSdsPLF0cEU8pRXw7vn3IycXddiDPk0PZQWH1iKJpU5/lzfKFP8cJYPYNB+W4Yye
SjOcnP50L+3vvYKnMYL5BOi56j2LFI+wnD1oUdLdO7AWtXg96k9Zl9dEqe1fWyKbmEtNcre3XxMl
3F5c4kW+4+E9aKLNHD+XGBfTfbdx/B9vLw3Pqa/d47QhR5oz1+D8m6uPa7pbbNvORS8o6PwLtpuw
pm4ZaAveZL0LLx7ZdP9MLdjgc2ARYGOdruHSHIeTk9ES+g94a62Ie/yug/ApwQeP3dUvfzaq/VkA
3QMrefaSeLU33xS9OajIwzXbAy2l9x/lk38Vqe3IxHYbhd1FsJTHWHy/y/KlggOzp5lu42VC3U8v
gAuihmCk6qx1GVsJ4Rd39s7P8NB7G3PVNUJpJ1nyUDX5ooFDaxRopId4hQ+8ln+cQpgJSAVGqx56
S2Os798m6Fyfd0WUu2BD+vYn0LEKNAqOMkP218fzgDeD9/7Pxb9oZBOMq1OON61NlZbQSE5DGdTS
MqIYTuCcCQfbh+nKpJX97j3FleWWZHivTHQvolnozCeLbb3N7k8hTiRp9eqHW2k11/5HIV9iUBel
xsnnGqzOD9LYNxxL5EHDwZQmS4dKyvl++4kmwF4iAu4KOqMpGVwjjPqo8I2o4s0XKngZnNDapl7l
l0OxbbEu9ud8Mx+R7XJqbRa482Sp6V0i428HMnLiN/ujIxYL++WsdDMD9i7QAU/GPESG8WX6FSNK
dh4L8lq5bbYKWuOifgOAahYZlvn6gOwzCOlMGnlozVa+Oop/2zCD5NVvd8SfTycjt3lz0Wv2je2j
cK+wHji7iEAZA6Yt/VWqsPHEcTrSKsBJmdj68yz+SVj1LnKr2oFMUA0IWswAVfyx2x5epZPCiL/e
zxUX0bj4T/qdNzDQOBhxL7HRJjr/ZoB/gE2mYYk+3l4PZH3vIQiIxc0c95Go+AO91p8zVxCOOvvb
bbX8kY736YM6wGN+uyxfpm/txRNjQp9TttDA+nQZY0VTcmlnWE++AUfJoOGsT97+NorOy7+8dDlM
L5xuuIKPQ0xzZCI2lPpK4bNoeoh+988gbANmsEn1pNCjMY+pYOe4dKd5o5jYH9xFvdo/1FOSh+T+
2QP4zxY729rHyddjCuQJ+5phkTyXFVA8EgBy0x1kGvzEFsWrC3QR3Hvb9iPyJEIcDNr9p3PazrQf
iR3OZQisYU3OIZJDgcxVRYKL3dJhbFXhh4yvC3xM9JdExYSNQGGrAnPyK/dywEO7o+PWCVM70kb+
elDdSnS9BawwroCfHwFb4vfq+STYP2ryod6ONd73hCAdKQl+0p1rJysfZVK1Sdps/t7W0neJsoEc
WMCovVw1dxFV4vzUtl+wa5YJmn0E797RnV6FerZx6udd1n6W61iIbupsj8pL4cG8OZZD984EEdvd
BFfQY37vTlDwWGPAzq0Xt+LXwiXdQr3Ydl6e+9w5iilGchxGWNE7B/+JByzg3aL7qSO1YUGMsXns
9sW3JF+Bekb/CnvkfF3MiGhRdo05TyhKo0IezP0O8dC15+QnabGrAfiV6EusRlyFCHdjB6V4mK1M
3TmkHK29eyUSIjCe3XVkgO/O67m5yBoqm/ydnlSelwU08diA6ztcumTt9CFrx6mKAGgn5MCkayOf
X6K1X65SKSttCAX53a+zvDhAYBK2EfXpQsXW99c3/TFmJHz6vgZbWtpSMQK/mkWowcevB1j49oPr
iIIBLIe1P0sYgzdD/5MVI4ltrylrvsJifkQm9j4pdYA0dtqA+90Pg+LJa6wTmwAHDf8IReqycUea
tJs5niQou2ysR/oMAZXFe/HJOj/08VKHYLDqHmB4eHT3c7pxwHAR2fz1isXZ8avM8nhAs0W4hrzF
sbC/J2cw1r8mGusFB5f5vZUqygMOp34eD7JKMIrRdJ7TWuPkz+eXbbz4+23dBAW+/3U5+s39WaW5
VuzgoBb7ok+ej9okXreN30zNk0T5OVEnDkjHX/wil4RxG5m19+wZq123U6flJWKOD2jYaY4xJcSU
3jPJSp6xJOicO7dgfkAkdCevK8526QiFmEYX5mDcSTBWFxudAS9TkDZPRuZpYdVGdJ3KQJqnb2mW
IPZROxMrQd83tUtg8REK5MbwrymGKrCJzP6N3UKSGcHguf/Q1LllxHK8imv/LKvAh3Axlwl6V7U7
lhzZMs/ZuAuVKkYG0oHKm7hxQfXTMVe5wUkG8L944XDRe20k/ITkR/2xggNFdPfSlzCl5uPJ1E6N
qqqiXjoe0HXthPdssJRYBDuH/Z7ixnTsFxb/H5rHJ4IUl3dN5kwFh9/iM6dV54Gm2FEjTvwywoFW
QNyQ9OGsc4FxV/Qw7PjV4z8jyYHshTWRflnAgoZOfQtjVGBjw7EYq2ZGdNcyZSx9rxPOfSkTYqB7
ahVvVMm/6BcopFax2dDLx+/bh8X/1g2v5lwANDuanKCag/CsoaW+moih8ZyvCmOsoEeSIMla55hr
9kKHvkC+dQdUa0QaNnD6RgQbbq6X0+z5yElb/6T51r3Oc9Jos3tFqbfme+erBKsNiTGVhQdC35yE
/O7YZGcuk4jnRbKpf0cFPVNpjvRFO0SIjW6nD8Xw82YbF1Dr7yD94rNzQYWeu72K5b9qVVo5kRx1
eWjTheCsUrcaV+VINRjEFDo4KwmsiXnxKo2wh1Eq0WyhIhzNQKt7loxi4UclOQRF316rE1NCZcnU
VNW1C2zb01WZEWcA0SR9sxRx0YkoUha29gDq3izJGpOqEQlZgjZ7FhIetfnc/n/4QyXXIHEIIKhL
LV9G3UE98204o28rSQWHoR8qdoVtZ6W8i6peEq4ZFAZguiNVbQ7qzj8sJ3kMwhlbtfhizz9w2vJk
MuJya2LJSNqm+PmobfXY8SFQZNMVmzlaAb3r22aIQbNWQ8mAO8FUVfSxcySJLC8Nqv7aVrWcorPk
sMdznKa95ldbCH3wiEQHMw/w490iMwtyjbovZNcfSoqUzzyabQzsc2HfeFlvg84x3yLvs6jSY6CA
vMygKrV1H9WoXE6lV0PsMZFn5J9QQxes1B1tEMnHW3hLZTf/kaYaZQZPgLczGybWaOTeQGaP5O+u
wiLkHQ+wMic5ZxIO3E8zfpKUKL0UjFc2z8V3yzdGpMEvn1/7LSceiSLCNNxRfmU8ExUNJ87EwMfV
WQ19/9eVRtrclcfURic4ZO4US38au4Z2Ygaxl28Tm9p1UuTMvsh06StoPUFlrFq7m6fCR56zev9L
imV2Ehpms0beNbV2J0Hug0qguNP7ZIetSVRVPqkPi4WKfUl2WxX5GyDmUZFuIyTm2ag67CBcDLPZ
iqiGULWn0XKMfNEq9064Ejpdeo2V6+9NJsf4RfMkLWlyBGiK9jXees2P2dsEAV9hFBYg756Oom5O
hpaLLY67Fs5lVSlcXE80AuufFmPjEQ1fvdokoLe6tmK4+6zn2Q1yfgybIScUDfGDi2LtZV33HQbS
EnH8HT2wOf/DPrr4JVHyoBqMI42qDUC1YxTyM9udZTgNY/tPVnoWa2psr9BDa4CyFLEmDddCvgc4
Lmvw7FXz6Loa90VNCTbTAORtNo0ilo+53BcAvKxQkkTVIRFzIBVejPtAM6vNy3fhG9V5QxZ/wncJ
nzP/5M8Fr/b8DYOy4PJSaJh2dBP/qXy0md0tfoJZsT2rjDFE67epKZ9FCCylZlA2Nhc2uRbb8Adc
oeysWvrUWdGddTwBLe+0qgRDcKUK2+TftWhSFV64e0mgDT67yPJf1ygRiWHqiHKdETPF4DP6uJ1D
ml3yPprWdkfIf/Gdwbz/O4LIWta5RAjNZuax4FuUYmgrbFjW2kMmfLTRae4AD5+nkpbK35//dydf
TwZWR2Tb/45m+7o/IlAz1TYRlrYRVEWcyvs0xmcDln3s4P2LPEP0ZxxcUDpfUWIrEBEa7ejXaOA9
1soma2hgTE8bDpi31cMjxex284spgQkPKwqAIy3PQT2io8/UD5o/bzGLeU+rJ9TsO1x/wGC+b4+w
6nKW7mG8KZAK01r2mxymMFv2sRF/WXuXhxqeUhuiqMJ5yaCpBP9gAybOMxRoQSqAnzQtrkebKRrL
J1/yGQ3P0UQwFJL51W3MkgixLC84StId3UiH6ia6/bP71gUnRi/W+5QjRUQJuXA3/vxd9xd7tN1f
HhEWISLmh7x/si1Gapk4I2tX3gRO5JLnSmtYs2jyU89E2mT7Bp8yR7f5W07gB8US0UTVGlPvR71I
Cx67+V51U4ap4mX001Tq3s1zrBWsGzi89sseVqpf64fCkNTOSxQmW2QQtDCBaHOmlYbwEKrD7BfX
eTK9EoB/i5z59ffSHgqyWniNOsWr/X2BG3E8nCYsVhO3wYtuNVpRXHSP1WkFQFqSZkCbPGh8mfTu
YFX3LThonfxgLGKV3G6DcWeMGbxMjmCcRCYcMbotV5qOf7MrjssFubnE8wkfcLk6vTHEB2KkAkcu
+M+zhQEppuuCPbyjWncsLFsjV0rJb4gBsxcGTgT9jchZrSxMLalqCQCDxyhIUm6BJiJfPIY/UMln
s9tnwBP9C4jIl8mmgmsPS/EfWEz8zQKB4Pe6NMFwYOTtmh0PMEercaIfK5WkdJ0YJ3ohzVymwQs1
2dwVsw0oahGHaWUIa1EfKUZ2IDfQgM4Ly8oMM8/zJNWUal8vQBzpesB4ylIlJwsl1bgJiYZmb3sK
IM7vJ+1KQ9YgtkUVFg2rDL7MQ2p5xw+vR/l/g+GlXKrl6WMOhqfMCk9yAvNo25FSaIb5TJumr4Is
bah7pEVBMdeM2+vwhiFou0tryKz8SQyTopsPLZvPYuZY98QVhJVOpnEabrIgXrowaVz475GUqjlS
JXrRJW6hxe/kraFyz00BTTBHWSXpPv28JbKd6FgHeTvK/zx8h1SIZegzogXNXSjQbffhOJvTm027
G9eTnh3p81kUGqTdTLtwx7slpNv2y7qe71wVHW0I9fDSZidG8tNGcKJgs99YSYhE5e2pSZ2zzEfg
SXpKwY88uxVfiCcN3MXzP5KUBiKWpAAlZ2xb9iz3yW2vCF0djHtqKfQVS/HRZ2MtCxnQEexnnw3A
H+5RGtibXM9infdZIGBj+nO/x+uceHhwNayDZJXJe6Zr8zpFrV/58S+KpHVjhI6fvGcdRAwAMxRm
5DUjRUtxgbAQFhuMJDtI8nU8FE+xOu2rLsimscsn3M0Yv0CTbsgzpdwG1ByaK0LpyQN7M3Hh/6ro
lXfhWp/xM+CBPgN8aiEQKEnJxaJ9F0CniJXvgg6B2WpaVg10/wKw51ml/OLnDIRyhydhnIGdngyi
sPShsR9SFqrFD8D+JorqoIfWu9I5r+ZpRbOqIX9Th7cVH4EVMEKJiHlIF6zufvuP05FMgt8KKQpg
Dm+J3rMe4veRMx9RxqkGwAAjUhwsZ7lZCBYKbWQF2E8DZGLhyA9tqvpxJsMUVYmCtlqtwL16+onK
NL7UTyT/HijocEeoKGd+FOPayGfuqYLv+OuV6P8VA8qe5oSLS10YjO/8EgdPw036bKqcl8kxOILD
4Op06OnIYelfrnYe3jqGb/aG14yOfh+crKD2rRZtpHMWjW8TPwiWycS1FrX9sYM9htdkm7Aul9cp
nGVBP769ARbCCf3yZ/fq4O0otphluSgArb4MT4NxquBTgbMBXihgAt/1QM8OGNubWd9zTZVTmK9O
y2kjIKBSbhmqEG1uVpQbBnadLRN5ld7CWR/LTKbQICcO3ByBE6mHUHg6NpxJh9t8eTtR7hgEVFCL
VEzHNWgoUD1j3iHhvxvK6zpqpHqcayCb20WO15UloJSUIbSwmPlX7LqtlAQUYxvs6ENrxb6t9gKm
DTybvHyclDetEovN/KMUV7AQsSiba651N2DFEk2mE7dxJxPgsKdI6Nk10hX1qu9OmiqfNVlhfsNj
FxN4rcbcuK+z2MeSAJYiDrNdfPVqVvSPYvIDZNQck8OaNaMEjzMjrEvxRnAi++jI196QHfLi3QFs
ye/6ZrEhIF5GsqDhTRM+oS05ZlcCqmGzj60LIhX6znGcybILhczsh7TEsUxQKF9yVu0BGrI6gSa+
l5z/Xsb59V2kFJJMYFrBO6fwHLUdvcxMAk8Y3cPnJc2w48H3VLSCdkfDVMtm1PiRpQCnXBnifkZn
AchoDCblo6IwjVQayMTCcWBxKVhO56jNVOIAZ9pe5aHZQkwkWywh+FwuBb25c8lqWVNtmui6GEH0
PDRfIZaI9570SwgXS1BX1O7fPF9x4JS7r16wBev9Pnol1hgLXndYp1jqV8c5/2NCXxKBW246wd5d
MU0TLTZznj6i2DPdaWVl3Fws3h9VAYbCduNVgaqjC1qf8xbYRfwxekw9kP1Eq5CCsaRYUZDsCAKG
SEvsBa+4aQNNvATVz8dcG/2TRI4E5odAW+7L9anFQ0U+BEwXDIH70LSSxf/S7asx8wpq365cFiEN
Qz706LIhDY5lQ0CJYDBJF9ZRhlmktE3Ja3FzvSINICYrHMgJ7qaMN0TLOLULeXc2zmxzq/YsuqHW
nUQ8SyXGq11xQlVEp239UEl+11awumxZmz8FsyInTsFmaH3irxmJJTAid2si04grdFlwH3hhn1u2
HuCSnAjlpGjbr6EIQmtLsuDifQH8bRPPwq+mbLEAHfJzEvDXLOTo28Vahak4BLBOf9WY/ZkPK2vW
dmIx/0Yek37Oc6dCXBfU5N7m1MqqNFU0Lun+yB/80ebS9sdr1sok8hKiGWB3Ef04Kt8i2nTcRnGH
d6f3iNtHPXf/lunKNAhcNcpodwg/k4Hhef2vcgdtaiEep3njjRzy9iO6Dm+pGvGVKw7HukXFKfXW
zOMg2uVH1jlJYq1jNtMF3gEde+Nm9YAmx2l84NZE5Y8uyngZEvQULWwr7hGU5ELlzD4LKgOY0uuE
+Qd+3KpJiyR/bnS9A1PeFwYNthZ4cSdSJ6a5qvYPLOjNcyTs7IGxZ91HILrdEe9/CXyYPgHQgKUp
zGTxUdTefiu6KLbMSH32euoGOOZCnxrhUdQDh6SEQDi82KE9gxDXTQFdDFhPY4aDUfIJfiDX9HRZ
rQxaYC7aCQ57K68n/axVOehIp7J+BEa/TdoWtTsHd8FPUbiztDc3pkbrm/7IQd+c1nKCcy8a90EI
BigD1SNZ+ZHBJU79x95yHkSKd5Rc1D6JmINtkyL/m/ze6GTmZuBcIlQFAfQBB2+CUeHh3spfxwZ6
kNxPbf7YevUPzCcBQkQedL66HknwIASryuXrmwgCNMVeIdvl861T5eT8B32cYYsL9CP3eMyOfM7j
WN7UqZ/6GLeephMFOHTGKA3iW7JMYj0ujZvAV4F2vvlsMrJ4D8Ei+X1DjJf24KjfNihVm2ldWRpv
xoReJZrXG715uEcwm1DJjkgEygGKu1fgvB4vkIjNpl2We4J6qS0oKkduyVKIYQtdin/KmSjTKuK5
5pXLOQZztCLFHfMMXqIuMjDOdFzSttb/g/H5USeBxKxTi2BNaiuozf1C7CE+JlhjFCEjT9Z9saJt
Zl6+k7jkpAwfONoY/pRQlhTRxZSME/bYi22++xETqt+E5XAyu7S+EsvFECYZ2BfFd11gA/SqJD6h
m+jXgN53e68NBelcqmVDWdZgD3rp2xC72PTOJpQ+chlKCqtMgm8PFqutNMaEQn4kYbEc+oGke8At
+ZxevYCxk7BDHPKGfNG1Xrx6JlpVe4bvSeaMTbZwB2y5lT4MbjCPl08IXBCzzuvg0Q5l+f9/6AVF
I5LzJ5Nqx5ag5UGueN1M8KewtLR3N1gRSKpUhWv8gFhYuBvUtKD192JhEKsMNj7ucksWRD6t2wbg
e9jiAxCbwrTpsotlqi6ZhpBCopByLE3XgXwQ6CtU08+HGfi5cj2o69wPUuw4iD1WhDYsoXcf/iX1
Pz6rdAaH1aD3celx6fwMb4t9PtNoT/BszLKuBFQN/iqGqbyZGyvr687c3yBN5rrX9FQBDXXrBxOT
rNbVq8UleYUFZsnBb+9E1eUHnFCi4p0mT3x+7lkkHcBK3bVZyqxM8qd+73wM0s2Z3BvriYz/ZcTc
fo3tJfpPTzL24BWY4MLs8MA3zjKKnQkl1pFwmv6dfVa2QriQ4lEzn11CJicKDOBKYsM5H3CFMxzq
QLZxOdo405L59aWRF4yNOwi+bZLATo4aCEy8/HQBrwn6nnPX1k3sR7QqrR0Y52yxhvpehJK2SulP
u3Ntaqtx8stmJbhGzJVz7km1c/YIkqCKGzfsE+5zvzJfSmMEWgHMGd3YILimQ09NHhvuQpANxNns
pMok7+XzBnvhx2MQnT/qa8fdT33yuWg1wISknMnyQzEJd15A0eFUZ1tlD1E9qUS5HNgPCQlI93fk
DrUvn/pCzoZtfxxR91lCxsfXpFZ1Q1NxYm+dZX9zJm7xVO6W+uO6w0Ted/a1k3t1lpbgYyQkEFYQ
L5GcVgvcGsCv5AZAxhfWyZ4RAssy1BQpevvFsYXix3oA3DRiMxHn1hNGb0I1cesmy6DqRB5QwqKV
kRWCCPEaKW4GjRYh9cI1+FS6qqMr1/sVsSQWc0zV4f/j+nbJYQ4POaUaBs4U/w4kbPzSasiLkFgO
UEOqaryq2X4NNFxQsAp3v3Mzw3SJCIvQMqdOTbl/8aD174ocbCBCyfZZBWpSgRabO6hxRhLulyVS
sEjA5TdSyi9vpMIu1UEgnltFyP86zB0Inr8MzkWe7W1dTkPrfBsokdW30oefGuNb4KqyuBPrmFbh
++rLI4FlTPFVejmDjd9AgpYxX1nxRjoTP5qAdarJ8Oc5ZtuC8S+dPvNSQ8hnyuCRbVHBr+bchrIi
IJoZQ81wei5gsdpnwrr3QehEWajJ6Tsb3dorTk99tySannpq4VvznGALUyHHxY66lYRDFyjWCIp1
qu9X/sOfipETTI3bubPxZmT3gZofdSbafGnmfDgWrSEl1nELP4IPvRxgbFj1uCa/MH9nqTm47a0G
ARcBk/65K7YI7pQ6gMzL81Exph5Ow84FA2iCGRQVmQni0U6b00tqT8hHpv9P+98tYqx0xLVpmw2j
epBbdzV4YsXSSid3//cZ1EFOtpXIG4J88BtqIARSR5r6DLi4VvFZn1T9teBrUNqWuYjFjvd0OxJW
9Yh/pJyZ0r41oykImuqhaRhnRDjX6WiSdukjihx6bJLGlmE6ELGzt9BlD14I8Rl3ceDxCw+IM17r
TrdYAJyrPtj9kqnyuat5RrqJ/eg+SR1KLRCyQ9ELFyAm6sXvhGkLtRazofOuSUT97lV95QiMHTs/
wl79fm7Lwi4I0sDK9TZAhowF1iy+8XdeHnyRDMHVx8Ex7QfZ0RaOwj0nSwXEEP9Lg9TyzM2fDLxV
Mp3ltR+0+wfR8uMbK4PFEFldOjWrefzzgkwmI21qU1tLKTQTWdOCOZh2MFj0wsdd7n2jLc393hH3
6nPk3KASM2d7QFMIliUDQxCle1lXrH+VGlSH/enD2G0wtpzneAs8Uz2iHvd0n5eu3Qu8myVovqV0
jqdOcgI0YVGqcHxqLDK1bFpnDb95v47iya0Ambvzw644lL8QHDr7FdCkNxOOZQmvkP0cxDyyC1id
9870GXFw8TcwAAXd9DGyLao0H8jzK65DZjUhgyoJstSTEy0NZLfLvZ9qI2ku/B/xbLl7BxSLxqGL
MtdMa+wgICi7OcowsRY0Sp93VwasNI1KV9LxgZUSXBPFFny35ilCOGxISpmdRKGyB0Fsp47CrLLN
nvdea6+SAYFpIXWfeLLaOkuXmVp2iAFOOjDB70GduVLoj8Pv8HoGcLkQVG5IQFeQL9fmDQ8WAUCg
2R6AXVyiT6vFt8QVVc4+820V2O01KuYXGQfSqguEimZGY0AxhRKLLFQ8ZgXV1Ykv0OT74lyLGOLZ
7ZAi1F/gIqD5kBsPy96yMku/DCh8HShxioNnmtV27pJmJIWPTFPkiuJuKVVVEA18YMXLxI6f0eLb
dmBexaXsxwtJZf5t+D+GFpp3OD9d3deVeHtUcty1iMg7rKrdT7lMkQGRgS44/F6rpfwN+72z/3Fe
6e1s0A71WOwjs3xj5h/eS0vlJiY2FMMtpLzTTrBa20XIT84UYRjdiwb8wHhlhr+x+rlkJbYIEOiF
8ZTkMNt008iiMDvMjIbz8WUAiHvrydX1e5pURV+J4O9Mb0o/57rVeSf+rZiyVteaEnNkiPuz73B3
v3HxD+JP+vrmO2HfCPjCCU6jHklJaquTiqOXFWZnJYqtUzazXxZMEYCdjhj26fGOpBVo/Y4xPGIA
FADk+i4vtj33R3bct9BotEerOMUFEV28C7eaSa3qKOJDmozZB6bb81D6dZnlLeLLKmuz+WHSVimT
06WusSG7y54IsXZq5DrFCeojjliIhSD8ExOlISWfKfoP9FiGo6eMIt+uGFplXG41LjH43fmQ33Nk
Qd7PT6zHWieEx3oXI+jxHOb8GCFzpUao1R6kefuZ5k8kzJTemwUVyesVHmEDJlUsbcl6D7UIzvB8
zaMl+CAA7aEYsA/gUiUsBnWZ54EGoyKbwcasEBnI5M2Wgs/GNF7/sDFWvdIZdK6kYAjd2bjeQyFt
olg6dY3u6yZ1CYM1kmctQ9huaE9KpnuO8rZ0fcFQwtNwzkSQ9x2wWS1LShiE7bZNBIonbGeWml3J
E/cndn64NTLI3xrLetwcsPqAjzg7FTvCwft3FviwguB9Red9xJQkVmYdVRZRjeGg7TfoC24BNNs6
soByfX7K2mkLobnIj9aGp2F5yJG16vF7UxJOIoIET1rXJzl2aLrnP76csxX45N2ShHtvp81GBdSm
5on06dNcLoNIppdRJDOqzZDjRcUjMxP5EwOk4fvzvYPg6LPTQWcMsxp+kq4h3VzrdSmMAzK1pwN3
oPIrfspfZ/WYqhRKTGgNCHvtgnu7ys+X677IaiRSBbDdnRrIBlN3ISNkJOcvYEBf6hdx9hrtHKI/
0Cv99mTmYfFrKCXsSuiz7mKLzPJ9KB1SkpD+QS55LTVi/xFTdx0TTKIFtIbx020bqhw9JEBsF7vY
1dOOHRLV5Tgv60AMlATcsyIUXvxe6inzD+5HDrdtXvkjEe4zzFRo8e1G15f4DCCMLpgtu6rKVP7B
OA02Jw4kFphgMDmrWnF/MMu3leN9BE8r8fNrw3eWLPbxK0Y3zvX62P9B9eA87qJn33YA8dGmovdw
s4WGoAPSh+LWvKw3u9/bTX8UaRgxhvcozeU0yUIqzar5EpFclWzftmjOSaWbG9WgsDqZNhI4pm2g
7CQ/z8004OJb6IVLj1rIs3nnVLHO6AM8I1P3+l69rmMNxPVh1OMLW8Zbjki82oLFqjemQ0Ix6elY
zaayHKuXtxh29ndZP7s0Wcig6rKnYfhtZFNM9w+wUNy4uZ6AwvxOOKwlUBeuJkxkvwnD+4nRGVBU
+qLqLIcIngdb7UABnNV044hQS0ds1BQfNbfHxSaesmAko6RZXIyrxyDa+PBX8CgAIu187YhJl5f6
aUIB4m6g8Oa47mcd4hQ5uMNVwtniktYUISJ2HJwu22rez6Ru55MSV7AunXUUUsI+2RAkog4EZel6
ZQw8phSPwPCGzWkIyu++WYaul1v+aGS79rJuuvIVkNQ3OswItROwOKPHTzr4jv4d9pUKttKcUIPq
TZGi4wxtGzoLEfXRKNtdfeRohrbKlBb2HOZoOSIjCS2+mRPsj9dP/PVmTnZv7xcel28zxGNhVvly
mVG9vSwxT+UjzbRTfQL4SLDlIk0KTXs0rXspEzHE/cQhlxoRJ4pIUmGJH6v6HpPsMZS2mWBOrlz5
Bw8B5KLt0wi0NiVbWCs89Im7fh1xylKXPxpBgrgGClIxRPakoU0S1JDzorYNjqsLQrOLlQ0R4oAz
C3S0RYCmTmTnmx+hUkNYcpWW5gt6FufxhTGi3ozBrA3jSasBaKpX2mPHEN/gLJmizbmgG1hnelwX
YeQ6ckPkVhU8xsjt3YBA6KPRbV3Q4HZ8rWZXW0Vb2/kBIqnWpJHgF02O5K2E4KsNwD9Rz+IfQFiC
JL3jS2R4J2SCMs3OszW46pQKVwtVNAP/qRLb3hd3xLpWANwOj7arG/1uETItKCI6/4NHd/+2rMhv
YvZDHPeotYC9/h/b5LK/GUsRAFqOYnDmY4nr94UfKWl+qEEaCIWUa24u23UCrzR8ZKYRIuWCLSwQ
XBBZYUcrF0YMu2euOBaHoy4RqtPz+6mWbxHp1mQ7hdcaOc1oU3t0wLO7MGjGue5wVvx8pol771it
vV4eb2k+HvoR8bEu/0AsrBGxDogudG6Cw2hgFeuyyla3GjwhDsTqUBUTECnRSMH6zK8IjwZmnlMf
wS46I+ViEd/BfDx2egFl8mCwcaz6HOfQflQgi52z5mYAtFlrdtObhAJo6twMN29nlXk82xWGsdQf
qWVbQT65pPGv6jMNszlc1TqpsbgnVpfC72yB5V6doC6p0flsEIe+ZZa+iMBxG59Bvhd4vENmL6vt
co43iY+bOm7B7h67IP6HLzciUIJ26J+mHjwtYq2bmXTai47YOKMKkUvX5cSPxfziakXagaCHxFYc
vbq2SorvYdWN6qjWCnlj/JbbewBftbWhSDXUn47AlpPIcWA3Y2wLfIQFWl3vZxM6lH4CkUyvt52h
JQEz85gTTWuzy7huVzXaAdNlLRQfx23Dc6z/hnku3fPuwsK+9E4CejGBzaTK/cmPmb6pfE0PqKra
9NXkKwdl7JTM8kPpLz9XVL7wg7Mf1r8OTXhKpJKGyJ7MKqPjRefPVyPX2unPG+3lFLSZv++yEAt6
u/Bdf7w9jaVP7KDq6PQQXBHvGYNsYcs4ZapXwGT+i+tuzHUa0EiuMiArDCz20cpR/1gSRIrUNbTG
D1+In4g2O1gKSjxpYUNk+7tb1MHU3agqWalpoXumolzlxquNPrGMQifAI+djXrKjQVlKFFXgITi3
i68W9SfBQ396GQMymc24Vfto/mrZZdTjeCkcU456kF0DYAaxqJgxtDg/1+0Le0enErGYOUDeeW4i
FVqxIt2qzvCYQSgvkS2XKOOYJq0RY5/x4c+RXInsz880xwXV+kEwsLNMkKSNvZF1UifIVT7kxRtK
+/ADnueBTtdvDfQLi2rlns5Pl3RiZ0d4KL7irwfme39wXp05k7mfpZYwQAAdeOnx05TC/kbRp7vq
2eovCH27O1LcMVxuNlXx0m+jyoHxAa0aWuuPvVabhhlto9/2kgcJfuVXH8bstj3fAL5MYB1Zn70+
5pxqNKmcySk6M9Paew6/LQ10zTzjhDbCzNiOoflzYP3HIhokXdgWyqMvna2uZMTCBc9+HzJ/85R5
IOzhZZPkNy80kGEqzvtPtszl4agCMd+o5OxTOi7jt71BSJUCbQR40+x70J2TK65yN2gGmNIjloCm
2eTLIeAKihWVhUH7uRW9JSZWdw==
`protect end_protected
