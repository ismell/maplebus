`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mjgAOmmqpUt1V+Rhx55PcsZFO50ANSJzUkq4iFT2ky0C1WINgCoS9aiI2Aoor0/FtBYKfc1lhyAC
A2yQaY0u8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gjwaSbcrNPL1CjiRK1olSBjrq4xEV61J1xGlt5XKQmKd32CsZVNRVqoIdIOQw5EEQ7uMTa7bpCef
/RRLmGjz/2hgGrgTwg5h2PJWHguc12Zs6C59vtsbmoplQOrftqG88iqVPmgqwLN+DTNOr5arrhn+
WjYZEBGst63L9iu3Khk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q5P6x1wYO7e2baBau0ec4MDS3ryR2YzQRaQhrf9aLeN+93m5ew7UeblmK6P8em0XD3V/frlrdjJr
vuNgfu7erA60Vrjdo6kExSAievijk93kh7MPyG1C7uDY1IKWawOPN0SnpTgnKNqgJWNP76YGs9dE
TN9mEgH2ADzwBzmsnM6NspqqEoZYVlXfQg9prMYa7vubVhbFy8YrYeUJcl/tvgZJjPwfOXGv+Ce9
6Lw3eVnbpPe/UcdW9doBauijqG3ME0OMECmmQVx3tDp7z92dYCehkqsqs9ChFA/rMqv7yoEeo0Tq
fYW2vFa8NzvhoAAn3MGMFPC05Hn9sO45pG9MOw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PhhRJ5ByvCD/sp7jeb/K7V07j0XnHI1QE90gfVDZlyBNRsnsijVbOgPrfQFzzQckBnxQRDgodqBT
UyEHG3baIJtqnx8S8FzCB+ms7FHJzH8qYiVcrBJbki9Cwu1coa+dV+gcYK/TykBXao/zKErqGGQe
o5y2fe4hLUiI94eeeb4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TAojQYz3bVMMZK9Nx5h3lda3DWpTQmZ9NPXuNw/InYDrG2TbGUzW6Wq6wdSILd3J4wAwg/M3zRal
0Okl56IhevBfwHBHR9xLcke5Q+fEjahGlIEiyHBXondVA3F5GQ343Sl6RxPF8lzUTfgXL7wJx8A2
SjgajF3hMQRocRSQ/AaGLTSAnfM8jJN9MMLQuNU2wvBRfbi8VZAqaKMgXz46LlEZJBasUpbtUHwL
r58zjjKIDHwYMrOB5SRbeeIszHIzYGbbXwuaGXoSgqoXST3hebuwdA7H0X6lL5AHQpXSqppzPZ6p
S9LM5cjn5dm06YUsC+fTFEUGkdx92p4gSMtILg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
hqWVuul9hWaPcg+Bmj71a5uWJgAz7ISsZeFhHHprOy3ttyKtQmt0NlGaWvBOwbbDSBGw/XDieEHj
cNaDEJid4luXvGZX7cDOVMGF2PDScXXbv3NVRiXO3prdT39xvWq1L7nDe11NLwMQ4rtE0WbjzrkX
QFacVNCry5HL6dz9TmcXk2aMvdB1kw2XUsFRy9W+VORpFO98vA4NZzMn/7zY5nHbBPhwWUUVDI6g
Zt9xeN2Mi4dsuCQSuGaKaGh3r0IZLwrehg/kYTqRNuBdAdIKnUzAj0HwNAL9gTtcQwdn72hTDkIc
vnGjFV61w6NUnj58Nz3c6clXOLZELvVW4y63Gw6zzIA7oBwpUMNobEANKn9rohFNkU0eXMIVKITe
vVXOTUOtcutuH/TeOTw3xhpBqicjAFt5YknGat9Sq+C91utsqoBRLHWo7L7cO7HHQdN9Uc8b/GXY
J/qjW0L5P927N9mAWNQt/ESywLjjKiCX9QVT8DU7gA5M5jVop1LZErBldRgI8sQ0KEcS9ep67WCl
wotHX8M/VKQOyJxEFHXEbq6YaHkM4MejHzoZQWYIqSRDbhou2Vz4Q+xrR8p9ax0kP4Au18WrwA10
hI4gA73RNxy4N1bGAGCkfwc15tNBVBOLsA+rYsH373AhbwBSJpzYIg1VUXFWV+UJ1fC3NaAZypqu
kRPFSbNPX3ZkwSLkH8adP42D12I54rgjXE0eh/F3pA4s4tPo9s6x7QAV47oJjz6wKHPRiF/JKCuQ
SOynBPmqvS5Z8JgHaSV2YwUbiYQvLb/m9Riz6SiNHVn/KbYGB9Kbu6FVQKbx4sWJyalzh2WRtrnf
g2krP+ZQviYrIQvjDDGAxRFOJYqAJZrKP/wxuZ8SJVl79/HUQvJXAxZumYruZSCJI7bFrJMFEuec
7b8V4R1ISCgHdqFVqv9jnsNpRkZLL40Xk7yY9KmBSWF22a7nzOBOuBFjspq9wlnZGgOCKk+Boyfq
I1gMz4w+kiq4pl7YGDKEJsiWA3SR9wjghNQ45JcernzBNmHKVPxj1xRBA70LX5tZeO8AVvVZp/Ob
Bx/T2OJZiNtLsyYYRzFxWvDm0Oow7l57blWAamPDx/507eMgHf8pgOp2UIByj6L+BwJu21mc91q7
Ftq5Kn59AFNw6ICKqJUBQcEThHxk9psVd67r8BqFA0kAUS/B1O1e643LW8r14TK7Ur49AGsLdqt4
+EW4lVxn1M01ATOKLYCH1+hM6QxowHgbYheBS+CZNZK30UtWyQrCe/ndOuU8LkePy93ASw3Eyflc
5MtKcKYw69CQyyN3e7qrCbZQkRnxulaFDlFNXeFqBHhTXBme966xVYhTf8Xe7ZscN9kMnuv+9Bcx
dmtYPLZhBQpBDZuZvu5GYj5xdnPU9UxAAuotziioooiHhj50HSulrsid5xFglblYUhyU8EgFsL0+
JScmOpcR85k2sQFycVoNDB8gogZISZk/svoT7DqcHeGeRYP2NcAXTsJo9qYylTUHGPdJFWoPlHQH
uuqM2qrJbFSrBHdWxuMUAZ4T/kEc5q55meNZBIhtl5pEobdndn+AfhRkcoyWEefDbf7OZvfwzdTH
wnipocvdvGFAXufIDO3sFU0U8IhRrhRJx5ALGhlDk8MScUNgNtb3WrmOugDOo2p/LtbHzXCaOAzT
QSHQ4VC78cT882hjYhIQWoAGv8qJE0Gk6UwWMKR+ncEkCghkXcV4b9zLTTunqdZdbjYF+Z0lmH4G
oGqePgdQOZcsnAwhS/9IZqDP3io706B6/kHBxRgtb6xaymC0U/86Vh2Mk+uMCK9Hd2fPF+adEBqa
+cpZy9YGyIxA6FIOX/49p9zb6Rfd0NVXlMlRLCzZEsgXzFbdEzkVZsgslDRWNL461AZqd+qaN43Q
OuOpebmWZTYCUDBPMpQzg9mdA/dfFZ2m8DJvx8BEXVi6XFR703bURrvvH3CSSJsilGRnCWc97pFo
Z2T6rPb1PSHwbZZL/svKGTtLhu4Flqi7ss3C2UfcUrqts8ZzJ8/oqM8cL4ujkK0HOIfzhlOh6ovW
9oB/DWPpHm179AcKqZ/F3Lv7ThBiDXzI+3w6+Gng+Zt8liHBWjJMJ5y9ZITMf0B/c+7gJxKUu9CP
/FnLacn/Uj2ohzdqwgZoFE2a89E/D/p2MfZ7P24/CwZqRxLpk/H4bkOewStrzOB2VeZL35rCUZL0
2Xomd0v1jPQtDD+nfTmKUgWUQ0sh51+2OLCG+USKjq1Lf+LHiSYM+TItM13lggi3sJxYNz4hbhwk
Vz50xvzSY6iQ48smhE162LaT0nv7Pnanc0BGotseTGHW/uxx+N90OhZc4XOJc2TMuTC5mhfwjhBK
smJz2/WhqFRIJGvq4BkMAu7wCEBCXzNLzOXA7dRw98by2lBoc1Nc5E3aen/W/qBM0fYxGbM1zRhs
tsjMDd6xYaTCs/8wbUUhEkc+F053gO72hYPrjrYNNwRz/hY+erPvRSM2TYWDuo3oN1DeqVmnkK9n
zWKEeClVgUq6k6Iixi7JyqZh+A8yLSc1NOemWdwahaLZ5mRCu1u7TRbPJVv0BTLIzT+fwj27X7Ag
b06VBTyeUc+IY3NuIRrh137n2R3EpSJOF0/uiZMQQIp7J/61h8jPk53tkcfHYvycVbGtm0bl4Oxw
MHm9fSFFUgSZJEkWKXlP/lmAZxh5fFWuXPf5oIzzMV9v0q9nXF7Y1DAuXqY2QnbpemVjW6bZM9kR
ypMp2YPA3pB+trwIL/VD+onqYgEzzVYi8qmqCe76OBgIMfWUwQX0hQ8WaWfCG48+4hUEneHU/laJ
tyrzdj3451EiUZbiZaFAWZLUGxZ00xtljEaa1d726Aq1RCl0CgY+zxh3KvFxnzPwdKm9m9JebIIm
09uZOhGOLXqd65dFfmH4JeyIgwJNSaKYgge94g2vSYikEQTbNPK1Q9/HsbetNJE+L6el/YnI3xi+
Nm3+/Xl+YKHPQ6uEkNhbc2eUgGYMuOVK4MH9rD7yVDQqLkIifO9PYxIwvafdCOH1U9qYS9coxzAf
KDgPSdWh/lMbttjbmg3nQPLgDf1R+XOqsbizO2u6HDgMWOVum6FxLjjb6cLTjIOmj8ou3VvYkWZD
C+SYR8qU6C8rWzNtbMXsdnx5MujaVdWry6xBTA7qW0u1ccx1cdtEI/HXsxETU/aO0xYxVT1EDCdw
3f1b7zOjxSVsklUDdei2shBubc7kKMLMszD4NCtyEf56XCI5NXlGqYD5K92D/e2rBuVP2Ab9cLIw
ZE8Crv8pBtb1E8gcouarxuejhd8WwtSEa+orb5CzdO7wealpl2sksDxUWH6LBtMn+xYOjxH1rLD9
Cm/SH5y/+mkbLL6LhUZKqei8eRI7cEpDfC4+IddRCZxEGPX1XZOt+keMMmNpkAxSlctkwNySCJfM
WxDDK7iX0Pu2aBUginIgYi6kmtpuMzc55NjPVt3utkVds8o18BtRKq2X0N4Nz5ZqHdqSLEhLxCVA
L5Te9Y+xv7Us/QiMvbYD+jAXTk7Ypcm7xKyfBvh8cokKt8ZaKtBMJ3oqNHvU+VgMN74pDa22zBKi
Ly/woXDMdgPLFYQtg8xY5vyizwWfSLwJj0p3YBFjRa3fKYyRboa+fKNk63RpRq7JK0+Gf0k5mBlT
338bseMdkxzpoYdb2YrMqhwgdb7fEUZcx4llDqq90Fgdw0zR8TqlJWwZWaOhzPHERZg11qDV6NUl
QF+g3PTM6ueXSHrzsXYcbc5a/mEVp8RpFEpNhqiZ1OehA1CHkjypowlJmMxe232hNDar2wsY9uB6
L+IkonEUyWcQgVjEG5yBeTQpInipglHo1U2AuxTAcoQJxWxcQzOdOBsiqgJezm74/8VPz6KeM9RF
gC61fSc8hA7fcaBaJ7/eu3kZgc7GVgbBvYuq0GOxyoGIT4ACfs2g0uZ4UQ8uCrLQNkUAu6kN9F1U
1EfIA9xFP8hRxg68Maehe84Dg3VG5Oql99kz8l0XUKLg8PjZ5p3a7HeEkbUdCMLCHWVDfvB8p6VA
XF+BIOj87diN4w71cmWYgBK1oUBznFXf9QMNwbsc6y23HVFnAFcPq2H3NjWiEOXE6IONbtVi7Q19
rTGS4S5bzPD4fR0eqOdsmoNEtBPk6KF6FqnfLjVpv9MGWtq3tmZVSb0uM64ZtZigo2jK52vxbG6n
p1pZdoJGufr9Nr+N2qSqaaaaibcMdX+mCFV1E1yc6Coqk3CRp/wTmG2snoa8oHgxGuN+TgndtYvR
wOYdKVWN+zfujAi0XW6iIjINt+edddiR5sKUgwSDaAybwoAqUf/xs3MRALnDxxAl9BjKBEexT1Q9
9r4x1BCrV8XX6ErsVm4TJwSuPDw1h5lxFRVZysp70GSF24Uf50T2jDJ3FdD2lNeYlerla/Z/PImI
Z/t6gqU/6Pwa2NCqfPJ4qrTfh+D1rbNz1zW88EAMKLfxw+/kbBokIgRQ07WdS0sNr53dQPq3QBxu
DZCscnf8Pvf98AIi/VzTxl39gv5seBkIpyCzb/RHPQXaJrf8lysx/LMGYBbmFS8JUUbimhvwuMUh
69cmVAzNUyBDm+xKUYX6Vjo1TGyeCBaHAvwdG3Zp8Yl8leAsDpWW2rim9DBBWs0NVknNrJscAKlS
yajUp085rjrWHJxJJ5rR81Leh9m1PBc85Z98Xn9IxDjVlMlWfDy+KJaHPQqQ/LNcWWTg1t5wiBB2
zCrSBSqv7HUo1ZKQ2mnaUVRoorLir2zqJCpAo3889yRKaTCQiDeogZlh6itzQXuiF7Bi5pdIOgYT
H5deZtGPT7Zol8feOlN9k+cTfFEvIgC9jhkCTrCYHHCK+oAGgPytOcNJYkBYeVk8zwlylFGnaLn2
RcrmijsPo/86hukXsUrij3DTL/hyIfZbojNSPeXMtmT7KPU8ceC35MAccqHzBl7O9MILeKeAuyLe
/InwxRiXDzG1JlHFhfU7prlpYVw2osJ7/CQZ5j4tC2YktZjW9Jl6ftYh91AoqJjgH7qDgKknjr3w
JDlYYUXKXig+JT2arc5/e1HOwoBu6gvynwIt8Ak3vTo1YBS8A5ZyBjEmXezixdNEe0/90zwG6plF
ciaYGlUqqo+Wy4KgF4+z4s0F1r4xyRsZp22x5Nv/XpZOJrYlWHA6MyGZUwf+YA7gyzchwsV1+wbF
9kAAT+ug7d7f1vn9pCFCZz4H46sThsDc4jB/6sdfJ0+pCARbsEOAV3DtKXG9MyIno5mmqD9opT0e
J+JmuRtC/mLrgNi+tOUoSFMiIG3PKB+Jh7z381HweqRcVRnlHkBQJouYs11cHG6c0TKsS8U4aTho
slp3scTX3qco2wQKJa6VLnbNEtad9pm9aRHrEZd2FhV6kUQTKe7SxxQMY8C9irr5mH+nwIgvZkEX
v+o4EdACVM/w1EaCgRP4QQoO/lqPGiFjL6vgQtf9sgHsftN4WTfbMmGEFijOx5EAi2Y98vxhsMmE
unjFpPiTxq6fDc7WPZGKPt08tlQoYhLyC0ndoMzzJDi1thUo81CL4DzHUugm8Dldfgg1CfU0IeYm
IFekTgKVCzsOwy0ZwLVN5Ad70cCZSyFkUwbSi4/OWMtveCA6+RctQQhtm5h9httep6Najgf6c3Lp
1R/so1xurCXbyeXH1lhzcYpPRT7lVO4PeKAj/jqUN6F0bnLH4DUkh3djkOf4DmOvJysL1P8AJ/yj
k7UR3+6h0bizHgHCz0nsONZsNwHgqF49RuMjP6hTm+e+wzyu//oW3hhadbGIWs33jzdMOFgQklyB
8iA/ShHBmryCMRvo1Ko7fYUMnE37+MOKuLwIgjwyYbBnBe9izlhZK7E10uPSLrm6YmKLrSxtDHMz
7gaBK/PfayVaB6tk0PwckuES34Railpu7THex2Ys0suQdRF4ZjhSdYpaY7s4BiNMt6x0v3VqnnOV
wf5PXoa8UN9CmwRdP/9doP5Co5xn4Sb85sBK7MsGXNwrk/8rign89ivZn+f5tzzhIcImiDALD4gv
qKwMIU8KGSI11ka49y1mbbtnJBoWPCZoqb3hHCsZJpgdCBO5IJCV6G5N2DFDas04SYPx5sJue3zj
FLPuWJpKb/EVSybfGGKgihJeJ8KjRlI/RYuZaLGttElFezj/HSR0sHlO2i65nUcx4Z3VUbJZzHJ9
1aCmdZATexEU4UEqDgvZbj0W/MZxu+zbUZM6lpePho4USkwLMbODlqJ8UtTMMlfrFvHeAHjtuzG8
Aw+N9bWHqSW0Ke7ugz/Kznj9lSo5oTEsxTsICTf965KueJaB+EXoVrcN6tq8FXjxuc37BNy6Rp9J
TMqMhtlovzINdllyTMXp3JJBF5Im3l57VZ6CEx+pwEFg7n10cSdVEjbXiDvOIKkcYPThrnRDP4CL
3ucjS94/h+mxpdyiZdCX+BEnhtfac1fAFe9z0ImmQlsujlMzjFcGsmfLZRduuYdepZCkK4tcdcAQ
7rxCv7/jMzaUjjItHbtYnfG1Pc2bqKHz/5AKtjVcOgk0eq6oLmCPoX0gNBlk6quoasTlyxY9Rj/H
GmxBLVnjAeuyHMAQdu1+s/dyfGwtub+wQU1DXQENe5DjvnNVpfYuj2sF8bAIOxXqLabuf0MfP9n5
yZaHqI3tjtLX12zupOMd4hZYAMBOj2SzrEKOWjnPqV/rs3goCdV0hcFmvgKN1S0udRYIxNjjtxIr
fNEJha9D6JLzqxgHKTpH4Y9Mz8DeLDu+NRuj42Cd7EHFRAkFaSPQBgQjf0RDrNKDi7sVYX8c2zda
JeRSWp1QfjCv0hZL9KQGG8O5J4iheiWvcHYD+9A9M7uwt89HU5tGFAGGrZNntpe2n8yGM/2a9c+d
dbiwRha2gidXTyxopnAxx9GZRXiZ/hxzo7TNm1rQzxDTzWvYHwDs7AlW57jUGe04DnCqNP8V00U7
w8EcPJ1Wy2tI9iyhdWa6PeYt7D9lbWR1aDCexeeo1pZEI4HAk/fOBxHFGJer5geaNimTXtxbcJcS
VGx2uJF09JkT39eR0MKwkOSJLr3e2KOJT3DC87HhL/TEZOshWMgJCBFQWsRT2pWaq7yVb4PcCjTf
8GhWSYzGAdmvzw4KiXq0jIKGZ1rnklKd7wF4DO+yrMjqgT6HXv+lOF5roveKTFa4vfOiFSB3NhwU
AFKaOXrG0Gtelrk8dCDTdlUguudvnvv+/A+ysv/RRIQAzviVnAnP+fgdsnj+PD3ZkRk0XKGZD0zg
srMaSMbUhOSqWNcAEIOaH8O7fJAAlBDAdj9LsnbLlAFA4OpwBKirfZgP6CYAxxCPsrESToS5GF8m
ljH3wfUvoMWmFtLqbPi7LLXfjbC6n9H6YWWIyxT8Jc+1cdi8E7tl4MI6ynazrywHsdtjWOnenXn0
sCS7kZy6eGO66VDJ4kbYmk0tJPt6hIU5VScuhRpKdJr4M6qzlcR/2KdiZQLy/wsHReK1mYpGCL27
7JT8uggrWXu11U+fFrRVivP2P0cp1dDM0I6bgLOYdXsdUMQWNbm4n18z8be0GxZ90hxn7AlfkE2p
0G9iYGhCOtmI0mIrhbK4bxkKYc/2fR6DJB+llk2NQT61AxIuBxbhIblEK80qrrpKP3uleU96GW95
bdWott4iIqfOYV56UiiSObeljwFYDkmWlARfQREv+KhPo+ezPWs665rf2fYzbDLgq9hMDtiOw7Ml
4Hh2p8RwIAeAKFQhmI4jlUU+pLn4VwnzN6eRZwOp7BWZa+mur97alQtIzr3eop0CRsQdYmn8Dec6
NPbGSF6OoXEkLfWL8kUjeoR4hFyyRE2Q8VFvRJZb8zmB6nksELgaCcOMwiFc6ReOw25o9uRCoo4p
2bS3HA/ZGzTUaXtAxb8sGLtZjN9aJJpOrTEC3wykH3Jac7dPYjAtl/6yefi6yi6HNL7vv2MBG3Sr
psV/dkIqQTOxJewTBHjUlPSsMeKPmEF9vBEX+FZl5rWlSf4KDHZ5bwizwb/OIu6Rs+aSk+XjHUDm
44gWXu+AX9mC+3GJ078bEIdDtiPsS0aNG92kEVHg/iasPRXd1dBHcZtS1RV/V3fTUCZyug4OgSfZ
4FvXLEkYR68JUqQ2pb1LVPbHTv7L679bltFkGIzmNN7wyUfqwJinII8iXTd+wLynBaQQ48EVznVc
PW+ngfTh2mX18TO7rs0Tg/HsTXJ2kKShf3QcHGnFj8TfExZi1eqcII4VXbhjnw3pE1Edy1AHFWHR
C1PRp97SVWkNZ73Ghauf/KljE9x264+LlmN1wW1M+eJkphMN1szZUZiVPpdmwkN4z4U3Fk6O0Y64
E6aQtngTCsgHw4DvMXDaf251ValGTA51hmXx5T/hAJwzejpbONVGY6z5xpN+AQisJSUCaMl+EOj6
oOPJQ1JRqJiJV3TMnEp415NdFuAi/X00S+GuZgVRUpR110A1xBoZ76uuNlbs1JkkR2nRXgZPgzR7
ei7/TwEo4vMzrxsJ/loZPBAgFl5BqmfSENxi1C/8ZfaAwUGykD7j8SSQYlQs6YecbgU0KUxr0w78
1kEuTpElqiHHHPaf79EGFqHt7uZdXTPavkMA4zRaSj7QJ6b2RS1X65LCOoWDdfVy5MXHdlhfB8Is
/A9as4a5UPTv0yXGMItV+ch7uR+V/hHg1uF6YONO01je/Io9J7bQCx844zNHoK0b3eCvIA1QffcP
mJqIaCUYc2qX5YviMS6LnI48rxAtGcNdTSC6lYoNQOj5rXwCPtLVmEy/k3NE5ECPDGEXcZHUO3iZ
k8M3ntUJfku68BAdviHBsuiff6vK1ypT4KHTMzkC3lAVZn0NDlUb/gceVnI1YnTnDms4JfrzD2bi
oYmCWOQsYrpA6lkfU6ncK7JhV//EGJRiAvXprKiON4aXG02ZUnZs70BxIiiTclY6HjqUzS2XeXsP
CCLkKsaz75qXV+gc8tW5OTWAPLXqr6OJVAzRKJY4bAfD+SNPDtTllg4BXrJsRKuuDlGr8oFe7f3s
mL8mYqrYq6wEKah/aLnablnWIjO325ML3IvnRgQ0uDY1OH4qrY9kCBTb0Pmz3MJR5bXLoikL5/w1
1aT65oC0qy6rY2zXTeD7v3mnUKONxY6gGygq7dPP8Mf79SOB0A0Aj+HkmPlIbtF+2IPSkMFHnxFy
PwMABh5rHYRsHVFIJ/vgjjThVGOPWOKSDdI1XUW/qTFbYXwF61EsBK+3xOxePbpL3uFGmIvnm6ud
6xFpagu9DANFpAnaNJs8fzAXMgLXLytl9BdeLdsIrOKymUh3+fR3f5K3Q0IAim2YuvUMnwBOYqrE
tUrNlG1VlrYV0z6TP9ycKuiEwjtBUlrcN2Qte4Ltya+IjDCGYD5k5cysbLHsddVMvxGv2zdwB7s2
JNkYuLVoyl0TwR8siqyfh9ppFVXQ22hQpHXjThSMnj9vC1ESn2esRvI+3VLQWkr7vTd3h8diPRrb
3PknZG+xHM/aHrNU06QaJ6i0lQe9vF8U2udEJc2C3p37XE1Rv96MHiHRwOJUa52Ml67ckf6hsM5g
MIEGR4FYe+cS7uhzZN/YQhH8QhThGQjfBPu3pKkZ1IAi5xIKuxhbjkAxN0wTQYlrO/8qNIljNwTH
qfswFgXkcGNoGe3hMO/VkboaL+NcHW1s1vPd7zAI0nYkKVl7L1tbtEqMm/d4kTcnJVJSTOPaKkna
Q+a71JnICL3f/eqrbvO9mY56KnqN1lrmFBWnJ4+db/KnGcsXdtD6I6z1dHjIqHnTyrpcfrGT6oob
x+Xzg5/JuU1wUZXprgiZ+xO9/LVntmKLmUrOWE47xO4aXIg4r7S9schkQew/AMEu31UXoo5HhxEM
ZDTfoyuq2NP3+RONgH6ecEtzTmRJRyTXAtoi8zisp6mBCHjjcBrRH52tM3D+77qWCW071LDdbEoY
AAXsDL2C+X9Ru+IMRCJlJXoqPX/hJyEEoSKJU1HxPTsBrCSA8PDXNO9LDEmkojBhDqGstMvouJsH
EAQ7KHTV3HsBwUGvrsUnk92FXQRcorQSwS8fKdjGZlgpjdGVgpIFEiX8y1/zjhKqJewdhtCgIPNy
Sdz8NlhTBdo39FC5fWCflj8U9VMCNBMwHUGUJfpPwSOST/yCZsn1p/49eQKuIugZXgaw9vvrH80M
YbFpXfcDuNOMnuPIf4f+gB31pd+Yl7w15rU/7iAQWLq9NjKB+xa2E2KbZi6QbvGZp5ZoGj48Z2wJ
wRnqF1Dut9uBgvyG5XAj4YGxTTgzMW5Dh0DvCkxLs0BfSUuVYxGR7y2eRg1kOvKZsAjHopIk4upr
DtzD14HDvkcQsE7kdFFNB0pnlRyhUr46qj/aaEmYjbvGPyrMPYfuUwYWFFGySp8Tc4e2kz7zdJD2
+qDjFRQlxdt/FWtNEw1xh48dMqMyXj1MC3DbnHwaIgWi05FgNsM+ORAn/DJFxPK+EklioG33NVlE
tTh/CWEXb5rFUSwcFsNDJp31wzSEHLMDMLAA/eqC1EAq+QijA5x5X2qTq7Zc7L7G721PNGmtys/O
jQzJhcf7JYLSeHGXbgerKt3Qqa+vnyI6TAknGg8Jz1284SR1U6POQp2lC+PpzdOb8QDRS0PyyBX9
TELdxVLMJRjqrPso6Cx0Gp9y+Crju5POI+mjFhgsYAQUKsLESrszXjUfRJBDV8JV27tZVoZLn/0z
4sFzsY/w2NEB6JLx7zhRYT+51Qz6Da1t7qr6R4PsdVVmYXohwolHw0FKS+NU2BfYteFw1FVJn2Iz
QhI5F7qk2VU7o8L1IKtFVo0l9rMctbrXW439ZzV815TIJBrOwpOrjjBv6EWw1OTjVLesgBGx5a3+
EIZVcfKR/YQD0S841wniDp3NqlJt4V6xjGzx9oYfptyqT5TGtQ2GyI/k1i8BIi5k8V00RgOxsQGU
B5hj/H+a8/po1TJn7a7FJ91Ri/AtC7WzrAHKyoq42c4+tbBKyXLqT7IuMAMPFoR/VhH3S722oTYg
ouIebz+WNmgFF92sa/VR9qdkpgXwsVxGT8CEGIuR2WEs/Esl8xJM29iXdYSykb96VZfiF+cfEysl
zkkZ6JpfG590facOSQvBOaQsh7zJdYAfbdxcQs6AKYuGdClt+CtbzfgEYqCnnlsqsw9z76W2FNEy
4L+pGEOKgy3M89UDPiNFsfbAzlxKxRzwzDBvMTnjjBIBO5oDK45Dvh7ku+3uCgj5C2nmj0U4PZ4Q
kTSqBtuar+UzTsUxBBvWnFZbvJX2ijr2/2d8rqB61arCBLoMVA2Y6NDJYhJMcOy2JNW1QRe9P6la
EPohhZYPijNT6wDfqKtKpBfFA0oPtOZKqtr/aua/Cisfriy2YBziN8ahVB8jLRnemiom+i+m2cLF
3eifk6LJ8cyR2O2RqP8qLCG5YGe+CVHdOdhUI6/0r4XHTFzbi65e8qaYVCMdNtJKcOLVKD42qTt8
paxKF+NoC1tMadmC5GACF30AHZbo9ie26ty57+GVAlDp4HonFFXXlc9u1Q9o89J7/LVqvMLC/L64
Uv4s7+A4yLP3nOdLkfJxKBw9ONZgLwVWa+sHUaLGM0NxTa8T9n0CsHFnN1MC0O2VSIHgyjfmpAq/
tGDRBrAmXEv75zgEMjI5RoTW7Uhh4zm5FAOLkwYm1VsSKcY5o5zbr497sP1HbqxyEKJX84FlYMCf
ZJ7RBodRnfa0MRffbcQWz+1DmcaZHkXCNMT+UA3oWTNiXXOW7t6l5fffB513qbXZv429OhVAm+me
Zxit95OE/JG/Srlw88cmgLfqMg0YAwLbk/MlabvilvMxZVtM73hw8l9uq+AIaXwGUIO2pHZALhFO
LQJqJyOzoxMXzB0ISkhnPyW8wTqA6Ecxrh5DFz0X/qyXs6W1cDTRgv/BWylCean0GHSLOTpxeXfb
a4Ts6pWanlYogYJcQ0YxcF5bY0rqzrT9E3gTAZ6PeFHQs9+eNh60rmR9N/Vy7ZbH5Rtp2LoC8jEF
ELVCxWzgyfgHplN+jasKo+fHQYf8Fylv3N0epZA4ktgOivaft8W/YrnDFd0YJs1Ha5gI+729KzSI
e/f/TN0SADzgRRZiA+NtY/oN+Xe1BVsXsK+e+P+UwVMXaUc7bM6ZKb9jVe1Am7laqF2ARKMGUFW6
oF3hQBwlPurjIUA8QA69jGJvRTGz2KUa6d9ghnKuZVAxEGhepsXpx9eFH3TN92G+xY3r/B7R2nOu
wnA6Lg71OgaA7wkqdFwxXFMaZgx6uoaBAD1XulCIvhJQtJOhBOwpZhLcGNVnPKS+TrgeohW4xYyu
C4ai020eAIinc8OPineNmbHA07T2uOBpxQY65g/za18kf3uiygcSYWij6azrtgM1LTVZoc46bEi8
5dNPYIYc51t+6YoftY+vQ30863Do7WUsu1s4WYzn0VZkM7bnrAvL1LakhKiDUtu9AOszHySyFv7G
0SohAl+H+VcNTxTCucB/DfTXvBnDkRsOMpWo/EbOCbkGnmOwn+oDiFRVi3hw+utpZOdE9VoFuPbF
SCppuAw1wMXl1x3DSFxK1KLIsWFy+Odcf58ROq00WsbtKas2phhDZ2tPjMJCnfLmxH4aYSfjniZ+
EVKtvs0bPFGBniVhrF02Lis7r2bcA3sA4OeHqNk15a92J1MvP4o3XxkYwxNpMbhvDfHFh3MENE9Y
SVPL4pZWZ0UElGJq1AqQcyO+xewgOdgmKfPjaCxRjv61siI4xP75A0/5Q+X/iWGulJJ0j12vWZ9q
v8BvkukmLFBb4BTEmd9/v7N3SaIYeb/1aT8BtobBA6jhPHvPv6ljZY/BS/WcGr0lCYX/XVceamTF
ISmKwv+b6SmLOBgPxvZi6O7qhAyCab6sZZscpRaJ4MWg35ooTliAxtZJm7DogNczoHqzw//6NbFH
wQMN8TyFbfkOTU9qr6pBOKNXoFXJT24zNkq5azn6ANKP/QUBXBEpG1anifMUz1DuEXnZh8xLbS52
TgOZL1VV1bANgPTSxZSZGP24Ags4shY5koaJWEZtrXi7YrmvWlSrR/82duEffOrvyB/rI1wG1W5e
v9tdWCsKHILOw4fgki/++CHA4PdaL8UuTVMzw/nQHiISNcNBJGdX0s8tb1WYZsLHkExsPK93HjWk
olLwqRg68JfO7UeAhqxmH9ITnOXyeYidOUTx9u+ayQ627tmPY3Wk4kP5wTIKCqR9ZWBitx0vjXgP
5hjGbZbvwM9Akh7gNk2XUE7WKfvKYD4eQdDt1Xd0z5VF5kl2zXHfY9p/s3asLhaB3jbTY1+sCFMM
nCx2kQUDS0jYd1cMu2KSNdyws81Bk3uv3GuFwgE+QB5D19EZtkwlcK/JSTeF1k1CP7dGarvIqMbo
y9hOwlgM2C/Sqwc9b+CaNYXSJUciLq82Fhy3c1/JfgsC/LuU6YV78EIkMM0i7L41osR1o4ABzXKr
zDVHUfUPGZe2q6TuuKBhzUymgTN5OskPs5SWUsFTyojo5u6/D6ddnDLa2S1/ORvNjqnwgxMbb5iE
AxVbrnWnNVSAMFb2xfafxGUQku56W3hC48vdB/NBx00HbiT87MxZQFbfT1jnHhrJY16lBj45bAkh
/dXDdYG0eRkblkTEy95Pk2ell/419UBWxKpABQHvMua24J74vMNv+o7tILFsj5EsLNv+qA2hyWtS
i4hFCE9+s1Dus3yvPu9YvRTtRXqZG1NTBNDx+Q2+pSJ+vU9q+/4eXP6SgcBBnVRkMYIqrgglIn4L
WwYN/0Y18fXBbNFmb8z6bkBcbCKI2WdcXjAmlD9BjaeH8f2yfALZICYonqotRMDdlh80HM05O5Fa
SEeCUYcT/zrK6vQAJTqZALMcCD79LdAjvjpjMhvTQwXWX+ynd/T3Gy9e15XtqVTdVFpGf+BnrCEN
Uyo3ylV7e8Fz3ASZn77x8kXv9bd5DWFRuCTHCnqYHapcBzbgjPeuTd0lmwOGhDiBIvjY3rzMofyM
Trs0tO9Z9YpXX+K3V00mU60W6KeTvmpUnmYGswMuLbnKLEIPT9wdzQWqandIJ817p1lLi1KqKR/7
fkE39SUkEjuZlCeoTpK7vbmqF7jAogGR81u9M4+xCmREl5FrV7etVZZfssaiaS0r0qd4sxrGCvu2
JEazfHheZnjTe2i3mDPytmeqO57YLWS2KYkegDIiXUBgYsXxsARcdchovY64p0SmQtV92rBmmmP5
beXs4cbaNa5hjo85yXfmvFXsBAZyGKv1XE6OP79MbqnscCanpK/yk25oNggvP7tKAo02CVL5ZKFY
su+g1pYHVYq50Ab5t3p6U89DKoy3/6I6dgEp01F0Uqd5jgoOT6dtAaVFLGdKs5mHF3pvUojPSaEH
2Wl3C8R5To33MKH+c8q0E7oYrDFcEYc3NVXpUaO1hIOiHlIW2IqYbcRCmHnD2ooXhJKKXaI6DRo0
UYK8akrPJXPbB75Xk0T4X09k5DWE2JfRzNWXhX+jL7I3kbdY9PiUmjOCk/ZZcwE4+NrMdpBOnMhw
aKCZi8VxwGPieK6Y9O6tHtWAeiWDs376MXITLMl85z7IMpmrwSEoIvs1v4ic/mDyeZ/I6q0o1xDh
SYT3LxapZ5Ps7MHHFTq1jMheGzGzZK+MEcjGMawouV0Y9s27ZUtD4uS4VWpT2Ed4Q+2lClxFyloi
r7AnPhHQOxO8y32q9Sz0gDG042CqDQGWmA5oACyJJPP3E9JLlg/V//f+X7lr2aRTRroCY9SrumH4
SX+2cIivG2XJvYoptCwp71EZMOCpn3ojx60KMrDXsWFbsIEHwvBo15W+h4OkLP9lQ2/IkwXpphmA
ou5i26KdysVWHH50HdujLOqoycbMH4DddQXiMVXvvbI1NVBvV2wsBqaqi6qJI5GZJuMTLHJBHloA
lbVaCqVA/o0MAzsO7Dsjoslu0gnWpB/P55kKd1zj2wKFMEWenOm7IREGJ2/3vE/ZVqE2LbL+UUIA
r1FVKNfUbxJfSoJFKA8dlorDB0vb9I337oPMtPR1z79+3qsZHsJAyhT3s1+HRqot7Z4AEAC8aJ86
SfYITbPstpz/Pmc1AntUgUzAVRIWkXqkrx2vc80QSfkVdTpvepJAz24c4TdUKfPNF0n/o64li/Nf
OZlPXrBJelendX8yoSs9SgWMlkRIgfUzTDQvBLrH6wLyxtmA1e2GCmvH8s1cDqJj0Af/HBhB7OEc
IlKiJz19zNqGtp9uz22cUVoyFLC61MppFuBu38Sjs03ho3A858QoO8wKPqMmn1xrH/UA9+AqCceD
pVWgbLYA3+o2JcHZ3sTtSzxuAccmcH5+hdIcx8u/DwIJ1/k0DXaZxapfxQyc+pQ5rKdXjsjC1aAY
OketRhHABF3RXQEtp89EZ5Pygb0uQP8ELvQfk2oUqP2p7b+/A0e3eLGwaWV0YdVvTVb6+pvzagZ/
itHegA8xAwfq+nhN2OX8gC0LT1oKkI1xoyIjRfv2Hfm2WbuWs+p2wC0dEKuhw6w098Z2Kdje96K+
GTSCEtLA7FCM8chaVwqSaOQVUJJOSb3T982NLO8L3dh++goIWaLOY670GJT6F2j4iTXLZ0BnO4XG
rnMifKEW4tBuD0+4fwOWSKbXEWsdeQW31c5NmEv/1lO6W62ECdqrn/OjKHiDDNs6YVxPp7e4cVWA
XcLUM9cA5IAA/R5IoiKNf042mpFnmhA6mSk12g1OR2EDivK1bd9YZYALshE1+TB9qCUnp3tzMeZX
inUEwrxxesfdgnGD/tSgsvBmyB4Hlc9zFjWEqlcmzVsSYhOPPbj8VLf6nQUE64kxHYcCoZ/frKz4
xI2FhbJ/jhj/pfpI763EkMYV/NlLld7um2XMpZ5bAentKtr5clYhKUyf87lH7xW3Sfc2m+vJKQmN
NGlgMol+VmRg+nUEK5NnpAd5WBouUxz1b5nvlHIN0IJr7S3i0XE60OrD9ksoI6WFbZlgySDrmyMm
SFpnx6SYYIg8w6zsY/MlCntWrRglUNkAciC8lH8Ib6vTq9tfuN3MEHpPetlE2NblYULFvi4j/Wrg
E298gmUXCIigpVMOrUXRcvTbRLbKJDYoNKqwxw5X9slnWIz05uAOwAhwCe3f4PEpBu7tGttW+izL
4jVBeSESssh6lYTxK4/XmvamnDT/ULKMPe4SghsUftjbTJru3ao0k3avhBNKVtC30XulRZ7opvco
sW26Fx+hcFuKSX1Zf43VMj+/jNjoiqQuX864SgZSEcWNDDBKvpcH3D3naQgcaKEJ8F4qK0xZjjNL
mEfZgo3ZWOe/gVotQ+6MqCSsrOEKfkbrGkhj1/E/oD0N3HsXVJSJf0JY8MHAQshDX+v3jBlgjk7l
kKOIo/csOzitOBEwiVFxe3933Az3zLrWFFLbrooleXPxPBaVVep7M1B+qbDLrP9qv8hwa3zt6c9a
eXkbZ4Cl51yS+02o2neF5XcoKIOHCFnsV48tFEZ/XXHO+gfKHHnLfSX6U4nfB6eYdrALRPEtSsJK
G4gE0Fad1MLB24Dw9kFkT5oPZgUEl4CcOyCU9NOICsz1VVdwwdngBa9bYYoMKiSzKlXXtD+Mc1Do
QtzNBzF4KT0Yo7w0PdXwHFr218JGPKxtcWkqZu/Z0tJ01KswHHcIOZu4/ZexADJPQVrg9FyMwWuQ
qjclgwSkcCe8GZYg/lKYuHYJ0zJEMSNwHQHRMANmRMuDt+rynhcSqdZrpdTbfUEoB5phZ3psDUWj
VQ1/iPMnH9aZNAHs6pepDmnQCx+TLoXVjvTiAwcxulKfBAkdMQmeJqJgV4KfyV5hWUWSerQmPZHq
FdwS7iZK5LA8gvQAWAhSOobdvr/bS0cldyysh5v4b9A4e/vZ9BqcdF04aA9pVTxGwbT1Ibft5Lmv
JHwesPq0aTmHqpaAzHwl4DxFFL0RsqnxjvVk2oBQ+++wcRfEwsJHtOxucmHpVJPQ8GmHFvQsLswK
ckzicKjnYFmEi7vCW5miC818BKwBmrqnC7nQxOpa5gvZNnINK8euJy/6O12NNGOQNms6JFHfOvqD
V3dI/2v4jWGq94RMY1VgoS+3B3oNlDtGeabZkpDqmXM4kpGcgGUBB+lzYnu/2bKswWcvCi6XdT43
TcgQZWh4D4D003db/ImKTZiWxBsg+GV1ajn3OSh07t6FvFUfja3da4oB70xhhT/9b6rvIdmOyvFD
bvg+CCWkG2doyg1RkubPlK3SvVpDzMO/Nib8qySgzwhu61cdzgiHEGyXXF6KwvyPXao75VrSe1f1
bZSFlgCL+2a+5pG8/9xBBQx34Num2Z91Pee0KLSvM91r8kaU2Z0XJYox0E9TETBDCoAQKwyN/OIv
L2JPY87boyEfB2zvNqL8sBroNSQozgn1jGI/CNZpJFCM4O6aCwFsKDRXjvr9KwtiTYksu22nFnY3
Jqez5hnOb0lu92b/xJzkMHZNd2HfqwtRWdZnjkYMqL+gavmGf0SQbhrvqBbD91ghQraXIRrR2e8N
1FhCGKI/+jEwdx1A5k4/QkH3fwVUWzE9uEkHcsMrfkWANBUmrfWEo55Pe5gSJNBKdmjd0kyN4KSy
019gSaxTJ6HGev/ljka387c/++fHxqA25LVGlHswuI8YSIJfRw2iZi92Ftb6MC6CvdtSGcBlFfs/
5YR8mAJNJeY3cIewlFrnYRec8/57j4JLtF/JHzKWySQP7FNIqp4jZczzHeZOGNszsdXLmJ2xvT3h
dczjlRxRnj3g58mnUuBchDzks12Hoi7VuqrtmTLvTInz5ZWIF+4HOA74nwwRhCHty+SgS+PMyAqI
wbcdnDMXjX8arKQzgUe1qczZDY6edf+KFUquBnwOGrcYtTVy2Wq2/DM08zgUwbAllJhmzv20euy1
EOW1abUnsB/FiZCVZ0sqrHLGK2ehDxM72VeIh/elpgCWRzO+2GZfJZA64OkYpXUevhq1boHFvdvF
1cT03UJiMd9ttlMFbXJGDQq6Ld2UMpaEnzhjzCzbo0zkASqbz0ZhFG0xS/78fugn8X7+VpTmqdcN
bygJIIdgUp1i2/qW/D0jEvs9zh91qPGjyejSu+1Aumfk3U5waqCCML69DOgfcF44wATFP6X6VLAy
EAuEqVAvY9IVi4ffHbUmo5K2eiqePBR/cO5U+AJC2acvO/tN3pt/BMJ0avaDVwdhRDygTKNYkQUG
roH/8/JA6tt5UtRVanzsHhhEGxkhbXdXquYCkpundbtik3jmrWaBmezAyahPTGAAbaXdr8kMemsk
YFEna1NvcaObSA1kX1mIEdeogXM4+9EZbAfDg4O/eGjm80FvTwmw+rBk4AlZWFHnY7Ilb174QmR4
KYZnBzZfByGSonmOUc/UCgL/bJxyonA9LUuyJNggxLvAjKl9oCK6XcklPMalU3zDsb7ev6kQjzUO
hfMboXnrXBn7dmkc9fIYIHLFP0CO+gqv36ZLePGO87nTLchhr37vfZtD47SDimm0flWiibPoiUHn
iXtaq+ELL7uUyyKa8S9j5mwRNLHAyI1iL7gHAOIdQ8qAqqOixpXeyg79CEPRxifyzYZve6aojewy
CnuEqG3BpzTbUw4Ou/TmM5JwjqC8GfwTW1Kf62CwwXkelSJq+8wm/haQstMdUCSg8jbz8OgMqsQO
G9ZZ5Vtvoo3dVhICBwGj5USNI6q+5OWtdz/azbc1Ccb/fL2hWeoHKc3fS3YPKl/ZzDYDSOUlh7Ll
8z3L7mmBPHWnK+kNqFDOYL83q1OffrBrUbF+NuE/FCnuIgPuC/TRdwscx5S/WK8DVf/o4ZI7Hn/i
4TDc6xt5pbfZgAhgrDRSFiTsn8VY9sd/hlFc1sEfbTEISMtphgFW6a4GkOAneVE5Bb9BA7L2lFG0
xrSYSMT689FGucNhBxP1xfdwsyhgqNCSB6E5b9sIcLhnzJ16Sh59H23q0PuIYzW1M2F/5k+FvVir
fRkEBkexT2jl3c/peJzjxaF7bEArEoH68GCOZAzBSH9FdOHyunRo04oNcUwe6VJwy3r68fsvRnYC
wWSGQZcbTKhFgVL6XWXDWdvCOE1hWQHH4RQM0RbZfzyIJXyt3Cjf5AyisjtyrPmvwaXEr7xyZfJm
dBMW1f73DsIazFfccrOp8jQmh6zgX+QrnQ1R/B0mUeNJ0S0T5rZBzcXWU5HiRUjmVK+DUX2oyUa7
KbbSY13nbBPZA/l2dtVZYNx7RlLLAXJ5vm1c5z2tonI8mKkswMD6p15RX1NoSH6y1gJzJZew6+we
GbwIOIJOToRCGutzJiQ/D/m5EjTnmlAgGEOrCGF+dHvI446sAPi3lwdkdoEzeSAefEM4URHnFWfj
PsZYq4PSfsSnBpFYNYYZD+Dnqiwe2FNQ85jNL5X63mo6PkYGQx7ULLtxM6ROU1eWkIdU0EypM2+Y
+DOFa6KsyjHpWbgalE0erCEifKHLhStbjUFNSoCrpKT8vgS5RCTCXGxCWpgPOTYiQwejBFSe6bEG
9wWoBxF4jecCagKZS3qwLwpOAgUynBs9crEmSbOZjsvXTu//Cfq/eXWQcY6slpStM2+4niOmeSI5
MgV/A08JW6mDDGWyQAQYHYtjfTDmWIIUKXzcoUoSwbWfXETI48oVzdQMYtw3YlQCu5mv0Cdl7wui
bSWWLFYM0RjVZ9Dx8TK2M4CpOdo8ouPaB+05aUCpk4FucQtZo5bdYMn/YiPFHtwE3YKlYqp0psxV
/TGHFi//Mp3P6D71eVCm9cjjvomsRqBdj80RfL0XLjmMix/gip7AcKl8/eU87ojzsWOv8Epb62wt
b6X7FniGMWuMMxS6mdyIq1Qv2zRasyXb+QOi0kjrviB0VsL+fwS6/gFm9vxUXaQvvlL0cuBD4sj5
uOmYKWNXTjKXTt685qXt4camm/P+z5HhuSLKhlKVDomRwnt8sCJVj4XNRhAr8akorUCPcDnVVAZF
2+yAn0NOFPVMdUf2tKUTCXTMNPdL2ywj4Qsr6x8SgmBmNHSnvlHCtokxCmoHqo1LBkjZQ3arGFTO
VErn+EYMi3xM8TXP//T2IY3MyRZTqNVrCy42gmsxNY0nsoItuOtEytvQ1RYKfMmWedUo6qBLvWGl
vOSl2MYeQs2EdI/QKFN1Y3NmvsY2XfZHCAFansWDxHfrmg/El3Tm/zh98DVyOPa6MYnrc0avivOI
uJBtpvxkC8PiNafo4Ys35fNjWvWV0+lZ4gIp8FfSJY6Zq6sUBN/JUrxVsy8AzPqPkVl0HL/xyMcW
VMMRZEx/sBfsuuajP9hUWMwj7IFUGhH14QioE9VvKwoKR5bsIKcjnm7jP9PQ/WftSqQ+luPGMNIa
edVcaZZ8H1gK6FyqqXd7+64MJpjAmoVpWmSsKXrI6QPw/dZvAYLMvxvH2/qO1x2xW6mIcHkrCrQ/
Le0KxY31iOQQvM7A7a8KhMHUp/mAJATsb+XL/cYiKoQNGONOvJB5NYYoWoSrk8aqevw3QIvsj9li
GFf6ASQgyu0VpLKWmctxdoYM1GMBZziW2Fhe5QdVMYMCVflBP33YTkw/KkX51btfStq0r3SDoM0f
mGQdcC4Ye2z9qvTp2IA4rUBnAqHhOzglCfOAjZ+4bqbADQm2HhxmT0FOncwrZQ34YKWNsloVyVFI
uUegGDFTSPbMCpd97OTeWU2FZ8AXeGFX5Ko2udf2wIZl8BS9k58PSfONO3WeZ1YwUQZqSGAlCk4v
7/yoNksNlFG6u2sFk5CcsfZvL7ekWN450FmwtzEAygD03dBeaQk4QAYfmAkZSiiE03VZgvl620w9
XJ4D6YGvlmxJ5/O3RU1Jux9DTYik6QOhx5sz4DOO0b5ZVxRQeIj0hZVb5yvA7Z/3dtCB7ZmjDB+5
f+1AA4BN0HXHStFT3lgx6s4qkXeM6Hrk7fJKaT/EnY24h/dB/z/D/hxyLA9MbLDX++wLVwnbTTn2
7i9g1lHLoKeoOvvN/BQe6XIKrx8myjt6wRbN/hdnGaW622AkWmy6YL087zyogAklNF2A+dxAg93N
YFiQvNAG/ukD0LXKvY1aKnKfTI5HlyuNQ16W5S7Azby3szma+RddedxgER0WGEjmgJYgs5x59k2r
irytYkUU5m1pc04FxBn6xnzhppnELhVStIjuj+XT00326ToYWe+uSSx6TmbBmEf5hnxtTDBrU3sd
Aohv/K1miY9FQAiaa9LoTpBvMhKUDlbVVqkL3H737joDVYBPJtXNVbvgYFkppSlw/CzPyMYXx9bb
gdksAM1TgU/FKo6mWYOCGEICqC+B8Acwk6LynX/Tpz7QTnKTYYkP0XQC7vz1+9+xe2nLjmLMlnp9
P8GnP+/ojJwGuHqr4TxJMpdMr2L3mtouqU/Gcc3NUQa1o/0S7q/EfSvQtduZzw+/lbf/JzUaPMvG
MZeD/phLpRe8hOLwW0MZ7X4OdqYYA9m6vqZjcAK/MJgIoRbgZcZOsuM7YK0n0Tf8qEtX9JObPY2J
z70fp0qg3fRLZayUomUcD6NrjlezDVCfV3AOqs3AtubGY64EGYjknAjK2/TT8dKNS9Yp1QQ4xa8T
D9ub/9MtETMZpbFI/Rm4x2Lfqyi1T+Lkj7858HR9xLzmcm3jIZtTyHRIe/Hfu0d88ouMNT/6Q1yV
BBSPQfJv5GcIf0hG2PlSES9lFZVDNJSJNIYoruOKN+8Dc+TcrmbvjkXRVZnRohJKY87gpMQWFgcC
1GbT3D9xfxwucYmbVWAU/BwwP9imunoMI7V3IHfzDBmw+wktXnVif7kr6rI5XWkAw1yM+Qyv3jx2
I91dQNTKyDvnRWEiLWnyqLnpmsk16vppqPbPNuMFi5EMjb2FJQawt7ujbYveSmGJsOFti2R/mf+S
Nksy13RXxMK3yIAudiXJIEw5xGJv7VKZ6HpqTkQaioAkXyEizbqTpXkw+XUcXrXshRtTXuMdNcvA
hixLVzdJzjgOdgouePAou7/MUkqPyDah35HxYHYnKgtUW1TOsgWAQZ25oW/Scidupm8qIqUU+fWb
4j4WRew86XDHnfBto7f0gYu2yjYSrTGWBFwnHnuDsuPrgPb51EjYVLYSA7/OgU7YFWVAsyyTFdAc
8s3vdNTsIpSVFpHFHMtX4nV8Ga9yavFd+7YPx11RrjTleVJEN0XxnkAA0C9na2jg3ah4Nx2YMiTx
6wq14kNpBQ3/645I/Iyel+1mA5sin8UDiY3GRs4sxcfR9nHuFV3Gzp5to76fWbyGzU3jcB6mFi5F
6FvTXdFDvaBHvmDc7fGneIj2Knmd/2g8pM7HKmub8Y6snsJoCUAFBDd1EdGCmNjaoIJuwRfvXyXJ
+zGsm4ryP9LNsqFMWbLIlB68SsTfr2JaNJvXEKeJut/aAkdyAYPg/uPpedl7NLfzzbH5ri+OdWm/
8HfO9q+14KQgkWOiCxoqXrZvXgbfOFCBRq2M3tDhB2DRe3O72RQeYQMhzghW5ocrtsM0MexvSF52
m+27o4SSF7s/h4QYQsslY0pGsBQatMa++5QsygZzwdXxfshe0Te0i0FbFjdxv/jdQGkxYyVsQp7+
+zE7Nb5n+RymWwczMzk9ji7ZzDaFs/2BCfLNGu394krSkvEgs1lcuzjiV43hGZqOUB/2RME6i42H
i9UNFmI6XMAmOb79rparUkb8LA3bCNj/GXJTqC/fcsJD6OBJTgjTMliJvS8WBOoVw+w1dMUi33wa
QG+RfBSDchbSLQuljH+tUrW9+EyWTVmI4bffBohkOlB2t74eBM941KjHivbhkj+iuEGRU3K+MsiF
pOZGsxA9MYpPvPajZ0u13yFUljuJjyFUbQKCorn93ZYvfpD7G0BRafGwJ1jHXAPxng1TjyzLjiOt
lsE1lGzq8srvRRKPXgg7Q/XeO7vo9KSEH/kvYB30m4ggqOzI5DVSpqFfEXLF2TFiVxaM26CwsoUc
hfB2cRbgGQrxCPDe7Pu5X7w+gC0pBikHdG/53wGvODvpCgSknDOzk7Fr+AUwIj1vnXiFh4S2bkq+
DVI2AYBjq9HkppswSi4+XsvxF7w+oni3LX/xBWXM1RGFzRniCp3/HpC+YHXiKtdW1E4t4mvrmzYO
+TElxKfJr7v1syh66dMQyZdxDrepq5qvVGyj6nWJOASMnAMdn0qCrrgzGgBj1vSEmv7Z3rjZmARh
PoJgN+BGmtmL6ra9bziAflo+mc1hAaRLRS4A2b3jrVKhgP3qpYS3NzfdQjMwmxF1sUepzoZDixjH
eBnMDZtKyECWpuu6POerRg0057lb8qnLnxMEc6jCV1anoeNtlMSokRNec4f60yqUKtYhbKhBHqyr
o3mQb0BRZ6rdXzRIc1AurchduQzoMvVgfgG8I/HyoaXScM8rQo44FgffSNHJhngdeWyasGkm8/5e
XED4nGO71RN04WfCTDBJwLn5q2kSunf5XnhwSJpk/waaPBpX2jlCguiIUncFAn23CbYX28TT7wvW
Z6m5pAXrGpXT+bfFwJGn9lPOSoUssOxI1WlKRz8ZbY0S/47pAGvBxkv24lVyqSAFR/yNDHE4uE81
LpxC3fbB515I3YilaVY9CPG+e7A3dWvOnaCzU8sZO1WrsgkaOYi3x9JYTgby39HXsZT/s0tGYWc+
qeqY4gc7Zt41OYB8OzA7y5ryPwdG1CTneJHxsHB7n4aNj/Lk+maTCvYpbYq6j3W+HMyDpMx5zWK/
LrfcYu5rVasPyxmq7Y33RXtp9moHwMXmwdJ5n5wTx99FIBlaBxq+5pO6wqBgHz9qh3YWKiVRirxM
IRMCKnUsEbwa9nV8IUhYeuh5yTdHEfz2iUXoB8dHvfEVvTqM1FnDj9HhveQdAgOjbfoI3sLg2NvV
meNLZM80dfXcfCpR/dmKJrFPHVy4OaQTbBPupWIchJw5D/nUU1vpyix64dDaNB4HHkfdJgSTM7yf
RP0PfMHOiv0A48Fda2TzwCQ4JEsQ0qW+ylVL7T2u06/rguwikVgAuHQv8T5VWtoe03gKCTb1V0Hb
USd11H6bB3en+qtiZMN/9SDU95ogceOxNb3Eor56n4o+OBliR2p+qkQO9AkOqhXIdgjFx7XNXESA
9gGMdfMioyesK4IjU2S4SAxVsx178O+zEpC7tcYmfGOh2Ycz/BhGcrxOJtFQTssAZWyjRAA1Hzb+
mKQJDvbbxcoj4+sxl0Zbf5kYfFGoT7M/BAs1wlVJtEm6Ra+/DjQyCiu4LP4/ys6RUwsvdBdv3FZ1
ZibYWfG56WgUidf7cnsJo3M9zK7mXYDzx3g3lS+Zqi3RgwuRmpPPryUtjAcG+FdWLIgLxfzFy4Vf
X7ZUtF6iXBQTDGnlr9y4/vthDB9b96wlqDDZJX4s7/l3VbD2AgT139AKnvXEZMrxiqMi6n7CZAyZ
e2N8U9vC6MFRFKnS7U8XCEHS2i6l2mVhUp1WNC18Kz9gND9A5unUTlghyPRZ+KJtTuhcYbSnGag3
HJdOVgNlXb/fQV+8KVQ1yn7r4T+LI7kwQwWKUcFAjsY7iUzW5sk3v5Gg5/pBI3Kf8WHqzlZjQ+aQ
TyOWqB5JZAlpJtJPdIgWo0RAayHFbiN4kCBf7I6H/F7+0IojuJbMPUSfyPCe39W3huBgCQFu6Gl7
3rv4eteBsqFIzaF4XfzETRTR80+bu7DoGnUPF+5HNVeh5IX7Jw57jedGhMkXBOJxyMwb+DPu4ea5
RrxUX4KcUi0fcIgPX+BNz8IXMd1LG4tdV1D6Yja/7iCuYLbbO3UYML5l4OyfKqOc7Qm+7yo1udkK
mIEqGdDbL3F/w2GDy1+3DaUOMSaHYhv1VLmUuWrYFnznbe7ea2y8Lo53XGyXCtPBX/tLpfR+upLg
c48DvTrgoXEjoaquMalBxHTPfELR7hSM2Hp3n2XmcImRpoZls09UhVgnc1pNxBJpYtyuF4c5U8+0
rAGTMGAoQxUYJmiTojR/JhVX8P9YRKR6CW6lkCSt5EsKfzjtHV+3Cp5L86nB6yfp2LNJidBlawct
5BJoN9ZHAE6dNvCDmVzBn7Prt5u3/Ftkh1dgIkLqqnDIrLh/dNpthV7xa+yvEKucFZX4xk67tck8
va6jbFVlMBBIqwyqk09+NlmhGKNoowLxQASX+TifrG7/72gezEw+DHWRSCq6ewfxipyflQd0D14r
KfjwoEx5N7D2h7FjHYkE8a7wxxBkUri+ZOsZGLV68q+S06Ed8gHXAYPjW7RjYmLy27lENOFOZb4e
X/IGG8v9AZ8Ym0LKIBclaQR8NgplehvjW7J9jRp2pjqN7CNtUkmMqiecSzsSeVYG0qlQ9TUfolPh
5yUT9HlY2nQEDGWD7AAVl1JMm2VvGg9OEi5jo2UwVAEfIR2t6RGVRVyh6MffU/8/mOuAmQCHrgoX
3ox9L/ZDgNFVTzD3xtXPKhcFthO50LCMh1FBRANFuQ/d/GNY3cKs9CpSRUz2SnT2gaybKj3EbJEE
ITADcqRPfBOx8ZXvaN6frn+rzpIZQJqtDiu+8HY9l5X5AgxvqIKuCsp7ylsAMsGnNKZm/h5FN/Gp
68vNdp2gNfyDifbEb3tPhDW/H43O8QIazqJfuQyKUhZc8YBfem+pYMDvvmn/dkZeZjtN7wxeNddM
xUxEM7ropesS9KnfLuJdBiDTPDQjcmUpRCjL/nKEkXzeaQqaCLtLGfIPo1X+KbC9cvd2Npqddfxw
qk+IFU2+sfHFpuh5shWO9hX+WtiIBv2f3zoxwUXYjBID7uaQ0Yqf1S8HpNrMFHp6oAtw02n0RLvV
nsofpdaXVffH/b30xgd5tWTtsE7RknyaZXrdTNx8UV9xzJtIrn6qH1yu2WC1CIaS9ZO41VOwCH5h
6Uplby1kewmb7g4GjKLpJYf50k8Kn6DcVPrrU4o2DQtPVh9GBG+1+EwAlHn9Xn1wdKmbyV/ti2Gn
5vk+Lo+5/fvYCfi4d/wwP+SWWmbPO1rXYcGhPQ0vWO/CZYTL7ZskP7fY349t4yI/o/Pdcp1Z8sfK
3BrDGbQi4wL3jJWWzugvmb4uHVpVkKmY6srcVMA2DEwgzZfGzG3WHIjoutrbcjnaDDKRhg2uGz8Y
FU5WqE4pGqBeeDGEE7IXPF2BWlROQNzfzr9p7n4Mmm9ZiQI6KjGNPWVaI4maj2FK1+uGWIOjwtos
gyt0yb0mRcly0TyyMRZ8u+zaYKozkptxjdow5scrDFNFyLfp5V8MRpUQi3DrvYkoIb6FsPEKKUjd
az48a+DWWwpO3ytmoZihQLbFG/R9uvyU4oHznsSqr1QFXg2FFp8RLGnbk6NDZtBHncL/RWrbMSCI
vkv/KZOT/lFosgFadlqd1wRK+BYtKosaIwnMykcATpT6ZV6bcTzR7167nrSxNKeYS815VumcKj04
gdwo2Zbb1MtYc2+Q05dJqXRb1TFFmDuO5sX3uG296KNsskXxrO0V3NAwTAQ/7mzRf/1hC6+W7eOf
MlUtFn+MAeQxUO6/6c4Z6Hh4GYSZ/XkiVfo0bMrDTDmLb2hRXIkl4cEKa1Jmnx2ChMKYQ/ug9RVQ
EyN1OJNaI+W65Nao5b36e9W+suPwFnf2ToJ2iKAYcwt8zBNSEKRfQU2udk3pIoBOGFEj36fnBja4
4362F2z5SJz+wxWvuCiyPH9xdBLQpY7WACcBqncEtOmZIfS0P0baO379yyVABUZTzL4a5swZcO3M
pL0YDph5uaNyN6jhnaoJGX/ATZj6zp9J79o3qgrL8rz6f2qHZLWkvPRMXLLEXA1srEG0fTtQ9XD0
25SKElC/5hkr5zHSKDLt6vZrVzYRVYhtvu6TgOrzysnamjy9mqiJGy2GFPucgqv4lMOCBy2zCdOS
7pBsWCWTrGxQRopvwPGhUP59MCfcIEcS1M6crwLbn/GjjntYIDxJS47cx/hbLy4nH7lYYEtkQHZP
aRiN4XWYexWnHyFBZXU9e/L2ed35LcXKsrJFfAlqX0IJ0d0HJDmLSy+nWLaShNVBAblfdWbKcu5t
RV2gUgNc6dEeBDPNf+Jb2PF2HTPqlLbwBph1e97Pj0QjhKb5tOX9oRFi3Wjz8B3znpXxv14pdxtv
UR+akgKtcwamrfo558uIMro7mvi5PZZUdllbv0kooy8tB9Tm2BHWhNlzALxJN1JORyzYye/GzAmA
KjUQtGJe37b2ERPxyVeUhfkBrU8RS+NkBlRThB70V68oCRluU/Mkq2nurTOBO4cSW3oGG4EJuO+W
OuwiwFMI0dkM85CFDWvRfxSCLAb+L4CptJ7wstfwKUC6oeGLOvwZCTfnQcIexyzr2v8+mubNU8ZO
jLJjt5Ix2346Vz6D+oWrE4rA1HDTAPR/el+RR6o4NHcY2EstJ3zKCsnSz3LvEl30PIPfcnsRXkBK
TITn6NNc6drwnFCDnm1Hsp+zQWuFnQixgO7rhwtIlVOd8U3sJX77dh9e8wgoR8k8X+PnQRBjTUgW
xZ+R5bZ7IwKGXOtIIztIcxzQWPn161hBOst3fXy6y77Ubdrd8eQhLQOa9q78aRmF9gsdaOppTE0C
FzUv/x+7+ChhKTRXNgwaYs0lsJzzpfJyyytHvw+5UdDMMdnkp1s6Ps1gPdqqXcnAzMMJlVjztHU2
ILGFFN30CWrz6yqBcR4pGaClpVBX52XhdzcUzuaGBZQY5Xi1L5XzTU4FjqbIhS+vF1RPg0OTQbAE
UZNtsyfpQR6PEtP/UqN0b2+2oAGAH8rsfa0t3ynTRcN110Omyezfc0MG6sIH3BU7uN1XDGS1Ymqi
wKhylcX+PPrReCoJZHovNOaUfA+blw/X8SkVQJ0ws3usHVCcQ01sYwAWCOZ6gzoQc96mQe/kkGPj
yKSBfJ1PK+vY4uvcbGBhmtQ5NGjZ6z7eelfPTRHwqGUt/MXgxS3eN9sYi314Gi3u7pjXNo1VfsAW
k+CkWokjXPk+/YHUuttA3NMvQ7um0vHsPrnpcTI7bZ2s/6cmtiP5XnxZcAq99YdnZUnXordG+D/L
yMgp3iBfOQ+Kh3in3WCIrmaZYk6AI/trAAvJO5/HoQLgNC0gCd/Cu5HPnPW7fzpw7ai7QdWyo8hX
BG+q89U7hRo717dhr4YFLT8tJzEDtaluPjpF/FcZMxJyvrSscCIMp6Vwp2dJYA5L+mUNGQVdQj3u
XZiHObJ11j4vdkWhQ98Dtpf2kFPe7NdoQ231KDRncj5Vys4T5Thyyk2LzgozJrWbFj5ImyngQutX
uMVHdifE1PaKhlYWisps1+Tnwp+FSB49yLyZnJ13hHTlFZd7RO8Zdm8LdcIoavCl3YRniCbGW/Jl
l7hOSbjDVqneiYv2XXtaGrduOAHC7451k7UI5j6Kx1gEy4zl3e8KrlvbJR/O+0TEl8SVkYw+JK/b
/MbkJJGuTc9HkRbaCOvxsIAg7YLX1hkKO1kAL/YJMepW5u54noj/7GOFChXa4SG1nc8+sEB9LXzI
5mGE4fjjusBu7mkarTqXOehSFvxZWmUZ+4WYFTBGs7jOYeV0H9mAFRw/rmPw25p2IsnVZtTfvrHX
ggCmYLCD8SylXe3H2POqr5QkD/YMplbBVdWa6DxzR3D+0QZKQCKOWGsPdjA+t0tgwKxC9raTZLU3
ChmmhFxc1yIRcCNEP+kjUqPs/t2OReq4iMKEGOZq2ktzK8bEpmDM5Uso+p0ZqeHXERgmlF8DFJb6
WBjbNWs8FaAxoeG6DKhFocgwXoNhOU0hDOwDi/3C4fIDO8NBpITG1FEcpmgaoU0SMm8hMwT/8PqN
DMsxGwC3t7k0cSj1jwaZkeayXIk+4hmL7b1GUbV3GJoLrQDujlMOAmq3qbR/cktx5BcpjK6dbWB2
jiU6PgNrTfHJXytH27kvA0bEAcHjZkQSYk3G/cvEFyBp5XQfr0IwqjE3QzznA0+T7pugASo0lBkQ
CQLwmiVXVWtkMNRIsf6+jlAUdiDUTgj+7eRVGkBYv1XhdflmZdejOz7w0Xq5SQEgfeD7sXOFs+EE
nmVPX3gaZj445mRbPCnH26wuFM50eK/Rz+nSyDtD9NXlHA510EbE00PLNU4oo5+UsGZ9yY8/XbYm
8lzgN2YT92EwPUHagGJqBJbd0/pnr5SvKm/HXjgd1sKogm2qc++MeJgB/lV3OFOOvApXtU72qyyf
d+sbodtZt7cSE60217cGSXo5mcRxKzrLvWYlwsVnzcFT73XBRw3RGu6KcEI1YqGSbluWXeI9K6qo
QJ7MEqrfa1KpDtCRd4llPybKAFkksYu2SzcmR8IkI/o0CTbw6LsNauH+TdH026zES1Ck1V8mDclC
5sdyT1aOH5NxbTtk3B1xisRkni2skWnh8bRAD78IsMW3xIA0zyfw1MdZQbdux7nhLY8UasD3Rq6Z
myg2hSgljGxtmIFK5YK2t5it0/YRjGx5oTBoAmiAzhOpgR+uQc3C1ZWi4Qf1jD+9LD/KvlMTBoZJ
12r+6QGzojSdjVRpOvbnpBAG827EDcss2m9uAFZy1vLPwcbINaBZCxhsu+lO69Dz6r5g/WgYpxuW
5hQi7qtXZ9jSENpgK/HDIH+j3HALTIUlfvKTxWxSLgztlRP0v/hl1ndZrf/Iv0hdAHnB91BS1Pd2
ASSnjcqaMwGIhYIiNj/+lAZgWu9K7CGFmJniDKVrvB45VBZBENquvguU+hLEiVCfQBznTY+OSE7+
5CAyHEbTWXOQgKMr2TuLROiotQSvmfFCjo6Uiv4YpQ22zYh69Sp0wFXdiufmlRBQrMtQfsVFT9oS
RaNFGLoLOrOvyzUWuK8TNSHDo0i2adQK4nILBLlpM2Qd+YKtiVtwoWDNP5BefklQuJnnC+NPU+m7
1bdZlzN8fcRK4dwHC3i4Jl+P0sUkcgIfwQxyqbGl8Fj4pS3N1WAPgRH7ZHh1d4WYMbOUAsJH8fyn
MQ0nNqTjnR4x7rfR8POTvr2G8MN1JNlbe4edGkc9CYPiHxxD3CROFMoRBTbdVSzLGu8655bf8ZeU
LNj6Ht0X6S78VS0Do5lOHcMjabQqzHG1RvFUW3/i22pfjhnkc47Zg3NenR7WwpKVOl5DBvhgBBE0
xCPDgGMmc7qxCjbseriZluNyy5vqlbb6Mc8uOYXtyRd2BHMxg8JwU1WFZCplummi6OCuD58dpHNu
uJa/rGSVyiJp+PmxY4tYvpgturcwibu3nEoLHJmIe86Kwx8TjFm9Njtk1TuCyTsdRNJisVq8SBK2
ajgsyyoJ4DMLbxOhn7hP53dhI0y0lpSK76SWmBak13iDxOrqo1Cnz7jhd8U2Zm62mNNnq2pBwOpF
8YbGYV1RZ3BfHNX6SBI6GdSsdvMgPif7EKUABOPgnx06qmCFjpjt0y2AEKY/i85OfHg/mEDbE8+w
Cynv5VnSUaAFucgB2iwPbrTAc85O0Bdpq4w8vHBTtnWk0IW8TDQtvULnfdBKpuUFA6SAGoY684w3
sI3bNWLrQBsKME1Y9clv5CVx+6aMNWVl7REqOXWlsOSx7Ltx4LvB6QewyC4O9M+/HqhpQLI+h19n
a7D3f4X59VpVwa3aRQXfQxNv8BZQF2eDlvYllGtZFbX78kemXc8/XdguGLA3c9cAae4qF3u47gKU
taRgrdIb615LItzmPcuWwpl5zCzx/+2wuhABmmluyzwvwPrVLlxE6NeJNuMlvSozbQGZJEXbfjNb
PLL0IbQnp/BQExL4RVVglOhE+3XogX7TTIGlpwBbRPMjetApej/7SnGIyADaP+kAXKl8AKHuF22P
GFqVh/S44epJmQfLbRWPYiJlQxEzQbr1W93Ka+E/EV1mvsBhVGS0/hxBdJ1GSVLTOBmvwU1boH0a
GvnDpSE3wy1pJ0gIBmNhyGfoRHEUAl0AvYUcBiLx/Qw1Vd6Eu44qzJ5wMyliPhDuGD3ECH9f/Srr
nD5SkTWPqOA9E1vmxJLg2/GoK+vcg4wreW38jk8/l1jDZEodc7fn08gOWreMVjSBv4DNtOLvGHYw
qt3bTj2wSwJwaU/tqLMJfQQOWJEmRidUijQaKFP7zBzYf9PQgUan033vVnZPHaAqCeNngN85wY1H
HrRDKzoio/oMz0bcaIoGNe7f4PKiJFMRXn/I+OnA/mC8DCLYVep3zPWGvLznrdaf3tc3rrNRNSJ+
a70tZxStrob0P9E0Ld+ksiXpQiYRikNsXRZUwVe291sSgC93rrSYNYuHcYpxArKDxCgBxrnBvnUi
D1m78rj5AsPwSKYgWrD2FlNnVDkL7/gVayTJZXxM/bgRt7DVBlZ3/ymdxz5xhJT1DmqlWzbCpkDm
M7ODXT7NM+6cBehF0SmhJkwC2srIEQLic+BsEsWKWuBxlBCwOpSjphEvm/8iYwcODYbygGZ8ip37
4H/Grlk1jJZNSeeqRgX23M74LZ0+NIwaMOxjHWmfEEwJe1/AZc64zVbsoUSMblx/LCB7l5TehQQk
yfX0caazNks2TDA/amdRYdc994YNQSuE8dtm8A4PKRsKQ3I/9y+5i0NU16HDR/CxLbyA7OZesZFB
vyQsZxed+za74B/1SmMtC8l/YUR/UPBj/eHtSIwMoH/u19oJm0Uil+2ln/sTduD+Q2Ky5lBHVzj3
tfc2e9MGasm+4OKQF1c1+JPjKbK6xjzkUxTbQB1Q4sih9Wx442/AcN1qUVMDENzzhyeMoyIR2IqU
Q3NC/hWq587J7yKOcblWk3SOlHEODALnb8QcyvpZezYrSRVwCF1swL2IILoJYHYT3x/FZj0PS9w5
N0+sRBY0MRCrypHLwjdLs/iFHmSXRfk9hSroa20tIF/JaBrLrn+CZTH9SQWqkh7I2bjYdvohQDP1
fVV6i/7OqUXZqfmNTAUj2EgQJZQq8CQERBPBpCjC7xKQeGXNhbP8CsBbkOdVBRVJd1epT5l7heIo
IJD5Lnfird337xnVF6+kpXE2AmO5ciPIjVmQ5XmOq6HPUUaG9ReSw3XNLK0bOYHaDrE1R7JaUWtK
lPJilW0/h/1B4dIH9WgcaKKv8ft62w0ybpTl5qu4h08K8uG+kdVDWecRkNFFZ+9GtX/tfe0LWazA
5rJvg1TOpsABiwygYQDM022bxOROWTUfa8IxaNvbHoCR563JGv21o1hnuJjWE5iz+c6/Vw6foy0C
PxUhS4TJ0/pWsGSOLFokqPtblFBoOY90jbHbSFNLdvLUEs9z1KYIuJAX2uQJMGFxmyQGqVd1QlG/
5Sdntd7F/e9zqS0eAfIIMpuDBDuc9i5k/Aw09IUxSi6qUnJr/b30tDLRxyiQwePsLEx+xREd4nur
K+6IWx9KXXq4tKPX35QK/QdSsGrKj2T2W+xVTHeTTOjndjBDluir/tRkkwmGbl0ZmR4QZOPM5AhN
DiyYFBxmjwabBBCB8gcHY/1r/uMLAGe7V53KiP/Zd9gn+dEn0gZktcQnz8mu4EcPKXMy9wmjlGpE
MCLEAxhRbfZSa92A06x5oo2gGt8ggMlc52zN53ZQ0EYJsU7k2u48IogycEuE7VpAxnYgKABypb05
0b6J4uMNe6p6cqBs8IEaziKI1U05IDM2CP3MqUxMM5Fd7WIki96PaFp+4+tRwc0UJtqK1FDxdRDQ
x2bPR0ki/hbrnvx0F3tsUxOTYF3xzyoobl4rAbGoUvP8ZWUaP69q90+QE2F6q2K1qhUFEhcozf80
b883igI+Ll/y4ErtvOsS8W2EDTvuMEk0SDr0P8rW+62TSe6Tdd06s2xzZf8eC9f06IS9BQZyzTo1
7agvfhMimMTvCC0VanqQO/TLo4xOxrxLRj9I3LHOB6Lh1bHLuTvKBP/7IpJGVN2oHmKP79M6nCTP
8elUTRzCyKZYAMW790/R3urJShPwLwi0RB7FonD6bfPlQ6jFZTseUiOLFPS5sQ+xmdfCjJI49n67
bfHXuGOx+TUdW4VUhKvCeNf3C5FUkCySIVLjOh2EKgRl004toMJsrXwCSSwRar95NCMgL45S4/06
LNLHs5q4eAJ+q3xGPxDDLZ/fHwjkP6vChve5IWZX+UyMMEpznWkQghkIAXLgaZVULUwBnyfsUVw9
fwbUVJgxZNZwZFuMx2W9H0yO+PEIz4IexrvEmlgM5ISiUaKdNWxXmbr0P9NpAISFoEWhwKCGWgNr
ovTif5rpLYaItin2fliLMWrISBfboX8hYtvKbcHvIeuRx8PxXFMIyU5/wpvySBYiIstDP31dJBUB
kpeKtNwqsIiPewLoceLSpudwL8Bi686mKG3ET1C4clGIaQeelssGfv72eW3kK7Imdr2R/H9P+wED
NImrlV2dyJGNIv8h8fBxAKHkP6vjXB0QdL96sm9g/l9+m2jXB6l6z1aRuYJrGOaXRaz4xl+L45RX
P0PIsbNrX2j0Fsg7cOXO8nlK5+QX/K3MMmxBPea+RSohgx8lfcP6s1bbG69IKKGK2SDir/4N1JDJ
6AMB3HKKWfPkXbt/zdSe+WiuXjyV8zW8vxg3DvUT702hkBuLwvH9tXVzqaTgRTINBdNyirIXrAbM
vCCOBGm590paLpLGxPI5NzwuaK2o3lLWfFn1gbDVnRx6N5HZz0sU5kkzbrt3AgCyU7W6UZ1LcTcu
9y2Vr8iOvmaUvypYCVMjifz7E/Wn8gTHpnz92wfec6hBNx2/fGEo88cSE4C/7MNZWmFxgaGoo3nd
+vGp3VHNNvut2ZGtrzk61YmfFK7w04UeRvCeKyzaVceek3Mp/9DQ0X1/6SBSyPktSTwWrvtidZGd
03uBQ7phFpioKgfvzCnRRshKNeYur6zUn5vl0j+co9aTN5AoiRwqngA+SLxmU3TEll+uzBTFuZxR
j5li1ANo1bkUWOn3zgPKn4rkJJWTNPlAJC+s9QvHD0q2406eFCCIhnWgz2oig/UnwTy1AJlhSL/D
Q5pH4YCSBX6drbhCSVC2WT3MnXCpuRtPkHSgNx5ySZpNiq4OrdiWfpfJi+2u1LcrCkUpAhSRBaYW
YHFdqbVeIxE4y1u4Mc5Q6mHEOeAY89PJgxjKJ4fLHf9aN9HY/A1c3c/K+j5bOI3vaorRxc5u5OiM
nLUUD8GTLbSlROB7KtgqEL5QTaAm+4uIVDZ0U8XKvFtBCeMSHR3pf5Ijo+ntMGYjNj/KZH5dsy6U
Yo0ZSg2uNz1ymYQpspCHi3dUyyNmwygNQeI4h0P43MxY5pGA20TZtqCYzJj34HHVKU3rBYpO4TeZ
KGlNWUCp+JdKfU7d4Otc0GC1vl2qWwbWGHyVEpoH90nNbrBb/HKaaH5jJVh8H3VmxMmYuLqW/Yp/
YQy8C+DIIoNZHPVZYM/JGx40OFGR6VJFziSReTPfDpIUJmvv+H1pDs0GfwHTAADmDHD7EnCO3R+Y
XYBpvEwqzZ6WNGoDp3LgFIFCgxiYFXfuSt6mS5N7Qs4Zsigk81pAsnIa5RaRQ0oF15JSk5LJynev
l1GLbdW0KFuDoWmzTFYroAlbnqvcgbyLMuM+A1QcR1FxIPLSg78cPtbYYrA4AcpEjRXL5xspIjCG
0hEMjCH7GpHh7cDYVrcP6P7lwZN/5iInIfi3bvrquXNzyBM+3gOgn70xUTBC3lUkpgwOAGsyQFER
4piT7dxLIrHqB2T+AeesmWhsel115ae87cggm55TGtOgG/QdzrK0zkBifEdTByuzcgifP4vj7SNE
H1kJ37COT8YZEoB4UO8/mZUu3yfRt7YgRfPzWuKUlhYWht7xTamH/bNRO7LfxL4xsSGTgOH30TSV
v05JEw5whnsrqAyeZS0t5o7M0fTQhVVWCmI2hYwIbT3Itlo+NErJhIc51wKtPUea0Ig+qLhm9ljs
rFbJ3jEtxraw3XxLjeAo+K+2RQUl0V03ISc411ySEBK6WFGD3QZRjEC9wA9fs5SBdOqDNw8eBC4A
OzNL3DPug4WGLkk4VUrOloFWrfNIWTrh8TX6pX4STCKGp/lHnGg8orbzewuwn+Ix9DTE4MgE5HoX
LJ8xvkbBelL87Sjsg8VWUXQcR8pst5h6JrFzkZluqlOGYsLjPlaU7yIKUFi9VYupJgyOZXvHmU90
rVbbxfCMEcwFAGNKes1XKB3Bjy7pAPaZoVs8NlDmkzH8649cZEDcPVv3KlvlKCizFxg0cGqxA3e0
auSkRL8V9VsPBrBH/iTwMOGiT9PEcXkYGVxnd1xReR/Bfg4boduf14kkJf6GzRH1c7EpeKCw/NZC
HntTwO5BJ+IO/5q8flKCSkFA+rtZv0IburkZ6bW18c3q73563Y73lcUQ3KNxULxj1lx6ZN6eneRz
MGD6NUaJ7P1DkqOtwwhmnhTsU1eNcimUku5dKdV6v9JkaajUZg6D3DgiksGNOasVWG8w7XZXZMVT
G2L3aDB2s3nDnVEs4s23LGMMWaYsruWsQfkJVxMyZSGtdYmCbhBh3rqD1nRrzCKOnaryA3MuAKz7
qAe39vk0enpNb+p7s3NlsWmmAKZRGjWUNY4UoxSkDlAkaGsYVjzdOApiCul1j0UY1VrmZJGKgMrU
Jgnj+QpINvmaCsTnoDEmKAviRJj0sps10Lvg3hFpIcuEuPHS9F9ZapfwyyLaRtmLXsK9gjGsQMnQ
y3DXWhzcduNDc30ThOGw0cm2/O59IrL/6UVBF/KAxQC38kGnlNNRiwdIMLddHo/4XTUD4JO+s+Tc
IFpa9S9fYadUuvMjcw0ReU0VrWGgR2VPlVxAh7cnpKDKY/COwa/RVKRYUmWdAopV4mto824jHuEc
lmRg4RJ59JsilW9DYAXxGsT+6p3LuszWAVeX2gnnUXtkK9aco1Fy+0YFJZ6aE3/FGF0o9r2FAXlI
rQ6Eu68V8ws4dQbfmB7rHM6lG4VlzbA9thtnVH4TCyJV019YWuddZlPFQ6waJMWzQ3PzwuFNEBxp
ULZyof3QhTWoe3sHAq3KlbIA7TjOqcDzPnXHw2FWt4rA26LpNgHgPhOEu4S4NM+V42sG+k1092ai
6SI2Y2dPeGM37vXCkp5um/h0xbgUzmGu8ODNJVjFAeakmq8bO8nTs45nFH7JQkSL6z5y8A8M18U8
BJocTcVkBFZcLWyvmjRxs1flIJl7GyWS75V2on2TFY7ut0vljtEn0pM7herz8Pl0u84FbIms5g0x
jZscD5uEY7LO0vOiCdylFWd9mpySjWlu+lk/M7bWMI3DPUM55q0v0152oeSEOnBF4nlWNXjnoZmc
fVePbItetoK+Ie2BU+ZiNQIXiO1ahKmgpf7SB4Hs6mBa95sIn/IxSplMzQG9g6Y5Fg4lR+3CUdSy
A5Vo1HtsQtA7zqyM0a/YTVI4TbIO5yPKpabm6RoIcmOcvOIk95NJ4Gi6iYj+sjiLSnlFxWb+mvkc
vrqF2iUURG5jM8ZCgKUR7QY5XIN/Wm77RJKxb3HIl6cpN1KEX4Cd90ef8h1wSx969VV+6QmNw+Lz
ehLNwENG3aG8kg5GcQ9TxJt+Rb8GMmUqANnu0Zk6t23Ui0r2DjDVgYjiCFuTcq/Qwqr3SeG1LIUU
IC/LXtXmqLrP82yPrgUcfIqsx1l3oD4RBGGPo011PfnefvKeNGa3nrHovZdHkVUjA+cE1nE0Bjg1
8EVskj/NL8K/YLzDeg0ea0v2JHxcCU3+U9LWPtSbk2/glmb3I+rtHMPr0WZlmt8ENoiZ6w+HhaEF
PXxdC+9ske92dydsf/2v5v3D5pU5wsA1muEiRGKE0qUdADsmChgZerpkqb/qyaJXzYv91y1447hM
DTGdrOgsameIP3OG3y+JqnoBHbIwFDouo2KkWgAVL/LOFQTLqnHrAAQj/hDwzdNLJtqSf53LZSGt
4CwEPo3VgtIeagY3kpjUYLKailze5xHv7LAJrfK6CUJ/K9z7eXCfcdWugbEpInGa6culAzPf9HFz
MKIJIbingc6Y17xM/ldkFJwiAuhsouupENOJYTH7x79DD56Vo/B3WI8fsd2ZtukEBBJRCzn/ywkQ
rliJYSmmgniIHa8Go1es6OjvSnrOX9QKIS5Ii/BROqUTxbr6DtsJeDrsoNR35UX1PztOSh/2eMbB
hsxJjYfkuL/xrgTT8XjAlX5Wee3QPxRj4EMWSsCMtO4knYtd9kP+1xAk4RST0vjKzKV8yXUnDysR
R+YaoaQ2NMXftxgk4RM4StrOXJBlqnq+ndT+S5O1HIusqW9cXy+J7WuItPMi+Vc7mHMD9771cZLK
gIQNm8VuH8xc5EwMG+gXKs5nt9Co/6kjXpzpNTcUkf9gz9F9D2VBFAc8niBbVZFHV0to1Em06huO
IJ+lfFLLmaArAvVPweiUZqXiwSZG1bJ0mMl1p8VluTmS3PMLI3+SgkxqI+IpW1RRExPqQPoVgS7B
acf6Dz82x4+l4ncvh27JnqJ7QxErE9uRQKPpI+ufoYln3DMtM6ws9UNRUcG/pGbKOJc+FFeM54jw
Av2gQhtF7ktQjXylNmMXIj7P0VyVNe9d5QVLxOvhher3J7R+0bBHjAYRIluBJRSpBksUx6Bd1LVT
3sImKY2NDC60ibo4h/rBAfEvKuquDEVczK/4gCEouwuItp4lwqBTtraJXskjKj6B7+Q3J8j7NFnv
iOn6UimP2unKmvCOSQMlai9Ou7A3d4q14tdIM/dnuzyQONRx6fdCpAEA1/Bal7GhyvGXrgJcKrQR
FYO2YH13rgWkLOAeUtoNpGGZzvUMv/nIjLgvoZ7WRF54W5gQhzIysZ8qiVEntGbGMv183kgea1VA
Tfplif7+OMpPPFaB4HNBTsJu2FVhYf1E+Oz6it/zzeGLAX9LieNjRxhNw4LSjrK/QpjJSA7vrcbA
nsAX5opkq3QdxY0aa99Io/smllr8KaiT8ydj07og7gi2gCCRNiE52l/UG61pNz9LUOmiT9SYaEVF
Sy6w2NeFXIPhjE3g2xoA+bUEqtHwQnk/iH+Qx2I3s6qtNb7alvtY0Dq1smcK/sSJvpeU2oxpKboX
eByHl3s+pgGe9Nhi8G2T4ITjVoP1Ic37472fUHHykcF0vk+BB9eIakjqbQUr75kov5SEFH3eSRSj
iF0uk1JznC5JGNN3JYrUUa3PEFZqkxnLmWGlduRoLrBicekuht3TPJOV6E6fTWen8mLREUKXDZa0
ed3373CFH2yVNzbGgA0dk6g6JsLwAYdcNSoJSlVAE30MikjpNA5yRU8w2Osp07RCngsjNhwvZdg6
bNcyWx7Dj5Gk5EdSZidta407C5a0L6Edh4wi114GlyQYwiCi8EpgbFVhAV6o/7ZpjU5luRfu1oG8
0DaqbstG/FzZoETzBgwFHn10gnfA2w7h23Ybboh4nj42tUTgdz8uJ33b2RlprjB3MPkhLCfNS7Ak
ZX4qf51TS5v326clTzMgft1/FGEx82sxRboOdmFZvkFidKXwDRIihQ2bQ3RFHVI4amR02dvnsLNm
kgqcvJlBDjE95Rup9DLxpJBqCYguX6yUyJC2NFCWmB6vzmuoxI8vGTraBceiFMrKA+A35t1o9kaR
5ZaoaYxI8/rktXaqqZW3dudMwO818AHTDVTgznxu26XHz8IbHxk7ttqhgTeVHWmIVpwK7Er+Q5hY
jqdaYWBP/qPbetbLhS8LrgcgBlQKhY1cbJanJDfsfaMQ1pzrpOhJr3gKRD6ZolqMOyXXhdKNbn3X
Li3S0kO8q/rkAaffH+Frang90k6WEcKnVdw+OB35XZSn2MHkbieWoH/pwzwes8dvSw7o9peFK5ao
Yj0uYNTgpmvpCs5UhrSnvPg2sTzFlUHc3noYpIPQuChlke3jM6fKHAV0jkbI8sQI892XqG0bo2Yl
0Q1JaUIda37mE3AdebcU5DQWQ9AmmlpQbschhgkcf0FUd6oc/gLCewCMszywJ+kWqn7KrbLg7j7k
3AnAr7SrF5jmNyi75WFBltdzTQ+XWFxpgAR4qFiOL2XAofzmFLvLRoHQDgYz1eXs7b1xMz+WDHUz
bL5BW1qLJLGBFnbyOBMrRP0rTt/7IlB/Ptw0kn//81PX8kUjAKIg3v2WfD19ysLrqkr9rIVNwMSV
Ifgm1p5kuw5IYrMLyDr90hSIFeS0nxaWtDt0860pnvtMM+OHgFrub55udD74q7XXTtJN7yM3Hm09
AMnzC/6OQFJ7D82DlkBQYRRCH9k3Za4l+fOlGWXoyuBEMv4iZ29dUmgWkGWE13YcVoh+/QTMGoFv
DqvgnPX3rBgz1/bp1vEqCVTnOb1lIxdFTP3182zM54GzO+04nF6EIwiVEQS66HKVYJq3wlA64rkl
Z5Q3YI5cn4scuwrf7sPoxUwZeIPe1eSLfzoIL+frc2wjRiQHwwmDVUbKmLEg+FIKVT7wjf2ks3uL
piowti/z7XFwhuxA+iVKXYtWMWrWhqXgKjMUGr+vLy5LYM3ZmI3KZcHX8czs0PfWZzr4bbcrnLcr
JWlw8vRvH1a6p5J6rHx/M8aNaAg1q9Yr91T5uJjCEChnOblyz/jn/fy1Cw+iUEUDb+7NtjAdzhe/
Ksejh+dkinwmEwXJ/EWb1Kee80jbOuaNf3li88N/NW0TmKt+v/7WDfqKEUyOTYl52xC/oipIBTNi
xCBoUzxY4VHsVKQDE9jPdO6HhOngB5SlhwxBoOXQVtzX6x+bgXJB3zaKga0VTUWzTfxZks9HkkxR
sNyXc0gt7q6CTIoBPyiHS5YWxFQDHPlXIhRgvWzHRkoMIAuHZEu+EcObKHsQs6AJGcM4J+3NFaCA
Zu1WZsrSfrS3usmoQKcjG1cJ9yOtXUuBNh7FoXXucW5vdmUxnC/n0X42LNDq8kYqYb6GW5c5Ct9U
Mf97PfERrfZdx9RRFVxtiUVNoGDpPLcEEve/RSMR5snuGCK5ZT1Ssl9k5hkESeLqIdKCPLffcsV4
drgIpciAFi/2nYnJHQwhp4GwQGe4zezSo4HjqXRiw4HYTBScMGCJqf4oosn3psCOg2CsrFbp9FQu
Ri96D5tUKg1MasTOn90SLICnQYVhBYh9lkG4eaBta/m3ysT8BxjlJX8J5aUNx8q43HNbJPOxV0Et
PLNy12TJnUbsRYVHdsOPdH4LRj6ARywaEN0HfTfkuZCiOJn1kGdfTwsEiAfPXnMqnz7GViH/XLzz
E1vCHKNtwzKZT+50F+xqlHxhTMQBmblYL4ZosGwPu7eaQSANhC9JoUnqNOtvlmdy4GYeV42LUZuT
UMLnF9Vm3LEN52ThZTr7I0eB83bLeaxiQj8zxcTQz+jmVAlS++Lkpem9R99o3iVc3NYpUK3HJK8T
30rlKv0b2dpPU6nqyS8CuhqxuuxFGpkk2+G8tYoTHmWAmsd1OZD1qYySR9Fv3Ux/dO7fRB2AI/RP
uydybEQqpeS0tDxooDrk8IiE21ZtKpHJDqN5ySWlrb/3NWg2++OeZAGVUEzbTHbHsd9TyFqdVPUo
b9NCw1EhV3p9mIJREx+hXwmap8zivTr4T4ni63ZWYJ0r393gEb2b3vqRICwX0/+o3GaDb3KyIdVF
DLDzmoyx1asFcBub+oeCfDrDi7vKnEidWJuTevC0HCpkEentbVzfh6tc6hnkL411/IqV808FkhZ3
GXU05HUIGxKsL5F9fIRFjGggFr59yVHbpWIGrxCvRyZQ1TfLnzUlYIe1e3IFyCyakVVaG86pm2OA
gxoxKOV1W/sCNmZeaHaOjpEuWfOZWB6s3t4t4hiqb0iblBRC2NUPmC4Sz2g1HfWrY+iGvs/ylNLi
jNUT2h0On71TZXUf1ic6fBOkDPC8vIjUW99B9RooaP35O8eveWOI6TAI8D0Z1chwW6+IMHsxMDTo
9x55hU2BSGOh26gqXLLICjK/hw5FRDaBH2ttVCgdmWwsx5thKM1RV50bM20Enm8ecYYpBhkD48Pk
wC6IrQnJJLyQG/CddHt0CJXaVDI/i0yIinM9tMrwnbCqJL5MGS97JoSt3i/X3iYm4HAlvYAYQKiz
kmBql9M982pCoJEyE2GEqRtNUizugq+ntbikxaxnl6SOf/Vbz6xAbKt45wGUMD+Ep9S49CItATTs
qoFt7vXD7uugmXQG1hqURS+bkcpmRFW+Wp3FRqr+uA3kmWR/OowrseToZIkmWiws+ZpyHZWEYfV4
1ji7pvNQEixCdNdl5QrxtkgYaxwEOgxDHhBef+BcvBMSjSYz60vjGmlsL8NZ3OhSvUMkfLiDcYHo
3HVVNz9cZZAiRxXjXNSE86PhGUBxOK5iD/AA59z4d4WRTLmSKQxbd3ZErTENjKcP/rZbzVcl+O3j
XKZLIj5Fv233j/Rx1sY6swLqIbwquBTRKk9FR475kX2ItnZ8p3j9K0/3zmcMsHACCbOXtK8SzVyW
gtB3OeAk1VnZynXUsyMkFTLrwG1DksiuPo+toEoV2H6uToaAXI4eM598cVGcTnuoNOWGaAJwbBFG
e3E21ABewKIJaNkykZc1eccImRhb9hX/FY7WAc0M8NM4wos9VpS0Jn0T+LSGQzIxZUEJOavByVhj
DR5ow8E2zuOkT3ndxHYXL7Jf4Om2PtCYoDK17CPXrhsC+pPYXztVDxni2Ffv08rPSiNkylZmKZOf
E6C3WbR+RDP/5l0VSacZoYPNurjzc16Ox/26kDH6oZ/MJMJi9qoh0Ahn+rj7w8zh+U5MhLKiQlHN
XAtKpntErx33Q45nG5+uZWeCGUziLwcUxYYaXLeJB74BpcSlzwI0yAtma8o19zqc46zHVZ4GrbjC
Xj9dw/RYCTP0JCTGU9AJVlLhNxzfKxe7LnkEGKiX57qIJXPwlTgBC1cDCbv+fAW8TVAmKLT0FhrX
nWcBjw4WekCFYoX21CTTLp5UyvV88Z7foU9ihuiyuaZZ1FdqXqr90XzJDGn2LDHW3txxGaSLO0aZ
oMKp33FHpfyE/WWCH3BryUHsJz8eMjnvLY6JPBWvAA6NkuDKpSQlw/V1qzxBe92hzH3YRHJFrHMK
rKx8D0TarH5udpQTmv7VpETup+lzqPLGKNNfkDQxMcP9IHHxGATaVcJaxslyiwTuRO3jwX45gpDj
yVtnDnDz4fle2VvmP+WlPEjVnLrgTAj7Xh+uoZaCO7HX5yugJZ7Uk9zHJtPDtVhaYs/MTQOAU7Ul
L/deHZoA68rIGvyjSyON9+sSQYfkJOLdxrc7aue8wK0Wl1R4n6v7BukxujjgC5ye1jF0cGNh7Y+5
fXIbuQRHY6Ec9tGPF37Tmau2z7rZCMkGSznHiICIiraXMBN0EvAXINcxn6uCp8GkSKgSGRFpMR1U
V9AG22aERLGsZrq4Xj5W3mpC7VhpC16TS1bYn2uJY9d2Z98ivVfyltyVtZh/aMUiRhbsc9nk8E4A
wa0AkTcBe7YevU8kaDTXiTsl8Yu7X01aRviuhKEoT77dvCRRBpGCpLW8BNRJ9GtQo4a9qvBCJuuy
pn7a9i6HmG+ReVx1yNzaPjhGkR7jbJJ5tgnU3uhQvJ8UTaXdngVkIK9IHMYXtUlKj94ZWHpcE+Iw
B5OJq8L616Qb8nWwWrolk8zu8dWSE0BVA3/U4TCMcG9L0TJ3lggjSBQ6qIKlWJjE1EEPFYrYvBCg
Y0MGAk2cIlIbpLQm21iWrWu2uwd8M/9R/oakNsImF1UHl+PrROduJJSP25dZ8/7ExZ+kIgkq+eom
8kgO8vng1BbsqCw4pd4dL00OhdmVrtrcmCWeecGIldgA1f8D55G1ilb+2Z/iVZ8nN3XSOVWLCwF1
lMOJQLYzsuOGSwPGEG05txSmKrwg/nX47dhIDcdaTQV4mzjBspz6dq+KePeoT8Bu6/S+4t/pxqfz
9s73Tt16lwRnhvnAH+kju1TF4UEyhkPKgc3g6Vbx2fHJLlFT3vdK/ZecXJSiDXRZPXwheLl+srnh
PqRmvd8J93HTFP8qiF4QxzZdJAAsiJwYlcnVYBnyPNzteKzJ98a8/5KOh2EyG+P7yZWsNcGKgTyW
30fg9TAOkN5J0uMZWvfX+KkfUzxtIYqrmxXF5E71OUVXWygOmsrRQTxj937eGP70hqoiS9sZGuUc
WgyNvYU528GcgvWgcvsBWVJINc+jVDfPAr2+KxlYQHfW0aJ0j9tqUDHrBpwOOm7fgh6n4OMW9ndB
Y7Br+AY4uhMxVJibT7SiJNWM05baDln0zL33UbyRFNbxw3zFPJgU7vCm1FLm8kMXUgvS7Xo2Chcu
umA9MW4pzVeD/fVVuFtEqiHO1qRZn6srj+VLzQWzFdsaBTWzZvbKTUfydi1o5tYu12KhU0/YamZG
PptDll1zTNIOW3yfscdgc926W2c62t5nYxSOHmNPvpUG8EHsFJqGtFCj8zCZ/bI+sWK+Tzp4Ks9y
zasbFLNtEOKU9f8A0aqF7gNQzfgzQGon59tsQ8GNgdyeBUFyZGJT4G3H4N6V1ZlLBoT5/HK3k7wd
vhme4jqy2bkkOpr3p2SXdS0i7tH4XJAqo0B4kPmPPyULeshmDKEriTcbeuekb3Yl+eMTXaSJpolu
59gKJ9PtBJKml2fIUrL5pX6CTQNyd7hMYXKCJa89t5HUzRtoVbQpUWM1HHx1NwWdfHwrzC8uaFaT
YfSxPQWI4zyMtki0mzX6lz6V3fHS8dLy/xSf22+c52l+49JqZMJOt4pW06QGWSrlCum/724hEMh5
0jNsPUhvfUxO88B47sF4bbosFlq9chM+9SImIhWiSrXNlBJHtc9i1uCS8cpHkvLzHawcBxpZGmHT
NlGZdSfbJRH+EB2nK+X8rZl6KmsCEFjwXTeMDHbP7sswyMG74DrKQKfEuaxG8cByou+8AhRyqRLD
tfkS0hVy/znh4wospJgXyZmwGp5gVvn8bs2CnbOGqU42MVTGEBURr6PgfQbjr99e8pvJaQelXAdw
FNrBPN4cDFWetJXfwkt5yEEjL/j+8iOMDhvMbPAwPZ5yRzBUS+whUQeo9zpOqnP0GDWUr5vLu2UQ
LKGkminsdNcsyu56frvrxXOFG8fyk/Ad+8jTZxedIQEZH81jKN/rr9lRfcZw32NMmrY0UF0MpumI
RnCQGaVonuP3pjbRRWUrnrzLQyB94vAV4COSByrkIIjyvUrdpQQ18sRoXHh82GYMc+xjEPc31XrJ
0Wv4QomjHv/1nBWSZHpje/8yHLLuJU409/3u/JiOtGyPh7z/BFNDnVue5CxkoxKylP8Vr2je53XL
1VeGjFU/a8kYTpw3HqeMfdaUaC60HaGFjjMJDg/EKTC41jzYA4MmAiD83sxmX6Sx7bG4otg4cyI+
+ZGTDPImRWVR7jIARnxmQnQ6VUYgu7s1L6JrGoSOK0wumya/RW+Po/+Xp1Mi6xf7KLb2l9iaIU8n
rI3phAKI1lHI2AibtKy9ZE7NjbS/Ksw0jAm0MPmtX1cUMF7SOOsPwvkr5cfiI7QhOoycPDSoAL5w
SUfa00KFYXZ65jsHQcS4WkLYvY8ogX02C8vkxUXYtzfxVccLMsLG9u1Qz+41NiaV6EZ7nQS94Q3Q
tNCHgXU1+K3jHwP+jEkJpm2pEFOoVqbfKSvzge3IQYX2bvhE3jhH3CiILhSkrMPximlCeEe5IC1p
RuA5VpuL2DXCgI1cvWuFC+tO1joXiwtNW2kFPkOkVagmKBFvsifrVNS98CLJfXtQbZFrZCqRxUSC
b+xUeAiPC1sCLCj7HDcUEQdkwIMMLB8DfKHIvjWlLy06vqs7ttF2iySqrkAXJbBXJvHXmCUYynmN
swkV5zFTfwqqcipFXTVTXQWSBBoOQu5JYV2CXnjIeej5wo+SF9L5Beun5zZXTkMQEO57YVsgsfNE
E/XGdzoIqMYoJb88u9xjzNkCSDLgyNE04uQluEky9I1kTffkTDeWj6DO2vYPVwpG0tGz9KGHTriR
cEnl6nkR7N4MSu3wpvT478qJHOVwdp/Hd4cMWYfovygSpNU5s/pxoiDc6wsqdvMzoyR5QVC+BMAW
5RCejqIqXgHFcEOEAWfxD8uHvCRySsuOzW2WgD89ctY6eb3IKY6deSKSR6ND2XBJ17oPrkXsE/WZ
UOf70a+XA2zdGCJuYaULHhNQaRhoB1fXiHD4NfVsQ6LG9rHH8gUpmJli+/VTv7FDxEunWVHMy8IP
4MsX9p6u7x6v6VcRkrSh9gAYZ4aNq6ZBhavrHEIPyo60l75z1golDEcE9znvgO07YV6zPlqJdXwE
1ozkSJR1FogBqRT7EqHplzA5OWRDRMtdGj+SWg4hxF7fLLzeqDGyYG6SyspqumJXEcGrAEZ1LOWO
g2uIW/gmpHTjdomv7MH/FvgZ+Is3iMqsO1o1IjYnwvakPNhiUfhcgdVivLXjaWRyAkZgVxBPwoMi
f9djDQnG06+VPuY433V+xN20X0UeSU/KsEOGf7ZUri7IoVItV0U48rAPljbvmxYyOBf5fI43z2nl
CKR/izHPSjs9FSBcOMEy3nnpkBCRr2bFKLdKwyGEb8gzPq04e9ZGL07w7CsvuYXSvGutYT/f/2qy
prmcLJ+9bpaNKbJCWkRsJNZmreWfgLqyE45vTadxZYtJVlpBmtO9qONaYYExLycXNT8Bzu5mMvxG
b7fQN3blxGZJ4ekgqBArXdjCfoayfMXplEd3Yuw+p6vQecdozVI21fbMrExgq92cWDWRWbL2bkKa
wuaiTlc0liHOgg3a9db0azqw8j1EXUA7PeK6b+y1hrHNQ5WJFb1/jAdCOJ00Z+x1FSZBLpeMH2LH
Qn36vBeih0juLTjHj8rWlxLRPqwcfdKO1MMoR78VtgMJGy6qc89lyXvGzTFsc66vKlVbP76YcZZ0
ruSOgtbTKS9+G2nN0N5lczd3WOcmqs2/3IYMDbfCzEGHTtXqGY9vjjd434WsRJ08lCl0QXicO8P2
bs20mzsDZu02L/yqj0X2u3thnLuMDZj/kMzGIO3SlPY4rx284sd+jIGETSCzLV6r8g+JHCHEI2A2
sSKqezXEhWkXQAVIlwoJ7Bl6Fetugb0utM8u7R+0c2MMxwLs439400gjrxOLGvNxrcgAyoTEU+S7
23u1SJALALwugU2KuUOU6mvHPzoAC+7bx0XM7RfMplpYECv9w1nlwLyq7yPbTLRqxdaoCKFSR5QG
mm9MGSj5ADfFAVK+NcEdGs3uhe/9s9/jERBzVJ9sA8+XyigEh3k4L6z5N5slneEUqkSkHHR7z1tD
tOGIiwr5KSWs5mMehYANJT7f0Sl+gBoQvszxfda23OAuB/y7a2u0jOGDQEkY1g9nr0q0j0J4/kwk
rq8hY/IW+GvbEK7YkNtGi247DqpJsr8cajPERKAVzlvX2Ru9Mu4i25/LpzQ17h9OOOx1GosSct10
dTDpXjhut1VEVh1xgY6UeDfIGSbmdXYkaiBt/dBG4AicnaOwmMU+LXuYq0f3NRnPTgZmUdnYInmO
cJX4icQQSkgeaa6GBhj0kcbZhCfB/z7TV8dHy9rTCpzJZVemYzrHwa7eV8wnl+MO1b4AQwCTyw0g
5yIHl8XErDUIFSw1lRmpIA8xxmimfd0SmDZbelizKwN3ovTx+UHoRANcNXFDHYFkMGxcI3VKpy9o
rPc1QD0Yw5pl2agn4wrJt9gwTYSz8aKcsDr8KVTIDmxcyQEGy7mrFjxPhyRCaQOvaBAbFMiusvrK
R+SwkpUPTwXJ2jno4aUFzoPRRQFSk0lijKDuLFlUttc0vHhzkykwo/j7No/KYXj4lh/LHQm+k7+D
bcKtsSTZVyWlFLxB7+Fi6GIMuIBeO67KKb6yry5Pzx4j4Fwbh/Sn26m/kN/YUbbHYRGEZSlqqMBg
62MeE5JEBkjIKFl9YBobsbRpUa93nwUsX62AEvTR3kSHEXS+yfw1CroTw9cAlm8SLZc1bQTcSg03
4engVD7twSAPqpSeiOrjLq+pHaBTlSviXLdTTNurQd8A0zteDHlX2z+jXtosrl5rwEghUjQqIwky
aRdoCXlLRmSNpJExW/KnOezFZyamJXhyJ24uD67KF8qNZzHmI6V/0pvzmXBr4o/dnkZwP4c/KF/M
nsf4B/f/hL5j8xVF4XUSZ4NDirdlleqvDNqjlpRWB2cLjIzxvMr3FfkHeEwSkRCPtCznQn6wbniV
y9IdFYZMQsbBEexRK6pXlPbRGuFKEOV0xaegADdvZXsY4vCozSZ5TMCozn9VjoHtgvOt6qZ+2OlW
cqnMitfwXcYZQD+Psye0W8d80fYeUZiTZo94ce1y92tw0hRFwRwxL9wdK3zkBmzNTHbJTq4V/bFd
2eovnisqIQfmxyg8tbkTD69r2dn8UbT6jIqWGAu4a8H7l5APUgnGIkK+54XJI9bTnTMQgqmao7h1
5yNIObnpH04CIY5tCMI/EwQA5DLnLQ8AdgkMmB2CGd69Or0TJhg7HMEotCWw2g1l4z2jVfUt1DOz
arze1HVwVjXreRYJcRsY77m4lE8gAMfbC8OVah74igevKaMp24KvsZnkapCrAy1zEvAZPozmYTui
5vVi0L8al3e2FM/8+ls/s6QVPUqkU/alWfu9FmxWxW4ILz2EkxbgpVooUV9V4tmSX3Ltqo5uX7Y5
OtHCAlIE1x1tVII+FcZ77JpaCTJ7hQELYvh7Epv1JFfKw9uSQyWzo0ZBmTIjb4qHCstzbhwYyhOW
efEhuwuxrG37OJBjF/NJi26b1cnZYzsnIottAFQ1j7GfHjoGsCV3VcwCFqXLBpPKUXFzRFngy409
MdLBlnBni1V7GWARA1BcSLkEJNIRO4vpWWl+67CK7g8N/sewc9VOj1eayg5xL8wiSoeYKEJiqk4A
CM9ZXdVbs/hwhYNDdfS/KhC4Alf+Y8Ug3cKItM18v0FkWdqD8kEYgDdoA7KWZW/DnMCJBzV20ISB
XJL1pnW3nKcDRj9cH8o66426aLrRn2YIMqZ3kwB4GVmnC6pk+0JIafhoWBvezlkItUHS9meyh5U7
kEW7CuBW8OX3yyVCjZZNDZoS32d88FLsvEjuteXo3hHy+N2ZgYWOvxURNDnVGzG1BlTfdjoszK1m
PDTu57++gG0RoCuScdS7A7fl4vE/np1zQ3+/B3q2cHinhdZkaa3cG0twUY99PTm5WlmLncw5KZiU
ShEx138nXzaKzqVYxL3W/hhVSdTKMSoq21O/hIA4+jM1aW41AjpuueKwI9Ggl+lzArsZoP8d/F92
VUzl47xkudHdhnxcioiFKpj8dcxDOZnpps551xRid3kzoRaZ3ZLTHvfQ2jBLIhayofYmzU9web0R
rpMn+7i73dlwAwc5LoovZNjp+TLS1qiHgMgb6TL/okd0v9NyBdT7UTPG4kUq+KZsE1SrXUKADnBo
1IKfkjU5Z9ie1ceE9a9uENI2ftslgPg+VgKV5rjuk+GsMvelZ+O8e/VM7rQ9/E3PFv+MEJKIGElM
JCif3JIDA06XXueJ+aARTMGn/7Ao2S7/gX+2pSg3cVE8wWu8QnvVVSndMRvuIW3KNyZ7C1uuCqSi
azPV5Vc7sCF4qL4Oh8zFGffsXAStm7kbM0K6TRI2sBpB6kX7Clu5ga742bQiXc2DxQBsv/ZsR98v
Qk222m29hQRAxJ4x0Je5Qe4n0Xv22jKIOWOqyFp/uYoqmn+9I2BwH6+fr/+Fgp9G5XTMjlQ1/bbQ
TXODaLgYsUKrzJMoWjZfa2WiFNgyJVxjWUUvjc2Qcyq6Zr778vLiwaMnbMQ6zCxkUNjsw3Y0dr6+
PU8ul8u3JAdir1ZcAGhYsCZgDP2EmewuVvVjeyuXO7QU0hbiRzm+IIpOsse4zLitJrPP5u8cK03D
1w34PsxR6aEGLdLkQImW+Vc7ACwl1+OpAb2jpP0bl7k7XatTVIugahjEynk+FU+BrxwRzVgwp5wg
EiGs8PgXzdi68Czqrtcg2r+7D96x0EZY1TQx79HkDxT3IimbZgdiJuYS0ulxCx1I840wN9WY8Djz
D7/b7oL/eRvlZqd6LJXjC2oCTTbotKNoyec6ddjn79eyYGvR4vRXPY1ZfppS86iID/luw5bAskWY
OoovUdol+50C25Bjz+i9P+zI6mhzly3H4o7HqxUpoC2v4P4W1xTmHSiZJO/JU3nWEejPNHY9Hp9S
idVVnbVq0/qYQ4wXo8dUJZVM/27b6uxY4ofgtmJDFwe9riJ3gIPq087Z3HvEYhyblFGdudDEVqdn
3jzWuVYE/AkiipgCLwjNRjSzZ7MRPTnBAKFOl2GrUn3GiLphcy1GNa3EpnJd32XgPRAOrK8+l1va
90mgk9r+MuuPmLDGXStGBsghgo5x8h8TYiJFKqbxQxCfHamY1trexi1zPqvN+lQ2VxtLDUWqMGww
kEVNUv3MwVHBvKetSHlHtgRfoaUfiLZ9+m+TBhXatEf/oyiyEToEYLDHWTxf8GpBDUuonyTtneLF
je8VROILLutlEe7SMxh59brOKj3ihZp6ALmxA86fjSQsGhibBCvM8qUsGRA3UFNOudYwefU4f6Bh
GQYq2kcHO4N39JAUWT51FaRW8zHUohWjwSWB/ejDxPMyIG4cLL4sMpPaziP/CJRbalsP/ghABdTL
zkVUmgRfo2nbOObdebM5xO3YwA6X6ALpuhC40GwZItW/ErfsFGWBkmMLpVPTg8QYoSfiSnkMcvyv
/r/4Ja0kH4Gxky1ucvE9ep239c7eg0M39GGE08oYK/q/OvdcG791o/DyZo3mis1TrdYq/rlZGdZS
i0cR5xTi6TT5fjuneFR0SVhHQ5Wx8MUUeBiiFEk2sycD1ouCdnJNxa6veAdclrbkKrKARpuV3iOZ
WDWoBN0JbKtdO+hiEMXERmFSZxiYl2kTjZw88x2eZvKMkTn7zA4uEyoS+HGY7tQr46vWOU9kBjKc
b2+ayGQQGSR7u3zUy8VpjmNCeVvuKxufXIGNsXPZE5HLKc/U8hQyb8T7+PO/ElZ/brogOiHXhiy+
lyvdMVE1uyEbllo0aFvnXWQikbQDBEY9OfT01p+dHuINVTfkb4G4In+1SCLiFv3GFPlkUiSAre9l
wtbK17kDisXwrwXi8tXfJ+JdJ48cfk14kvCF8cslhHVL+YSSWh9zKBItMZ4qjMSQ8/36l1gmNnUE
GvHeozdBUKU4VL9iAHPL9Zc8HOONPoCkPQqEYCyhP7uRb9mVpyB2PqdmHXE5kQXsOYxJAo1jSPee
A3RYSybbHezDFbDAVEaeXbhINFnN9Wu0yC58tBej6FsR8cSMFPh/1fMU6RR4rDOYr8p7NB+dm/pe
RssqYygxjWbOZelRx7Zl7FQPKsTyUyMjVvkowwlbOhTARW3IDZBF9HSxixd8UHAb25zJFlVz3Hms
PP4k9dFrdbqEGOZcROi9Ome7LVFq+5ORNRPYD/lD/vVlhX67yEoBzQmcGTQ8Lv8F1oeLz0drqEVq
QM9shits3lTuah6QAO2xyzqRldts0uF3xazpZbWPky0y0HynVvSKjSqHd9t2K9LN66wMKTF8RN66
uGTPDJYVD6AeNsSTke9MJ86Dr6yR12sjjs6oMc4vwM82FU40MpP/tbjUz2zE/NoU0QQ/ci7vH9x7
m/wivzpeKSuIMGxIcYD3eLz78uApEUvn+HBCrSfQsjUGfdce2xoyWDx0zzVBPWcXTFKE0ZOIVwwW
WmHhZLFajH9E/+hUVnavp694KJMcprSlWSXfn6g0DcPN2uMVNYpVRe2TmWXtZ2ajEsvWPLOMUB3S
KxBko7IqNW6BdXsMzZxolcoAHp7fx8tv0/KSwSZ4cwl4bp6yERG/lpJLG3/JsDRYHsrRQvFZmyEt
sKaqJ0AwD4XgFLI+2jnvt5KNeiabugdVije4jj/2nnUuBdrKXMfInB1f5RiNxXG33ziuuZ1CL3X8
Yx466RCtn4rYdYCZAK6e7SVp18zTEXMqV1guHgstwK2cTvjOp8us6385Cuckl6/Rw6lqtQRcrh3A
rn0LWjFWQojgDsR+J52i/TtXE4yMD5fg0/QhpYq1saDsVs3QHQ5mENqURKlQJnL9s+QVictPVoS8
2Rlhc7QXd7TrVNJriACSN3SD5Nh08aCdES0zCAJ9eqnOLDn8XYsfwGrm09hbGuCHBFYa//sMMapr
9zT4D6wnNRQtF1/fRY7efMfjVVjaC2fouj16BirlVNCyldBfygvjpoaUQ/mS8fWoc9TYaCIBkLdS
3TWPlGq68RR3x1Vi+CvkSmfKsEJaI7c/0ggNAE6xHJvI7aG6QHDBNAdRjBFwuNLVBhMuVtM5GzLC
nGJj5TJ+thcMbC1M9cBNb2MhRywE0gAFq71Xj0bLAzPpxvAyKutNIC1dyRZ0o+JTrZdhRLqWgZoD
q9GBy6EgH28CWHIJh1YKeM6fdyt8F3H09FyQ8j5qsZqGFFAjrPerXg1bE4RkzGy/EuDOwBqGtEJm
yxhwc8V4uAEcDRpNjk81HDM3P70KmsME7TKvH3kMgNPG5+lIaxAay6oLs9IQbUuUVExr0bz1sI7s
q0/VwLtwY6UKjhQttD/Q1//1gF75fiwT1+W7yrhops6zzpq0nysDjxcGr54nO8yYpLXKYBS1inAF
rWyKNvRSKBlahZKN71uPUl9sTvF2tj7/7fpyOxULQkT+Dj1D/PYQGv8MxCdMZfoRUZqem5qymy3U
egXiQdgHI9tfxEQ3vnPxaEj+stR45shMJvxp27Re9OcVHGp4yd+EA1JSDezWaZyCdnGGIbqigQjH
nmLJd/cMO/p4E8mXmguJS67S7+2baTU/KCVONMPXAGudSvv0Btp2X7Mx8DKcppNsZ3NySxv5hO/N
CDfqLneAz+1BrcjaWPqKH0FDgNJQpGjVatG83XR8zwQlQK8XVRbETJbMvOyYhm5XFB5KRiWTDhxb
7lvha2gXIv94IASY+/BFrBBBMKNYihSSVb3rYNKw3UrFwHGkThqb5LhQ5guiTdWg/zJ3CsF/cHQI
FLYaTUZYj76m0uv5qwLwk8VWVuj4KzVMJHqR/I6LgVDEtAIXGJIay+ovKvlCFrOLhLdm+OKCeihr
P9KsUUhID4chExyrNnk2rZFekU4LSpA5eR6HfgTBwg0iAUqJs2Hcq+NBtGNXrdZDWu3F4bGKDOT6
lGYGYbhUcU54RH3laLMQ0B+/cq8qRFH76XwGh9TU6m+eTFcHqb0sXkUcgTRXLBMgAhKk9VJwJfNk
vSDwgsyGM/lXJ+rnBWlNhxWj9gUv0vfgHBDBCdvRZbh71pu+2zjcZHOcZ0YdJZQKmybsI9JzQREY
5ghQ2WXyKybECeQCvOnCxzBFbsfF8/mIFOSzW86LnehwfySzpP9YJHvsRy8axSTFSUu8tV41WdFJ
5i3AjgfCqFljhWTRDYUh+t0pJgJ3KfAzDDUlPVpBQ4k7+EwDhAVfirOX+I+oOFZOHLgwxhKpCoNs
c8AGU01pFrNxZiyQMPVLsTVlIwSGgi8fikO0f/5FUEuHzQ5NeoEa+64+1eK9IyZxAAFoYV6aXHkI
1tubKacHtZQA53O58S2ELaegXkU5PhCWFejhK4L16765C8vz2AsZcr+iZKj+ZFqGXRZFjm9P+k0r
yru4vVKARFMS4V3B56PfmmCMo295O8ALfWRFz1fRJEjOiDEnLjQahPvPcGcUxXIooxm+9oTKz84D
EBAdzUmEwUKUtj4C0v5usHaaR7NyjrJ+1pN+iLK0tbo/0oBqgFjXltBlDVoNHQaMWs8c1H2w3Qqs
pERZWt+ngZfv0PVB2cegOgyODt0bsRdBSYYZXMMhYI8Sz/do/BW92zyZonsjWtMRPALYWGuqw6GA
5iB4dXBteH46TAoFOIJ6I+Cf5QSKMnJ27GrwpBiFkbiTbSbAE7C9v0QABjTQbzLqcRygRzIB65AC
IkVdIl3PmK2BnTOw301eRM/uGVhXlqn0YpswktNLZOm9hSnScojwR0dkyy19gJU6WFu3Cx2eaBhd
rnWJFpfNC9avMs0JgjCd/eRdowQnqGRbdUMTSprfni4Oc4Y2gh6GFJGbm5BPvez8Fdj2hh2Z2GBn
GJKk1ZpUiclE5tIxuYcFXhhapGxL+ajPcEEz5oqLiSqj+h5jwO72DmwmzC9KMMQa6qxqCWnuvlXJ
/prJErLKQFlmfPRi82OM2yKksL+gO94wfCFmfxVBg/2Q6QTjVPfYOSdEGpWgwwM97iOYE+2aLnW2
hn/qZz1eqUuKoihBa7pwjzk6A8HoVwPTrmcmljkbqxaAXRnJ3TvvBGNkZTheCBQLFElIkJHV1hWw
zi3VAeNI25VC+KLcSh6k2y7UGK4HjULwi+OZNXjwjzB5XokmPfmrhlJFI3nCFNUWjRwDtcueYTyl
p9D2musXzMENym2TZaxg3FhvK1F3FsHnvTaRb6pvMG0nHcs0G6vmFB2gF2lH+cxz+9iZabBJ40yx
HEyzQvz2nNVpeLG/QWCk3B/+tHRB42ZQG6REtsssF2Obt7ggywOVRWo1vIMufzCbh3MAuljBOBzi
+AmceU2PQPmoh6XDmjv407dKN4zGDOaTraOx9KgWmwQOIHznjM2wU1E3G2xaPiIlU/uTFF5iqmrw
mV1S9JaPGE38vFzspwqd/uyLXWsobNOkJuUtbWmOFbVEkOS25xYH4N506rBT3dwy8uuvAp+NAR1W
pQ4lE74pwNCECIGp0xNxLQxQTOFwMGgkXB6KyndWF6au/xeoJxrZgnf4v4RqDCl3z7HkCVMv76XX
ODFRc7CX2v3QYUf57YyurXECgRrYhXu//picfTiqvgQP3sSIsFudDDRdY4XcqjkVXfD1CYGrQ7kB
jHHMyaALPQjP4ao01W0Nh7rUUEGQPpdE6y/7YB55fUIv08NHsw74bKf/Ffju8p2IdDTKSqxjnpZ0
VtUNHq0sWmlJHXQNVcI/2gvHiEeo9eFTpuO3+ENomgCyKSJDfJsANjOUK2NaMZ3OlM5nx9RBPa8o
i+gETiDWbd8/xBi+w/lwNE46HcxezN2yrkj01ouWkKrJMM8yo3CRlJKHlscNbvt5q/i1y+i+K4x0
ec2sj+Fo13CSQI98wYIKYlERDqY+ykzFzHASKL9UL5/TwLtMm83JVGt7JOgXNM9Hx/89Gx6GZXAx
N5Ms14FVaEPUUXI1bmp1HT6xesbPEqXcMPqp6tsIC/b9nIzN/T94yZHQWBO1paVxFQhfdBSscTUj
x+OwyzAvsri11D+Q6yPsJPs+eUOV1TvIkVNK+/CvFnyY6lJbY1hR+uZsnrT2e9Q4vpWkSZl9EMpu
4JHLbZ7cjAKTDZVRZWwWT2RS4BCRURSOIH3o7LDvWxMVhPktCLO33TIyDwoxiS2BeZA/eCmvDrWC
aFAlcrKFDZY3xl85v8m8tp9sQgWJCyRySWhyNsDp178NA0vgJzNxf6oCxDOytQlFp5xmSQd6mcnC
/hs2kXALVkdU9eF379XP2hB0CtBMYe7PlNgBA02T6FsWycLPg/TwdYtRM5Q0RhVncUL5BWqll8A8
FzRUTDAY/xRx6qj+GVwPbHREDUL1BmES/3x1T7GgUXl5Yxe2X4yNl3q4IaSY1Z8MAwqG+x/DVvRb
XN+sUmRlKihks+8rK1/fkh7yfrHLwUqv6HvwpFFssYUQLCJtzVlqCNK+hNTAmr+y/AJe8WIlyl7B
hl/HqenRJgWZl3725j2v/0CdnFz0tAjKmIMJNVU/2ehx8dQBIfr3k+C8BeMIW3N8ozaTmDM1VVkw
/jvEDUrYkUH7ox+2Jmsw58ig53o10uSoAKfC3+sQQEv9I58XmRVe57rah7bmohNv4f53duYH+xUz
e+Zda1YqDjM/8lO9kDy9orTPE7NS50Vzh6xY/yNuTaPmOZvM989juz1UFtIGPlmRUAvCL6J1dyEG
Pxpz829bTLwio6HRxwj84tLyQak/ISoVSfzj7i1Kq62cL/uEjaa2MGRMQF3PdTZHWjsLl2ayyF0o
538QDTCvwFQY3rxrWXA5LhCBv2IYL4rau/XIAgChb44cQAgPYTR0ZdPWUcA55zvuM0JENvUu2plE
2cQOGMzWnZFMuKzDeTdqyctFb1ZnIAawxPTOjGB8QBPrU75ptie10LImBiT+AGYcr0SWImDWbmsd
vkHbYJDi9wNUJuSvStCR4scmVWhQ2tqOUUztfpOCBXHOPwR/gYSgOvYa79hKTE17UuFO8dT2B4w6
GDEQ0lCOCc8o3F481/0qzx8AEOuvsepSH6caHR0hKkQK0baEXAP2rwMp6rkT5p8Nj2fPLIz+jKlZ
2c6l4pgmGMcihtPAVKqlZnDu/44UJ3GrAPP9NEQVP+41OxZSMQoMzyWkfWUTlI1DODJaYG5oBf05
WyrkyoLitfYq6tBDmkLY+S+DIJrwUMi9o1CEsXl66e+BlvmtcbV7QcKDfngfhbT5RRZqQbFLgwTS
eOnAx+ahnTaRQGZ5g1r04o0JvZPj8awqTkxaQq6SWnOht42XiehKmwzma6rCT2W5JXyfV99CBUYG
tt2Ae2DlNETBC4pq811oXUu8C2CJqjs5ul/UuUkjLriQzyXuPFivOL39YMg18lrWPXX9yToXl2Zr
z8OeUSuB8neN6pIYc8y4SMgkAmoMXuoVl5bJvW16crKq72pQ8168mJam6uqPjgbiB1kfOk0KgXGG
lDCIQk+Z6WFIJDBZT9j5LjVLs++Jc7Skjg/7pOYslAwJNI09orp28J4Zw3qnV+CrMc/NxlXIgH9R
8G0RmqCoLJTg6NsjsmucgJfzj6Wl290EJVbOqbfJtSceMPKktEkJkl4nC6Gsf4Pzr5fzGR0hY6RD
F/ufQ/ojJsj0FGMWyslxvqU6Thr2NJ3LFxvfl7lcRMxBeRDqIHO0szbsyWsrAu9KZsib7eU+tkNm
828kB6EQF2UfEpBFeeJ1Slb5TN2P+786sBdsE7ZtzIbcSnqBL9bN8SGdxCZddRgRnpUDWSL6JSlA
uemb+FyPtXOcxzZuxZyxRWXrYcjz8hngKMNZU+tsnO8cJTO2WXDIoD9ci9TYWzQD/d4lvIGqp8PX
8hrdSoaZ7bQXezXrUpiD2GFLFc7D4s96KL/tgXLzuniXoLo+uF8GHonZWi5V3V3OWX1qbd0R3dnr
x2KLlnfXQnSIssvNEzPvdLKmYz86oV9rg5RH9X3eLnj24QrcDrKWistUgUDHv1imNZXC9Yh3gC49
YoEGL934AiNs8kRpUKOvQyOez+f6t7cQNCxxYGzD2ld2Pv/rn7SyzM0aHV/pOt8yDjU9tqdsJOTw
ZVYGlDzfJddgD5zpTJYk+MvjYtYemQDkZECiJRT9o6PkRgNi1o/8IYIdWfzdlO2tdR+3dwKvlNDg
MMXwKskdeNTHVhIKup/o4WWbByavw7qlLPNeu9RHlS6b4YskDyme5UAq8PEGevjFInRnW3FBeUWg
xe5cpWL8Yho3mMs39brPE3/sv8FOrwRU6m2YbDWWf1uRY6QI12rhjT59lNs06SAepV4+rPW8esvu
FE4bz2VMefOWRPXCrJbuEvNxXwCeJLtvRm1ak+MHk2vHuh+IP7LN3cY6NgSWeq4+ahhJQrGb5BBi
fj+pggNA9/UDckLI+0GLLtiWk4xVypJuB9qWRSq9KBWLTHvsFbVhjOkHD6j6d3wV8xXCW851sd3+
NUFwlYbwWoqWmOOwzgcEp14HONc4Gl6rsRcbhwSWoDxqsegS5yHtlU+FgR5E6Lpww5M/IsLN4hp6
/tlbxLGTj9PYInqhZSdAf7lqOUC+t+mbY/CyUBFmNyjnuzSTivPB40VcCx1loUSuh+lO2Wz8EjMo
JKDftcCXlMSmH4HXA7y59pr4cHZ52kBNmuVBxkt4Ky1V0WNETar1jXlALbIA9U1lV+7IZ+e1tUuU
H7glSsVnxGxVDaVm4vKwUul0HJ12Dkjm6xbNYJHFOklYNwZ00z9/6P0ko3FiNsIiVfwSrmHzUEas
VzgvRoPk+MgHgT5pVPXzvC5BsWJ4uA+CMmwJQukwl85a5UGPIbpTNVrCDA1KwCAYdMuWgUeAtnY6
0Xars9QluANbCHSbh9gbtRR8FG2G4uPHYbztcLguAbF6ivub+Lcm0aJma3N4NWjmzi+eqLSJvh2s
jYCPpYcCJAq00wiMnGKicnorexT7aHz1T0MxbAr5qfRrYtWWzXqAco3U2VLyJQXEUCAurva/uKUL
vSQbrSz8LyJzSHZhhMlh3EispqOQyUrTUJ/Mxq6sZNHBUQE95zhw3fCf/NJTINOecpwUh82tfzTu
8G1mcCsy7TJmj12C/DvTj9xN3XOvyLILJkx1lHeyqNyXSR3OzAKZQmAZsVZZajjVt9kzgXG5EyiL
SRgoXhvWye4mnIn2m+WjAv4XpeFYLWBMZJZHglPFky8RyXldfOLDVbY0vcQ90u2s5CFkhIciSanu
w2pgTDniIJFOSL09AvHDteC4dLuz5UtdSO3lhnFC0J2QPM+guuuuF737NOFET9th2h41vrNtMwUW
5iURgOnkjEMiiFRyLvk/DWAWDCszHTqL0Mp0CSooJpK6EYf1Fq0jhy8WdIOPl55Ygw+uI74DQwbm
iMq5psBoLYR2pcReR6d78hyhi6LBEKxnd45gnIxyhWBzqjhs4hOof5MZiGZmNLV/RqDc8bXeSwpY
Nf+4WvPEPiHBHw8ETkToyWfNa5W4q1Oy+RdYmQdm2nMGHbY35w2svhwZ41sOU5HMZ+z8FVVd4EX1
6I08ZSXt47Iv6EsEN+vrWd6sBJftXhwqBKILf/fS4S3CCw0P3jDZlJV6HjBAc1dNPa6KgchkJdZT
Hqka/jIbVAxS6zem7l6GEaP/gCC7lRwuY2+158sk1/iuLogZZKnLa3fJxGsW/5BuyrlLN5vayYib
8ezwFoJmBkjuPXgo/AmHHSvSPUewzNvbdKxwdkrhCABj6dEL3gVaMZ0CuHsbN9+F2YE7ISOeKInK
lxaHvycTGa9skKx5faVC6rmnmw2exaOCMiANJJZ6cXr04ST5JN7ZUtkob0Hnpm3NgWAm68Lo8q2d
Qgp/PMzjYQhr55ZePmxRnG6admEUY0obv8F4uRMsBcXj0o8nnUjDkV2Ly8G861e3/YyPBt2FXpp0
lgmmxZ0QEolIXyMDZJcqxdQmH75ZFRrNf8aApBlnNmAebhw3wstlVsEJ2Q2DnG4c8nGvQgoIx9tm
A42T3QIWDFHXiwCkTrO/vFOsrtrHC+aDOkNBof4WlZBk72KhxvZPj486ENLB5ylySVniZ6k2j9OG
qM32k2FpxPpGkA1r6/9868/EgNT2qmmJJr0LFws0cdeKKtQbMYIDl1c/otwwtBltua0iXj4A3TvY
Qs6FUXxGqux5ZF2QKXd1Awv+rxNyklRBkMKKitVsWnjqOKtzWUUeL3MigxLqquUCpYhJjL2CoCiT
lrOv00mSfMtg52xF2BNi4RWApFfzlxEX33UyzkB1sQc9k3QSumo60cIMiNDP4ROoS52djBKA92ne
so/ht4hpl8qMWuJUPxXvPqe+lw1XQWcB8RbkvM9NljvDQyqvgDknmZWxgS226SK1nmH0ZXLdXAXH
cHdqWQ/4GF079DtAWQNxUDBHc2/xkng1y+Yr30rnIw3NR0JjgW8w/nJKEVKQY+nt5jkDwnLrRzKD
02ETXHoSiC/XtmTsRkrOxw7NJhgMLnrK4enQktI2Lhsam/XjWCrNub3fr9wpD2JN5q13rusA+I/g
+OXyKAL18bS4hM2bW4BsPQylaYaAHZrdY4WgWdWuHMJbPfp3OIMoWJpPd4QHhUAgiflSr7TWb3oO
oTwrzqK9DSCznO5NwQZPNw62pQS1LhuADWQMfjoTXoJsToULzulobPCec4liqcZ5+di5E8JcfKJs
Dv64/fRW/AlSh8jl1HKGn/Q/7ocHMdv1+BOzpxzKS/Ob1q8mxYYkO8y+GxjOtpNmD5xI3dnzp+Qd
o4I7tuEnkjnUF+J8X6CibXlkpPrvIDokJMbpSCOK9uu4iT541ICW0yQUKmjfLzPiOwP2m1BI6z0H
f1jjQE1P5Oe2F4kvOgKobyAhrZQtzJ2ypblWFINujlXNuVcnje2yPkEKy4VygfYp4sM71kHRT1tY
YDZJMwXxaX5ac/DMKTxZr6U780R6uHXhRP7gdaJXjLCNBPZqyCrDj2QHGC1XUbs3o2Mz0DIJ+E99
9Fxe5x+k2g3b85HvHqAZug8oSDEzxaj24iU3P5IkX+jERC4LnSsDjl2nffaeXan5rCecZqHYE2Sd
iEA+6cv6nESG2feLQHR63S2AWeQPkkcHaSLpmkEuazyXzf3jWCn6i444gGsTLVaJHzOpPaZJKI/H
vRhnrckvMjK7A+HWxI6/2oeBQYocI9xEr3SZP9wT1abBox6IcymEDdmx6w6E37mitnGNzxtuEQAm
v8lUjfxO4B0oAIsrnVkcFtOnU5U0gdy+9YAWOyB9u3XgCoBwuFbtQNMLGFJ810s6YU5IqhEKDK8y
tueD1dWmSqZFZcveXIRT8Ew8d/gk5l3f4MiZM+5h+qirYM4sLw9gUsFSnqw4vOhsI+S/VhIycjTW
hze2rdUI/UAe/EfRDUxBtLmxrF5qC7R7FRM0DPkxly4ygCaO6OhA8uzOsVBg3BM34hjRIHUye4sb
M/3kOVvFQq15DVKrsBPuLVzvOuuC0seqARt6INSbn5gJkcGCTkWGK9Qtg3yOqAq6JXDFKTZjl2Rc
MtoLAAGC7S3YJW0m/QQeaDZ113xglIC/rRe0eGDH1Sjovs6P0cvL9xff/7ZbYcZuPE2gx1tjoWd2
bs50Hz3zat4Uj39rA4El/oNuLK9FpZm6y4RoeZl8eZw7+5I9AAdk5ZmNDXP+fXncd6WV9dyD4xVF
+SifCw8OoCoksKYh6+WGuI8Dt+4kKQB3KomGE5YLBwBWPnUmZRPNoMWMWl7fTs6RfSLX56Cjfcvv
wIkxvr9FJcEx2dPpssMX8qsMeVxNBiuwrobk60qukt6HtOIBL13bP75XKwxhip9anO2X2kfHOOWy
zMSjpCCLSE7Hg6JrdfE7vrhAPALwwO+c/Bb+C7JQdSwBCxCYvc+e0qPuxqmLl/Ui7s635X2SZ1T2
N3bdOmSrowhWueerVGoO74bOFjvaZFw/bcuRxQhOMuyizE2Loa2NetqBHjUrEKmSTmFELOWbEZoJ
NZgErgxoBRU0Lr6PZOqB/3MX+yti4MG7Q38Ktw0Tupq5Ajke14SergLaRDPPQO+SeoWRmWc3gFYo
gfBtUPtw812+yVOgbXZrzo+IjRKs/iIoNIvbmL+CJ+denVt6LUX+iVVaPiesUjmHAYXc8XT7Th96
BFlMewL5vIJxq2eYys+M/AZQkfqtkX6CrFPEfKyVghI7HLaPDWYKsUQsXKeQd3h5pW/3FpromVRG
UnC7iTdp7kgNl9yThVJHUIRigWjOZqSJ2Jm7jWpWrA77kS3JzJzbi/gTWVKYu0r/2XTltA/E6dQh
qNmhnOLjtbBVSeUMCj9b87FToDtjvP4JgEkxWmgGz0WzgKFJpVWrLhhofN/UekiNWYHsbpLbURoU
7lsemdNDiYnuG2tYcONYmQVndvIL2xedxWp88LEl0GcTwaYY6WMxtKfuWNGwzMKO0hVrfTEZPeSn
m7lMZmw2YbqUNY0i7SpCTvXOUOWg2Rbu7s7yzIR866d4Fy7wj+aKGbIViBnUOdvyDKgKdMyqvcaK
ynujiS7/9a5o/hxMb2xlOAKDBlfYPd0z0KSGHA2TsF1DmjKIp78dwwstB40/Z7DXTCT+um/lL4GL
gOUMSY6hhEWwVtsV/M3ts7jgtTCh2rm5H7OVPrJO+CPyGjMOfOCLcPr7WSROYLBgI/RvqHhpScpg
4Vqtl8hDfesxPBncQV7H5u6seS6TujjgPph9R3VcP3ZlSThJCddR8qDgehzWU1xQHg+EdWv1EiHg
xE3nZiDH62xqpyhkyBocRJlq/6S6227NRhhRwiBZ7XB6wBHP4jvRJuQSE1sHBxaLfEmSSZphpluO
5NPQoAwMo52RG7U0Uga/kQ6is7WC0hmAG6AhW8i1qjl3wy9LGIOJcbTq3yLKm8a2Mq17rPYARiBB
VXDWYRgl3w+g3Si6uK8ghaOr09nYesknxPYLBsZlVlwAlEFkzR/2LZqTJAt8kQppclj6dNr0vVme
MbRh9JBpIRMfdF6UMUN7I6wPVe5r71kq6vXIN/mwq3fBYA4mfMk8jsEDb876Wb0N4Kmj/6w1HcOq
1gTz8dxuwZnXwlZfi2YpnHpybQxhvaOG/jxmIfkSFI1mvIdaPxQrg5Yw4pJEEDEj5Na9iQgZTc3h
P7TQwmobL9ytIVBXFYqMrwEbYw83Hhm8XpqOamsH4eZ/eiAOGd2+/wQH2fP7NhbxeXunNuprxNwI
y0KU68BLxzfDeDlQSfVKeBIPSfGiL167rVg43vRvZQ6Wr8GHp0YvZoDA9ivyLhHGl20dIIKS6DNO
Ykxz0wJmf4M7GghjPwERC1vwdTFBvLQuCMW9oz71N8iXJ0ZJl74svmRlU6+AYuH8E1oMEKZU+CJD
hhyUS1gLBgZ4nEIpAS1phTt1u4ZlTvb4S81L21xu1P4AW5Px41zqhlEHS7WkdZHdCKLHA8yfY2yw
ud6Yk/1uhMdY1GyzOkMZ3sjHIA594k9TenGXqjnp/otrzxceND+BJy6u0JtXKyDWU1NEUsNhKzZs
y+8MSV3qH0ncIMLOx1beHweAPx1RtjnJApgy7cvNXqY5prsQkGqaoCaaXw+SJg4MxNYGUz/x45zy
UaPIxvMdisYY6GnLnYlRnHaZswIZm91GbJ/46BL0qMTNXWtRuEuWVbtXmpUr1DmKB1ZDKer8OfjJ
weSqV0MS1Tf+90IHW8EEmQsY/vtzwifyOToMZQWWdX+a1S+NUqnmGy832nax9ofvN2zHb/f/fFcK
l1qTC2MC7DNldM0fHU3eS6Kr6XF8rO1Sr3R6YU/geOTVlmXEHgOAGW9zSFiyKXSLEb8JPa/x8G/1
z6gd0C+EPiSaPLc9N4ALMZcAtm0aviRwTTR24V2HAVpNPG/CnlKWoPsSn0TwCdA0tXMq8rOMfikl
lWKjKIQOJt9c9V1RNe/o35m+9HWM6q23OqIOfRizZclzV0qtt59+By+TaaU0NLDQ7C0o0a+yxczl
jgi3Al/ctEwzfj7K6gBhf/Ss9wYFRYEIndWSCTrSZAcoUsX6IjpyOLp4OrwgB4V4jEe68SSXXLPK
fz8kIZVpd1o34G/Je7TJQFFpGZeR4M3xqngb8baYTU58qT5X5rlFiMtvqFGuC0KwohMn04pqqsIe
eL4Hhg3IZoVzG52qKDoWb6uNN/ame4utyeTZXv/PPs9Y2Un04/82tTaXp60DKlXjXFmUOeH2AVVa
atN2X14k+gkvfxzzNotg9nYC6OZVpcv2JdD5ia0i+uO4iq8Sf5Ss1R3+bB6HthLltH1vf69bmBBB
PmTGkVRusbZBrl4EujlMw6dHFmmADbRI5ReotpfQ62cZI4s10+LtsZY2iPpxzz7PNVPTe+Gaks3r
iwub8dIv968xe4FOV7N/MidOc5V9w5QtI/aH8/ZiqnjPcOkSwMyJ3hEazx8CB7WzQbWovzX8y7Wi
m8Fnt3A60GokKUlAx5j8fsTqgkGXCmMnMRSFnwzo7mErvgrLqEU7xvk7eLm9Y/KWVYm1ef/IFWaT
XU9wkT3NnC5i9+4HJxfx5/EuP02QtngY55wTFpsVJEQDb5cQ9zFrtvXU7rQ6fPN4MY5K/6m0CfNY
WlP/vxTr8fXBnMWO2Qhz8oz994l8UsvAd6d2+ohH4PZGh0RHxsGiMII03uplqF7bXjE16tZT6Q6n
MLJIhwonrs86ipX5PbG1XwvNOBbhSeO8CScfGO1PLvV5HhZlPKKBM2+XJcMh+cRHEpvQo1a2YTRi
ZnPoVw6WDT0evoYjRB2osrl1s0QbJID/1mehUzgga5EZZ/9b43YNmySMLRT/tzh47PXgHiXMGQIZ
87VoRcDkG1sxqZeFXV0XwpqBV6EwwXSAgZ0c3tfeFRSkO0oSHabcgHG09cNgjMTQbMMGQzTxWZ2f
nbpb8RFrLyOsiVpyZ8f1H/bvo2I8XAc/4f8mo8vdwxWs0nl9X8to7zWb/vkZmgd8f5mGiSbMcQEE
jMdaqM+02/FUmajKM8zs7Mm7UXQFFDeylVZGOFmBXHt01RWOnQzjFDS2CiYGvPgrEstwfYj37QE/
t3rhu6vT+pTmNmV6O2eTz9Whq0UTvF5FkpIGPgOzt3wUI5nkMLlNhs02VRZCXMbDxOU4Bvd/3Pwe
naL2FJnZLcisgmebdhW1PP3nZFLWcEVhSBRBXFLm/OVs4nTh/AyyHS7mcWOUgTaTDI01SFnGBksN
f5n0lBA/uLQnlvLxFXDpiuTW5cF4C2FR4VqR01R0W33IVFee33q68MlVlvwfGh6pPQVQPz4/7jOV
T/Sc65JhjrbTVPzEgt2jv+xmZXQnbjh4/vD01/NNDHQLyeqjmex1YGxDEk+9OGYYiUf+wdZJlkYa
j5qImKw3GHVANVIdhegeSGzvmXrltDUC5mLH5TZhUZ5l2rJIHbfzNXOuOtxqGabmjsr9Dr+DWxd+
JqlxQUD155xAygiqY40iXs6ljgt8Lvc+p6rc8xeFg3rdfP75LAfNCJ1KV8YUSB7g7TbfZwoD/UFC
cH6A8ZQaI9w/jfPvhejD6h6E7yOFDRKOPQMgRmdrQoKwpQvKgg2izDPPPdKXNIgd/GpyRXoYRxCn
jbNpu86TAjMk7NIR9gY5tsyLsGlUv9Ht5Y/ytv1CYA6Rq77XLD6fWlZmuawiVV5YPC2IJefca1Tm
3/RIj63/3fkyPE6kNLlaqq6E1Up5dk/RI71I9isP65Rlocus4iGHw5HjLSJqK/9T9LPvhHq1vPf/
zsZo7GCa0WZiYepM1TzSXzrxqe/jdYhEOH5u5nFw1XO1k/q8mgfGy2GGF9AtoNZoizoxNBbotJpF
kKRFtZ+UxOPvVGV02+kMnL8+q6SGJlu7gm0+iZtRsLvrzBUUoBNSxItFBloYUuu+v3ila/v/y7mN
5x4jIQS8KF0u8O0DVonlckl2Irpgg3EJWbQEVh0MnScjvvpAabcKaP5Nh7szGmF/K/K8hhTMIrlt
FTDQjOiAjSaX9zGO3g94MZoIgwNe9ZBIALpF4LC9ttnBFgQzFgwd9r24WUSEoPXY/zkpw+3G26Jg
/THCVeTfirg0ZzpBMn43uA0FA65AHnxNIB70H5P4mNZQ6DPRvP/Lkj9/QfrCix6rD9CAteR7YMtd
zWfOqtQ0mSr7hZe20nRr9OEZaPPBe7TeaQNBs2zSA3cosx6Xu8lfegRQmeVQxMwqUTEbs6+GJF6J
0Dc3+ZFLFM7va5izr63fTuKlCxslgGTY9BTs3CIrm2htP07IbKLX1LaQlIgPNaucmaENaytEdco3
Uu0casope21Bg7uNQ+BTd5KtTXbJdGqJl2W2ZTDuUV8z5ytmJzfccf4ZBrUxnT3Icdgo1zmfhFyV
0kUc+CYt2aty79kewhIXFAjMZin4QSEIAGiFm9yVgiZKSZqOXr6Gj66Q9reppOQQ8BoJOQKDA0Ha
mj1fpAgDmHVe1Y2pUM/3+zGoHZ/VIW6AIMWVNx67x6Xs0CKhztxyoRepT89YjyNl9TC9pG/bPPKT
CFAX9Ht4egeUo4slg6gb13GZOgSi5uVdSsKPzueT9XnVFHEjRWtYBBmlBpoIM1OXhYrJTWMeGGyd
G6MMSpDmTpV+VSFzSVK63K5UzCRnobiVavYLw9GrCQkuqokO/8JV03XRLbrZ+l2hRGgHADSKYb0c
TTY1lJcB9k35QI8ptMBPOe1utry7d+Kr8RpJ4XucSY3atNPb3eYydjs1D3N5qpJpkeQNRsw8TZCO
5OiE/hjuwKGYN8cTabU6RWX2Yaf42fvQjjFtxAklGpJc8gQVeUJpyOjBl3XSuTqpKM2fXGvahP1U
ii/TG3/6IaJ3DTLHCVUfuCuV+msplbcTE2X7W9ogFfwKqAXMnJoUZwy4qKmomczd2wqnH7+yoWFL
wiJhF8wtLYMfw8z4++eCqtT8IUpLQBJJzWD1DfsLjTFcGbb0QIyTmuSiKROGk6w+UYHqlQJfb7E4
eZ5FoMdk8ApjDyOz1ecrzJ+/s8gLyuVEq0tLs0OlrV6dutEhobrg+5kRihla7LdOISl5uK7Owda5
Ru/SsMUwH9E0uE2sCsPSo7l2ON1IEAJ0zfVO0OY+fSf0KQTB2J3z4PE/c6vRrlvzPn4VTsrtjq5Q
QQVmPaSZx5e1Ty3anVOPawLerGRH4gGCi4M+NzKTnOCDHUd/mEo2GSf00lwFreF/JPRiV2/55WnE
8U7yLHhO10r9g/ZtLj8Z5Z3G8hYN2dXY38HRpraCJCrTqSqDG7v0MF8U4IunnJVD9RNe8WwFiKL9
hdp/4Tq4M1uihblS35QCyPf4kCGDq/poyqh1KTQPoucZDxCe+WQXcSqCOCvYRvkshTgy/QPj7wAG
AI60n4zp/QgqXLBsrIqaDW0J+iaXN4RXXagF6nwRtgR6hXiCzTOPncVDjnF9HID9IZIufNlEmbth
U1Y4NKJNMeSvX1QyV/2zYqjLwqwsqWfD0QERNLzIoU/x9udkcFlVf/9llW/blP4ja8/zof8MDuCW
jwvIr5kB3dtqzVrisrwdGyja9Mse/h/Bxxi3OiCw/BXGQmPY+XcSy/xE9aiW2t7sllEOUY61OzFi
4txPUKAXi2vFhhzkMMKG5ZicFgNUcWleXVhpc2zhVgz6LXN4EAkyXhj22ay3ZJp7CPbp8EloqAFO
sI1zTUzyCfFQ3vl9Gurbn/3gg3tDm4MAlQ8tD2GallSNBiStNWC0JeUwDDxq3es7hJAP+m4wfxg+
MGFRsbSREHr8u8ls7b5tdA83fW+K2Mj5pvI1oigLERW+HjLMBFPpXChGsSexUmMkdPlBuMHHhiPk
gLD0LI7a4Fp8/xPx7mH3uW3EPQ0yseJ3ctZjP7yRS8Y4RvghdbVXy5zXe+K6PRiJYQqZiR8Q39/U
FxymBM6djK16EVDR3SzODYmQ8Xps0dsOKFqhr0gsLAUapCnR7/JfJb9EY2DfuXxRqAG9PmDLUwQL
7nVO8x3qIZyQuHYrtEdKxW5Jyfjqb5OFPGswVtmVlIrRgca/+0ohQYdI5ZzaiD0a0O+8XHYwkRpH
e2VqR2Sii+f6lumCYqzxNvGmXAa5UapWACsMgk0Oh9IQHoILNEUq9oIEdCIJTqUN4H3r4I6jCkNu
uOML4WnjlqZdx0D1Qr1HeaBW9FzjRxeLQTJQ9sxXYDfXyZKQ0z4mE2Vqjj42ddpDPdKoVWXioFMl
QpUrPP3E+F2ZXHIJW1V6EPDIGGaOBzGPEtKv8bPPNsLhVmuzHkDBv4mqvLXYUPOaZWJ3WH7ZMuGk
8cjAIOMQZBb5tsBAQy4DUowUneKntwnDKtc0f6zHh+tjewaYywXn3D+aObuX4frmJMZ0Pc+0TDGs
izb8oo9wK1X8L4LKy2CUCTAEWyDMeH/b3HkTJx/SUqCJZ4m11DRmEitfRaiuY9VOr4ngT1GtkXtY
U0bsBxr9Mz7UYuEaJJiAv5LJDtZSCaFYm0/2ySbbvarIyaodWKMj8jfdjPyqA4GAi55aDZkzzWGu
2jSJYoL8JFqp88p3guLiR/wnyPpQERZouJkw0JsE/bsV+NkTvSGrBqQDwGFs9Op51+PFtgfEZhB+
P6Zowx7eKk7dfY2rLlgWabBpKPTZDkYGEn2HRjAA+YmZL+Ian5aDSb7oLa4ff9/TPG8OrZ4Ca9mw
HMMB2wKyzIEptLi4Qmr7Nvw+XNkTVjtBalmnPHljHk5lysQLOl1YAbFFheQQR3fjsWPwZK89DwlS
hncivARx8hwqC/+e3Z8+uE5sT5EmIK6den0ysRmPJ/qbvfoFBM+39K+Ay5sKKjNGn6B7cDQsmjXs
nBs1Irl+76+1BLB1135k3z/RbcmbUKrGwDeETpLgHjaqVpl3IHtMgSMxqO1Kc/NtqvF1XidOiX73
MbVnKcjTd1tjs/8dTcvpd6/6xPFkOo6V8kDcWuM2O4dwI0u7Q7HW3Uv4P47SBU2/xBDpp6mk3/JU
IRpEt0dXU25aH0g6yWmqf3abyQfNyvRn2ikqXLrSROy2AoyP5roBZ0Ty3zA0eYhBYYE5A169gp8B
29UDuBsSkN7dKYrxhpqN2JOu74tfMv7u0A6nFf9SOpZi6kW/aqj0+3gzG6nxLawxWdEf0Nwcy8LT
+ubj1b/y9L8m/bQLX503BSM1AVEo0iqKqcGEFyqCneHR7421GoYWAVd7pxcdfSCyuqvzlmYfn+eE
fq9eYb5kxMeNYewsIcyrVD/dl6dqsU3Kb5pJwQVCmGKLx5YGw+k1UchZxLz1gYagzN2+u2kurTbE
JGe/BefBEgYjrgLyPIZBbYKSgMinYVTkE/4ZYZJUWXW1iw5LnslrNDqxtXgAN7TyDFA4L+2ZG/Gr
bp1AjgZEz+yyLZCQFtIod3QgHzbG0QJKUwPIDXVIYz4zA16naiCcZ3Cpx+IlT8KUUHqwd7EV4d4a
LGMzx5GBjUzKrFYBKvWMwmfmWnZvlt3U2detu8Nw2exIAumoN40CdC6n8qyFvzsYQ/xAtvV+8yDy
NdHF3uTJhuuJt1mAE1MSp/GNtRHR8PaBBbPlPAwlbsW3yUeCwQFJvAOig57B0qwzEBHNx3r3vlo1
hvtZ+mGyJSfL4fJNNIcYc1vdVuw6oZY94z2SVT0KQA3RDnSjRy/1nL35e7ZZnFIooBY5QFfmYNET
2ML2qCxQFJiVQTMUGQ717v8MreoSq9cYnN9y+YALzWMCkqF0bh64Tk5uShEnn0OpzFyIsoyDB4hn
6Nif/+gpucQ2MVOnD0KsWtm7cLHDqUgMEAhqFNnJ3D933Uzisbmkm0VUEWdAI/7KC3g/I03Fx24O
KBClL2CWG4vtQ/yoceX2vP/TSvViS5LCtzPtY9Z4bh5SrqKaQs5gyDEvsll7NB0Sgt2ueTI+XFQc
HYp0LngR4HdT0+0w/sMB0fJULznzlqaUYjWQfXYM8cHjW+wjWJ6KEd3wJO9EAsROw2WPvIkFwlDf
v4wJnEmtVJKheYcHq/yDndDiLZdkkiKqCyA25raf7sDLTqLfk1t/LTRbOBRq2pi2NvSK4DTzD+LS
rLwmoU5gfME+925GzxxB6TScvV04ad3bVc3rd0KkuQdCq3Ndpg2FWs0cFJ0pXtRq7+6Z4zk6qRx+
hJzMC+19uAhzSnneqprqKM5TJhFPxhFa0fHLnbqzzHXq7XBOvKL2jQFJ03TkTYBhs0EE2cu7a7I9
2oixN7RWZjP6UvlDt17NavdGMicGu8tXsUyYd4g3eZn8NusbII9ujz8O3YOUfpxJMSYV8q3C+lvv
t5MuavBAUNwb85Avn78lFQIDv8npsVCEEPtwu4ZaSnX63Zf1eis7v3LOPOh52+xUhT1BDhnQl8wf
IPL25QMMUxvL5+tUDvkaVGxMWD1Yp5B0VETaaZIsrJ9PWrK/NIfrB4heI4Glte2chgEisX84ialy
YBcFD/qedZhcX3FtEXHgzJzcB9NxW7PYgoSigDeofNieuzTbzBuCLZYE761uh45ewm3raPlxj2l+
FQlL53Vd50/hUxbxI/skgMOqm3BZyYIs+obj55DwZSI1rTBBlqfCc3Show8b08iXJSMQNR9MOBld
mSqAeNBl44i+b/LBbSJpig2DCAg7TpPkwNhhn6Hsy/2rJK7TGQeatEgyCHdfVUq0pH7wZ3xsmnsU
/NsXGO0a0TjnxUIf+4fD+kGplhcXTlGh3DofeQzR6isM4R/9SBqpPefX4oJkqfKAsm4/Pr8JdWp7
Du2sH2LMwFt0GZCXI83P8hvVnrLGRrWM/xD8ezgWT0c0vmPlsH0BfIjLl4KQs8KjV9+0PRtYkI2R
kNtk5N0vPWvsq4y5wKWgAn3t2/z5YNXmO0fuSo/Uc72kX10yCOkgywiomkifdfY685cmnhfNUM4M
pZOcgywyThz0ALm9qnm1XALFJaIMlUiBFs36PK7rbW5xE1tH/QZ37fgM/7n6NBEYll9B/unr3z2V
Lf01D0dfNpSkakihvlWlUWFQOrUHI/62c5OAPbruL5+jDKFzpAL0AXtPO8IC41lNYb5vzscoYVsk
ahalPLWtG34m9EidWhptnOUxFpvJd/osCqIBLUj0ljwCNPS9t0b64xBIYUU9I+wfU/ydrUsgGcaK
ex6S2975cNXf2DHoor4zEuPQu9ZVKjIDrKI9dMa0SqdRtOae668qBnpxm+bts6seBLqkzg3EvPpW
qXY545BWRE2dnZQhZdzlVHlZKKt4ltRhYu2ukDWihF0Yg0+MJdPnCtYhrORKLfrJXJGASxGp+q4D
F81dZTwS7gIBSQiRjsMBI6rnwC1Bw3R5nUpoaKHJZx/g6UaxgWjQnvB4zKD3ExnrEcCuHlRCQnRk
SFuPGbcHfQMM9lferuys9RmIzohgej+xOi2kypPYDEoWNgkLEwE7mMgxQY+rmdNwgLvpe5c62b8O
JmMY9jY4vJfs2Wmxo2Uc1u5azdukRdCpqL5woq9115xAg7Jr0tfHEWnYHXpnR55/Abr8i6rFUpVE
gmI/57hy++7OfAxWmu191lx5GvxcxWcOM7AbGxDDddD1lEdyrOXWmGQHlH+llqfrBnSxO99BdF5C
SdchQlzPW/PHGdrze1mJ7SSfhkT3DoRsJyF938MFMqcimp+WAEXcTvMRRXaPRbHkm0MaAUMazrox
Z0TuK6bQatobNeHCZ75QaHd+FGv9K2CJ0WLZz+R0ecKNUbl4hcBBU/7Yq5PPBUFUVP1xh7qt6ttL
pO3Kf3kV00rlLWlZESBtY0sjbwI88KY2qTFjxXZbsCw2E7QX+MV5oIVRZ5Zt3MH3vTPRb1iXP82f
6AzmbIjHDQKOOfPEwlCCxujsx4Q2zodN43wIVx5ZsiHNXNOj+EVw1KQX8mL/p7i9r8p+fBNM1oCe
k/TaSjeVMAxhXEvpy6cSMUKkAwZs3I2LqNjxnaU5ArR1qCR7nKg2P7ynv5DzrhobL9kMQeRyd0p0
V3fEcgYTU9B6hoq1S+O+nU61IeNmoOJFlr7/idgyX2T7hJuXm6cif6fUL2SgXu+5LG+SL6Ps0gBh
u+woRSKTDXJ62U3q4qHnJ1tgfwgKmBUz95IGLijCIWXrlW462KRJYTsM9r4Z+LH1bIXb41Cb6Xsg
O7lMU4y8MfPqRio8jGayrHTLhm7wl0MtliUxXNRd2ujN/dwpEQXIKd51Vc4FcxhpKbF6zpGrRG9T
qN8ByAwtQzXKV8y4/5WEUTV/KyQDFnlaX5zx/ULwYuUvqYGw+9vsHZGin9ltfTXl3Qzb3dWAR7Bg
kJ1STP6BZ1hDmlVD4g6USz9q1LZ66inYRiAT8ChkEuaTAmE29b4Z1VcqcTjDbDXhjebuph77AsDL
uAtsouTHxmPq5pdBv6ksu6JgX95txFgeAM/bt0SU3EpAs6qJZM/RMZbtb9RCT3pNkcDL5V4ZV/Th
xLkEWZji8yMYBBzXs8Fg7gGZDG9UQD0jvnKYttdvUNZ32kGmDu8xM5ocwagJjxOzDEXtDH41MfC5
CHbdF8qJFBbkWydLCfE4lfelwa+LfdFW+Jq2fvf8ePxACI+lp6voL+XkOTC0fr30izGXRKOS8nqp
VzAqUIxKM0T1DuOeQUO6uqu4k2NQUKmTvEsd+myo31lL6CSNgS8XlLseEq7uw+ffp+9H3xS0CY0G
rj32pgbYF+5mO4auqMekU/0UPVGOSo5lxn+F9jrKn05zJNyZ2i/aMdbCFJg6+1euGADrfS9k7au9
oeDZtJGPilWb2iU5I+Gmde9FAd/CWcXQDV9IT5TXKDiU5n0ytGE9bWP7DOF7cicV7f0zjfIHReQc
JHvWAliqDzn/b2cqnZZHCqO1AoRIFHrL0BmYVBSYHIz/TlUNPUtttJ+OlYPph/E+Z1q69SFPDgvX
QyQhiCtGNBSMZy46TMz153fM60Zv2Crx+yReqB7oy/sTy21UC2vTDx+X9VPUx5qqjVfxptQROZ+U
JpGEl4aNHoOMU7LnoTxT0D3z7HV+XuFHr92NhcYAy12782TJRI7H+avLDodqnjEC1zDLdCxGgJ4p
nX+PaD45EkmArpf+1Pvbsqgqd+LFvO4tjxQEFvH6EUjF3WtpjMp0mp3zMakTvRcq7b+jbztlxsN8
4Se3xYgr5A+RMJL0adjXCH3uRlFCBsyC7maw9lbUoQNcOz5HCNoDwjxTmFHtNdWGRDse2dSeGpnf
i+h0P4it5JgAwMrDEzQPuJrxQIHso3sLZz/bELIUseC232fhh+2dL1+MhR55bunpF8jKvW6XvG8a
XAtLm6spX/NklGPQBbAmVfWHLv0C4SYEpCQ7FqypmM1HC/ZiQoG7DuA0gRVf2mjoK9UJ/G8cIiNb
Ozpt4g+HXN3ciG+MBlP4DctRG7lOWSj7EQY9p9aqrEcOpMzreioKOyJ7XEHv2hgRezJnsJyQLJdh
19p0gPUX4+klCFojsw5rAkkvwh4Akk2scywf7ygqnaUjfJSmDxsaKD4LHwsLxdzbNQ4ubIBYcdCb
sdrosBCktOBAgmIMFvaxpgZk4hpzMxCun+mLXr/SHUAPjM/x22Aaa2iet8uV+OKwfAHZC6ePeAB/
RrCPrDXDwZeXUTDl2ECuDxbmVU14kXWNuj8AnJZylyaQtznynwFcuuXUQLY5z3NmC0UTkzcShD4p
2pf9XApfYMWKDMy8NziZo3uxcSgo4S83MgcfjewW7wjuVkvktjYIfoQcufuoHnt9sP5mamohH02u
bjKX+DHgDde1OUj0uPlzDDoGR6dycYZi2zUX/ZvGmTHbJjGnBlB51wMh5GTnwAN1rGGy5G6jhU0C
zBNUB1NRsd7gPABTgIknlGpORXYa+PI5TsWrDHdCkU6QSYxXZb1NR2Eh3bKcl5/8rdTIt9sFuJNC
crqcdaUXBHT5v96xZKYKWAQ9K9a4PhaHtHgY1SLbnxfgDjxDFk9ihXu4j50B42T03AQxQeTZxEI6
QjTC1II1rWZrCym19kSEXVGdMGp32prfN18V1ho6FbVKtTAmZ2mbQzGAgA9kx0djmpGaSFm5pqT2
8QoY9CzJltSj63Nn76Y6Dv6WtMn/XXP4FpJnNpCTG5aFTR8MAWbMHsvQQwpC7ID5crpT9F+OD0lX
c6y/BVdbV4SFupXEbjs3j6kWlkwNEfUjSCakFIzgLJdVBKRRZtpUAoraPv3qjdfxopDuJZInBl1+
1cbX8smxlRXXHyu8w+MpmT8SYFibI34OhGQF+ZdDFX7wOr/DACtnOQ4NwtHSYcmlL83JxOT/Q+S6
c9hrFWp7dgRKgUvNFljSZtWy4qNXdZjKOhbhJ7ucZP3KJ+WpeEfzKWq9cpSrLZcrqOqGNGUZiKih
nllVC2j6VKP4EshjhRXn5/pIZRSPbF8nqvV32ecZ9RzK7OvqAH5oFKzPsQrGUa3CCKZ6QsEEZ3qe
4OE77AJs7WMdk8qX03fsVTbDAERIf4KrihEtVZ2HIO5x2/J9GW5VFu6EN9OyM8dyqydXbUikLQM9
XzQON+PmzWrXxr1zsgA5YKYerbac8YvOQbGhabaqWr0GE6nfi3OQhpomdbj6DUoKTGkgxs6pl+RB
wSKz3FuQxGrozNbSbqyFm5xx1Sf6S9HNkNKIAnNOi4cexqyL53RfYEpt5HAtu6LoXiNtNWyXFhFc
D2oq2wbNj4+H1JW0imz+wjhJVKymr+6VI6J+/fEBiHaTMScGWglYV21cG49+lluM8M9IUHiDaYL3
c/WY35oFEh6bPSZZOce5tMA/wmIObyRfvxysNmcZqddRiXMDTVYuMyiyGXEHp65TvTBkI9ilfi92
AyLzDBmaF9dg2JdKnH2M/Tz/4EjZV1VyeovF3evUPkH4GWOULB2nhz2OjxihxTQ5hmNCgq6XdwKQ
ByNku98IRI9HtPnoAUs/I+PeKIqEnAPczbBEogiTXuVK5ixGjNfX32KhAfzHq0k16MW2zOUSx265
IMQD1kZdrbaiwRV9oQM7CIb9+ChxE+jQRDc6HU9Cj4TRkaRlpcUwGP9iNUvVVt0lXTZSKegwrrrr
JxFHiLlItr/+uvzLSSM7NAG3z+o5fkg1LQOXPf39xOHcS8JlRGQ7rGJKN99h4/CPOCmq69BxXHNn
9lmJt6g3lEL+10uK7399z3N9XLUoUsVF5fdJ7HF77VU8PHZ92Knq4rn1bOS97NSBEDttXycsglkK
N0GNJsf3YjFa2yjygEoPShVrA0Y1sLEkOVNskFsF1aX5ND5FQ5iiQMIP0irLENaUs7BnHmvqhe1a
xZVuRC/qTSna1CyApEbLHEHTuAfNSXgg+kbuRqWeaSf+aq7NPlgUPGkuA11+3VsksCT8urFK61M0
EVQgwE/3CziBSiZnok5MJxTB2H9n/5GXmYq2zQXdItbEp9z0AhzrjHT/z8avLfGpSJYFG4S3Ub3F
btrUWoK1dp67SS1sQMI/6uaou4SCY9GYoe5hoAwbFmEooZ0sGhYpaFAh1sF+brmOJsw2c4v402TF
IQNdTZ9ouGIki9CQ+AhQTa8lrT9LcSJuY8NVo4fz6GnLqK29ycBgNUP31ZQF1b7Tpy8Xkb8wviX5
3bjWYpZhr8Suw/uFOfu4dKFjJfUYbFyNJ2R/h4l6UY2BZowYJBP85nv026WrmF3SntU9f03B6/Y9
GR2EwMfptNHibOxtcdg+g++xN2gYwgUELupLbcBBrGFi/d0JJQD5+LTxXdsg0oCpf8gliiQh+eX7
HoN2mAxO8qtYh/xbidFqymPC5JHlcZj9FVoeEWC93s6gtghRbypaozeFqQcLuFObWu3eEKHqMK+W
NMrwC1+qauJtSjMAwO7fnb10QntM3Gqf6bL/A3uDSoujTpm6vfj60EQ+lgOvWYmp24f6EeF4VY5E
mY7EYeU7WPWHAy9dghGz8Xl5LIYIlDKDmu1++75VsoOn7IjHScc3pvNf9jqbdjnQkoHzvJyXu3mO
dgrXLrATsK19SSjJCKAWsGwBQiBvFl9sxEp1xm00u1a4JzYwaF+6iELuC9gcKyZfl/vtaWjbqRuY
MP+0sppdWRIUxHaEq9DBtPSlyVXnCbyzP1ZoluNqEVjK9+8I5ZfUOK4oXD/JHY04apMvlF+jAFd/
XnpVr4zUNJI0r7EgO45SuiZEvptAHF2TYcD/E2lwhRhCzGqJmgNTE3NliPpZv0pESTYk1Obb5aFq
mNKGumm2TKpMhGwPbNDFx9mS/aWPRvBe3yDqG0kPW2dz9mbqGklCoYgAUrYnC6kY1meFlvg/9024
JZzfeXQqclsyaIDSE0e7kQFh4PeXXlHeC0KHvsgXWrwk3d16mayNNhsp9sK/ZmQh086H02HPELl+
lL13bRuuUKMntiRqwbN6ILSsSdNtPSkTdxC/kketwmJRPSS5kppzlPoifmcaCaKjbv4Q4zrEF7a1
CmugF9l90Y/flD/jtN2rrceRpQf6d+rg/t5vQn7vO2D2ZVqLZsJEPgOP91WUpEQPflc3165ui7/m
chMASU8dQi1xMAU6QWRtQy8MoR6UUTruaR5hMrR6KJyu6wwPMoAY25vT5vDBq6BeDxolPO08aR8o
jqoMguRgBPHxWh6R55JmMBKTNqkHA/6GkSZpzu9cvMpcNjbbQQ1X8EyjJR6IUmddfZAXqOLOca7X
DQrlnNSGVVsF7MAhfDsOFJDVeJ5IIWmQjknEWLng/M3L+L5NnRkFzi+dyA0bARpIeBYlYl3VZ8R9
ulvWFihbYvFw52N0hFtRhSvanEVpXQ9bnkWUSf9raZb7+3sXr/+itsz4ikSYdj+NtAiIvCD0t7FR
QTNVu8ScRtLVtHrV7DQVvRrw+JMGvwXIUwllDkB6KloQ21npGTEdPZu3SWjtfznDEZ0BBCUFi6uE
XTWcB6hM/6BEMbz0hilPpNatyntcV1+4LQikTQCs09XqJ5+xR0kKBOwud9nyz/pFw2J6ChuxCqSc
bl/smK3sJuxV1oHEVPNjDAXQM7AD1c1SASREcLocyc8vqeORhxRRKZG0BSm3TPZpanzTTX+4BrHU
T1yTffod57jNjXN8COTwngX/8odN7fn1GhZzeRk7iRCo4kFrLHsvC12CihQuSje64bNOCi0wthDu
b+qY39htowCiI0l0teBKrqOc7zYqmZWlLdkBHy+u6ob1KUcVQR57V7DGKMnvds3/xqvD+7ewFu3B
hxhs/MoGcoOnFAAzBSaPWBgcim0KXpG/Wa/K8vPecgInDYMHU4ME4rXS52M+H1DnSkhZ+XGrxV76
hR36B72rIUnymVOaeT0au6YwEMZuEYl3JR35epBdX0of6jTZXC8mwAYtK8nSIxUJZiZtSVWpXknZ
yVxoLI9ScVPe6C78aXFIIFJvNOlCKKHKdu0z/8L18EpaFHQhmA0pArueV8mlQz0OK27ia4XP2SrS
RyvvaULk3SmfNVKbJKa5BtOwkJO5AHVJ2ereMAz9I8KKes81TJQOp/Y0gbSOoPgT2d2GEanKYke4
gXN+DFDrVAAVs0zsMGmQM4PIT8pP74Gh4GVZPW+yB186qFVDZjhT42CI7o68YzASM3QV1vunbFVa
saekuJlVDspJlhGAY2ybVsHNIEXNJqX4nBM1giicOsTlS6wGfVbDKMl71VmiHsLXftAPQ4ywOK5r
seHw3khoBRT6FWr42i14Q+gVbhxdTFmqslvP9wntCLfkzzTZhc5u97UJW8UbmXrpOsLvonU04ChO
8eH2QjfbrOhzd1yAa4iGxaqHql0kjIidAUKCrnDmyC/W49BWZYtMwqxX9fVsgBtIXnyFvCyI6T0h
1qfbnLGaGyWZUZccKm8lWeGcNbifSLVgnlfaCBbHOQKpGCkQicfKJ12ZS4XnF2IiXi2Wli3tl0n7
GatK0NCFsH5pP67j4n+pU7dhcDTQ1juNnr1vUKHgL/SsNfAuZyoNXqKHSs4QM7IY97qMDVMWmn8g
oIMSmLFBplpeZElvq5iU4mlM23Z63mAGxYhIMp297A0fFLoFNV/NXqOeTK17rpfhx0n4SPBUa6d6
AJz4z1gXWVqeKtXi7v4/8yVVYgkHrH2ldYEqYHr4X4c2/RexZ/6DBSs+y+HURr3607g23+dl6Vjp
fadO6x2d/JHP8QAa9L2jDQtE+DNViIU8bzdd5ME+kbn+o5p9Cdj/sItbakSAjydtnCSeXuEBC5/4
4EQPC/GcV8O9eCQ5dv4ZkUmWeUiXzpBnV8OYSPGiyaEehqwdXXqjxKRL6Dit+lFo93qzZvftLu1S
8azWBsVsvisyKJF52izRYfnAppNqPQHKcM/H7YStRMfCtiMxHbk8uaNO8NgH1eFMhBUHP6uf/+T4
mIxpfpZU9pDGEpvSrUqbnxUTEVlMr3YJ8ghzEDRaJrM5IHA6DcYv6fDuXwH+nxsomVtHs7IWKNtV
K83jSeNvvR2CyF16WS81b12WbfTSIPizwHdCa7e152UTf83eMBS3Zeao56jBZH/K/Uk9bkMtO43H
eBG4IKzJkeuQVs7+/uclXeltmx1G7wJ2kJu0FOhU7G1QZ/zLOWBxdikMNBfEs2QITIK5gLU+Hoab
w2KnseMVhJWX1oIpYZIIOtKBsJxONHB0zEWaLow8DWxfMLrTbGijsHSrM8xKAoSd7sX8h7c5HL/A
6gHYxBWq0Nj/0Vr+qiGVaqphxUh5VLKJuT+Oo6f2P+LzTUtUOlqQ66myex2yCrXtZcmmBNUSGkvo
KsLur1P/N/KS5Vt9pu4pjWoClELZF6/GMiioJBIuMQUwPKsLJorP7ryKC6hNqFMr/iy/08FKQgvx
Hgj1u1nHDKRd+oFmuzOWcydM2SXtQSrXmvAxI10i+/Oa+bUUzmIqK0Giqo+VO1Zk+4+8s7sD4E05
Q69hRPEXKG1gHzCzi2VjfpK9MkXR0mvqNY3cG6ye0OPZRZrcsbHnOi0edPQU+kOuJUxdC+ocnEVN
hFL5TwYCm345mIEcIW9zaVoeJROMrG19TTeQhWo+ycnNKK2nhWSf40w5dUQZucxAsnc8pnpW0qQA
OW5M8bfwDlKbVoYAqsrcCETWmHo7MhuGV4moGqLaB8yrSloB1gIH19dsB9xEPW/EDnzCQR+UbiWH
QlOuJ4atTixnp1+i8W66pcNKh3r5PCOpHEna3y6dj9lOJjE0zGmsEUMEpr4ucn15d9jeJBauRm99
bCGorzNoakH0gCPQSlOHCGDf2GulYZDLs8ViCqlX8v6yXQRAHfXhZv7dRWEAE7XdmL/I5svkXkHs
yvr8frEvsIBb7zoaY5pgWfVLjh6Xj4qAVg8CoZR3Iq8MX7v12n3VBQwfeOJPulJ5SBzbLR9gZE1g
/CvP2Pq4lj+62iM7rVO4Vj6aR1W0O50WuN0FaeD4RaN4BnDYDZkSSRVsAAYcijqtrDl+0/JYC3+v
PvQZX7I2LmHPc/U9CPBsoQBHgCrEXqH2pl5hSoJ5tRtyOyr4RSz0DkWCx0mBZZVOpMy4ERqk05Vm
Lq5LshD7Sx+uW+rQaTOMqsln8vABHOe+xCTr74K5mWT3JLUcDA1B4I1s2i1ME299RfD7k4gKxIAn
JkQQa8LLDpETyMo9O7Kj6j2y9FKGa9FzQnYefHtr5L7Raq9/1MxtZ2f6jfaLNhc7+x2t4m1C/hDh
JcbfL4t7rKbZSjBiLlvrWviox3+F0h20LEfBobML8cc/iQ2wncYz57TzQ0c4Bb6XSDbIjF5sakEV
aH3peOFCKSPZt6BVUbaBnDkyx7eyt5u5BREXvJp7oVMOX2g8hdLQw19B3jroJ5sU6rmmh6DtbVFD
kabaVB1DawKzy53KnLg53j0pE8f6afBoM78cNQ03oYNV7RXv2ecTLlB7xQFVNzbznP7GcK4BI3j/
PcLB/T9tXpsYOme/ap5Evk975zScoLrNfmXI4KS5GjzGBUkqEDhgWiKMU4tN2l2PdfoX/5ASRKfE
ueD4YKnXG3G6xJBTmUXh2MNbiIzDOEkidPe7ryGVDbYQXhUQbp1WgXXnFG3kFiSIzod4BAnRaQeP
q+TwLq7U0fsyPgKF7jWBlYchfcZiMTBFI74aPrruAd8GAI+oSPPouKLY08tz4DThQY3OF/aCM8PN
2wds902iM0M2BP0XzTruxlIYZby4khSeKZ335SOh71//TwLypDBbncjJ1aOg1MT/Uz85RgJ2kYCy
KBZuG7fLMAniHCORyAF62tyF1S1K6sQswOEOS8KwvTrjnkWeeQSjxxLKeF1+KFjWD7Yq3jKKqw+3
V6uAMu8BwRzg0x4tifOkIvvyLsJjfjDg7JQ+RLPUd17mx/mQdIS5QaCXimsTGlq1OF9/9fciO+Iy
A1xIb5OoAq1OsN9PkWH8qOUG6aZ70/dPOKotNg5UOkguEeaPgTO97on0TBTjqfxTLq8birw2pjVe
+psuU18hIc9RLe3kVDfFIduSrcbO/NN1E3lTzaGiO5j/eRNYWiVDi38+9TybJaHbHXdvU8qkVKi6
PAjaF2rKYbYEvgHhArBWE2SEGcSBfjPS5+6koE2QY7zl0YEEw/4vbeU1q23C3rampXVlaENxXfGQ
JhsWAxrNgB4NEhVCxPwybUubw6YaGBe9gEsbl37r1RnUPWW54/1FRSjJg6/faHSIh5yzKYKqr9ir
UKo6xCLJDHb5y0lvBS/bkhsfhVg6SiOzkdjExh0FdgvXOZsmUr1Tshw82aMPal8CSp1EkWlRYwHy
IUnThVoDGPhqjqcQ+wjOKfmOrYAkkAAII1T5w0bDYmx+1mmHi9OjAaIWs1TY5wVMQxFmRlCBpdjQ
Vf/52lBm4FJ6Cc4XEKLS353CiqABIvGtgRBySbGVJvrrjP2p0Sy0mvBsPzb1Stjv0altLcP0zZae
SrFcHRSqxBWV+Oc8ohm5I/udfuCksx+O4/9NMqfS3PsdnKlzeq2AfXpF/J/uiG7NG2BeB6VQHjZS
ps/7L7Z6T5jXZrDkxYgDsg2T3ctey3y5jPzJiMGochd6Rm9QsZ97dXw3w+i/ueHLqmrUB/TYyJUj
KctlPdEq4IVB45A9jC3F0S/1TEeIZrthT/NXaPmPpQj8si8X8T8nXnQJEshPz7YUIf2Q4D/PnVlc
CkIQOdtlZ2wThh7RhoBlbYOKCc6fTPwR1t10dX2b006dP0jRrLq0z2C4K/IMk/ArjXvFAk2PA0Y3
zLi20UCoHrXFB1t1UB4S7krmKXkFtjwjoUZ2t0yxgA/FRDDQcmU6DMJzq1HYL0DErKkC2NAR55vd
Pwd8pHnv9TYFaYleBuRHYq1w5retLXJ0gEi6CSJcDYImB8WPGJw8iOn+YX1MQSoeM70uWbS1nBYU
9u6iHnOtIXGcawe5etToWBrZOjhsALbqKptzYg95yYy8AgEDT9AkWmqIjKnfVMBWQCfq8+tYoXMU
y8NzhaBDVW3/y6C3ULcGDhV7OgXjiZ8M13c69gqDCjmfUTy+Ho1XnkH4Y8TT6kk9ZCfy7zgya40f
a2eiHjT5QbhuQYuctSh174i7e7DzSeQcWTBtqDJkF3rSl8D/AO0qRboFC4a6VfC04ctE+W7nb8GP
ha7INPc6lamFc0j17qUsgHgfeKyxRKS4Vlb1+KV/a2lbusV9gmE4y6P+Sv/imI1l2Dh+LohRG/QD
gciZe7lzt9eLFQPDRQjfmA5tRXhtP6MYVS90tZ1u/V+zwtscWNKG1RVsQQ9qjKz7K+/R9XPE92+X
GKec0FFPQwBg0XcRW80GE8NbxVW2uwTgrbf4K6WV7QSdO2LyuqTQK0fh9ZYARcleH7MydRk6Agn3
axb2TxfjyUUPk60TJttRidm0x462jNG+0RfWHKTUcX2mUexZyas2VAovbNi/Jae63oNk3GbuNu8c
BrglAyhSY99LCKs9Jv4utoqZHMqPH6qx9saQe4ycsNt3Gyc+T18f/H4an4G8dI1xI0EsrqOYADHJ
JPgXHiV6JRUPMdUfGQPzNlnlhDQT9eM2lBNISxuAU366B8+SDCZzLhd0wSiQmjEpfDO/nsRWPSET
0MigC2xaORzt6jfkkWUE+KdVxVJnsyL34orDRQ7btNylUCVA0o7ukEZJ1jhhOfDRVJjXb70sHkJm
qSdmxYR78mXKF1/UHtwgu98F6IKP58cfny9fX4T5LSEakuSE/K2yeiQZnMrqxJRnVSsPG78dElkr
amfh3ez3IuKrsdvXnH7p6uB9BKpdMPhKgnk0P1DLMnWd4nU4sN1KSzT8K6sIP1v5Pk7Qg4f8D8XY
Hf5xS0LeRlSlIVKs6brGhuVJxuuayS6WenK0z2cffxLJn9saP7e/AzsfeF/HIqHQqfi2hquX4zek
9kWh9hvKQ2bM3HZVnK3UQbxyXbZ1g/dKNZNekIaiPNBdOmFcG8vPkIskFWGu31P0da8lB4cCej14
lqW5pS7g+3Ef494l4xjYDVTqmBIy7q8fwHsnXRRp2l7/TfznBX0aY0+7y99Iu+5f4WEzh3nU51Bc
TNwJfRrM64XcCVr19vAD9B1PTTRtHYUCXkynfo2HeliDbH8Xl+AoeHc+zeqfsM3vFHk+gtH8Wpka
KOCob2a1H6vWlwMi4h4Ooi1+g9NBsZOO2OuCLaTzObqc3uPMzGN2M8KV6fIYgHCO179L+3yaW46Y
dO162F8/+2L62ceIS4D2rbdFJ3wP6wM3tLxSCeL0ekNHQWvg/MLThHpyTHCnUxaPXW1DknW8gZuF
PkDhgPFr+Hw6fV+PdJHbtKWKyPR2SYZW29ldzgh36FVk+eh0JEtRdkenyE+KtGg8UEYGXCgl0xum
Vdzal8HKoPt5PXpeIBdbWf0Vz5sMWTaGBWra0+vjrJaw9Ci29l/M4lWxVvgg/dypczZpnCXWfmAO
CbBnajo6s9HEAgugjlKAK2dHwXnJmnDFsWuBSHWcuWI4B7l82tECy58rfvi9mSCR4hUCZOigVBxo
Z2egef4K87y6/quNboDag6HSgKqJOb+MiPJFtj6p+e2kOl4xZ9DKBkO42JzUlrAvzgzqMjHGiJbh
3qoGK+g=
`protect end_protected
