`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Z6BHU2DpKswXqZYCFbHbs6a8d1sMlEerj8R5p7Q4uroQXoAm/ziSLPHXFPy+m2ZJ146Y2Lfr/BMZ
5nVerCq7Yg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bd0FLQRO1CM4cxLq8qAPSICBO5PIFgH74KkIqfoCaND+HNeiRPEc+zyr+szFQE6psJUwUQbU3aaR
wiPNvDP1qVUmWouryD9w5kFYtEcSVOesfRo1lLaaopl5xXJiF8Is8J+0U6DCv9DFWRHzurRsSGDn
6KlB8TsTP2X5WTsJL44=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OD2PLZMCm8mYqjpsOPbZ+fUR1/mwKOTLNHDzPuOokE8UCgBAEcqONYgcSOr3spaM/XVjCFYmAuv3
lGlHbmrxPz70MTtXrZB+fG3ehJ+MN/Lmh49BKKDcYLg909bHsGc3hlOC8PaX34MFYVDcuCOnprV0
2abBmLaHFysESVGtsFlwxwwC2FB6CAs7LqndGSBxptzLAK96zx0rIbEsERRyjgn6XgPL70cz8bSy
1/DXbkVXMjrRMigx3p4/rCglfBZddLABuRCXwIBIIq0FoKpYLtybYDnX0o8haXN8fbTHXszVV5NN
SbfgQJiIZY7+NmZ+9DyTQrGdJxl6ozqPLRxZ0Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PCGFe9q7siwFqzekcSvOanqLjpn6mQJgh2ORUjjCXYYSP3cd0+4zUU6fhAeIm4UxVtdXIWsKC/6T
R3e8pUrnLUbrRSa41Z4v5oHK7aYhrQePZVoIL/P6IzIxxiuLfM7fp+fdw2Gdg87hO5Gl/BDuZ/j0
PjwMYHOfnT8P85jZdwA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nW7WFpjBPnqrXIIVZi2xrjN9+OwED1jPwXqw2SJp5Ol0BVn8NTTSzt8wFMR8lCkQuuelBkSQ+EiU
x1hjDEIdL3yyBgJJi9Ulv01Z07MmJvkQ67k0VXiU+g96nXA6efVXR1PTfbU4vEcSIvUB/ctDclYY
fkS5gg7lnoiOBMq4uUgtwYkSCdUbkH7G2Rm1vviE1PSBZpOcKHxoAZY/8cNS0tmm/Pgi1IIBaku8
hRb6Pna4V3CcliCvJ13AT1gn3WDgbLO67RDFv9lQaXZ0Xw2/laf0otSPWdl9/I5X/MW+o+h4EfiW
HEBnCJjhVU0/gg0cP+xgr5ndm6dEx3XNg6F1XQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16560)
`protect data_block
TB7MW8Bm1bUm2QgDxPjKoRYk2JIohhiSCuQ1hse6vuejol39U/ElymzSw0/e/pBQk0bl328apIun
i8UrjPRGqiUJUsilj6gOGCL5IV3UmIPvyqCunh4EsBh1SdruIRvHYq1ypL8MzEA5JxsoE6MFByhf
DwKDjMddWAQOs7cZuikV+ddv8r5qv4nJ0koYqT2vE0lQwXxF5b5Dej59H2vq26zmSBFvLX/E6gEK
PpFdtPXZHI9h3k539Vlxh1POp2haNW50CJLal+dKpI6/RVII0NSxwl7xhtHmzrUSEQScicJ7699u
fEA54xnpbbR7Lm98fRILH/rpCeWbOekWs0DoWlYmpklCEaB+yp/gb+ywrwlm7W+9WCT/qkzwGxBE
zXo8LWvnoVI4nDnqPBtrdDJ1ORGhEdRuoZdoJVQNtF1y+8HZPBldElIaKDEUlCwktCwaWfa0sTo8
4AQm+V4tj6WvFrdmo7djOvoGlsItsLWlB5Z8V4nDjx6g25pGmL4qsAROskNOg0hpqYPOsK4IB1sB
Acu63XEt62DUVb+ij8NnhwfAk5ky+USdMr/v3S0nnPKaLCJHyq4TM1htPVHl7jmM5yqsbGVKaae0
uWr+U12VFOHfcxcYIL0cPyuFgN5CBMezkVNh8Eafy+h2gaLt7gZvY8wUr5LASm9d3qyBkqjATYSx
3bRqVRmjPw7DPe/WXfUGkJZPryxAjiUxKs93gFQovcvcW36JmtVpYKDtLoPps/uyew3u/LJAC7oA
76GztniZVFkkMYwCCIr0RmlMAvByNoCEKlnP0g0jHO2Ca2vywfiadEAF64BZg6xLYWNwpxfNn9Uo
3YBxpeD8PLvYF+G4OhBWUKCtBedkt5feIyx3Sr5UKVP0czIS3ErW3wd164HJiQt39SS2KleC9Vt1
JoTeHJqtK7t1o2+NGu1tDKrVvxbkIt1tycrlGaF4ZqxDe4wPausgu9lMfUasIpYcKDlBA1sbNP4j
RJ0tUVENY2jON2OGuMGI1j4/4JLLyHbItXfbT09nAMJ77gv/jC4h5Ym+yThPEPTxAwnvvA8ikF62
wUTOtrO1IaeUhYm6lqIubG/iZXVkFOEJ4UjBSCKLaucFK3cLhe3K4pGz9Q/NZyW6LkqgsIJNfykv
LuHdmQgNsNAJ0HDGlf+SYUNmWoiBG+H9DG857zSIDBa7u42hfGz3sgm2BM4PMWDOiT9l1rVq7PHa
1PokskUcZRwPkNMtwpOme4eXJ2LUs0+r3dKhTkauDfuZrR99C7MZEOaMq8V22d9AYzTjoX8hksl1
w/DqGOFLPMJ970UNgzX9R7wJNEiG/UPHoMuduBOwRp4kLDbPlhKeCfgq7z4nHwqSIyPt4xYvpu82
rD69kJ++tOcLf8YRaAWQp1rSbkFNMpFX+8l6CceFJcwjbvSpWHFFsbo7HelxahY1cwltqjKQxbk/
FBa5Th204MT+ra2RBgddstT4OlhVpAUYgB7wa0kDeC/wrIb0yKaVzmQzqp2T3rgFVncmg82AmFc/
9oXDtz8KwRitPXWqrneE7Zi7l4YvxFVvSJ1zBGL616cDgbnYsuKinXMOPYSh8uH7gA6Qmj5OrrTK
uCtJ3KZJx45f93G3djy+KT6Onuu3QptATLqtrtE/hel85N6PpW+aq+dUB1K8JmJAqB2xAmfxUDXq
B7whGbYdkhLudNWATyaj2S9FrFUeg9uOeziMYzfaTzy4G79PoWxgjVwAhjSQnlymBKZJ0Dyi7USD
sjDr14vKT2J/cYNlrBolpOmlo0vTflQJ8umFNRc8jMAULjjhVgJTXW77YwoXm2nHNVQ7hxwZC52C
6Kzqo/aAYI9wJlkUvlbKAOQpwzuX1BtiT5hN+cqEWcZ2HOI23NdIJ9a0jbFgfQvsKd5AotCKu02c
S9S8Gp6vngWgpNk6n18tzBtdegYNm94iX+4VEMLbrRqGejQkuH553WU7zJNt/m1bc8igzyq3HGHb
oX50TrWr0OLxVTtrc1qEurI7UsVayxaVem4QV5h+y/51KAY8WG1JLnus20y1W3i8/pGJmgZ0s6kp
3ZkoeTP9XEU4DKe6NAPCyJlYgizgnjlfLQJESbZWCkLjROjU7C9ATzkqqdzpTRpscn08w9pRchJx
EIBSy9zR1OQn9H/vKOCAocqS+M07ZVXOzMY/RB+WldXgSAH+ICkNilnHOL+p7py+owRF/u6LGawv
hWSK6kUAjkhjV1EoRtTx0i0xOhi/rR//ZpYVfyTCIuiHcoCFEKL2Td4A7dlAde65dHOMFQFIUdRU
jdMBIZGnN9X86SL8/Uy/oEbPoM4ZAq+Esq0p3CcHimj+z9NQpaQExbss7f22iZALDDf8rIVJuBuE
iRBzlqq7MHJ1pgVpvzA/B7lHUdLloftM42Xd8qFfZvqw46iYNfypE+yYJrOO8/+foTwOOUP0QAnr
FLVadvyWp5Xbsf9s46fUGbtz8n+KJ/s6P60NqUWr0Cf77m18hb1EWn2sUb6N64xoOH6mqXSrgx3W
YbhNMm1YkXbw77BgTb2rk8zqkykFmt3Ou5ZxHgyapcAvm9kToNvMPMe+7+pGAyTsg4pPyCilMWCn
uesUiCOumg2gwJHV/u93O4jTxZUAesjo6FSDVA3blXWyb51nwlupzYSxf7JjUZy0/PAEQblvje7y
/iFZJN1fdeBKo2NcEKEvg1oE1KfUCyIPuI1LgAdth3whnGVLfD5GKajKnaStfIVfhhlG7CvOfR5m
vsqIy9qFsHcYNFPPTHdbCRzqxzHz8ZpCLoW0lTjL1GLkdJ+36C3Y6x3bntd+umDCSZ1u2qqheKhy
P/JHPqKSWuFNzQ8Qlw3nG82PbRusHrHl5wyN22HtWZ92LBjvlaYs1r7+c/e+cuSSCDyGJTVNLc7p
VceD8cHXX2JYV29/Vz80/zXDdIGMUZ6sNK0QVEMxRpcbJg8p0pCCig4TbEgtmSnKIvFuT14lyH2C
/0kssAGP6OyBw0LQL7rkhaZfWgrDcPy4jxs9/bg6+qGAbsi580qG0XghZCayBVOUgGOW74DI+Wvn
bCwOMYyKgbLSMr+72vhvFcTMZRM754STwToDZAIZaEwCPQFO7cEqZQR57y5Oh63iz0x+VJguDE+H
EGfuIGfwR7avYfsKUH40zHHRYADnaJ8A2ymS/r+stFSl5EV6Qg2tf6kHY+KO3yqZDrRtBuLw3yM4
0GVLT96VLZdUiqM6HA7vfpRuWzbyGaGBAzn/1fZ6xrujtdO1e7ozSvO1n1ZlFieLciBs7pwb1d6W
9BSck1YkyHbmCccwX0jkAlR3Xupn6mzg0New4Ew9+Eeo1XdFUsBXy+PtSwNMgdLaTrBecNvgpHed
8U2VEeL1WcOenCkdFSL+NvGMLkLFCkw8GB45DmaXPkVPPWwFwK2W3J9n8Ee5tz47/NeTSIDklnHU
cEgKsX8sA1H9VBX1hnGYXYYbEDNc2EfbmofYC+J+O4+h50EzpEy1tBa8V6cjf/tyeUYi/y0c1Nwq
OMKjI6jWJ75LFo4tIFqDSnSI5inyapyntq9zGkf7kIplsGFoQ4IUetDwRvo4RYFoaGH7J9qZaqE3
ivJPpJ/1bsBfWOC2SP/53e+sOWeXTmIHcc8TUeHB3x93TBhfEy4y3JmxFb34GWOnZNwbFiobdytN
w3IoHFp+gFp6NKVRm+xuxqiFXDuTv73oPR35nz5kirVsUwZW063DehXXkUeT6EX36ewBK4tmy3cg
SG3Z+A4AlSIyPN82HuQ2tjdEliSnLQCSvPbv+dWSgP384qIVuplDZ4G1aSE24vLknSC90W5LIwp7
YKAlOh8q6ZWZKINmRXnIDIWm+tLX/7lcq2jAU4UjSki2gVFkcBJiuRDEOKK2F2Yw3ZuVWqifZ3FO
KVrq6chfEzH7Ym9G5ci4eM7Uv1b7RdERY2bUIUlWf/j4p5z/Y8mSLhECirHHfxT2PG0cmpOAHdr4
ao2oftjNKEmrbMuTwtZ1qc/DXABpg/X+PnC2lAPFZDhHeKFyTVB28ckdX3tS4rRc7U9f5M5s+XmR
9ULlzucFzxNj9KRnb4tKbioxxu1Ch5t/49KtDgd0XDYdfvtZI1zycOAozFG1QqXJtPrYgLRv5+U8
PT2Q7i2XUqKufXGtlppElZZJ8Bxk1vSMk24/zG0dGZ9v3E9dBsbiu67ZbL9fbRvyNok0CcRifiZ7
rQXomPZJAzhHHNWv/Nx6K+qF3y5WqRaQqQ0aRU0LFlu95ax4YUr5+QZ44+IdnBshKcUw0rjHFU56
iI9dU2IOkhBOnRQSV0hgo+x2oMOTFHkBELSSIUvfmJwYQ0vth7CKgsHQHSXJbzWXHt9eWgOMJfO+
O47OVIcCouIBC/CGUXfKxpIA2a3Sgl8OV/u0wHdQEeYGqdLQLif7X/i/LXCwuwHeSji2Gc0XDfyl
Jd9nU6w5t5/t5EcJxZCM9WRbrBIHZs9hQdp71Y57aen6H03mARdRWQ8sZIXVAbRkKwLRbvJWDGYK
c9eWBKAtriMmmPf+pnlzOTtHDCJLZUZCV8U+Gfu5/v5oPSNhxAguz2a6YEvAqJVw13kibd4Bzbkh
fWp0zkCxc+igVbcK/HgfmqRiWz/CzUnWZYHFLE/AowIjub0Rl0LnCoN/DPX3ZuH/orfuqgr76GGu
T5dglUaDmz8WEeK28n5mxH2y8Wc/c5w+pQMaN4JL9K7zBNwRB0BZz9TvmzOX+Xvyhz3ESaTYN0sp
K8SO/a+/XowSIhhMZYSR0kYu8VSEkTHe8hGK7+ioO6Sd2UlENlqM39/E3L5B2XLK48bbojKyqZVM
aasIttuGxwBG7dRgXtXoMNYRAebBcJtxWCCqpzhhOznAE7rjz0R6yxUoGUFt5USw2/bOmTtbHS27
odI9gE7SiM+oHTSxh2rgPnuHHQbDQ6UnLvmN22tKYAsUgOf/g3UeeMNjuWFDdmjRdFUXe09JCs2E
wk6iPjklLNsaF8u/RFEFa3gC8qbQEfQulgAUI9+TL7WaO3gxNUAQEE1rDw+dfMLwUG4lyXPF4plh
EDvZGAVmLhmN01/7/IBf3xLvVSqe8ZD/37jhMA7GPcEe6GlkttLalqAbMfa2anHGxh42hI9gFuRz
J6ss0JEu9kX0xWGce2EQeuVU7iZWQb9cDorkvsYpbUXqaNyjPjVkc9sphQ1/qWvKtwzm64R9TN+f
zZoFmk5XQDcPyc/dX9hm2RG90lLICs1ZvMauf7fA0lmS6f5yExhs5QoIGNRl/2RH37EOsk2NIt9g
CnViD3KIcpmhbw5igqwM6SOvicyvM0QL1O9pZwijETHPiGUyvkPUWhn9YlFvPKzCKGQ1EGIN+y88
eGa5DuCXHBY+MkvcyZzKDH7N6PLXyz/Op4AXZnCtaR8Cdwn216gTAEqNbUv4K0olrA6mk6m+k2js
lw/yF/JypeVjbnArRDNxHI4r3XIEPbRh7w/BYcdk7Uzan8P6E5wTG+ARn2ZXILxIi6ICqKmiqYNN
DhDyeRCT1a/hn0Sc+OP+wbUCR+o2b/DWZK7h5DJGjfjAsMqhcLmlMWv8IkjueX7gph62P+PqL+fl
7Y9Rj1J3ft0NAwrfwd4gsmDRez16EkQ0Fmz93mm7Kh30j+/L1AK44/cuGhnyxDb1rRk/Goz19Ins
f6pyUUGNQcK5zWbADv7RJtAimPnl0/ihuzPw+iy213h3W7DaPDwmhOwdAsUc8GWm0vD5242txiA4
6Jg4mYtGMJNfpDB92QcxgBqX26CUR4IbCALOdMN7MeHZfIdZ61/f0CgvbRHpXJTJlnOn0g5hFbIA
Z59pRuN1yslvZn2VfP3TRxRPcz7RrdjXUu9+GjNlUg5Hu8QguLKVMkks2BCGENzsGzMVUf+MPSUR
VM+rC0W2QOJ62kfOaOXpdO+GiV06BwnKkrKY1I7ZMEaUTisP2tW5nMBc2UICnefOJgg5JatuUfDA
Q85dj8zmrN0oa0jQ9rXdjMFN1RhH84lx4NMfyqnGGlpzEJWw72DRKgViDsXG1rHH9xFlNCcgbkzi
ZNQA9pFPqpaS+Nu5fqGytkNnf98V/TOH8q24CoSFBNx4za0JXM90iTTTClp8ZPBoh6WgSou1L2Y9
g6zZSwI2DpCN2BFqpafnlmNY72zHeVf89MJLM+mVA9IXO2f1VFyejTehB+RwtmtvcsiYJMQiuAlu
yvjJI1RGZVnz68YoxJL9ZlRFV12mudIdr0n2xhlf0XwTfkLRZCz2q0i93F4eHkdW/78ybQ65ufzO
Dw1RDtl0sVGBlP3w2dq24/6RJMSsDrqm8ieLU1XMkkuohJgvHT0bYmjDYO56N0KXAi5u8O1HAV1h
hT4MQ+qL+TJZay3d/WotnSb2+G3f3bIXzNMyiBA/ywHP5eM8ecOyMHYzjhCfOAu/fboikXnMF7XL
MgGpGmomMn1c32l+HmLuScK8qoOCkgpE6+F8FyyhkhfeYC7V4YkV5ienonSfekVu86k5ydlgHKF6
nT4GJi/a7yZZLJRvNmRVrT6juZiSc//+Eyyv7V4OIt3MW+QdDQC/ly/dm9FlUuNv/N3J4I6Qybae
sjA+IqDeDf6ErfFDuzd+Z5aKUk3Nv/mhZFl7rXw842q/HgAMjPiQHQyhnXBzvxdNlwyZvEJSsQNL
byp/g9YVsIAwoVzvnaEoBcBIRF89QY4xm5ascAVLkySmLALO55jisJp60f0BPbu8dpHEkAWBTIHl
cikWwJctatwIFjCGmVVUSkFkcp/WBKMEdg3BGZJ7S6hiBCUrB6FAWNROnHnsM3ESpBXN6kRx6XP3
meo4Bt0UciLuUdL1C3Wgs4qo1xEqejjT1A4d7071+j7VDkozLv/gHgaA6PmVVYvbeqvOUyJhDq0R
wS35pu/zWRsVpFfKd3I1TNR7smEEQhfABDeMzWvnDb+ZeTXZISmf9DEsjO6WKsm2ijYpQ7cvuWhZ
GPj+6UAvtw4iw0kKLwJXPBdHX+9i8u3ixvG3NfvyFbqNRkcuV9W+oBSUitp3Pqakhy0gKaPbnHii
eYHTmlwGB7UCSFvZPKUzEEm5r4H6DSPoahSnFyxaNpHUJLjceigL4xUUaZ7tB7+hLRJMjbIxHDDc
79dHxc54szn2jlyIEn23wuSgyJLbDEMML8Myvwfy29Zi02Oqv6vUaPKnMy0crR7gOK1H7ukOlpvM
AQdzj7cun6+D7vm26f15i5t7ZSCmwhQ3vif9mqEmlR6E4tPaSPo5CziQLDHbjiHP0Xz9TkGMT6Io
lEyQXul6yLYebk7uyMvM2jCHlrDRmvBUyGtYQ2oKZoTOY/gdJwmd2QRPBfusRK0RpuvfESBv0IBz
dpZTWmzucX8hXEkrocr9Ry8OcpSVgd5nkg2zt7Dg+b0AiyubCl/KJ9+n7+xGrgF7nVHD5gH7TO6Q
/eyROZUJ98naXZzV+pjFdukz0RRZK85iDDls29QDUgFTznXkHuNM5rElTsGzQDGMYgJuy5xISoT0
tQBbpi2vIzy6yXZYqretIKHqHgyvg9MQ+UkFaT9dHNT8Asy121keWIasacVXEvxi9GYZEKmUCauE
TlJpPpl3w1ZDzE80XQIgkFb7hiqlntkCiT/Z5jCdb9XnOzzg4YXTde8v6kKQA1QBWVJQSzpGWxi5
j+oYJQigiZriBAA0tQVH1li7R+I77gZOOL/emcQYSX5p3sISbNzUmv4y1zKdEwzOQ4mEkrbt7FwP
fwMrtPRouhT9GlKGM1EF/zg9CZay2VCexIl+U2ty8PkPKJ9CM/C5QkZ6ozmH6fVcLa3DOjeCMKPX
FsQgccBgXJr6zmOBehU7kRNjmdtw8w2wSdP5VimuEt5a23Hmk0mYrKEWtOhTKuVF8SUWA5IOJ+e8
kHt9U6o+MBVMbL9r/IPUMj/qyC9td6zOLgnfSM68uQVUpJSsUjBdH+imdlL8dENqs4Th9cDyfN3T
s82EHdsZViDjhoXtLcTS4tWQdmWBS5XO9CqQWZw/m/rCzkgPng9tM+OWtHyBRGrp7Sp4IfJxqOLV
e6KncR0VZ1Wz5NInGBYq4sZ2v8gCSY16cpNl3eb2iW/eGCv3oXzU4wMuZQTyu76Zmmt5p+LWmOL3
RT+6qYIlwZGaIblQZ7xfXslV/S+ZIelzZwluHKsgM/rXqqAkUz1NlEdMXXA7M/unewrANs0s6mVX
X+QvB7GaQN29lX8QEVBf/NsILhEfFn8J/Qj8iOiGp7+oA4/4VDKWoiwGYJcyTuW9IwxRGE1ktk/C
HOZx1S0CFWN+AUs65WONCObpGQ63ywp2a+jw2w7FLv6kNB4agk2Z1XFwSyhxhvbVwL1YLYTzB34y
pQ808UArYSXPtfQeI5aiR7q7Nrn6W1PkVqEiopMothMcDbSdEf39g/Ssbf+r1VV5khxGc7uRHJ7t
n+eXAoCpb+O/fTUr+TCP4/gK40TqZhtosNZpZ3aagrNAsVF2QAR6gk45Cq6nkJQl9YUpLX3L7Ydt
8KfAprrrbwQd0BWSIv+BFeOjWS7UULdVY9ec9guU754SWyRBOlKOZi5uDlpFLRWsprUFjGRNPhWa
OeDYEc/RpcFRvOVay66rON6beRZOrlUycvYH/kLGGXnj0eqqphinp+mmQg4aO76TxMSfG8MszaQb
Kbpm4odajK/BjX3XVXJL140RZLqV/VfehSTvIJZE+IPdFxellrQFI6n1wXHyNqS0EZyofi2kwX3q
XjtD2CXwGEaxjSAJU0a7xk0VWx2wHVXa+JnLRjtdpirwk9wHtoc2zcPcOR10eMlgLsyf7F/hr79Q
ejGwZya5+C8luj6S04GFWvTRzTAWwn+JQwBZxCn4JoeKGV5HfFept2WjbhNttH4VO/94au0nM13U
xYBGIyXtPZjK7Udt93fnrcHPTyxS0qKOu9JC7Lc5J3B+oZdenYxNNjNx+Me7ulD6DOGnlXLsTDig
QhrY1V5iobtZeMh4gFVEfDErbq9nYF/U7oqosHsf/8k2/KHqvFk5hZWnSSJRRuTTVBlp5y9ySuK0
Ou4iCy0J20AdBto5ekMTNo/49OFWHDY/mQTZw6FrJHhh3/oCr0t8h66omIHUiBgjo/QNpC30V9TJ
dvF6tQf5VX334gv8eR4oHnPyY3VsiH5q2s1CVLnBA8YoFvXNSRjgNvVWoLwJmU9RyAtmlSjYpSf/
5+kkiH9mbqGkjzNf/l4IEQxwX1h/mLNY+F6wweXCkwJ1wuY5nw03MnMzAn1lMGSU6eJK8nAa8stm
280O8xH77MR/oj/21Xia/dzU6seSXmXRREx57DS1f4BZEjr2MDNOgMbWJxpE7yVa8Kb3SP/v9aAg
DcsB+XKAVlkuLo7eNiCb5gvNMLVKGzuIa02ekucHIJdR8LzWG3PkTfiOv6Ze+DXd1rA7MLRcVJLt
4aYKDk0EoEEzh3zGePWAVECM9uxh1S61GyVKBNIEzDBmO/P8lKdwr4NEI7Gm+E5QuSTt2haQge19
tHf/5bfvkXd6qBdxampzSVF/lzRe/wnV7XwV6vrahTaN80+s00hR18jCqXhdZ9R4G2rP0vIHoeDc
IcsaVGW0b4oh5OSBiPDythh3nt6BSsXzCsLFx4Ol6aOXTguRTYXUfPKC5AlLj+458vmvR0cAR/Si
uVCV/FAsSj/fPKGa1sY5OtfYpOoq1LO25JEkNRSKO6mtjlifdyGsaP/4YHZO6E9E3edJ43CrBGAr
PJ0RPr7wNCDtLP6JovP7e1RTbDh9w4xLgR3H6f6Hk8+oQTwELwFq86sLM+avHDZPm+KwkqiV/p5t
C6vh9MMjU/W4bs8Uk/MDIjxhlkEEMREaVVcyjMfjJFnnEk1dPvEst1eBvhblZgx78dosx963JnNL
vmSiLsGg8z86GdtYRSo3E6VG2sRmfSXaMyjFSgK/+8XvpaTn2J7aTI74hKALLTfTGy2IU0zsbOQQ
y2/RrTvpDEjrEXZdSbmaJQ1ObLBeyxjowNwe+4G2vqKy2ipaCR24u1stbIlUbRHzXtk+BdjvYUx3
s+nj3mie4inJRGibbHbzDEaIyeg6ZqTvJdLh3wq9joCkd5rA0gtdBHQNas4AmPP965wB/qWKNQE2
t2VeLpiwx+2bSyFMcIuupBqpanaug+DN/fwdVhSurVGAHmPLnRMwig6UzaHfTfZU8LngBSw0SIzc
zeZpqGrF7+AwvR03eWekHKghVFAvzW1/2eb4adNZYqNeka8rEsy7thSdRYfwOaA24Yp8wij3zLUi
huoPo0pZ8YpGLr9JW8xFsrP+p7skhY6JClBJqdEM2DlKqVPbikm4PZMVlTy3sad+VeIIJKiwKs40
mcCXjo6Avz5P+vc0pRZLUlc/2IugdG8N9+f5TD9vbwKLnYaTCWxMFKZDj3o2KIdREkxDv5xlg3vG
VXm5uVQr/tFxX9sH9CAZ3elUBegmWtBIeaMHvcqR0inx0+IQMG4SAK3FV2XYPK9IeOfJ7Lg5oc8N
Kh7vGzGJWn2pecs+/M6TgHWXqUHjBbWJHqXf9lNciv5K+N7YNyKN+oSI6VFMXIOCNFWIU5SoqZr3
r0+RUkcRDLBgVBomzAgUGSGdICrEHs27hfeIHgxoLs61AHCFvkGYaHICqV81+lmS2AEN6XeMvCEF
znCQBaAVEGtuumc5e7SoevSk7tWBl4mTt6YE/hFL+auLWeJCALF/UUQ1Ec/ZnUILAiMaFDFxBpIs
KnykxBdUFjjarg0Pr+4nenwoiHWNcKTZrQQyXIJM5K7bjfuU3KuM8urtiUI/VU1S9g2vHVPT76zT
KdX48Um2GOYIFSDotk1HmoYdInY9QMq9yt6kPpaDWqsHv/Y+5eb6xDOYuFuxG+T+sL91Dt5VgbiN
8mUzJKHJgfC1mGkHB86SQEzfQIhTgR9mbb0IO0dJVHOZBPqumDK48LJq+vUv8dT/kppm2njwIOm1
c/rr2Hu9v/ZAdQqL8sr0FFwd2Wf8PO0bKb3c5fx4O1ju0XJjTxIHe6gXyS8hUMRJpciUMFP8+wBV
Zt3wAh4sCWQ6BGhtQJPAbwJsk93tS/d0/GoZg0IKBIpViLB3BneQ/vCL+wqzKLBDjrGq+Vr9chJL
zKpxIe6YPbNE9bufMEIyZWDM+F1xwUDEOZEtVr7zQ+H1Mh2tTAZwvBhH9jXTNuaRwxbv8qXQLQxX
cqw8OUx9s5uafmKRbRzjZrfw6u2vIFdQ7SFfPhjmPyxL123GzJHLUfbGsgCcPd0LxPX+wWNoEmtO
LxU0ogpYLXGaZaWcKgYrC/Vrg0ZMa6DM19I1C/x+ak3Hn1eUYCMILDuYaNo+XjhNxYhW7Dz7YNzu
IvyVLruJ+NIu3ax3iaNS38SaUhOPMONq1RxRkOxWKDyPOfQ0cgkoYY7hcrnPmnE+a5TWU744YVm0
0mztNz1SyVcS4jnkEgZROFOm5pMLugW0fNhyp/HFlySUTrZJX+1ChnVQbnleUNuaqh7EKSQiPcUw
Nb3AaLTD/lKHVXqiruuPrSRpGGq7KPw3wwJ8uPyMUl1p7LvsOPFifU9H+i5Bva/N72RSROrGOzDU
BT89WOQTIApGz5IasX3S5VBpP6oqMGVt1OqK4iHOWg7c9Upf8y5QbUUzFT5QHw2ZtLX3eJu8Tj7r
oSf4y18e9CysBc3GMR5vvKwz3FC52iPK15AOcZ7z8u1WxoSdQiFyf2o9t2tDf4fTgIeNVbXDmhbM
jRKntcANON4fSe+xf+At2Orp/bdiTlbuEgzlHgxMhMtqeRjx4btTkMzbRvhrlUc/5bMLvB65yQT8
zC+AyeBAtu7zi1+vFG9Vjw+YKkYVk4ICOPHbVRcquC1zazwMggkennfgYIjuPq9XLyuhrPvpbqiN
VNBO9bh9UU8m4qt07e4gP9dibuXEZIDu+4vzqrtGYna3bO/0W9uEIZpiPNxGWDhbH4bMRqQ/kuQy
Gl4vRJI764CtHwe5FAHMAtW0gIgy+TNu+4askjYIVKrJUddpyeO9fX7CKvs4/0hMmEYRbSaGElCL
N8iRPcbgQUVlBdhditqqMSQihqVOQG2YS+243vbGr/SJSlPbfdttA4MetYEiqMjj/Rc2uVrbhbxk
Wx6Gi8q1vAEjZoRx2UWsMS0paEX1uowPKbM5gcT02oJoPxQEbJ4hK9A7PJN/tXWtDdH58qDekb+M
CSJh0k9PAWcFsHyRt8IoQQZzzjV7V0PW+dV5wAy8V7Vk4w6ssyMqtbOT6WSCfPYIfTzNTH3O3w6A
isTQXGUaFyscgC0udWAPr4eto1uBHOoG0zFGAuqaFcnL9xFrHBnnked5/DhrJYhJXxy8CWuAYZLa
5i4wIiE6Gj5M1dW8HDR8aYYcXc0rTNIt6PvmR1QTslaxaw90jPwOzJFb8JPEeOmZ7lVF8P4YIB8C
7I4N3LZBy747V7+t/HnB7IdTo8F2yLl8SPBjzslz8EWs6UQ7MbnJx6IEM90X29K9fHOFw1ftm5KZ
C0IOBVBXAp13IEVZDmM3CM9jZDAnWkyv9uhvz8BIBhP3HDZ0gyE6Vi5PEvKwS3uh8+Bxq7a2SLDa
GctK58BPGAm4HMetUZzgATDiBzAf/t+fjDbtkSUpHl7ccgxN2F+nKbQhHNowACPbC6IIVsieMDR+
c4HJXwlPfBmRYJZS7Mw2HflxE1ynHzkNu8Y/NYhuYZLFIe85Co0sF0LUQ1NnPxOaRn4hmH3NyPpN
50oAApfC70s7A9iSFg2P/qUa1oets3ulfeTkqrFt0w0zynAlMF5iy4P+5DuYTeKotVyPX+83FGHs
S36mCRTCgfHZQxXhbEMe0FLKa7FyI2R3kc5BfJ+fk1ytfrCP9MwVZUiL+BnKPau3G29aMTuY9ZMC
6OxeHT9YXJInaxGw1eMpbP9iiS94yAtxGNAwjtEmm4IRb6x1dgQi89Q/NHjjiHBDJQKH1TC96zIB
sv1dCqBZ7xJA4mhStJH/wPD7XFYL6Vu5yho4tyb8efPQwMmjBC3CBP4QNuVOsnwHbacQ9QG4PUJq
MbEsZcdGXzhmyA072rrxUEwQDR54tt8LNLdaeI9Qbwn0hygKOH7jVc7ciw7P6ARHeJhWqAEqKrwh
77pjRM4GZFh7aoOc+pisWtfpiZqzyuKuIPhdf3vNeaihVhhp04+JOzHuGcaUDtbVorZyLi6XHniz
HkgWeQ5HAfYaJk5mPwwSYkfu8A3iMY4ZRYQ1I6ycQwBdmXq1sVS0kg6WNPtfhEqgOfkOyb3sOgCS
higBKvu6rJNFYteOmJEEg8rJ2G60QnD/XU75GyScOPNwXaSoQ5iif6JxxBKu1H4VJr0SCQwIghEr
3QiS2j3YetDrbqvhMWl1hb3gCdUDmqAtcZCOmyZ7HpC1vkn1OFsr3G2f1wUPRrsn1SMA3i4HA1sx
uSDDRp1ld24TEJdxhCQV0K+op/39BaHOC5oSi+ubKUgV+XKHWgTkxsKefozem6MlYqzkxJSAzlK3
tntb4NwA3eJbhMiiQyBbtSdXxH6DLeCogUSzP/f4p49AeO4kMEzV+tR1Rgleycz15VbmxAHTTAdF
1XbzkDcaAahhZiJs6c4KluLzXx8S/uHVjU0+yYFIcTqvhDxwpxfQD6tIela37YcFvuWLYu0L/TKW
wZRm/PSMfMjw8gxPjpeJyHOXUbSb66b710Fse/5wtj4Gb01xUHH1T3IoSmdj0XOsoYPlKcCuvitV
cXmeQOhe8xvnHSEspXGdcjn+NXh27W7ZktS3pjJB77ezdAS7fH5lw9HJSpwFhiTHTLrUpD6UZ8pL
kiNSJsmC3wpGPm1gAgNM0D/3hGGU9R9tkHXW7QbU1y0C9dy0lkg/q14nmEQbMD8FuRgwS82wKJzO
dOtLW3UagT/IhnNsvlsQQ/yMI1o10a5KjpDlkuTL0TcHdU/deEdNS6uSpbhQlvt24rR8glJ+SfZR
/Pn5ky/eXn4q831fbUQtg5p5sE3nFjWDQjsDKrJvu+14RW24t2jgkDc7bIQw59f8gmIg4Prh/Il5
TJS6XKMi2riZeVsoJsloI4kLrKTdPSB41Io0zv/Fz+OzbzdB2U0okttt1XM0JcNeIHdxt6WJydDk
4hOsc8Yjk/cyaAYcErnwq2FBFDYs1iRiWc9AC1elJptXBvz4V6paAMWsv7+ZlTJExOGCuVXfGZVR
IaKAHCDA2hCtDz0SXkp86I8G/hV1SPXaxTzrOCv4dPSHGMD8JGqwJcibQkJEKmhOR5ZYtiFMecV6
C4zmHXGilPy95FSooBJ+FFc1bBw2TvBK47DpxAH+e9ABQd3vCpsRWrExmBfGV9GfGgZ+DPqPB6Sv
90cK92Tsbm1WUg0wUXU5+sNjdiUhzEp97sUgmca+aG9ylCkvp53BMYPzn9gesi9Chvm7wJYfgZZX
lXsLT2jzrhfLODclV0eMPJrtNPULchn44r5Nvmb/jkQxxS2qNSbmo6bMfx2w54U1TX6z3XrhngBp
8qCZetQpd0RgbgJ8GypPFDCQWMgqtcqNl6JIeKO815FcSLymnEWSb69+URnm12OZNdDDnerbut7R
nvfUokrl6mgAHexC/ZEL5aQKQ0f7RTXcUPauG0HI9XFYLnFcOsRiMqHTWGhkb+RVj0nVhUFm6pdX
g2jwP6J/G/MTSOlDMNQGTPr10pT70sA8ENuYXqoZdgokJLTcH3xMFhQcjgZYIKUkA2GrFk5dulbG
tVVf/+369VXwHC71yPegZKT84WYmyeJ5XqGpjuyjlqTZ4EMbygnNVLd8yy2ZRGPtPipBXvF2gE8k
7JmUcwiEYAFEvcYZTxgky1Rg7a4GwWuM0ZId86PDgf9adj1C3VMaGbOJIjAwvK1HA98sBnaWVQUq
0g4Q+lqGwTsHzDh/Ub6+GeHCeIZTyiiLnN+NC9iwmPLqvI3y6tkxfIxT6KGYRtOavOk9oCvS6IA+
RbbJDmfN7TlcBkT85lrZMzfkg5I4Gb9oxnyPdxlmJxXohzhsVcslHWBuryEbGbpPGUQKx3i6Pxgd
LW2M9bwBMD7131/ypgurijogu4r9im1dlpEYjNkTv7f0u3efJXUOhg9oguCpGVWFlZL2M3zNi8wO
CqqTy2AFgIyhBhwmk/Jb6qKlURxej4ue0QC5NFFVYZ7D9e5wx3JXnMNVEDw3kv+PPto6XvMvXnn6
E2Ls+e6adXe6fpAwG6hxCnQ947G8GeEVO5EXw6QxAhwbMBvz5wevjkG4ZqFChheZv5M9LVZgN4ma
EnlYVh7UjriScUUgNo3EdOG1Yd1rJwfCHBnoToyk6BQ83G8tG5xgSYMEGSrRDO7cWF0XBtoGoseo
OdQjF7W7fm88PrLBPwyu0jzVNsxP5fNEvYwxkhs+wS/kYtYyZptSIq3DSVfcAtB5wDLHv8SakIeq
ltVwzbAdmwDscMIUZKaEv7oNdybiLzGmCZYR3emkh9PfGJ33qe9W7prIhPfVjLK4q0AI0BxheKfi
t6Gzx4K6Tivs8BYAuRMScOHLgHKmd0ZQc0FKBvdJIuG4TFBV232zNYyh861vtQ4W8Yd/keQU0qqB
naXOXjEyJ3mKkrNU4DRkqUsJqc0VFtTmFe13CttKGCKqhKAqaHC5iwifdcAmqEfENPU+qU3L1nyr
/uJSxmc7zj+00FZnLqV4sjTbqA8S6ePCbqRVuQTPXegCvAZiWhZOCz9EOyi+xpq1rU02FOhE/rMY
KYeF2sUkl6Nae9c9agrcEjcaHVkcoMKZytfM5a+gHdQ/IZ0Elyjp0up/ReNqd9rj7NHRoR18jdcV
y1FqqIgEimd/FpZSeSv6BmXzqFDuOHGdH5pmFwUepkyf6c6LhRAufWOAbujEw+IRzmDuZ84Hi2Pd
QEtTK1l8QMDucLfDJxDDzNv1zyxkRFIzTzsx8lOcztjQp6zr3ISGzsqNh9Ogi1r5EASQhtsqZDCm
7IvAHu+b5bD2cmV6KriLaz0G36BcpAUO/MY2FPj3ma9ZK/ZjWzPgbRKWY93KB534EpUp3LvKh+LS
9JgpRmCbJ6dMdQCGRElR06Yis/zPxtgdGBtvFJMMsUOecpuprJvmYGQbVJeIdbbwDQEHErEaXuSN
1TRUNd1fzle4iR92UXNLc0ljx4sU1c1YqHFUuKcBwL/Qo2IhsxeA30NzkQkZA0z8n6tOXVnGqd8b
sx2gyxviatPAWJMeaaBcm+hLofpODg6PIYG8fTgPew5tzYiJD7NTywPEGoaLrMCYKmh8q/nRZNVP
JmzvtgmSma4qtFv9LdpTl6z1Ovtx4PSzJdfoZ+MumzaBkEaWY6ja1ysZ3dp65elUMMctR/0YaY5B
l3rKHg8/rz3rlyiMkSBfMVsnXGnGG71uQl5Z4DwIVd/oqr4ZT3izxblFdXFDzJWLtTik2LoVRnKH
ackzFq5gnMYnHIr8WzBtMhaDnGh/l7QUzqFnMyknQ9FyfvYIZ8m1EnJLeOYjhndarKSaJrhuzYse
uPyYLleA4zC3uwydkxnpxX8TAIhY+xo5mDNd50CUpx/EzQbNIBpWbW0W3nlUvsHQV0i/b638aRT5
q3jhQz7Ypq98VHjnyed+j7XjkZWc+mRArTu9Y7/19t6Kp6bZxQgdgEDlC6ZWGBo8VNTj/pK+wjr1
39kLphGmBTcoCNmuMJiuYkS/YKv7StpF4Hk2fiqyVH4kjqvxlP46bDmQwX4cMRHmy1ILDy4Y4urH
XiqBnlmOZvKA12QWiaWmAO+5zxBNgEfcgDU69Imq9qjphYeK980gKHM9ha3HIpsXmoNsiX1nXahd
n04teHJjFTIoWoZ7u0yM1aKxKKB2K+T2Pew4iabBbb6e1VcDpcScTQzT/iJndEsVzVyfKHnV4r5r
L+ztMZcx8O6ja/F9Q7Gi0g25Sd1XfOiDhakUksirngiluyitXRzZOmoY81fZAx24mr9eZkhUpb5I
+OA7YStwFWv+7bCgbVvRjYoHegRofgwgb+KSt3Te5eqWg3IGxOdgx85LAo/cCQZ3ecKYsY8WLi3t
mh+AG0rKKbCo0Vf8uqsprPGSUt/hSjlxWNjZieH30LZ0IcwTEqpjlWs5k+/xaf9qKNkw9D6bjoCW
Sx0vYd53rI9uEnHAzrmvadyQbKwuI/Twvkzm3Tx8ZLV4remXG9CqX2tZi7fXJxqpq95RyzTp2jC4
JJ3nB2qWh9iNdPXy8VxhLqTtI6zuG/A2HKS0zDkP0lpPTFTB9nLJiK5WkdgQ306OnJJZTXywPsD/
bwCt5qQPU48I0GbDekoGdWlrDYhm+0R1+sg+wzbcBEK4hoFAOwvURVantjD5+8FoloIkUvhgiMVI
KgIk3/T1VPovQuuMIKmbQRCBbzMvyImpWoy5qrV40XkY8QowXOeL2BCXh/HfHld5owb5HdcxTZyD
Pr8Ec+/RqSYxu41X20EJUYSyvtvq4pV8w2RKVd7y1e8na7O75rNpzi8LxcAq8RkXzNxZ+MoTCVaM
yu721SHSF0XB2L+SZusdUt6Eya21DDZS3hjujYWprYDfX7wRgJDZqDxRJvwTMQ+gDzEdATBJssYK
U0w3zbvrAx3PmlI7gi6EtrbvtbL0QbysSl+GN0YxAyaocus1kY4RbR8tohdtfvUkhsEaWZTEhk3g
npZkS8DHu+TG7ueE8DJrcoaQkst0NyApqWaOKveavMnm40r1Gos7Xyvfixe+wFFN+B5uEb//TI2a
BnK5LZyu0q2cygNnj3BSGAGEeoSrTY2HASl9h9HkzcHAKmnJv26700ZtCP1XsCcxL9BzrzIuz4Ao
c3zv5bLQdGkBMfOwE+CdfTIgyXREPkBuPPRCE1WxLqGmcnbcUB4Pw3gxZdabNQQu9Vju1UBFYF52
hwWIXCJJsljY+6eQZCrukuL+bmjuoot29+LUa6vYp7qrxVJWMXhEHtH71PBFwH9WmGnR3OGIPriw
x2qg+I0TW6rIcWyLtnr9NT2jkN8AXuUiEefIy3oigX/0/emDKuLS4uc5BJSH3TuclxqzKMzFoLQh
CvqJZUpxfepxxi/q3VF5+c3OpweASoXvcJmZT/oK5aQQlifSarTgQm6tdPq3/WBoQpsAWpFx6/xx
/Oy3MIK8R7UwU/pYjNeu/t+HVL2dOq5e+eCjIhLsYlnvOFkr5wU+fE14Nfu6rzwJJJ1mEu7ERJEg
6timF7kWzyiQQbIHh4bU6ImzVLMjTjSOHHLTuT5jtUEnfxojlkN+Vki6ghkP7AjcDOVg5vM53K4J
Xwoy4B/QeBHd77Lt79wQk/4mo0IzXs9khRyZ5xr5rICzq9TJeQSzw8IaBWE/jEFaHwdlQMP5mFef
Rl5eV9QNq2EiR+yI/FcxsBhgavIwDXxmGesUK02o3nBEV5liFkWJNhkOL0FwCV8sjW0HEk/p9zpD
b21j20Gxxvza+J0tB2CaufLXGvCyWFbURjptRD9wd4ecTaVlcsd6gXEVYee4yxzgM3tRuvzKT4OZ
dfVZYrR6acqENeulmF1XoORCpU+3eLFpH8hxaTxqt9rgxDX2MGgOZl/LXphNyHeADqwQzVAGO2uB
Tz2x8OtN3+/KFbJ7VO7GC7/GRruZpc73a6b83CgL9xoZcKl9gul4PXyKe+qSep0rTIoq6OAxOIur
CYUtolZKBHPPjT3xGMAzPK+nwmksswME/ct0a3HzXSJtJBdT0u+HlypERpo1twp2sDKryP6gbfpm
ZgytaZ4ZMpdcZTUCF+57kO+BiPOKdaEGzK7OU/eoUb1dbEyDl6Mbcru/j5rfTZFGWJUrkMrr4BLm
5KCvGOmWTwqCWzeg4p0sWtYzeku8yoqxBx/OrxKOFKMW6FmKX+nzTZQhZENsbJ7V93DwywZi10kK
OGkiNEmSULRUSOmwCsO9KaLxX79wlbKfB8nxNCN6gBUnWPvKewcUmARQsQI4jvDo1eoZiR2JRihm
16RKTZYDavrTeYMMP+5vgB7VBa+oeGxbXHhuQc0SXR+1Hz/j8xLR4Ez+pzqgTY4cQjAnyWfYEdLP
scu6VcZ0JS3kUT6LJGTi6DBDq2/5sCUAVkU9EDEy8WxD8XVKlclJx1zdnCViti2+iSwrNRCWrFrh
AyUL1eRgXcSoKuTvclwuKypa4z1vEiqFRoHVnUWKls0O0CMMEJ9CzYtLfWOSml2KQwsgIQ8a7C0C
oILuK6Lilll5ZrdOPNxJt27SDDE6n5YOfkqKi41PvsLA3RgmHd9BjOhdyLDkSHGltxiRCNGdCVAZ
z2GjjGBJD/rxQOtEf9Ho8bNCjJ7dZ2CxEjQcxF+vQKpSkFA7vbLl4cl1xCMo4YASnyOn7am5r1SP
Ggdp5CDwmNG6tv1kovkaU1kSfyfOFRdtcgPp0bmWei+KReWbjlpS42LPHhtLS6gekoXBXD7A7HoE
gBzxCVHjZ8QBI0ySmQwFcwN2nCt07h1fetUNXj9vsBl6YTIcauw+09KuWG7aWHqPNtv89C92kgDY
a625Xb9K8xmdfd1uifV3polnlvZQY1r5MEKtkzOraEm2wY6BvbNmlJVnF7lNCL0nXI+jDAMumjjO
rEXMSMBaat7AFoELHPbraKixL/qOFwmqihKXkMbhtv7LR58QopvQFTDR4lCfFQmpx/FOoh0pVn7E
MphuoUqehxN0GJYIVb9Kvl2rfYIuDXGwDTimF+OJC/qpExwzO6oaLx9+KA0Ah/reKi31yXtrgdMB
/ra4qDiXuTNso4tPe7qIWHK+2oFTjc0Ws7TzHezepNd1m2CQTa6q4WR00qBdwfP8MMbE3b2ZdGTn
b6VByvG6JhzzzoGU6hdHkxQU4eyIiiFqRKotLv5CIWmN1Z7cZ2HL6isf3rhEs26yzOI9F/wxB2Wq
vEDUCVWsB6jqk6oOcVlu9IgEt/YpPOIc9s2SiJJsIZ4Xz06FDXq71qKpEbheXmrk/gKNmCC4c8GU
dlZgxyNwRmz05OpwXXekCydMW3X9oU0d39Mryw4sCbqwT3IfobIGt+N2LDqG8Vu+O8tv/lh8LQa1
CAMjrIegjvD5FEpYJgOSFtZMDRDEVAYaOV/sN0+VcA9g3nJSDAMlJxHWIlo9bpCJAWjpVDe+Z7Ob
KR6N/xUk7J/40xbfA2ba3cICcRvO7LzzzupBkSv/noaaarA2WFI1A7JC71p0QyZf61RTa1O4Owrr
L/64fepW4Au4K2F+Oby6lxzHzJB8fwD5Jgahva5xzPxJJgomc9j/yZR3BkL/rzn/W0DaqGbssJfK
G6AB9GkOtoQzuvtzhTvuLrjBQ9SWAPJCWr4Ztdr6UMnXhMfgoS7/r+ruHbLUJIw1CdvMsApGPwUf
UCNcdBGcMbMC/cxXRNjc2K2hhJGUY1PL1L3ufKiGCxnLxy0NolIiOoDPE22qTRd7uCetrRht6kNY
Boko08PdhAMsK3hyTZgu0ceRWDM6ATmCwScr0iXIT/gUzuZzFq9xqAUDUqDgj64YMFPF23HzkWN1
E5cniRAE1dILo5gn6mss8QN60Tuo0dydC8m+lBXh2yER5du8Cy1j0arUCK8vXqlds2D5r0JCJcJJ
qPnVJcz2/wLC+mueuDbrqrkfSW+ONkeB7ftS0xYcmM27E6rxraDPjsnqDFBhO6iEfOh+JQ6Efk/e
GFTPC7rIohjLX0RJmlyvtoz7oDtU5Mt3HkfKhh3MfHOGGcdU9zjlKYao450CK0iSAGUbM/gXCMdQ
wBgOJIIsC2BBrRVMDhn5EN5NQkF3a434ZfsjB9hYFFlgg/xMZm5Vp2MMmTefJtXdkkEdhvWtEXYX
lgmpWlRsOH6jgYBgZedSwavycxa6TFUHEnj4srmilf89wuOav/EpFblR9D6pC3Ar9Wf16c+ScG2y
KHR1J8eMxXbONjrnmUw8+UX3xXHOcklMdpFCcwXjaP5/JSs7OcFcfOzvLsKLUTdPVbgXhgLnbPFv
R9KLjaSUM8trgyhfZUa/amAlXrrIcYxfQIJdI3NK5/rx3yG5QinqETaH6/1yARFpgOrmaOdF7m4+
OQP0q8L/T1XtFdBB1f6Ekj8iB0oH5zmyiWGl6W9oZWqJAhoXtQBh3dCrP+yIA8UXa5KxdlwBcyVR
oD3U7HUKs5xD3jLwNT6qxnB6G1hqnhdLwzFm7LMkGm8/1YYzLgwYp9ljREKZ5IdsGjys1mKVo5Wx
2urQ7OH3TdUl4WUWVfZrRwtI9VOTRKCNLOZZ3OYp2avc9V/jTdavl8ohfVdek6kOqKp9gVNgrK01
ou0dHpCyVzjoLxDKsiiEifI8cWyLAHiijwwjbcpcNEmlBefRYdaiZvGCQUi3EaOnRt1lDw1biqxm
gxJbiFJxnRRerk+4ZnVrth6ZAPtOYDtI8gek/AavDrS/ljQN1JLXxfippjVFhX54bg5NTVGjbKfz
ATxXXwQuFfLPLMpvR16oCc9/cH4eShQUaOQcM4Do4o5Bnbc/W32faC3utxOG2lwvyQ5pisH96dZV
9N8lLok6w5K5MULpcANhGFamCHndGZlnoUVAxH1oSpaGt0tNEQPB1KBDGUDzR5pBVxwZGSib0eBj
AqY1VLq/CIHMtz21RP8iTDu1eqpD+j2pxmjvMNHImMdLt6rlhR37F6IqZNADQdJieQgitV69Xrd0
w32XdaArNpoNMZK4NQ7h5Lg6oJdFHTU2vKfz+Q8fvNttXVPHk7Dpnym2/N/95t+x6sTzp9SpuJL/
wteBADLy8DpQ4osFgfJnN1jW13hvTCK/am8bZ3EcGc8UQ7JqeMQ7qibJpXAuC3fCNYL1WxEmCVDy
JR9a5AwGuIIMD4LfTfiIAz6790e1+p40hzK+Zjie5IliQycZWzOl1JJM/tysHaBBAVxjv51ILS3r
0CTd34kcwbzg6qh2FlPyMABtHNQKmZ9QAwF56goiZpYhZ1lNdlT6GIpgONqi2mM0o2xVlqk6PpJ7
ndESx88ukKGqa9PDu3xN3lbtVRF4Et6Qq5pGXrYXrib9q1yLtOIYex3pPmNX4F21IY0qACXI7oY5
/zV7enWMFMkSCeUPssk0EUt8iesnGrjYZ5FGv03qL+Vimw/TyPekeq7g6oXm+j2R6/9M4jngdcWa
Ln8GJA/cDvKoYVqRXk0Vw4GdAas+LJcudfoPajIb7stpNQm3tpJoiEr5P75Le1mE2+L71maPUS4C
ZwK0LICyvLBAfxEH5XknzldnfcVwsOyQS+F5vX/vBQOLz2sFIivoTz8Ceef7bgu5I0qocgMQQX3C
JJmBCcQelQEvDX9yFqMaBuv/Pu/36Er46vDWRhKF
`protect end_protected
