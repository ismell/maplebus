`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZXRWDLkqcwei7g2aXJ6gpee67Mcuv4YxaFJpGb/KlrUC+tNGJZI9+bAL5C2O3n9sxUilqldWdCaX
76bcgq4rtw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bIX7p5W0I/Dj6HKJsQQV2A4WE7INKqL/CDQ34jxRNZL49Elv4FSz9I+/XqAO57jVcknS8kQ8Zk7h
XMbvTVpgniAnpTjl0S/2OeEd9OTrlQFveviS6zr4qc+mDwtGCytVPzUIoAZmv2IEGp9udC9KG200
Tdi0mpponsB4LTj0EM4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lkeb9OfU+oB+VihKXbOT1EUypxzPnDUvCiRAB7abHy5b3bhU8yaiw2Llfh8I2DJ6+zd1H2Ca83TT
Jjv5xSEI+YFjUXExP46RZfUM80A3Wo9Uf7XXexhkiyBoSgcDmYFHOoqZLaQtGnT9DtmvpkJ1Zrmy
VR5vapP5v7BIEdpaW4bfkpH/2X6gJiUYrsRRv9p5wm6iEHODTsn5qjk5RQld+1f0XjGjHig5FMrt
ho1R5DcYxeBhUvYqc6JYXzu38eh1tFDPqNTasXQLCCVM5MOuh7tR1wP9W1yv7WDWNvaWFYgaXUnM
VcUcNHrXSBhZwyDUG04ggRKca7T73OUCxwi6Mw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EM/nhmn0u0CaU82Y1a/YlSGWI0cx8Ig7gbT09AiORzyGGIaYovQMwBcZwBYuKUo1HtXIyDCKTzwm
05/1R76hxOJWMnwMEUZlb9y8PDAl7+rWLT6vsUtlMK0bisdPJO6ho9qJiS+vW+RU38HM0EOvTBIR
IGN3Si1tvJRH5NZBLjs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h+HI/g8gdGVB+qszmHp4/4taDR5pSlN+V4dLt7laC8AiHF3mzb7VpWQvlK6xgsNzRaqYSeDKjPNs
Kybh0qPbPa9pJjzu+8Xolt94/92CMQIhAHfCVV6Ftj5tjGAACqL7orzWkRoIqkIM4WJgfObOYs6p
6/HfDGVTWr6RSFMcBd8HGzGXHRkcBg3txkFwMfvCDA1TZpGfVf8ZTPYWfU2PDUCLvRLgLcE8n9Bi
af7wdkW/JBc9UXh5olTdH+F3s0q/gVtxUWVHDyH13hNDTDhxP35jnN5y93y/UiDCaZkzzVt6mJWC
WfcVfZgnlDIZW9YN0ux6k1fMOdsdPWm2FPKnfg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
ox0ymm7zJbqKwGNNOTb7sKPBVaIvx1SNVkPCYG2sbHyYCJpCMmCYD+HgrKKhzbdHW/32Ip9O0RAD
4LCe5SaqVRDXUaZ+NV8Ffwt4u9yMEeZ7gGLcMyxY6Qgunt/DQQyy4Qv+yKOiOMVseItamZ70qE2T
J5aFM8MxmGd/mnNXAP2X29W8oYi6/xGc6blY99LLJrDhY1za6I/HBGFx4WPgfina5F4cf/NiuPH+
wKK8VXXufIz+xdZ3+7cVD8eZVFkmr6GphrenYlFl/IvpLLQy/2P4rStLTe7+MPkQ8ThO87delJAr
pkeT5dxrAZ0pG8TRsRY1V7uhMHAeWSCV1IEyfl1Akpu3KeNf3e4GBqQlvU0fdbhz184BsLf5Ry5z
vdg86Lf9GbRgz6Tm6IAiWAotHxR6iaosUt4BzCt8KNXUD/7WZiF6RA+W/nEwoBh+TwAB+D0ucYO/
Vvr14kY4bX9Ju00rzXbLMgzhKSeRx1QYBmIheVDf2j+QTitdVHPrXc3Cu4t7HJv5AjYt3uA6R1Ir
HjLayOGR4nwVEoHfU71hyrRyPO1J+Qi1aesm8tprpbhJQ70BhLMrag/JmsPoBrhHX4K4g7TxvYEF
kixGclUtcIg/9GBIo3+e3azUdk+MlAGLEr/oD659duFLY1WW0tqstiqThRONdpJiU9tm52o73Spg
+flGmZrcrhw9WpaOOA/VLp1u4pldhCf3/JBIViUhfcAOskpzCQqvMxBB9RCfpTP5/nu+c01dbhh8
ASJlgR//IKkYsFogvpQQFy9+u3cym34o0Qg9eIa+7jwH2JycclYh7sl6HEwlatC0fsO9la4SNvoN
kXsXwpm2727hGv3ze5NGc4iLkhwWpNriFJTSIiq9LJSrqwRwTN3auqVcu9pZFXKpvy4SBmzrlxeF
ErZUskptDttdiUuGqp/0tYEyV09A9fK8DmNoIpj4wlPOhtkmeibcnItQqo1aSHSDo31yIUqRJfbp
oJ0VB6QTkfwcRvBFIkhalm4LPherAWRnzpc3+b30uYatHZvpwWHI6RK6ISGY5YtXl6wluC2fv9VI
coTZqJ7aGy57gJbyCDoyTu9cdpab41Isfj0sS0KBj9UQH5cN/xg0AVqdOIHI3uPjIizFuXKuDBKj
XkyxyAP/5ZvRNcbxdeI4TX5cE5m0fWB35cNdZe7BVDVEMk33cOxeortDebBxwZrICmd9AGXtrWrL
pxU0Nsrt2aGRQOMFj3wOfxWF4vBqKoExWMrWT4UG07ZEuDm83KpC6RAfWlWueycEMSEElc7IgH9z
9exTFZwVXnDr+1JMY03SugK99WTlp6KWMzDFJ0ngxFOYqsIvzgK35t3sPQoutWGE19xSMvo+jGv/
MpWcmi9USJTNvTFLWEfSFp4ZEcQ2Fzwcy4W8UjGM7vpYEv8wTk0zm7bAHGj37XJC7VNo3VtAK1+q
XxQUBSvET+LBAjOTxgN3Vf0wVw6fytbPHhURTRcElsHSZg8O3K1EtDeMWm1j2oqkMmdJsbOo8mRA
CAuOcEu7amt0JLADJSo9q8BbOTQaJasQ2SixmBaTBVAUEn9CJm80RLArAd8licLLBnYWXsYAKV0M
RTVy0rrJu7Mrdk/QMj8s+oHHcFKuujuYXLRs26gUquCw3s3RsDr+CuGFF4ibMOWsQ3FrOZW2Lt9i
NTAQj1IE0k6q3tgrOXwMCOKfae2WmDaSw+CuQruJd4U/21iCe0cjwQUjABkBWm9nzUHTcSaMDJrX
mJifh45vPi87XpxxgfsSU708NWksTmZljSKVBFW7PRNv2JvdNlMdQBddEsH6cXqTQqP8c5ZXO6Av
PJeWs4D9QcwzMEx7y2+yqIObsP7dermGUalmtsDHnIOhqe/Hjd80hKTOPi3PrfG+cderolOQijgc
C+tlhrhhTAjU1sYU1wJlv0y3wGMOEsP+ZQlTPIvsIjVJeg0d3a59iguBqPgyOizBTQnBvxLQ1IIn
JrBx5WCChBAi8Hh3eQeO0fGuMQlyNQuhzR+egMOgIPLJWGYueHaNxe71BEu2rSZ5mdQRB9hPrFyU
9DwFttrvi5QUmaWRkaPNXAzck7SgxFM77OHq1aId8vxt7577RrRF+x9o+SshIYrIjik5cKVU8H0g
EpErWijkkXH4498GE0waJTv+bFVcKMKhtIsGVQ7tEkpPDdVugnUUywy+7t1z8PfMVN0MypWb7Reu
TYhfyIWjHjhbdo8rJ8q9atmENW3rCfLfL2ibY0ykyvQ5YWlYA4b76iSDeAMQoQ4SQKaLd03DW58p
oGdzMHfz0I3j85Y5QWZ7SYYki+5V+jl537GmTJuHzM2870geAK8yVMC7VOiSPwrWkakMOcaWgQkw
9FRAO+Pw9x7CQWJ/5/esWrL9ZCPvf+b9fGxuNSDecV9Q+D5SaNcu37doeOo2+l4JpZI83Iofsfrw
4MY8BikkNPEco1HTOn4oNSKTwksf8elmXheP5gSZOdjzXFdAUksES3Bi4iJ6hEd7UcpoGCYP23MA
hl8Sf1Kh7xVj4KS6N/jlxQTFcZCzWWPrRqJn4Jy5WLEEj9owKYgYjcyumG6iV+no1nUdt8MV4cfg
0DTLXL+XN9S5alluPd05KbPW8qJ9ldIR1beXnww4Sf9M3+JVEdRplCWxbzg/WJElCNFDJUIKlecZ
IIvvgw2ZhtSsK5229uPPqTi83WHauTiI10cXhL+uPM//lJVL1467GkYwiLNahHxfTY2zLr5V2+SC
1VWvEKb9rPjo2mkE458+tfWUDMxZENhn9Ou5sJz/GqTyyLVUgfCWyW17hvTw3uwgq9Sk322rKBlA
8HVKvgew5z6J5rvoJ+ccAA9RuOm4iopS9TV0iIT13aurj9gdxmf+jUC7Y7NHTpbm8ksJm2rCacX4
aXED5mZY3Nn4Ddpro1Xm/uqeftKm219+NVkVrjouPWHl83lAhOsYqQnYpLeQW74wFWgoNaazYkCy
O2jfuxXfO+i3fk/HQ7QmY7VAcHqX1Ic0bYnih7MCDZm5HAoySyYEikvCxunDLpxH2XjSZs+KY04Y
QNUL3+kS5Gbo9krjRWzhb7LTWukfO17BCIrQYhkk4GJxcBeLgWtUsD94s35+zU/6i/APae1pgnTP
slKM+nZ5kYuo2AQXYxDgQ8XUWGsuLLMW1ZCg5Jh4maKeiyT+RHdrmmliv5OsWB8DTh8MN3RYAoHd
k3DknL3+Wc9hpJbLN74o7BM0H3B35QdYnvvs4LB/YjaKkH8yy++C95vdwto3C9d7F6JFoRh1IMN2
HFphCwAmf4BbvK5Uc4l8+S68H3GjdVLAxHnFNB/SNSZlSQhRj42ugAt3WLT+nZmgsLN2THheSSzv
c83RrnFga8J0NPQjfT3vErhRFnYR+lYPlmaOlpwdkm5T7LVsP0R0blBd/mtS1m5VEIGiaCCfNaDn
zWnTXUdSFNCUXnLLO4bEx3AFGGlrG2AzJYdxOerkdgvZ3kQp5sTAfMeLuXIEYQueuy1VSTAxIANP
uDpjhdGGn7WJ7HIeXt+UY5gcPIwxR1+K6+jSPR2uFrl/OPMJDU6ic0Ac0HYmPH9hg+oAdAV+bMSE
adPphE8W4MhzZy0/auO0viwJPM9fwCFmR08A7vFSyllp8rSHTgau/bkndOnXBjL/9nf6+sYo4ssy
bqw+U6o4qt+t0gEm5pl8/YausRcLgq4gAu3KUmJM7/DbZKlJPb4y4jZIzJ/tmrV7c75Jpbi6GfwE
kwScdZsrsZ8L4Er46vPH4oP8zUXIYQMVhtmF6J7z5ToU9/7PCrVMU8FU80u9ElytBXlSNsCznHBs
tjY8NZ+Ems/+yn3RGD7HkFa+pb4EubV++XepwuN9sZuyHpGlICUgN6pqxswz/zL8QRpOzg7AzbVR
oQseyeBwrWIhwjIl2dyzRNkEJJrtSzUFNZ3FCG37zB9VDBAD4Jxm2zocE6jhz+dKAbJuoEQ/Jk1G
XaEjKmaN7agQzSj9IaMc/CKdDZWcgVDB+INuIkqGpC8M5+YCehHKqYdSnI0qKoyGyyOfis6P1glL
sN2uMMydGqs1jO9EgoYG5t7tz63e84j2+/IEogtoUmMUG8kzmasel8SGNS82KARQA5mLkFbFpYDo
XtU4yB4/c51Jowov6cCliVSFl7QKd1eiQTeI7nhh63kTjMchcbOT5Fk5cYi1TDDW/Ep0K8OBVg0t
NCTyduJ7xy/X8lTOPlwtDA5YQRqN4AfRGU9z/F+AX00Kc+uNrAhAOn9wBArxFUfDHV7EniFEY2cM
Ve7mgbt2TK+MEWgyha2/g/kAeHQYC/DCYE1u9BuihuAtPA9GNaEGT6vGt11iA0BEp5+NYg7fpn7V
onnGg2NFVsO0GvsvyLTLghxdjC7PHhBMCraNV/ORkACsYGnCnUEoxP8FpUhgVE0CGNbInvvhD4zX
/X4kh0uesW9KTNXq1jo9j7z3dxemLuKEmnV3xuDC5VklNaxVSodgren/xctCMKjEM9wJlGcNoeUr
WjF9jkki9m/b0PIpwdMa1HREYfc7ps87OXZ+aRaAaVTmvzeh9hPupD20S0Q6ClpxWUwOgHKsaF3f
rcZe0VMac0pv2nEApY/WaP6EH6aL1M6JJzdKHZi8B5bAV1n84Pe7t2tsb2fiZQboj9Rbmk9hYzFH
jgAGhPYwuQgdNokGDtiF+jNCVLEGNaR/a0s2n5LxGrYIAKa7Qv6BfUgx3cmgLjZ7Z3gQlo95HUOG
Xb7Mv8Ig6kZilR4b3jzyg7jd1ItJFf0RD7OFTRLOvWGoi7FDk+FxUkIqaNve2simIEH9wXlGTlQV
kgiXV9InhBhtJ5KmkvkO35hG8avaX3SuTENvWmvutBfSnmPA6nRfSQAgqVc66pe2wnBbvW8olaKy
QeqmOAtxyxCXTI7dvJ/p8gD3ZcrRnRHHw/KiB3g9hxvkbOl62DlN2ulDPbEqJ+kggGx/8yM5I3m0
+6t284IWtShnHTiOMC44Iar6mtY+vuCugqbjatuIABtIPYwEFLJRIDHQBaXXGhDh9B8dnUTQLfwP
JwhOTirClPrbGQ2IEdugE0eTLeO8KQCgILPDoVfiXpQjjtvVWAMbwDYgLBFDRrpesOC/yDj5nKSY
L5Et3lodGWItLyDruWyYX0drvhHjrqrt0dUlEYVVI2KtjFAE5HQs11/OHaE64ZgM07KHV8hckaKR
7k0VZnZHxYY3q1XcjSwbCzwZv5jA2jPRFFEJkl67ay/kUy1Hk5/OaYQJ8GRsJ3+nl4/IeO6TA7YP
xne5Rj2GGG4PkfCl7K9+CB4Q++SRsCs5Eq1n/nRJkVNTxhwsWNaahhkZpUlOYKpF/eOuqNTJE+Yw
10biUOVexG6PUFC7TvYlCLNkdxz7fMaLWO84swF/4aggj188pKJIgzSORY3FRLoFvFiUxHr86gdj
twBU/Q3ayeTDvFFPblRH0JH7OSYEr+m6MzvhUgJ44HEzqaIK2yWqAp3Lw6ypILbjfLC5Kf99Rx4J
hlT4u3vAHrist8RRkEEvXE7fNNl1gB360MCTLLjJ2IdXCZDq2lhi3o2bGycyMv5kxdtdlTnkO0VE
MeLUMMEIm1Ja9dP7O1c9XkyoEmq5OBZ+6An4Ph08GhmzD66qvB7b3h1fHPZ9Si2v3Kfqy0uggdKj
blWysoHDrLjUuvrFNRXp/spSzRWc5uwKbeiD03/HxAxHv+RyrQyNxDkM3nmxEmF+YCv8/iKa2Qx8
XsSl0n+FX0424wk9k/DHEvYEf8WOjnYfJwO769MlDBu4M7n1OIMFoWiXv7l/A0uC8FXhSUsh0kXP
rW1X4zBUyQjt/1pZxsSdwAeOu1REu0Vb1N1sD74v+AfGgO7FnQWrz0cv6Cm2WVDD8KCuP1Zw4h7e
kTmH5am3Tf5qHgoBvV/SLLVL0V2Hyv/i6zTp5x3M3AFOREtMH8jRyjMTgTW1mIcx6vHfNYCttatL
y2haLczrkSJImmFfTj6COHNMEVRPVvJ8N8gY+Ii15EoqFHRvt8xkbQopXCybgnbktj1xVGtpIUIs
ZcUcKkmfOouFKlhmQCR7vJzV9hLYZEI6vamW+ll0OgCPzRxdSj3ENT5NNkDWz64l+G7Tt2V1qjdG
uoiedakN1BwmIdkRtKhduvnPCiVQ/Qf1bjR0dCRJjp09teRJuo2DLIGIaI38TuPZk/CcdpYxU9A2
1N0pg8G6QHntLIjt05LWO1qh03k75taxACucM8TmxDysAxaaB0C8Y3s0CldCfTk1MT4XW5pSwX4K
1hXoGomH5uvrPi6yGK2Ke8briff0T8CgUXuIZHKBCdolrIiKBUCCJiOs0kWfr6aGMIz7gj0LwPsK
Rs2t2mcC/Q4nWJP7zKifRyJNEVi8x757GHzYUPkc8QGfh+3lF18n3UfMkbrfZk04F92/5g+2059t
oFiIve4Urg6y70SrtSZ22294q3b4QGJzmz6v/D8azGnMnX/JcbS8+pNFyBC1bhdKWX4vTspn18Nu
w09ldXuGGyL3hi2Y89Zh0OZev/PyK1sEVcgRSr7C3W4Hxo0CmzltYiv+ffRSRU3UbSCj9wf8qcyu
rtRkW19bkb2D9KAdPcAx/VQqkaR1eeGJyAKM6HDd++s0m45e5N9QRm1qwu2mETgYqh6FS2/vQ/ME
newTwGsx1UG8K+g9lJyCRsQ3m8Q92eTAsbm5ULNLf2i+DqngnoIp1QWHPxs6qbx8/m1+T2s0jOrE
U3YYPRtaqEViCaw3LIVKAzw1I0yr+TkPghCREdim0t0L/0r3bJknute40fimnKu1XG8N33708lTu
Haa3xJT6O9p5SU2Yp8urPu/GezuIq+NMN8EMBenfiYtGqFN30mgF8oaVbiQ8djAe0GgtofNf0TC0
k15CUBOU3axarWM4pXBX7Vm4RpLVsCuZtgtrK4TcioBgnt4J3yz/z78vEL4jnKoNRPsTMZo5IPnk
c04blhPM4no1TK4BZYnus2LfQ9/ui1AxAeVc8H7QLpugTgjh9jZISQ2k2fXgxJdzAgtoSOlP+91h
Ok7Y8KIrOZSSQQwABzp46eXPxbC+VRvTVOXhuK6u8oD3m1CwzP0MDJwzGYcbvIB8OtbZk6LAvck1
3TJ6ptUkBklzcIy2+YCwtm151TbH1W//c7l4vdbqb7q5FVaHrRb4kpOPYtGi+NfhCOxCYKX6hv1y
7S5A7WStyGoqj+8g3aMNFrS4RioyEbCdH/qvMN7H8EDLLx4v8j5X0eKCV7bnv6ZWwEkepb5DQ/v4
Poo6CNaOiQj0SQ61RBG/upDwUWt+3I8xX/CHsYRiy2Bu05Zsd+aqQDlugVJdBWRs5gvDb2VIFcWE
Dk6ljzdLdZskf31yIOERjy2zUZXRHcFJWSXKr83t5IJ1jVZyaCpgRCQTb12Xd4hsMRVGocy9p9gr
PB4aF/e/lY1tyarOrD8eSh60xjU0iMU4WOiD9VsgakmKEa+08jtodUTKTyJfYuNUBimCnki9kdsC
e2JA7fKe2mf8dwC6K1Qkt6Z9OEBRbatetD8H1LuyP/Kmzuu49wZQFj7zR2t3qKY+XObjZ5IlYldd
Nf8ztVFeWtRSFBKoTIud7VQl8rxNum6rrn+6tB8YTjskpDtuhAcBi4CdBaQC3U4CYVh7uGW+vhoR
K5UnJ0Ido8hvelLWOTPL7uwM2IMNI248L0YoSOoijCUsjAtR6MJmGZwpZa0UFWN5XZoK/uibHP5E
I8mGSr1dt3Rqr/1kntuCylbhEhLwZV2InXA4xY4JLnl7BItWWTGqEVt3FNuQOLpnSzj76oh38q6g
u1/VNtEiJmLi89rOLPQeBRqsCzSyqZvDn2yvYzIk4DDIsGCrVuvP2UIooEPknTGmaOEVCUMHEhbr
049Kq0DR6xOTawwCVDU0B7xm3mmwtuntjedhJ7vyTqn3EMZjVXltZs0e0PZy4L93+3+EY5947oP2
II9d1spc5apsOhS17F2Au7rJ/QLFuSgacDl+REdhzp03ZfguxLXUkQrg/ur8eSkcXUxVtg39Cio6
l1qpulqeB/3llxmbElbVvpsSxMC9isAvDdXbNVjMckz0vN4ewpsMzR/sE4Q9tGn4n/qn0aqTTRWj
3whT7U1wetB6nAVxE40lycok/zpwpShiaP/GO3F+3Of0Z8GKtWBF63hs8J+eC4sVTVcuAiAkfzjx
jwaIHXETnpySVPueJldiUzKdijLUFezvosgyIPVO0JN6RHYAzee4GqknUcAgrLgr0v62+3TA5Pm4
PdeQkiryUUVHztqc2BXZqw9hKk+Iqe9S5sijsffYavS6eRzd2UsGT2axLyT0PU1C0FgGpY2gU7Jj
Vv7oHy440iI2vrwPf3iN58pvazFnGK8pigRyJqzmiqotSpfp3qqeKVeo3lD82L7JPk2g9VuxRbM6
4auibEMJuJRpm19wi3pnvusgj7RdBuP+loXf/Ult/IAjH55LugjI8vAn62vMEdRafM/gRvAh5zva
jL/EZXWAgd4/zGw6yQ7JpgaVQc2dj7YCt/k+SUqDfA9M/pLzJcfQqDAjxvBFs2wHUN3knEzspFHa
x2P8xc2T2c/a4ZWqJM3IyGX4rgu8NZaf8/Z4+B6PWgC3uPwdCuGBKuLraGc4Qgl9UObsWHMOldPT
K/WBUVRhTexEt9xBFaqsviArGybI813vFQvuwucdN5fVkoxQHGOyZLQ6iLqYXSSiVYReVVvqMQ9Y
U1k8LMlhdBS72QtZuIqcuaqDefJDCUkzzDYei5NAY/+J18ZmkIMpmb/jV98cdhYONhAi1E4bUlr+
UfdLlbs7/5wMhNcHwWSaiZIjVyNVP1ZiuDEHIekAyO90SE9hw1h4iU1oz1BY5LJ/AAjZdK0zDz7T
FNzrDEWAGggsH5JdCIQWEfa51ZwN+MPb+FTiSGGR5Rtd8mcgl9E00uk4aSYSLBmgJpbB5jGx8F79
wjs4b+Y89Vaeitoydz10bpZqDJDZDIJ8V6Olr4vkn0WnhHosunZDQqElkKnunbAmt50LFIA4VRFe
hfJQeo3c7SKft6c1Gy09lk5MNl9rwLRkaBkmq8QM+MF0vpw3ycZugUhH1fVuDfO4sA1OmX25khur
m1Z4UEFbp6RcErrBcGBOzjvVvRtiPNHj8KkUWJNsTDC0NssGywXavPA5c0qNDpOt3SNpeptV81yD
k1SsE5Sokz2+qyg0TMUC/PYzK8zE8oRK8SRZEIshYmRIsRb2BnWEFr3btd+LCdgN+EdoHR5mMEUo
3pukpgsA5e1rIYO4duKEscfiGRH4SGaq5FAlQaQiZ5vHd/LCFGKzJMWek8Onx8MsyKgIfljYH/4n
I94uXKFca+lMSR2gb0tGqiU+Px3smlOxWfjmiXHYlMtz4rb7C6f7xJJBVKpL5VgzSKvVNjJwo+u3
Gl3ae0Tgc0d1wxLT5hby/z4HIr8s48tvQ00g+ZF+GQfm8SXTmESiOfNqxpQHbAAk9LUGZCN15cOr
4168zDyo2eTGtt5VNLSXimEgCnm7/6LpeGJXMrS6MBdDxENvi5hLvZZVbGAr5ZFCWElZL/CvL24i
zbs1mPt8ItwNYLVY5VzCn3nF9Mg3EeH20g1/k/hAGj51xhTYQMEsWtpkeCk6YHxmecxqg9pCLLY1
+exyaUKSjBfY6zvMIBzvaWOFdjgC70tCEbPrWgBgIe2C/0ad+AECfzSBk4Lr2xsQLkTciEDISfg5
ydh2ZlpXAtVY/kqEQLsCCH94XHPcOsRwNLOCwbHuGxg2xFXtvTEqe0+KUl/UWQWKRSEd2z99xUJf
4RB+0ZCMmKEUgpek9R189RBCt8QC8PV5GKBGmQqR59xo/Adik0LIDMisg/GaDlZ2EDeVB45benCk
lGNtHV/zziRsd1umGN9NjCRmLxrvOVW4oH8W2EzUqlwk41nJ/hRCvDUs39n6hj8y+mO3HVWKTGwV
sx0sCDFcuLGUKouA2JI4wiU4u19OoK2RWMLqcyODkrqpoHhJFsmxr8Bcf7+Ebi8vfNzaYk7uJHOj
sAEdeuabr3vDFELBZ16IWfKP/vaskRzKypif6Ie2fx0ubJGRG6EQibjWgkFX40E/4YV1nF54nx4O
DYWr82A9sq+eSzkYmQ5pGTZX1YsFdVocofvup2Jz9uDie/VOXtgn4C5pUF8P96Vs85i3sJv2cUGF
wsmU8HykRnrkQNRQ8fzmRsMk8gPYbCUTFbd2RIG9InRATDLy2bOU3sSVp8ws4vCH1Zdmq/Hyffwj
fli9eBlA1YitS+jCdA2TjBqUuPlX+RTiujCTHs2h4/OSxd7i/QoIwQJdF7QPy7XF4ZBp3C8Sf9hl
4r8NyHBZIYkAIRzczcq/vhru4N11RXdwii3VUnQ4xZiL0/4Cca/jZlaK/kKHxWRl5BMAjhZStFqo
U1EyFYWn0Q78ZTGk7wjpUQyxpIAwv6olBPQeUYN4CsB6octMWjax1moPeN+qYz6JUz2t2czapR8T
82QPVc5rfralLigkmVoOMBLme2t2wTQM1kSEADqqU7OhK/BRtlB6d2mijYiAKtodLEHZoouIEhkM
nR0kylQWldQn2XMhL+otn1rkqhETfJdMLkjhReBx/cY4B2pyxSlB97RYGY6KEc+czGW4m0iQ5Dt/
/lyQMFOqmHWBgpvvhCJXyzuPPcsTThRIVojVznk+ccQWZUTzxIeUT0BjFNtqznggj/tzMauZidOt
ekd57GRyJuaJVdz8ejJpdjSxuihz93rbAY24oBRxdRJdnxHNU+iutBSLlTXTUepb+hIoaTvfTvs0
LcaGvhY1Z2WjPhrj+2m3aAMOM3L/4tjFXuVL+jyrB8jaEpADWTHKuaXoAzqEABhk6WlOq9EcwxEr
H8SCxn1MR/Nxm0nqs0DVxwiTQSRyvJtGuayN8GeM6bCPjgOwYXs9DPCi7oee541W5wZn/CER8N8I
d6GeoC6j86Ijcj632NuA1fBqi1Vx3pjm4bayAEBFQqFqk8errEYWWlxR351rR0pvz183Al0xutie
9YKmenggEH/UEnjxvSuLRE/asUje34Dg/akW/IPPJNFjGFJIxe755fEwU8MrppUsCnuyZrm/JVze
jKloT8h6W4vjWEPI40l00zOcn+5Sj/RJ4/XCvrTyhp8vROifSFpWY5XkXJrgLJXei1vnPpko9slX
SSGlOv4sP2yznxbpXqYz8kxJfvYYg9XoN2iefN2S
`protect end_protected
