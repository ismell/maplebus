`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aZ51O0d+KtGKSavz1Awv/c7ZYyjj3asZjppg5CKu14DJI8ku6S+K53KQWUtoEcZv1hgj/uC6Saq6
Dyq68Z0n4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WdX3+cWn/4z6l2oj8kJE5ESEpA4DP0Mx0mmWyavie/cFz8kHzLl/Qfy3AecGPerCGyHqOxjTHGgO
3iSZtSt60dw670649ZURQUB1e5D4AFED+SLDPUZK5Sw0Xl0ew7bMuTwyooaaO2El0XZeDDWZVCKI
YARDA5WTDfJYYxDul0c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ikaNepJ16Lhc58KeoOscyDqJ9qeE6CQzvUSYvm2KTjXG0oJYuIA44daPbLNY/NLxDa+zo4S70RaZ
MofDwcpSc6tvftFlOcE8Ls2sVj4J7s27d+K6oFnBEyrV3/6LCCopNM0rNbDueGl0rbzJQm2IDKFv
l+eT7aUEo2sA+4PjITEhQzs0p+7HqHmG0LnihStnWziT05db1Kcym7CS73qDHUp9wXYBCoKdpFlX
K8qo9mVpij2F1SDMHdYw9FytzqUqLZ2c6zc2R7BB3sIcSy05zy5knr+HhErpCl+0ZHDHagOl11n7
214omig3GMP1DlreuEs0+Oz+XOkVwf5FS9S01A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YgShRiLn2QNDQ3M/X88wH81YSgWwqJdgvj61P7byKtlszvjW/1Ls/bz+yuF1Tw2enJYB7pyZqPRA
8W7178E1N5UvcOkSHHX9ljee3LjzalD1dfxvEU9J3JYXPmgOx9VC1hDeGtmaFTWTgJCl6MzVV8QL
q2ZAih3XkHZ90+WBcpM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WJUpgYEmimgCKQZWN5HshcITVPkd9NT2vdloof0CVlSYpei/rucu7JmMcTKY1YYs2NQO6TqPdMZc
OTdd3C6F/8jPZpNtSBo6i6NrH/m8slcNpcUBuzFlz17CPLJwoU1hf1sz0BaBO0n4W7TFU3VTecwE
VgwTsVJA9r+zKO2arW5NadMONjQF33Cq7tywrI1T/5CZELQB7oeLfCM+xnjMJZ+TDNQMBv7Q1GoS
mIqb3U/gJmZ5YdRKlFB0XgfJMu9oGFTqAksPcatOVEkouQBbX1yYKtfDYs2IwNqJtSc56gzZbjXn
LlFbftiFAQxmRnLdMHxJB54hIudPFuXG21000Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54480)
`protect data_block
IFWAMX8woG0LhcjIrT4M0Bj9XWm97mHeGUfujx/tPjxezL4iy9FdTVlXFlOgLyodqID4fNr60DFh
biYAcuXL2MM2e8B/sL+mSbO3QCwdSdPGX1kWHhZRoHnUtWwkTiLMzXdg2CVx3tsL6PH3/nhgaYWb
APKS6+568IJ79A9U6vpOGh6oPOvUZT5sjPMOWP3O0tIL3XE3xNzsVFN3k3sVW3g6/x1aUqx7PFZG
qYeeiHDozZ7o0P5i8pKoc3c7KRZFwwYhsNoenM3Ai4II08cm3Jt1fbNWOJBQoKW7jpPWPB3E75Yv
Cn3btp+1s1lnBXW65Omuk91qbTLd7bq2QJWpN1D1HZMIxo8QAdVjzNmQxGwMRpHa6kCcSsuFM1It
trX0vvE+JAqHgPYyy+VCmKh4ZFMbNj7D4Zkh37ugb7NP4BD8Y3yLGBHW+CXkKVDC1ga2exFq6yG4
8LlyFRB2+XmNdaPAlwlVJuEzoTCXLDAyA+7uTl2s+0rPCnut73DypNmNRmt9iK8Y3BRVEf4o1D8S
dio6OUANzdEdwdC7REDVSGEi4MTP7gHtjgKKphJY7uw470iG0Gf+811T7IqH+VZCrgSS7/Fuacu0
VAS5n5sCSZjW0P45mIeEyKbA+yNeY4WlOSiUPboI9ga5UOhKflDdRXRHkoXWuXvv1UE6ojb0mmAh
yuUhPEZUt/ykRkK3+pBciO5CFlg4pYS17IKwg6xkdqNUBefj3zHjAKUk8E5FTU0y7SeLsKeD+j+w
khE+gcu44b5TAr7CqxSj6VMm7lQLupTqNXTi09aNUNYwk7+UXAfeu46TvsV6sbApEhG7OAmFR236
baDPyQPkckjWjfGwQ895skm1ULPxJ0tw2QRUD3TRKfS2LcNe1g83AAtRETharwQbsu9vj4PfGPOb
29CE7gLdeTXdkJHC3WoDPlEAgo80W7s0nyLSJo/D4OG3Taoxe2TFR9+ADiFZ3bjoQYJdKFefpIzG
p0nWI7ztsOkGzCAJjaFPKtsw+8e9Tqr4Ru/N6rz4C7GWC0xY3rhgG2bAUb9fi8BEM2FHIq4NyDHg
rqjUa4xmJu5nrKVtkuRrHOvAoMOpq4y2hDWGmW/3KD2HH+pDt4ieOaoQsFL/TxxZBBPH3NAvD2SW
r7qaQwyN65vdn0Maznsbh9Rvzfq7ZUUZS23g3mxHPgjpLEEnk3sl+mtY2AFDokBzVX3INctoYpTK
0+7IFXatLgJtda5EQeCe6b4mCeugfnl1iifn/opvtT7SdiMOIJvoHm4bR/Ch4pBovo0rtIWtXBII
uMufdPgY+xRbaLMvM4KcsonNrJGQrMNvHQD/H9gOMb4pzffOn0xrU46Ud2DaBk4smeZNYZbXHVav
yNiEzE3J1CSSe5W5I6PCUoi4IPnCs3oyJ/Q+yvOEcjqpwqEpfYo1EJt4tsFfPirHYNxoCygl+MaY
HnqSGszRfvD4lNb4ZkROQMLbeG8uEkZmkzGbd6vId4BjRKyaPuSvuwxpjF/pbvGRlrU4K0RPl9hw
wn3levmTIR8O9MFAQzIZqOzbkZXiMwaNbmcjoCLHVl9/N4zA1WjUnVlvovA5wem5YcwlxGzon4Yr
qwgTCyHJKToUfWQS/+DpTAMkX5MvUzrsL/L2+Hr3/e7OW/JbmKCKlQHYVW7nYc4HRovP+VMxfOGO
3B1gldIEPVML0MW8nq+mB5kczZuT4fP0id3y+7LHtyr9+Zfk90cK37aFdd0bweHs66FE6kl6C0fW
9ruf5NyLcFlaMBG+R09OQhrh6PAMdUgGm70MjHjYU8+IS2zUBiwYZaKkUzSNii/mVc2OFrYfTxpY
TDdrayg0d3mjvxyPFzu0FSH6SLnn5GvKDVbczVcAqiwmDuHwQ/xJ4WaC32xNnHKMNIwkcEhHciez
+EqToObZnveCuh31upiYMw14Pe6W2hFT6L8C+ZKXzd6E4+lpWe7syGVKBJTEQ4sVs4Ky6eoyaVm5
5l03LM0IlJm4lB/USLXiKou9lavWMwv6y8ZyTwDzThc3Av0d2ZaIFJb0dSUWT0qW5A37zA+rO3VE
Iqhog6nuUZQqqnEmJ2jG7al49f+d1Z/vMKYvXRAxgryFc3GV0I7JCs59ADThTvFttIPjwYxWtqNa
tjRM3DhMRLriytdxMf+1pdKqI9QflYgWptP4MaTMQixNXUByi9paVyBz1OD3VNVodT4ijQll1fgd
7s7PPliEGS7OutXwp7LRrfyn4dirkZb3/0Gejek1nIY4TMiI+3ZFrBGNOGJ0wqJriUDS0CGPlgYS
8Kw4b5UjPnP+mMbjSRIXYJRXI0Tj69gjZE7obBsIxb1YhGc7Rpt0Xc2+yW/QBoX/SxIat6VyA/JU
+dflstp4k5NTp7IF2+fDvTAfMLVuiMpWXOPy/rTZEx7X4IKAiS8N8gGjRSAG1oqYK3J6Va9aEkqZ
yniVp4KYl+Jr2WLvpjTcHeTiK749N5Bls/s72Ckejq+pj74VroZt3vfGndOQciSrAdvtWXvzPkiU
15ZYIwj6zHz7frYBf8abYh5xuS0zFqRNJxYmjbE/bqDTe/MSH0eqYkmpqnAxfrXFiwMSk++eaIxR
iJsgpNmM+K05tJdDclNYyi3f1wHpvwcZyQ3d8BfAPk4OBLEJqBbsApqh7S/6olG5a2u3uY/eX5sT
HSF6A12vvGgFymWk+kbZaFJdy9EjNvQ2X+9uzRMc0NR7gXReUHOR1fYwrJHtKJGGhNf1Mwx2ah6a
TJQ3v8kULqpRGhyl4LRetjfgIYcAaaW23KAFf3fxEDuUX6q3NocDNzQt5xNQNRmrFu/ZT7mWRv7j
66dM12PyfxCcVga+o93ePnrscTSIBe0TSse9wTt+OzcL2BVHedgkB5wXDhFgPgIm9eFgRucvQfDG
71YeRWwFJc7WXgThZU/lCljYzvX6SCvmR5oypnVV1fTp9BSFHhtDzHbCdKoXibTwSSzInLhn9tmD
8eK0XBEB6vEVl+eFtXN9Azt3BkAsAqda1Baqbvda0xzLDA8q8LCUmmxS9/BgK9WQEEX1zhSJKlkJ
wtJG79azpbgP1Xwhm0J04GcUZxYoo9/beJY6Jm4/2MjtG3/QCBL1WudXLzcMHKIGU/ZsxUmsbokP
qJQfjKi9HkfW1xPldkZHkXK3mko4zr4onAiMrtTaW0uij09MNFzw1hTUKS+/VpvfGiHU8GpSRa6u
CdZ0+HQjWyFpXMyVCgLsXgN2N9SZ1gyS5KYD4LoRSk8kw3t3bAUPBL6I6OeD/Vkb9x8UImrqPFqP
qoiuVkGA+6X94KesR6JU7OstZC2nl3b3/IygCwKbS500iErBO8pa8fgCdOS2Y7MIukzfxLC4WhUE
vwbVB5+/4XHsXw+jtCKYlsIZtWY3TrdGt8LStkRdn97Uks9jEm4hvuXtheTpl5ERNw9FYt/MEEpd
lYCECzyD7iWuAAuWVpYUojvmQAUTWFIpuo6MvIkNE4QYFrdK5O+PV+AqpxBYn87+cpRya504gFuC
FYe+fVDowNP/chGLiGdbasXIjkPl64ZHvHUEO+CcsDSz5N/y2Tc6gPuLeOTMD8ZxqBC2Y2JXNywx
LuZziQEtevTJv5N71ukJ2CDzbZDu5O0HF8she4tuxpl33DnNFZOFt7px/uP4vCRaGcp1dQLUkOL/
/R6Jhs7VcoFERInkfhcdPiBv1u112gRUPBtLFJIb7AeEOv+gb9yrqY3we8euRCyxAyhr/mc6K2nF
xKEAMBzr8lHDJ7EcBWAw2y0HD70QP6H0LMtVVEQ6Zbp4Io9upXwKRpUhP6zYIWkQ6k2tvZWXdm4H
kHaZpIlPF9SR2qd4azCn1tYtTka8kjuxf+M77r6t6AlFZcd3I0weZeUmQ9PK7ewaE2sgFSAziqyG
3AOf/4iH2nZ+G+RTkv/xHAQLj6KlXQenQP14OyMEnd8KwJT2ICvMX06gzE7vMerV/Y0US0xWwyqy
KWoBiNKXqxbTCJqtNZi9r9KzL/fWiLn0JFGZdh1B5FtUXFrDVZakRGp5IcQUQb7m0WwRqROTYyJM
7yHTmYEbJaHILC/iX+XeHGNip4lyvwYC3GZGftRq/FDKujGmC/F7yeKWiuqjVRzOv8sSbiD7BW8k
M57+FWVtHKiDHgfuUsH5MuvyA4oGy6EZVPAyc+aeYXMSW9j396ZQfiHyvs7rOBsJ+ntdUG/TNrZd
fZo8UBHdUEVDrX947Ekwd4IIj3IJr6JekMZy2FShlLn+6oBbko+vY8pnze8HpSMWE4Uz9F9AtyR7
rikjR1y5JLzqbcqy7EHhU92BcYecURIszNwUfxXncQc90bl90Me6J/bRIwQHOEkPAo9vKhybTj+f
o7oJoyKN6qQPlNzy9S3qbDWNu1FhzYjbEJdF9lL7b6HYRMLXxAC/azf31TqCbXZePi6b+voe8v02
ylZM8Ik2WgagP32DqDaUFrhYR0GMNTnmLHmT0GIuC/yD10FX90GnVWEgDluZE2m9qRpF+I0aO6zQ
n5BBaj01wdaC78Ufu0BfGQ696LUMi4RzJmEtqwc3dYNyexiQymDRbAbdGT0dyFF86j8n9CLfABSj
QprLm4KrQaLaNGocw598u7Ni39WD2YgAgQPV4X3fqAXIN6CzH7vv46LGWfB1s8HOoZ49KBOye6bS
D0w4vA1VyUyma+kZQcfuHDYqloFt2ED2n1z0VaaY0LxIDIdwYiq8/3jzemfZ5xjdLF696IB0UoP4
E5foRJWqQ7QZY40CTV09nhK7YePiIHg3apfL+joRy/ZDwod6KmTjtSFmD54BlX4SGSjCStV68rwv
NyB9ik5Lc5cXQcr/0RoVWGj0IBwx5gRijMmZ0pBV/Vr5DRHuu10gw+dPRwX+39zfZ8FajdQAAfmn
+vwowxSW5x5i288GWrlXmqFXazahsUouCWrhQ7vXcBjhwpnz0c5H565FEXjSvNok0bMEa8sk3wBg
FJhMZh7Kfbx6w86rSfaDB7wvNFZ/PPTYc0x5rL/hRfica423Nv4F74DpLU9AZKx3ohdcyC5vgN7r
T3+N8QyCkeVghOp2YTX4ybJh6HJaPIwkMlTwp3eSkzK9/PMxc+kbUBDuvfH8U5Qj5vRlosz9elAI
gYKqvl3yISpO6uvXuxm6/uzBCd1d1sqFzP7aKAXGUZN4YGTgqWSmL3r8klKiS2TlW5ZJRgjI7/jW
rOmn5SUKYEyNSFUzE4qgKMCIRUiQuSPGVNDCyRI6ViqeeNPPQlkdte1pVyYNvKV803lfUz69gzZw
bdpYv0S1W1maFGHEDxvZz89Z2OfshkDjSNm06zJckhg2+NtwZFs5DbZTdYbutF8yC4lL7iZDXRw+
22NE036jxuP8cLtgnr8r68jB+xPX23hfM3LwN6Nh59P2kQuDexU1A09369s8+bmaTwm8mH6EYb9z
cMyLs4TLVU3CGuFR7SX1K5D2MI89H6ib4s9mlWknwyif7LMSGFj/ydbNBPDkx7ploVmZtoFw37q0
QiImiBjbZzxq7HuJfTble5rhhktXHVIbSegOee3/HnMcOsMUAdU0pbFWDxk7eE6vWC0YV5LEq3Wo
O7Fza6EkB5zjvJ+D5pDi7/YC4FIkCLJzruXmoliFL0x64ohQtBuaqjerDviJSEa1deBjgNo6aScH
bxhzNic3ejtkaYvr6F7xwRPGaxkTW6COXjadxor7FQZ2sz0SRTkaSz5UbjTPR3wA1RR30JgZN9hv
DSrPgvUZPuAdl5M6SjqZDkoUW2y+I5xMnEXiJtdSfsrQdne30vCn24lMcm+Ot/VRl7X2y9xdTKir
X5Cw2JF9n4hXWoAhKJMVxDIbP2PW5T8OhklNvIQi8VTrJz/UEAEYgRl40vohtb8kOoJWOXdZ9V8v
lPRp5qQZFTrm1EWr5h0ba99V7doOc8uIy1hFQ+R/4gIX90goswUKTcBQ2YrCsPqz6/0wPsvJm5Js
jKcL2+mHF98DzgmYfI5GTT6Nw0L2y+wmcl60sLEC69B/CHXX53uju4e/p7btu7nzP+mbP4FmsS2S
dD4sAUcAy4aQCbP1ziGL7nE6AxxIVin5nbkI5G54sFtR+vzUpUpvgTjcfj1Kjalwy6IU4+j+Xtjy
XQqRwx392QREmpnQ2eCKPEgcEEf344gJNLAC1JO69VYzry0Y2FAgwKCgJxQL+X3o/aGG4B6jssB8
O8ZnK39oskGAkyF7B3cWgtTkATxjO9Zs4YYN4dzDMCfjyStGlv3qRhTDzU3v3k8dVaG6/8M09ugV
wt96/MikAgKRgU0+AqVrb25isioG0jNEKOXHcF9VgFFDm2unWpPznghD78HuEtuJjbjPnASATQEY
wBFsfUYjpS6soDwExWHrF8xlZFd1U3t68eYGD81aaqRYQi6esjYOOPFmaJvctyt3OPc1Mi15+VuV
dg5WG3xS8JDvdmCbdhOykAAQTl+hBeNpXuPwstxG7hR5AjpudaHROFFXKIVPRxCoHE1Wc3vUQBPC
MKw+cQaaXl8Sf5Qk+ABGexrtz0/1HdoDTR/F8jMguGj4/MkLCzofXJwZGED9bScy1DwHXxgPXDg7
njLan7N7vIiEqIvo9TK7/QIOtpT4htMsMGGxagXZf+B0CbLulrqAhdkpONm37zDB+/dVdR5vzgiU
a3FwU85lLvFz5f/n9yrwUkX2DHEW6ZLGefPZ70G7o/Rsu6W/yoiE+FR27GXpyuaNTW1wYtT3PRkp
A7Oiebjn6k+XS7CcW+gsZZD1piD3MdCrGCi8XsijcVBk0hlWnP/yyG711OnyyjDtJkqXgHEBDaV4
KEbUnMvpdoODPdTV/LdZvhlRz5P2Pk3gOPXB97gZ00SvyKAS+dWprAguZQ+RAXrHKbyrg30oo+RZ
tQ5S8l+9M66MCggWiPd6IXih83wd8CJdB5TJTFf+tgbMdz7xX8IxTpSPCyODvskDiav3AeQKo3s5
bRpqwpAmb7i9UrV/T+gKe9nddNzIkVW78XGCC3/4CiOvdkQjcmK5uXF4UMj7jGrUgBotC25Qgoc4
ERpaM0ecVpBAKPqbtB6A92TTNt5grxXkWfHBpq5XjVn/6251WFPDfzzBnV9JtkigQSa9hpMdyxxu
wVj1T0gQelgtWssG/X1ans5hxXd2p6mO67DBSzdolLxgS01qy10m//PyHvRdw7jYtSlDKzdtl2R/
v4InRmB6HOePzsP8G6TcrWY9XxB9JVqIGFwhzPKGN3V2E9Pw2iu08mH0bnjbUbJie375rT5Eq6vP
pXJ7JjiVFM3qLOUAjlYtUzcVpcm9aIDZgJs9HBSbAcQtbyZHzG3cWN7ERxNg8FUqqMateDtgJ8N6
T/O02xg4Sn7VRl1+aR+O0fvi9DREQmBGjfavqyH314kjFcynfB6b0JumxJInomQPIpxorSSoFpnR
GaKCysLeakoCV0tj0xcfUcqPjwxC26i5D9ciYT60LdnUpGNsHUV1bUDW5Mw5TBP6qpBb/zQWI8EH
Z7K76atWCHDrIurG9HYs2VsSgrj/ldwixFYCtW+aQZ9x9oFRGe2v+jJl9B7AxzO0h6rUYghhndmp
sTGK6x/VghuuuK/m9Xxq1WCRBe+wjZbZNKWOrBTDZbIH28Eo5RYOIxkdOw8jyRYA8hWaB79ZVLwS
b/+TaWUCNBvFBg0T4ss0/iWckfHjiHBvOwfbtOqnljNLOwAuwufnP53cTAlVBelABeCVnGtVjtv/
ciJTcDGJnp2d6XnD35hWgCjRhXDpUwCik876oF+jHWhrPLPFjHhHXRctrbDD0xTBW3OU/WTH9o1K
9TOX6US8gaT0hgmE1B/OenkJ3N9UXAG7a5dwsmKAQkNUZ0QeEyKqtsOV66ew7AWtUdyGKL2yfAYO
Jm7UbBi5S717TvwYSc1nyJbWuh3apNA2nUO4B2HYcTVnea+Q+N5TjsV9zXIWg6QyuHuJu684mkZr
VZ63TU3sONpJzbbXJvsLFxOCdQ8TosaVhiI5n9gzuqm3L0hKdbaP2XTCs64ZKPMAHW1jFzzaoxLk
/dTWA7fuAm3M0BluxyFQ9pEhTZgMVuZ+cl6Q0M8gxwEgrFh6soEknXVHsDDuA3b+AlaQUWmorzeQ
ekUoJ436CQm2W1Vs04j7GZQBd+4NXPsoeA4dPixGmvz7Tomn1fnq5T7Ae4O5MKYt2sQ6YCdn58Bb
kFTM0ll/BdFeuSbpmY+UZXKJe1pV+dqH7gjNEW8ZFOLgO01yUDeKrUHdK7Zf0p30LMT3V3DxoOeC
UgY0gfgNDKHJGjzy0QoMXnXIQsBSgDlRU4p3GtFF+/CutKLCkUS5p6GvSUqZiEyUmXBB0K9706an
jDwC5EFr/qm1dT4rG9W2AVZOmcfvwYk1jQcByEsDtGav6DfmxBHw+S6OvPLuOBuJvjJynidCpPHD
pnGLNb+iH7l9GP4nSS3lPLon8PZ1nFYrTdhfkIERNQzhzW1XLHD9vSyWAaIor5SauWXEX0TCpy+G
nCOhU/WLfuw2c8D1yaW8xflDdlMdeYwoqLQvJJsawIR5BFR+NT7OTsblc7PILBh9tCyKCnjbfLgP
0RKlrd6fJX94vNWMP9UWqkWGPEVdHrlK+/+xaseiNzHXYfznp1dO9JPtH5uJSqj362a+2T60HhPe
mRw5HstCFKYpHpLBZkxJH4bct3tVhURl4njXqqo0pHyVpPrFPisIli+zdHkzSUqBPYR/TMvSZjWj
GecBBu8fJi/7HQqLQjthnIuutGdQIUG40AFoaaAEcQm6G/IQX731nFen76z42czJfSYehqlBPesf
Me/rhZbeHYAdIVLauhwpkTGrwOmx0VTAeVWKnTM3KZejz+ShXJYRrjTPGo+9KAa/kVlg73IrP98c
DOwDj65h8FWkhX01Tkkxuju7RvCjgUdtTDmUwDP8DI0fN+tcCus7lqmIwB2+jszbWgauswN1/Zf5
DGPBr7bP2fFISWa87K1M4dNz7YIfsdZgck4uK5PRmfmLmquwiPM/8mWm2GiZy7gTBltGQ5WwpcWB
E3+AN9wMMDFfuVj4XEb+8QgfW/T5JN4yv61XVrlUpovH9Z6TyZvl3jh+TZRP7ELI+TaiI5YsXc7b
n1LR33DIGg2h81epm93JGRVQdjg90sJgIdsKDcMjmxgeUJp944kCZud+Ey3aM91pHFM6U9ruDC1Q
qAoY7KMSPOJzcGebUkRgLm+XxRAJ3OIQofcYJzhvpKXzHQXQo4d0HmF1Pv5ZCqUUoQuwlp8Fz+sO
FJ77VDVLB+e2Z4NohHrRoc7n38xwEdJORKcV+ZPzfb6yg/gwgCsVWjC6TGUqmtuFgwtMCWjsILSO
kM18oj7zhuM2cuWBT7XG1El/9K8TXgx3bfgFq+a4Asp3Islro6dR2UPui3/CaMds1IKMWAAeIbKm
xW27TFZEWpNPrF0vQnwYKOpEFiVm23ZE/xEAZQBCGwyIF6q1yiSvDZHVcjzC39lmtj9u9WfWKJGT
uIs2sDbEpMlW/Np5RKfTfebdaE9zIJc2mM2b6ntTKQxXndwQm38Y2N2ibKecHR2KHsuPEwlAJrBy
smRFFUYUiSlEsc29/2YSzcVnHAx6tNDSgPVktP9307d1p69xv/Olt1Co+xVhmDVKbLpqAkF9rxVE
ZueJzK9gc1tvt0CEa2olmEOthIhSpt8EvqmagJc0klzDbx8yGLWMDymxiBaN0mWYZ651QeZK+Am1
v/VaxD+VQ9fbQVNt0XMp69/pMpSkdGADvfr2pq/4sgEBwAL1xGSCib4GI8csN1YfuVj5liN68Iu9
RqISZ9xO4uHon2K6DWA1QDz7+EwfSdKjCmpD+4GY8DgT/FGWyz+gn9uJ4l/tsjfOtu+L0FIA5Za7
Dod8Uon/L52BmgW/39keqVFb4n1xIcpHFuWcvnyYrbVNBC/HtL7KOMaXpyodFZUKVz0XkFIyMzDF
XYyTYIowoh+5vjcmLMgolnqAOlTfFeeLBvmmBEERVP0BDWjnIKSd/LrshbMb+XI1fnxM9HOxQDya
AQXOf7sJCXuCYI05F3SSWuwx8bqosyTnGdksgAWwUwbsHheTx4SJpt2aUZQqrMRgRwsDWk6NPxJr
KqGe1akl+D6n13U90TsBafdgI5NpHT8380ldj1HJQDf2BsVkco4SUrXUmm72ZJONYbgbqgQ1iQIl
9yjNyNLhRewcdw+RMsaQq/D/OAFidGyw/o3+xSICJK7/akSq4stcc/LsROV11Va2Bt7BdOAaEBAB
roUoD6IA6jyI4NhJsrDi/catFqZnvXc/+3VJUz2Ay7O+nSNYIMnzydkGwvPv9yJCH0IRNafqqaig
1Rwty5EMJlwp0gCiC54/z3WcZxTjGGMreDDSY2wp1s0sxzRJOR/+HIG8xc7DbhRy/zTqoCbDXwwM
gH5g/5pJv6/hWjOtIE549xbN26EW8iUZwuo/Rrmb80j4NoS/C4elqDPYJgvNUBbeTgGoNFDdBs5P
nBWfg0vePt1NunzCKvzzsZP5GZtYhKH5JdfJHlrft7gdVqA34aboqMl+wlXB7q7VKfIhsuM6Dz6g
tLg5aUt5wwlRm8piUbATYfstaJ3/a3LD6wFB1kqD9tw290O8pSJbIk9XbmNvlAHh0+J98pWGmIQb
OIvfkh1kYHV9+hnE5o3zn5JtIzp30/2DNolKl/nYUgSr+5Fmsp2nssWFDxnjQWuixvHbhwmmLNhV
mHX9GRq1ICPgWcG5OOr90MNvvLoGwJU9/ygJ34spo8z+Nu3z2c40EBUUvPtWX95MDPz9gMzBB1JM
Cl1KrUKWWYlmD2m4PeXwGhgMmoO5P3/yTPXwtw/QiAc9pZaT4vHPoBKNIXw+UIpUM7SDcleGAAjX
zDWBAJjeC5xd2RMfKwLuNHNF4rswCLDQH364FiZLVGFjjQPzrZu/hdkZZ0eS7coCMGLO7tyn0jA9
0fkhhMuzV8CN2sidh7bPp7nrwz4OjAWlAnfBy51/5VFffN8d07aT00ZGvPEurMbtPbQDOnI/6cBw
s/QjrloNOP6/99X7+jw0esiK0FYSHaJoF7o234arSEvO/2E+hhtOWITyw4LzBEBb8HxLE6mOblU3
T1pseGhxR4jOtnniKFWYEpYE8icx11DYhyTpwstTwIRgPZXcWLyht6fio6IcEOcVP585E4KFNzWF
4NeCBpiToqEJOIIOEniFPCcr7M10pY4vmF1wESfpjJO3NzbuJ0QlS14pGdfkkv8FniBKT0tJ+JrV
pSNbY0O2DvnnzilwHFk8eSG3HfNOAeZGDncIxboEUc92yPSwBJQK6mB0NBjKOtJ/P9I4ivRta5x3
SmhdxoOQ8YfOg1+ccj6tpF8nWtukH7nL3vAm00FMisGK6belA6ug2n4OduQA/e5+V8Q2jk08UNLN
QuumDcEwxFCReb2jsK1LrRBwoove+aG2nWlt+4ITzLwjfam5ZCGQ4uXDEDiuaT47asW+wGsVAy6z
zpaWjILjhMslyMxU5CQEgwI8fKGEhiu6F4ZT86tWv2FfbJAtZ2zNhn5YaPSJ9uRpokLpEsOVU0kA
wa9qGmqvNNokUI586tS9J/xhksve8h88PIXpIyV8GQkmse2QL0d8LqfcCHI8WHy6xDwYJOAPN7sI
PXl6h+BPlzE08OXWvTFlyofAxOXniNmIJLgi8tMjSSHDRzXoEzmRT7qWyt22uiEJo0fNFUHrnZsp
2gYznA0UBJfnrn8sal/snc0bbu2RaJH5aV6MBED+TdMHUnjjzDUV1VFtNumq+mptGbxdYm4uMp4N
vk9fxZ5evIl3lI9UjS6josEUCyuhJ0jhIysFFKB1fUDQUfQQFAtv0PzDuCCXCWCIhIOjcNZKcAfe
72gxM9g6fvpC0B61ZE+8CdSYy6UDPbk/Ho9zjDixc8V2czqY3KCEdcwGaVCbPFAsIG+X+rxSwZQg
U9r7onE/Rk7GwLN0a0MfSNdvOuxnufG0G4Io25xyDz65UekEYw9795mDjOw4+jLUqyaOSfmgHq6L
t3t3u4M3XRUGnSMO92vASekSX3xRmmx/xqWk055I/iCZH2GKcHUiwUNDNO3CvqVbEaXC7kCiaxQf
5ZstiKHrg4kwBEFdcfnFYLpJuNagTo1ZJnaMG/+uMKe32Iu8JqkV+m5ItXH1iWIroSz+HYc4x71i
41lVcMQBn5Gtoaq4nPePk8echL92OL9jyx6L2hgebL/Nypj8uxVowROD/GJg0DRl+cRS528gQSEs
++1tTrIYtChQeHzzfMEU7pbzFgS64oNh8BNRirX1ZP9lKJTVN7HMFvsNz/kkkc2flChLHFFh7tXf
uZxgswbCkjvkO3DoZOcNi4ezg04RVFX7NFpIEdrLu6Qzv5SVPEmH6Qyhyi5OF7u5fdWRw9xumQ8s
TRMpX6A5uKORlHpgUpypxMPusKCaw2u7EUhiIPy4UkHwm9d+xmdPi7IhfUQxVcjhLFSpYX79rKpb
bEtUv6wZHkiUh4P4l52tfBpAi4BkQTJbiRMRvr1+YPIIPbqOfA5cDSA5Vz5ZRF9c40wZNdrQxxAv
tLIfRfbI6KtRbc1ZLQqtU1SajIXHxH4iqK5oqiNAw+qgzCYx9+5o25Oe+bctXefCJabhFyLbF/ol
G5Z/KmlwXHPyAGAafqaB4jX692hNE/TnwRlW1f/kNI4ttj9XJ4Iq0BYGjbxpSrF2XNJi4BhfvQc2
1RQh9+yaf5FeB7z/BiFWKJDrCUTNI1Fpn7tkicmIHx0qb7/HonyCulHrOZH6M2585kuks4IiLzdg
KOPBAE/C9QpOlTskrhX/gpa7Idu5Kgcbs5rAifno17ob0RHxOqCSMQpsmdkWApgX65lyJecI1VlD
mPniIglVvKlIbxIzysjsJcco7ANHwVenh7LkIIXhMrC3yDBRyC9wtE6VIh+8WYdfjkraS5U0cjRc
MEDoEouzDqArGvLdoOz20WouL1dd1+h1ZoNLLOAKtVuiX2jEvTH370YnrwQoafuZbjzJjv3ZeuWS
ontXzQqqeSxR70Sj+/cTBqvfpZ+OZhrKsPYt22TPFuFygvg8uQ38nm/0NQqaLR9AfL9R5IhUDlpt
GG4RwsdQ2/F0jmRawJFv3OQ9GD4uUq3tfckfJLNmEe0O7jWsYA+Rl0oDfJBg54ms9KQiEaIt7JZt
mkOv02JxT2AxWc3+UbCuf/cGOZJ/bpyQ5JeYCHxMBuheV41eONM6X3FLKs71jzOGl9u1P8MFe8mA
afc0bpDjIb7xoTo9ez+pXBzUEdMozOyPvH5yvDQaWvZYhQQy/5WPsZN77iP6VUwp/tAY1kK6G98i
6wWrSPxQdAUTXDxX+1qI7jVqnknmDIAmQsCTd8mIa9pwKrxQcxR74Qtc5t7qIFIA/2r9cle8mf3r
71xhvxDe/ZD7BqrEDdFYlGk4SAL6yCrFvPS77FxasZSw8p2KzK8ifjwdC2NRZpRA3HUBx7APQxFN
dwyrqPSvm1ThVdrfVi+pQBTnKLeFzBEKusZOuF/76k5aFeE1Yqrx0GL745gh2I9OFCj5g2Ati9z4
5NjZ/CCFxwJ7/aXlLJtHuUh4d2cDNvnpnsWyMlxLJjom1ht7ER2CI0ihgI41+/iJImT766b1TPHa
nn8FSvhuqH6Xlt5p9ux+eCYrA2nn64PEB89zSe7I0O9VshtoDYIApxOnDGRGa8LKjQ9Y11B7vG0/
Jx5VbmKpulyhQ1OxludkUH/C47Uyzsm02hfALm5EAJnbiZtaMewfyvCDw92jR6ek7isYf2hz5zRX
KDBjByB2xX8OijGMBEdkE5IOaJmG1wXjnlKlb7R1fLZIdepyJL9SiseU+ASvKXt2DrQNIG/SstCy
u4fomnp2f6+vygAqkiX9Huoez485ZzCNPbZnKMow6H1K3CVZgreVhOyxUFdsDa3hMUF9+GrtOSr9
4YMluj29EpPikoVDhDVxMjiukCUI0PF6pEgkeTlHEDrXGXK02/LXE/JWphWlHeam3Iuy7H443TlB
5kGqyxPNhkY8SAYabEk+K3FkZlKFqUCsMVhryvf5Ydi01VMQ5uC0CutczTh1L5QvROSBKvkkrmwl
K4pPwkW74oQZz54HxtTxw7W/tBdXczcnFdOC5nrfMPN2sg1gT6fJIPXKT7pJ3lZhAblpyaYLp0bO
+TFkhBTSmySH3PwI5RkwHgP2E/kM+lzWKt5gHkqqm53BfJTIe1G7KlMF4o3GObfMtJEyu24s2kK7
rE8gszSRaK/DpcEcKbnpdhRv7BDakwFm0/u0VSXX0AQ1WtKU0rsVfmmQYPRc4v/qarC4JUi4b8rb
SLaWpAszuVtZ59nl9ISysl02gh/BWQg/8V4ezxHUXJsOQNSDtl+AhNgAzQSVF9DoxJCz0IWpZFQ4
zTvo+TiseCilr41yxVQ0R8bHgCB83UQs7JFnu0hC7E0UKtc5snEnyI5i5awn6qL6kTijqUtxL3MF
XT6wQ1myL09cWQH4Dzn50jhJrOUwU7BAoU7iVDH3FC+LeX2sHGapcswx5GKDMFBLQwayGYFrSZUJ
rBwBEERSHVumQsTvzA1Cow4E70TRGJWWwkpg9+C3mzJCeYiXB04QPTQlDR7GAeeCRJeb520aenTB
yR5CWLfLgD7Hr7y+T/Nyq9sSDPOVvS6IG737SE6M7+ZK0BpLslBN/Z+8IKa0NBBKhqEnnO+gdjkm
Ik0dKkodNkDVaOlElbutDrLqoJ25Vjun8coh6CKkiGU94491QCYvp+yrkRMF7EfALk5PS9I2L3LS
wJ66606gRZbCWbRIsx6ajc7INXxYdx8l5fWAowpo1NJGLYavJ729HICltyPIXCUj8j+vJKXpfGah
59XGuOv8yzU7VkshIGpKfBA10aZQnMj8gVvmw69MEjhAriAFHWFzHGGC+sNhcSfBGel4CupYYyMc
utWYXEWT7tP09MgylbT/hYibYWHi3gRXrd+OwxJTVXtze+pY7NGK+aGSJk2nJsGpgfYdMjUaTbOI
BUkhrsFIEOK180aRoovwSWmdxUCtq4/mf1Pz75d10uQT2Ac12Osew6nraE7MyC29JJ6JOXDtjDeO
2w2I7f1vc0ZwrZYDWcNR5zc15VUcLWK6dTdnUFQAnGZ0wWwEohyM2FLYnIWYy0H4oGQukF4o4TML
uAAWzUUyg5lybtQOZ9eDZhwoBS9FuJ+hDNw+U+7SAIafqx/RF+dB2Ypt5eZaWxCjge1Q+sVOiwZy
2jyVcdL5wKEiKXAW4zvJv29zf4XbbNjhVYmgV6Qklg6v1ZIm3movOIMpa5SkMRVc3K637tAn0TJs
CDho1TP+i65vlsgLV+BAO7W0HVzNZxDzG+mdRtNvCn5T5O0a/cU7ltGCT27S1CnUoW2MscoV9Xhl
MbvqLcYLj1UYtOhiZ5XByfZQwsHilj0CUuN/dd4SXe055OiDuUiRtPX7xdCg52vL+I7p7l9YXAvI
lqY4FqB8ZeR2LdIOYTcF8apH8f2VJJ11oEuP4iGMMGjwC5qUdPS0kUTnEoMDijySAxGofXGcqbuP
rc/6LSj+j3kv7YhqG5eZAmBXspP+g5Duf1+GmAAwE60DKMbMfMRQduY48eJLxf9drWeTxxH4Z3EN
D4fM/YSyuwhR/dDXZjk5VCjuDYssEIDWtRuVnoIO1W0pInfM3Zqy5pFnQyc9X1LB5omSM4Vhl7GB
WrO+ROJTZKVOfLj8oPGHlUJzjF1CKSbV/q5afj8BpnY+OE3Bf0X6TQ6kMFVPLYgK2SUxihouB4Pm
/4BUomk+0z/OINyVZKkvrcZuEh2WP85TcE1jOs/dC+EHcxvp9XUCfViezcyjyvPY16MjuUzOBMT9
ylLNBeGhO64JGhxsbF2b0Z1YnJUeSLpL698xHHzA5nnbkVDfpu7U1HEa5UbIOfQU+rkAcLLCFJmi
Yns656pdXecOw5n+TtuwQuaKPpAx6iKmDAOODz+7C7IEwhFRgIm4GvNpkTTOxCFJZkgGwTft9eNQ
PhxjGlIMPCxkVgIjwERcCDdgxt1Tzj3GO6f5ONfCvDcYMAV/NM9806H9k7pOwWaWDLv9nk057riF
2T4AS/6Qmp0n6wbrIzS2pdq9m20Ptfp0Jl6FWPnQ/a3W0j8HGqwdpGA7QkEycv6CprIDnGS2WyM/
34Hff2W9wzmlNipm1QZy9gMrzgTgdcJmgLf3D+HM5vsf0nRe6/Q8KDS8oe8YLZ7OTgaNi1qiRP6q
qGr4SFc5C9UlPDpXgHNv+x2pma7USJsfcltzUXx08u5oxiUqtRS8a/xqEmJ7lXPW+9BIdFnGq7Z7
tIRBY5SmlkKXikZ54x1WvGSImfuqrzGMl4RO8SA+fWY5hzlFwwsHjj8x9/1Ii05MYNYXLSt+J/D6
y3rSs7xzerfF7+R7IEqe2xvr3hLxgcnWT/EtHU55My/Er97d0DmuNIwRQhPm/xmRaEVSQvTjHmu8
q6SRpowzsyTweu1su6EDaIp8xMp1HzzvkauOQU/DAxs7KDoXjr9HmVXfj14TbBaO9pqfBFmsZWYs
leEYTLYKmOCgYZpNCvZMwdTQQq4NHgA6O9hkVqsdGBM3pltf7MjHpWIWOdU23eweTM1JxqTl3stm
NxtKmpgDeObmAL/JoTSVnjQTGSRcexEu4X+fq/QNhmopeNNNhsVzRbYt5sK8Ny4rTRjSAuivvUmE
rp9Stgg6mSP4Ep2tLzgHICMiuXV+na9nSRyXUwHpdbbhsziCKUBmUQ8P0GQMGEgcAsP6BxIJXlnv
/y3Fp/vtX113Ee4NmvA+Q0cLR+A74KBZeFpb7i8Qthg3efoCL5xK2oMTBPfjYz1t9QgxWJKLs4is
xrkeoCQ2FRa+RswfKq2S1gtvrXwbng96aRA/I3IqJl7sd347TEQ7WrfznSfUuAsxmmWjopsek3nP
AZPPnCa+k1CUuBSlzmiKiuSIUzwbAYQONx67W3zI9J4GLQxeTB8gsKgs5rMBkZmJ9t0iAb9yJl+0
DqmZgCWDnSJkSkddEnqwjkHaQUMIGZoWCHy++uFFMkFsP4Y6I2+EQfz/dReztafEaJunq4hLY9n2
DObKZDhmAdQCUiK2PF+NLdtWTcbxH98qtBlaWmnI5/eH3K0RbntkbB5AJE3fqXx7Hi/xYndcHctX
c6kKoPXUH3ua2vqbOnpLtoxKsEi/8vnGYBrWyYdrzATMEWHdk4q80XqgEADWuqrjaap5zhpGOOh0
JQuP10C1tLK0FhQmc3LwP+DFtgXTn9OWyoX2hVpHelZrh3S6lPJ/ZwP37tyfUX8nwUeM0ulXMGwS
XqEGtkf+Jdc04Q+L2KeAj/UF1ku9MOFevtv/p8+Yef4SWXbI9bbi6XM/DKJLbTmTd7w9JPETSyJs
806cDaQITwg4rn1WV6h+C8+eyzLrZZ9We1iHyJyGq6lAjFLrPmv5J1MvpJl5Kgw2GbzbpTR07dZP
Fs3VKHk0/DhE7OWypOb3dTQ0DR+p2hRtlBZv0bksYdeuDmAo2vIohH5ZOv5RylwjBpr44sSbX/8o
8Qo6ZgbA5DHGHZiMhS75uHlMMzzYx70Mgi9luuA7VcjSNaLpTJg8Af7XYN6GnxeeB/KSp8utUjm8
GTYK5XQ4GwcBkbEjSK1yUisXK5uhGMROWdoYup4p5oiF1C++IuN+GneYDIyF4n4GR5SWgXLCrkCc
JO3GAK/XZ1dNF5SrOcr4MTZrLRhsNHTknUPRyoFy0X9z++4qeqNYA037IfYI7r3zEQPUK3PZcRXJ
+eo8BAEKR9LesAZkS5Tiy+37bCxvqBO4FZGgQVxH6QGyvtLtn9AI8bepAv4rPVyxh2KNrdIpYPfI
naQSk7yTjrh5QSUHB6wDTrYCNl1t6GusNQsVBkgIHVlNpQ87g0BOWg9W/S1maxgNOd1CQ5ms4PBd
PdmlZiLhvJYMiZDxIRQnsFsK3bjI6RlnJ8xLk3XKgkvjVAO3tkTbVGqQuAd9+zCadpX8Mt093xZt
ugPvPdnickyCz2XSRcU4aq9VLyne0xYqk0NIc1HCkTm7y3mUU5itx5MOArqC7+HpEMtGaP+MCrCs
AnSUqjPrIxzhb6wQijeMWMvyXCtPAOB5bxOujJLd2oGUx5fC3WR/HL4ewuAPK1QmfoPCIAjhpMfs
0NwIBWhiS5ic+LqNjUcM/AXbG0+kp7jo4dpG4zVfMUtbawxAbb5SK5xvMPSjyPxi1vYfzE8NC5Fw
w/Zt88S5Qy3Dnbuc9FK7tynIGMh2VdKA7zwZzAUR4hM/kMQV5BLrmhcYVAQDeP93lcVpY6C28r6y
4ucpWKDxHCDhwQFn+UXyRCOcIpZb+lGlxgU4E26r4YQ0K/uNHiaGzYeJ9IFQPAeW0c10Rob6zYx5
+7+3tvaqeCex3s3g/ONkqbdyOY6dbbW+aHg7RwCUK27tCWtvqS1ztaE6mHSbE4j3hBpd9waIQA+R
Lt+RN7r9vhLhTqdmtZlUCtApNUigM/Jvk/fYT1+AeT8jiY6YiPn1W5TedR22LkAu/7GzzqitfxSr
bN9R0/bgENGVrlkPKry8A3QlJzj1FvllskGb0X5rNuyGXVgmdazKlrCJB26hcfv2hVreJvgTXm8p
1+Mzp/N13EjOfGjy07jUk/IRkdzgJhgQiyN3ta+7epwdxoGdVMDGOdwBGPXDtM7PeqsPv8gW/E2B
kAwTD+gEb6R/l3ZKcdRq3BmaP1lgk2FkMR4N22tYqQJq4DslefrJuIQiPD2kMGGYPpx+wiQQR7ik
aGWm8+isYfzogLStG/6eQlITuwqv2Ibr7vpv68o01hsBCnb3i4Vfov3krvTrqwStVxUWufg3g1d3
yw127wD5YqMwCFavdiDsDKrc4TGSNA+ep25ZidAG6N3es2bbbTUOLjyP4jUHemxBC+5k7Do3W78+
TsuG0GBPe5QJ/9Fe1tcqAMGat7li79hzlT4cn5fmiAVBCt8AWaSxDgpHJJfFnfeT0xebtBcFwyWz
tT//l3OGpTFYV8TGFLGAuzLgWbjXF8yvqHxUmhcF5KGpQ42sSqZqNUTf9KbS9lgMHRijDHhxC/6i
fEVeq+72MRHt0Td4UaFtlrqMsIs7PJ/OzvwnVwc2AOHHRBGKRa+sWnzkCdP/Y+wPR3HC4YQv7oES
VPtPpIeqG75JP2w1KBW1RCWEcn1eeND2kgQeuyGioegN12qY07iNrYKxneDwZAM2FnlQZEbQjpln
cpH1OvoGe94q5D/0Z/ia7gDTbTkOIYd48q4imPL7kCVP9sEBVe58HqceiwAtvzIFU8pcQix9TpJh
yrrEhktVIOsTCTR6/IV888VEk/XpH0aNqVSJIA5M2F7z25G3ZJR4nSaj8NboVMTUawsnaOgpytHq
/bg/awAr4sp+xK9q7okKPMGhpr4S87WIjsinAS7Ih1TR1cj0lpwfgcF+5LjflqsfZipprwVlQUuA
BNociazp7XXpvkGEyYaVZtcrbCLfOecbNSd8dgWZE9AuRVoUT/7XxZcspJL4qApje+/xjv8LZhd5
nHG3nbq7nPAjzOjAogaNHsaiat+8UqQsXiPLIySScbPY0ybZwppe3JvBPSd8fmaNLP154ovm9GSc
0GO8QR7hBzoG0OgYQf8uNklZTm+4Az+eYdEJTOM1gqlI3DlLHIBHVKTZOLpzrwtYaKyVeoANcB3t
eq8mBPhisZqWiiWUKmJxsoN7cXk1pJEDY/NRWw0MiVNzxbZmY/TKMvZJq6x02r+veMUV1SdGYMbm
1NEA37CS106VPJH9uh1cdhK5DrklhJWgXAbDjeJj8e4VCt6118kNEilBxEXM1oi8cSehTz4yBijo
StcZ1pjcBmDEKjYNmHPjXiXVxTFsNyW3NMUt6VF+FBebi2f2ESA5AmWwCO5t/8dCijEJMgmRAiDt
gQdQS5JGH/Yeasxg0Ba9Ba3i9m5RIBE34LpMDLteCZRPGLlFVHAPciaG8i3J9E5M0pchkmbpU8wc
tY3/BKXYDzfekEWdX8FYxX4otw7WGsXeX4mVUTYsq1vnKsajyQvOFdDlT44g0+0A9eGCv5hmVMch
4gehOEvFTuWuFn4VE0Dll9BDkPDC+4SY1xYyDRcdjJwq4mbeVC5oRoGZscVtzu38XRTbxj4cosMP
qQA0cOcsQpe5ROApf4bHJQgy7aHBXmDKHnaIstGxc9Lmd/PGqsiBwNS3eUfVX7FkXl8qHJfmkvPl
buFeMvWVzaUiCzSrLBfCuN37rkVFt2XcFKuNoSSAZko/xQFYGU/Omv2jqCexNJAkEu0xFaoebC5E
M9B1YfZ1d9o6h1W6PXfdD9ueOZrbUSVncHUC6SQ0SyfTwRqsseamx+FhVdCKaVWBeuLoPqnXGhC1
vV6oKkr03srM8ByC14lHsD7wJbrMj3+qAu1DB4ViQyVgAl30KLls6XE8v9Dpd0TTMuAjRzOKLvZy
ldoNd6i5KFgtSp+s/wBiqa7auUEjkJn6PZRtyRWvhU/HOT52IIyXVnJxgw9YUMFlE3Tf7Bgwj2/7
TkoBfLv0ZCcLmp93DCCGuM3suk2R45yo/BiXkJ+/XD8i8DdShi4+34McPF0iRCMKWNLSOKQLIhrH
2u8SPBuQ3qBLYxTL4/P7YOyv5CsbUIsSgusu/khTafhmOL608AEpvqBPFcvLat1RqLR5CpdsOC89
Av8GDtoxjK6w0HaamhhgtJHOlTPpNyT39Beauq0u5NnsTlOQiHlEIlzOL1TfVALC+/lswXeRxML/
CxWlcJ3dfx61pwy221U52K043p0AhJKv8/zzUnoPVDWEI0/3IVyzAeINBJqfMG5G+7Nurtp5m5Km
Wpk1zAyp2M4htw+aqJTssWxXAjxg2YOYZAILSOQj++P8O615hr3zCLDhFmX6HCYvGDayiB5vu+cc
8vjG99+Cntkj7JEUrS2IYHpBiaf2g5eMpak0gCgQ8h/09zekX9wCbYrIMaYtnbHqk3D6wAqobdSZ
gPWlhLrfzDG0Q0ZNWqzrW5PNQ0mqk6Wm1BjsRSeEGrOwWZ/fLNk4wDsIzo1Wv8hmdmDhqtimNyvL
j6pnvaRLM2OuVHQ4/YD+bZOMcUDCvO5VVHAWqo4eB2hk/pkcj/F+7flgmUiQBV3OrfyrgnPzoHAv
gTSSIKYquP3yMYZ68KPpWMh9dSsnqOzXPEUBcl1qtb3b8DKuVP6RTTAqZdaaT841yGEdMqNVcQHw
qMHnnG77gEK96Az8DVcfqYGYf9YRchL0TQM8D4Qik2QXE5ZIr7B8BoBK3MUIQ7DZojNrsQ1Dh35S
3iMl7ILRC0cQX/gyJ+OyyzapAHCi+zqso5NkV+mPlahJck9vzp5czdWcYmurDR0q40wVnnN8QAnd
BNkBabkrZmMPUhiOxSjHSPdXB6w6NxRNrWKNlmHQKGbB3xw/TvPNUwRuAhkTwb277G2PS2X6ths2
nEFbPKV+F1nTihyDvMu78PKEKUZBHGZD2ysiILeyhOtW95LTC3To6VX6pWijXgoXIrYCbS4kVXsG
d/X3z+N2jWyjZyVaRYKFekpNvyDXJIv9skO5XLSUpE8OTXY6g9SDCI+Feg9ZlKmKgBVPodZ+kgDj
dY92mcX1ZVf0KOO6luhbznIhrsHCfNqdXmLi+FsxkSBLDarfmw2oJxgmIdvuOIWwOLK3FPuMZufU
ljwd/aBlHXACfcRPO4AlWTF0ZGWwm8+xm8nbbLicrNaxE8LuRv0mKJ9WaKLIZJpyzM3rMxZpUf/Q
b6AReNkemeIugjCObdPn/TNQxJJBmIMR0vR88Kk9aH6c1SGYTLLRGMfDVy/yn3UenkL6gc0LJo5O
IxAa5Hjrdp9A2IzOb25qFjXCu1P/E+5U4jUSW9fooLdyUMGTGsDPG+Wvrg/9N5GmezyVAZmOdUL8
dCOA1B65IAHMzicotrBhojkPZx6N+AJCFIHwDdDeLJl6rkeGumjG7vXzfG2g7byEZFG4Ht3TPBM4
/O/AZoOZM2774C5KElP7+5z8v7kkGYmOOleTIVxr8NPrkeCRgZxU0+kqLRNmByokQjoZKPVEP1pI
NkO4KFXPenJzm8bvSSE3MEENDNJoHq4dxecoykGNAbdFBkw+7LFx9ru5AuMGDLOz4IvN5hwZ5pbj
pqnVraDQnHoL2capvSjmpO3KBQED6BbMSczBQ/VrN+Ey3QSATl0Vc+31fOL9r3K7TEL7wD5yjXLE
Z2bmyAuNxZ4aA7RUqT8FpdklsZqhIlfqeT69v6rfbbytO8HoAdVc0VkjorpNVe/TS4Xc/9ynw7FW
bldFxFngBPNTsRE7wciCtdvcvl3jzZ3JR6QS0rXOjT8qnUSNXZMZ7fkMnATYzckpYKydBiJJtaPs
wPAz1vGRnkYMG0UoT7Z+HBnDZ4xU+tMA0LBSKxSCxeF6NgpdkxPex5KdHTaL0DArGzrEGCgDdGbZ
UDwadm4H+sNiMFbOvswd72msQ66UE+uMV52GJ4JjhiAnRGyTMJdytKmuNrlObettnmL4kEHbwlwp
4LVZ/n1G7Uc+52rsDuFaH0IqMHJQS1nA7DWf8u2Bm1scXaSutaP2Li9JC2bJjnhcBxxPfM676nlF
r1IhM9PMYZ6ZuTYCSsBPTfy1BcdXQsWK6IoUwF4sifpf94aV4zs8Ne4VWq0zSYQZl+ADba1yJbPe
ZCyW4YaLL8Si6QxlSNiR9CalQkoHZE8VMLi2tRaCwcK72wAhuirY53TpkcqlyiBHe64fGiGHT3/m
HuS/7sJsaJ0UBip5IhRCOl7XcWUpK5dbC1RceC57TVyURL03vcoCYx4nKVOoBuwgMRKe+bZMKwpo
iPeRumYDFbYMWxDyNcNQQgGIKtC/Tj2HOKzrx5RXeiOn4bfpsO3dyqhbUbkZwMfRKBx5/fFE5aHS
lTXIKS/FE2pWWQ8WIHg57/gIOWiDmEAciTpwZ4rCy5tAlT2t0VsxqBw3vg8Kg38PI4ZCyb9byq0c
mbXlDNAngXC21rvKMoQOxp4O/mfQ8FSuWvcrwCydc8sGOV0UBykg1w8K8IxzkDGRB0GnbUPdzCVL
wAMnVONQOEY8Zddn63B/TBcQ1Cc/IaiqFur1henjpLuFQv2cNGyify+Wfga0N+NIjnrBJGvKJzfj
F+RIwUp/F28h4b9uPEu3QZ1ewXRNdKZ3h34ce7wTP81ibxsKBkPi0aYGdhXu+uaxDMYzQUWTpDKc
aUbecMPlePdp6in9hr8o4YScBOYdPEKnA8lrHVFNJCAddJK0moIEAo0xWnyjk24/HfXq8zU6cOY3
f9PfyZP639fzgmWkr68bw9loLqBJ6a91Z2VpBmd0PcpjHREyTSYg6jXJStOK1VwsTjkkZtzH61nG
vRnQRsKZ/zcQFmC8sODV5y9avJCLDUNmoQTCaaf6CRSfuTbHA446nC6D/MgyEavZW/SOUaV//biq
UL+aOhwN7cakp0/UKwEj3m8pWkuc90hiKJl2G7HOiRzlFyL8eVQ68pQTjiEuKYIx3mYET+ljSEGj
oUXSzWfjE6kyxH6+XdOiMWy8pMa4hDHYY32dFXZpnel4Q73tx0pQw2Z1oKUFJ2Nnzx5ZsAeBBhXe
9zyBLD1KIurrh6Z90Y7crpdMWADrsYyrgKmGR+UpAd4lm9agU+DBq9bca26OFDjx9hW2VvXfc2DV
ejLoXczDSBMGTo53KnkEEjd3jLPnVU3Ajbf2Y5Fwb/7v24lIUQcf+Xf5ZNn3+DSb6SIUfzSA+hKF
2W6zUiUrtjcZFXhuq2TdF1X4yi5PK62pQvolJ4iY1+5NBEsCy5Gj824c/QLOa2UfGa3qMyFuq48b
NUeilqbRkNMJV99TznvAbJhOcnb2fqWr++wZpgd5FKfULK0zRw7RQwmUdaU/Vqed70W4/H9c5Imo
wSRACe2GbvZhy2F6HfclE6p4LVqbABxJ0T22wWOVSoUhCAndWTk6PIyREUMQfVpVOkRdNKzeC4Re
TEIgHNvoF3e0SDVRUv4GX1YT5mfZvv8AwiJYIQOLfaKlUq338vRIFrmFnzO2oYsNFU+gpb7tMUX3
vtMr4qVhQzovtLh+Zo7TL4h8gVln2ilPVAosi+2lDoS/DDcl4VStiYB55oc4pz3Jkb2xKdm7m/y7
kwKrKjwlPG6zkPyUPCDvbefYoOxZZXok3fxYSVQF3+OYNX9T/gT0hjF24Ue1PGqmQeFOiiQ+or4E
Bevd9MdXJg7rxW6zmkSr90/U+R8EgBvbrjOl79MYE6UirD+7vwubSoNv42I9l11nalltP2jmR/+R
y7uKf8yCESgRUJxoPSYieXDYShL8nLh1SbMVBZjfC3rbI3zFzU7lpwjuOYwzpttZTB2xREx8dLEA
GeUHrsnt2li24ACPTLRwQyC7g/Hc7qOdyJz26khM30eFNBjH/9r8Asmb/0WSUNX99EfXoAiaTMuX
RvOeUGh4NbHbgXBrvHusjDxNUYpuG3ExNf/7Zx3TJ6DWial3JynhKbHX/9/aejIJsadzzk77Rigj
1jksjaQJ3So+0UwT1JRka7QNRv2yTMnPbcWB0pV3OBnKzIwXTpE8iODl6bEZfdaUYJYnC8s0RPna
9RG4/jcA/V2+gnY+zRzszEITBcq3U0uQ51lQzzkOP+aJDwsspZG02fYmrcG0+2s9HV0aeU2f2PdZ
VWimBeSsnHOgS1AJNpTnYr0woyv2t/E//hBXwHc0i1iznrfGnZ673hBeSyXjHh5I9zoeuWCTJEkK
WzzKsPDyhx/WBBy1C+HaHl9GSDROVTYgP2FqNcwkfwRapAzD5jbDiTzmiWgZ/GH42dmaG8ZPKI62
0PGr3eeaku8TeSw/+kRpkGOruWMIIIm+sh0Ocb2+ZohnJ5xt99w1188XaNiEHlKhDQX2FQeyDavO
rRqYlfKB3TpmKxO9GPv/8UNiC12dDQaCOt1QEXn6JIe8/QQbsyjtU1sUbosmz10kw6G1TBt/vfFA
XAQXJ3/tvR7Lwoacg1idERmybtJ7VI+Y4hl25mVjwhMorN1pISbCSYvlDAAuM05xJSRR/SeWSEj4
+fL/GusQMXrQOEQd1CDTPZCRF8ADz1A1QP8CturwEBdappfdvSnT/TuMt8w4/v9FUaUUOIIg0esn
54QSOhdtfv8f9F1jADNdUKDzB14WP5Qii/nkn05fIegfu+jsAgCirWOPZpxarDaP9X7bAEMEqOPm
P5hImexM8dM1S6gwHzJ3WSN7kBIP1EJW6/vBb1MgNwrT+SEEjPrr/lJ+Cb5utdla5gykHbOStIZA
exR8oS5pp84VUHF3Zv182XRCQSv+RvNlyDDetD3qohXdJ87+CzmAbVUmfAZ0rF2LzifYijWdvV0Y
ScgN1cFDdifr86zfloSejNWTvyUSM2UWOZls+If0jqmNY8wh2ALfmJbNtZhebG1KfuMWCJQX1rq3
vW9zf+vC7wQpDLVpROARyu61k2sxWCQa7ujb6Gysqs15/Sf8cbbQqcOEHAgiu/apBYvrJFfI3s/6
3r0r5HGrXX2cnywnmH7Xwx2vZNK9QxufjGErdpDI3XlAnmstQFLqrfhElWc0r5HItNLqBquxNSnc
NVht04U6vMR9cn6juBYLFWeTWaMsjv2Kfla9z199FFRDBex/MEKHcNvMu87JEEk8jjjlLoV/xKUa
xFipb+bUV3GijnKhThP1P1NWOAbOCL4/FirDnLHyigXFqeOYOUKGlAfO2C3oW1bgyHGvYHSksljF
VcLoqXJBRtIIXD2+5L++lDwbVLfZMsGkLL6LvAnTaZ5mIEEkg9PEbHhrI/6IpVpi/fJxeB03bn72
59gCX0Ite1bNIB6jVNcNwiltiJ1oYCemE/dS8+Vb5jB+NlfXCdnhSHFkYU7lEqFvXBm0roW8zhFo
EKGLA3FuSxic+w4wtZwnR5Liix7xD76MACwvXHwBWBkKkTdWIWkR94FoUpZrBbAi4RapKSCUzKXN
mUbISBpZUPaGvR1wDo73mAS6OUhwlB+2qcNAt6w+PqsTMUQaqaKuEaGuSbOx3EzT0fUIy6tKyJi8
bhbJjd2nvVoxca5kZrMid+epC/7W9ItHR3oDxUZ/zIUeXulbQQgpUnieiklAl8vtgDC2PzGHkMiB
T7do0M+H50X2apG+ZX4YuvCXIlYdf5pqxI/DPLn8zG5K2zWDHcMZxjavDTbR9/596dE59QNoztyn
QqAaODZ9vVLgV3H8xbo9VB0u8DPpjnG0P+wKBX9xnI7U8iIlcIYVkdA8XZEQrAxbhxmn9xf9Hx+B
kLZ2nMFpUj0zyO8/YQkB7ASxSQgvIO8qam4MNnUqywynr9VEYXMXk047u2mBK3ufs4EfOWas/ycZ
Jd0xOVxtz6QN3KyBFY2KE0vpJH6zKJX4i3GR3pMVt1zgC/b73nMPo1S3cv/q2GploG3sbIn78XFJ
TEJajvQXYbtzhtedA1Ma8yHbByWglaoQWSiMw0SuUzHsz3ZO8Qvz2h6SfFkKyfk0mr61XS1Q3Y06
MlYrxEnFWtiZxWmNgsuxYrFBFkb+IUZlXtRXGn2wSzJsPosp+O412Y32UcQjGY2R7/b0oifzc6BQ
0Ov6dxjAcoNiQnYqjwMZBtih3+jEYKFwW5+r7HpLekqM8NxlX9gIGPqld9DlremZWEW1bVLllTsE
dM+PPYmkuadMJyFLb85kp9Zt6InuFIzA4r8SRnPa8WjgyyiT26AXSIwgh2jc6nCLGx9DvsemMVTK
E8PWWJExZOdobrdpHY6B9xIBhci0JEYYgKsW1EjJSdfXX45PitQmIa+kJ5TXOndq+rvwAnyZ3UWa
/ickmWot02mMeQDU/itU39sItCw9KSoImeOVkPFnpOdFaH3jj+myA64F+O9XI3yA6ass02h/TyZK
5H6W3078OvJfFoGvEq3y/dwQhAE65mXw12+io1f+dmzF3WUGUYTkJIuyG0Geafm1XkeRxhowVFyc
ZLcAuAIUf+9wPkv8l1UusCjLAcQZe/OC+DfLvy9Nyn6aU6T8q7g2i5s8ZsrmHeOteNxUpFTWetvy
t7ixS0wNM6zELWaXjNlbQlkNZxcBxYBNw6kjouMLd64Y6TwtqqCbHbwpgCQL4uyCOU5lD2ABmHOh
+dw1LWAufNsj+wScvia9qR55VTEpkwGTyMM+UY/k8ocsEP8xdpKDGENmsI95ga39FGrTVBdV4mfh
9dsbYUzuptnv/GkFe6CpGbm/4dImQDTHfYLsDLb11B1WPlWw7s91eIlbE50oeMBRWJ+KzEFelD5P
Xy/RCa9uJ8UbfwjPT1wXgGOn4pcibOcM+Gb0CNPTCJzEGKUhlY2NvWXXBnnEogSaArxLKwOM8O8M
fGQ45LxIMEscQqJPwIOdUpRRwCLXXnW8ZL2ETvJfF70zpWHfnlsQdaEsWgxj3pMwkfXOeDcuOF44
3iGq3DAb9pQtEhq9Ag2B4bxLQKus76TD5x91O+K2pOZzIhcNh6iV+j1NxNydj/Z5jfS3PdkEqdl8
EvKBsJcQdCnrAdzell9Q8xV0ylC2zzFICqsO93C1/lsPqx05RJ0nrMqvHEcGGfNulqvmrb4TXzwH
azB73C8nwE2kh2BjA1QcSt84Z1nfSLCvi7mIt+urAvKRuee0Af2MXYePo4ns9kcHAmd2ygHUgWYp
DDjDaMgkFykDXwvfxlfvReR8RLndAl6oEMtjFG0nE6fZvGWEbGr0jXUyDzuMdbeSf/2MXiCX+hVG
2zWUoHzu6FdGtt5nEpx9GvLJNhbTPAgQmCVGP8uf7YS1wpYdnrzar4clSAe37cMqNbMjfYV9qCpB
0SH+DkkIjABAJ9Sg+edZ3LvCnnO0VV3LZbnynC/FLC+2WRwT7V2UhYMfqdDPgusJwUy6R4+H3fRQ
F1t0SkQ9G86cKhOyqzvJNz8/eLhCp5Ay4xPkdhnv+LL5GKqbt+a7eIW1cvfags34360FMdo2rpZq
4sy+Nya2WqCgyyWzPKlWUb680RrxWpOadxXzJsPJcNpTh8Gz0BZ9blFycRzlwOG2ZATCKoSqyF/k
EhK4xmbSlMdQb7cF2RSXz9k3Ip+gtOW74XRroAgWjmjVg7hfGZtZycu/miveUHABvoUTHkmcLbHp
ePZd3SATQQNs+76AzB/pdHuYixCmPx0TpyGoI3kB37FxzYR/RGRgvGMyRiS9D3LoKHIxzptHxlxM
i21u6GpEcBdDMDr8Tb5Inxmc1hQZRGpmhiKyNcRixz/fPiryWTWe1wbvZaRTQ5wy13zzSxb+YAZX
2D1I3ariCHBy9eXdYSW/f2LCn0ldoyvUDmp/XHH6M0pHthIn/TNWESUkNiB4kIptOWWdcK4ZdAxE
KB6vw1rcQevwUacyj0MeDWc5bFwk5s52lrdNMoS9jD+ioYbkWH8XN9q58il/ZneNhQhcrKGScEeT
6A58F80m81NaJMVadVvoj8BfEYFODIXCslVK2odfUXCvE++jOUFKXXHx9Ds8vwG0QAfzjV28YsZE
VcbKX9yksvnBONAMoPNYSc+a/TKukgnqANDAPb++72qdS2GaJQBD/Bic/m1wEi39PHtNRVwHolSO
nscAunJuJVLxy02YfIvb5A+9l4bAm66dIzDpqGLizVfRPzyU0T3wyO8wvWMO9wfKByHwJ2bNDVFl
CPenU6AeoZ6ORLu5lBTh6dGcGFfBKSmeX1pHot1Qng7V5GmNzT3aiXOf4EoLlsO2zH58vpwZXYU7
vUmpMp+Ll+gOsMblKdJo4z2PZC8geuUa97wUmCPtgeV6fdEtVx28X1YuS80m0qpfhcfQpv1RqE7S
0IfiKQ0WOxOZSVvs7Efh9zlkASTt7bXbs9543lQVIXlYcyEJlrpYff0UQspZ3VIVamibvmDWKaAx
fHYimrQUyhFhLHmlCWTlzByCYZ3UHvPiR3M6Z1KCv3W59xJ4apXsCpLM3USbfRoZYbVC27/TqBUG
BbRmSGFbfHZ2fX6d8YASwmIyFlRwM6USShUynaaxasQI3duye2X2wskk12pBraoJiQnCwQDeNdxR
O5H8vKfNSmWBNkUzuKjCKTSNvx2B/lo0VaojmalURmonjP6gR8jgPCmuFwk4ASzYO3+V4MDgkFBU
bzY1NgUbThI/d3QXDO0SAd73V/PgcpDWxTklh9mnH14A7q0QYBDAwvbd7ri33Y8RtoCWOFL4tA/S
Kier4xCXGgsWSVRdEHoVYxxO+K2YqfzIKhwIigwRCJMj5aO0uYBdWoMxmA4Y42t7ALnuoIVz8Nas
0EB6XPog56b99mQTbnmvfrPlJxFMgbyXBkBoTmaT+IdtijKzNelL0LaeaL35T2NX/Vtb7VHQhKjb
StrkojMOKpA5zN9eJdgNCjdcyYfKSOOIvEMDdIC9vaT09hROpAAmK6TOg5sxrQXR7sgMwN4ZfO1V
XDGUVIYPfTdXUnZIvHUqQVuXLCxI3Vzi9EAfhsOIjkfSrOEcf1heQtjbOAn+Jim5q9nQIYq/G2OE
NQgiLzd1fGlKoPMjtpYtWVqKs4gLERL4eHfTjOjWOxs+A0NNsGjMnqJIdccaqZs3yCd13jpNzY8h
fNIcuidQX+aT+p1yJWXlxkumIpOKGwyXbEwHhNtvxuR7/Ij1wBWi8IT7KqwGZCYC4Q9pGvpg569g
gaOl1w/v1Qj3ieQzq4rwvp/qgZWqaBAd60FESzny5xbemFMjYMIENtIC13USYmZBsvqcFE27N3IA
+qEW6IhL+d5ynIeycZqBhl6kNYFO5GD9RAzkDCztcSZKQbZVISG0nBBtiyJOb1WMNqpTG2jPtsam
ob3g/PS8Q+85BSGYRfdjUfAJLf6XkvL+fLzulBvMdOzTDT8xdVRpdwPIWCRuwROyjrDka3A+fPEm
uw/yuDTiwCuCDbZ/haKILyEbdxqyv84bLbdaswq2ATNLm1j+Ko9zqejJiPVko0zoGvdESGBzTHA3
YkduP6GzsZjOowJyRDc9VTOoudjU6kNL7ISR1NiBIgS/2I4dFuE8m48BrICtMzhPpOwZ/J2CRRje
A09/wbqLCPFluOaobo+GINXyKk63/ZIIWdTyNaXQ8oD7hIsYSI3iZv3pqAb/bPazSK41JgYk2WRK
M1XJFmyiR6D+I2ga0O4h5rDEn5nZBnUgjOuSdmKqhF426UMXf7g67SwHk6orUNI+/1I1938j0jGA
QTCyWwlUEf3lUm7iOkDhK7myTgFpudV43BD1B1y/2rUtalVr7LAVc2XDDQCYdVRZj9mHI5vxK/rc
AAFWaEJvepSe7ETx+q/VvcHgD2bbbT+FxWfJHg1c8lIpNDX1ulFjAegVwvPIZ+MaFSuz6KjbXpiN
gC0yCF1LheUGHENsiSsZmu+FKEs6RHsAkhKFqXyUATEQcVPP3hamdSq6w8nckNwGR+RqN/X71rFe
tXBbQdiirEUMKpZ7fO3kkFz4CS2fh9rpatgAqRyfbnqbAeFt/Ex3mRLQI9RYslYG5X1Wy5j1ly02
ucmqskBTx8l1bkduTd/4b8V7uOIaev+cVGrhilaVteuisew1TlTGkq4cTfJxXbyPVORaHV5KQ679
EDWo2rg0zAcWQBtzKBY8IiAWaC4AUay9rEuwoEPYyGlSp+FZ3dD0asBXHcdsYLwB5U9yge1SjE5P
NYwdudNn+dI42SXMs6FJRY8GmhUt7DwvijKSFKeagPw9djmxyXdwy2nQAM08p1Zs1xuQrEqF8Du/
3riH5lyU2B7DfXdOn453Ck5VPEx+DXPFr5yUA53aqb8mDXM+cmy3QA6wN1ioAMH/7hFZntfBzJkS
bM2AWdQlOrFlZOGTEC6xu23Zv1YN8HqSfZmNwO9mX8wPNsvASBgyYytkNc3FB2rJcVn9bmvKdPJE
4WqBy4PQr8zUE//lk7KN2ZLz/GeZl+DXTSoG4d7RyDxCfw1BkmnEtYInlbsWqxAHsKLAt0wgXH3O
uScp0xbbDbIP1hDmg1vzjdej6bzc8fG1ltmmvehhsNZHvsUe8S2lm1a3KwGBzMr1Gn2u5XzTGatj
0rYpGQRjF/MpZUaYxOJdp+IrDAbfePs8ImgmV6rCxDGm2+ByXKg5merc9CykLLsvbnRjnWdSJ+Ge
KhiGFL+XUh8jGKzYymiwzWc2XDLse2rHzhskIPC9qnBBwMnfQOESzYFlFMbKfw/RDv4++HksJsJq
z96m3s0BY7KQjI9VZvpR11K65vPVkAwamK4AzgjZUs7Isetzy1WjhedbEQfWI/XI07P+BRcyt8yc
p5ybE7YRiH1feRG1tsEYl2fC9OA+AyEUqrPk3/udLHvd2k7kbDrk6HbHf9RvgPk84dtFa4u1oQ+K
Zp++NjbvC3FYQAOthfGOxb1HPvLvT8MQkMv0jfezAlBx/5PSxGSZFT6jaru4QK3S8okauoTif9Vg
RcXlS75PGTGZT4BcygehIyjBaLcpffZyS3u36UIOjl4O/qhSXs9EaVAK9SsVdhE11ezqIB/Qosnw
gUOzpRQn7ZZlSOqfkJa1DKXNc2535o3/+wGjbjvXERx+dfF8JGdM1JgV1j1qRJxgspzmu7sMiDsz
feNOc30eLEaO9ibuCqTTuv7jZAkAHIT92U6zOj/BygDRlXJqlBrxX26DEjbWpswb5JJyLP6wRo14
OHA3+NJcQy6Y/5m1JtdKC3VcbyyImHh0tgiovGi6MUoxnLMn1HNb+4Awf7po62BMtiAFtLzCjnXo
B7mFG0yWAJ0TVJjOYLzE9TtlyBrMSm9L23CNdzTyRzX/yAaiR42I3HqVNcD1h7wfju8tr/cQ8I/+
h39aRF7+jUvtbWkWA+VzQ/T+X3as7UF5NrO/bsczZfWjH50oi9AiSFJUzZyF//hp/PL1zbemkqa3
rSAzTulvw1CllOIqgWdP9M0JVbuaLWiVXcloaV5YGdrRKyB/DzFAOiQKQBhYULYTQEwQ0a4nG3wk
OPFF3vkAH1Olekc5hn6Bjsz04V7Gq6JI/d9O2g9K9K/4C4WyhKCzPTSbk38Es6QCDFrr+gpFtKZO
Xdn25Zf8oFaFDycbwx6wu/TW24RVIoy+bkTk0c0c+swIgiXgnJra0CX2mAh5zjOE/fV2Vzek8XK6
C4WNc3LCa7pVptApHMb0CVIkiQ1nW51d8QxOsvLloc7JQPrmrtFf2Qrqakmuj8R5Iu46de/4YzGk
QzKw067JeJS7vxy6pw426ZIxQW/Ok1ky5vEaKobV89Gwcy6AgpFBGTtqI7ffHuii9Im3G+wipI8J
rJmqsrfy7SPgjUGeMJGGqGbu3LkZWVZJUTwGgmJD928fYzDxksTpaoWEaM3g0VcEzD23MGb78MWa
5fOrcYmqXkR1xZHxaENboH+FO+QuKQebnuu1SzgyftKqSMOwYeHrIOk8n9irM0RlA8uTk2q6cP5m
m2J4s0O83t9b0aGy8G/BZfnlbBD/uqR4xjbKJNL/MQ+YLet9e3TQSUhw4ktDtZvoz6DAH0mM0Tmw
NU8Qb5InRy/ep5ZDlBSSAlnTryNO6MXoEbAj499N7IlM/f3AxSiLi6X9WkDh6OBIob1iIw8KOViR
KQgWRObjqAqQY9dvAMLP4s4YpLAAC2D9EdN7pUORW1CiRz+06GrIrWN+OjdCEpwPAslmZ4vRaRWZ
aehOlNezrT8jQUl9F4Nb4voQvOuuxDNePhEO27SQRtiLG9fOafHTBjhSQpnIFKR1nYkateEzk9QP
eUJ7TbJ20j664sSqMvRU/geWgANcfu0jCJYI7cG83XmIOvHfhRiQHV3QuRFOdn68kS3KKeapElIh
0tDHTi8eMOm8I3Vgofcm1qHKEJqnguVOsWV7A5YuEUHYZQSjcQKPNNPQ+6OiPzhvVm3flz0aHLcQ
l+sbydu+oUofJfEJzxCQ0SJJ/VYBBdzzMfbBFziYulX57tOJC24DBzxcvJ/doYN27lPkBbaCF4Vf
HRcmCn/Cq5TIp3QWY9Ai3ydnTLGrPkYrzMwk6aPigyPK4VkNkTfZDyIjEZtbkKQuB8W80YNEAKTY
7q5oHyJJva3sEwFkJrdiI1BlfnMhGxgpQwCATka7+yUR0xiVJHmxj1Q/XWp+G4gQjwm6OJQkzNiL
Okh1ChfoNKrdRoT9V11clv3oOTQPU506kQUrAAAUMbKF3SYw+1Y7vY4AZn0KKXyWJIL1Q1Y3pKqP
QZpQTDvqdE2x9X+PI2xyLECLt+cLHWoAaG3J5pHBrM2Ri9Clixqlw/SvYEvHztwUY93xu0gSH4cL
dTjyRg6Vg7KIkL4jQ2FmpZ1LpU1p59kZNit+b0ioO3sSJgWBlW8PVg/rdR0vwsn+Du3JttADIbNd
oDjwgbUQenAd3/2RnZLvwGaMivRevlR7GvAbi+YK1FUxI5iwq/DN6IQv4UGErFw5oZrRGtkL4Mr/
RfkYIEWwVK78XRgqoRwG+QsErIuNsal6zzetQ/vzIB0UmaDHcnJREWk3bR13MdazSxQz/zKmqZR0
vOmNq4/CCL7glrwegS7h8XWf3jsBoGKgftBuilWWIhgIIs14JC+1U6wPEVpC0GQSKq5zsEJuUuLw
4AVxlibShmOTJeCx3Rin5XLTCnhUAGxcwtToDeFFeobUI1BNhzcDaDGtfCF0TGGA3+TwjLYqu6Op
8RbROZyuFbCqAbJ57olD+KCaNLlMDX/GB2O6sJE/p8Y/G/h4KobqNqIoHkZg8hizuFOBHc91aEVP
/0fuCfi+tKCURhfsMBzMGTh8m6Zb5HjkFPi5ztJUdZIKQy5hus++GQ8cIsCxXza5rLQbbzoDZYdT
GScq23k7rZC1zBFU2qkAd6ba5G0EYNzQFJTkDMIOUpg9i8VUfDuswSUDTBONcwcO7SqNFdrvs7G4
9JFC3LnSY0DTFEkGPT8hYLnFvYf6/9rwTKaWnIPJEdsUs5AcIIrxCPhhXPr8bGn6ninEbhkRV5OH
sdCeez5R46BWgyEFclltPiVpVIqZ6fWRkKZ3i2dKAfVTVttoizxLswZXq21D0cUZxVahNurEHlp5
D0QRW2CDEV8u6zpuCK2ChdWljRdZA2OVIW9ek+Y6LaO+Pmqm73e0GolVM3Pn1PmmHGxVcZ7lhJAN
lxiQMj3qQ7WdNr5IcZB0S7ypjXF5Nw+uEKvEHDRw+hkhe7smHibCmVfbPkROg9uqAGb0PP4YhFbG
i9z/44FD17peCRWidqwEJY2uj394eXBedbsssUpBcbnQbGxV93wqFhtt1+x6azJ+NruwSa9gIXZa
PEzZyybNEmuM0aBEOn9T+sX12A/jE4P2eEsLifu1x30MD7x22KN+C6Y6Tdas6b0ohBLasFo1B4XO
XfR3koGKb2OW93ANjF1p6JO33dS4SfUD4p/DVJCB4T1gSSyurBHrdoN+Q4JLKJRVX4lxdKCATOzv
F+rnvwToeKHj4fac2JYoMLC3GqOoLFb/t473pKzNCovBxeVS5wbu7Jt/gyscOfKavyU2XWcuYEr2
GElYWQXzEguQldFrn+/VXWPd2FkkagL4L0MQepB1kadW22Zbyahxnnssza654lPTuG0iKpUmfA9+
PMVdvM8kz+3KI08zQ6U58TQ4SdpH0SkLDQxS4JfBrC9IKsOHb11jQoDA9AFurU16ssyNVJ7bpIU7
O/foKSmLK0c2Cmox/FCJK11ZTFBxJE3+lriQAzEx148MqO6wK15bpflAIolB/Tt7+tk4BoFzfzqK
Z7W+0Xg+K9Gera5maCvo3efTgMBUu7Mi0rnrFLudejtKfSGofIhpvigwzSpkkYKcjBiqlmKzqCR0
XmSp+H8IaaurrEaY2a2yMGa8/Ed803zB5+bUd0+MwU/ujM8JVsjvxSf28c1pPru5BHwujibYFAez
AGrY3g5rKxWpNW3krQU2jXz2ixSfhqhRbHcT9WuOqe4I5MDN5WUlgLIsY4M3C1bleWxeOijHAH0e
aEeJVFGoEyO3W/IFKGJTv5KwwekFgtjYSr0lvzaAiwesP84TADJ6ek+DYAYquXBBTK2GvaSgNzKz
cY/6ePDJvCTRQuQvOM3r5vZboBYv8mT1wQHPCNU1nVDeT9rSO1iRg3Q5q+yl+SFszW0AK8Fujlkt
0ttEGdf9TuqqV400aC0M+1IDaig04rb6STRYzlKJo1E3z+wvIzmS6eBHX3H1UdW0ZrsKBcDr5S/s
OdFt1PXPPsZ3dCIPLrcbuzxOV8yke5rQaz4JnV52YjfMhNJkrMtfo3FkiJcrBPoVjKH62ccB4D41
vdOTUxFZ39ZeqP0pGHfTHRtzQfKq1EtoGL7Yc1iScnvv6Zl4XUclSIXypK44WJD/xUhThuJs/scS
VmnERZ/xD0ieHpnvdt5oi8qICATyAsKGuf/jHlHZ7B7QpyFAp4ZJ4IN6lYpJ4IPkbQy6w+J1H0qK
JiYLWCesbg233U0pFxopZY/KxOMyAlrKr9e0EUGtPCbu2JUmopV5TFKG7/sN6u9tG1Y2vOt3x1t+
kz41e6fl22eS9q2BguH3pw3Qr7STDMYaEl4lnBobMbuYolaip4h5AFx8UcV2UYUthUiOWNj+gaXy
qTnAqgJQpFXQdA4PXaA0zUwSYihWq+FSgZ/USlVi09ya3ImnamsPMNsvfpXczNUh53J4wn72a318
FjPRaiIxcN0dFBqhJKUGYLno8yGz8ioJa12fUqJF675/cnT1HGA3kuEHb/b+85k3qYwxO8ttfabM
YVzdBnk6+temHzHyaXF5NMl1aB6y7IhWiltMbHNXbfS7HCWY+kAufMIPergp8iqpFFLMChC0Eh1Y
j5s4Zk7IvucDT4O5wh2GdhMtNnuFoEX5VORqc6viDpLp9aXbAUFMGC5vuEeJx3t/p/VZP9wqkVRX
qrPK9Nsllr8ndzqF8gVZuURAUTj3XqHV7CCt3fMaiUqphtbRJiUDTVj+9YZn8Eib6H8qcYLwx+HW
DcuTxykj0L2c1MWDsFrWbD3uHR+725wrBg8+FOs12M5vkaeVLfGRR4kJvFdrItW3uX1ICOkjnBkY
NlIjSOrZZ/Z5myfc6O+WB9nxODF5ZNdEdFRzwb/B702VDGWNW5oIJND4z1iuobz9rfbWip6DXR+R
I12Jm0uzocggdolSXYsSj3opytzvHBeX368OgV3C3+5NA4wKkBz5av/cudm0uudPhlXCqVvV2n8b
SUl5rBXveEAge3Z8IbNU1Y7q583UzdTC5c0ugDS1tywb5qP79oKkAoQQbQ8lYcKlQTilEDe4B/jO
1uop2kT95grRWGUXITaKVYv25b4+/KGfYRTlr6B4Vm4qQNFAhqVE61xhaPjAdDUjWkaffDPzO1iR
yWIbFHMi7akS8M2u3yBYRbSoogMv/6ECKv7HKvS7UW5xmcBUJs+kumMbdcXvJFYoeEM9OiRGSCrf
t5irljKDk0gh/2XeilzCjR5t3ltZlEnqYyRaRKqO06oy+pShMFPhCmrTpZsVLaKXixUGATuLjwrg
0U28J1Ua6N+pk+ZjD3p19QCzAskfuLDrTXqZebQzMkx2SEFOLgv/PT3BRI9HlMa0c0sX3WDrNCR4
j7S7LDvmEXJZCTlOLBLRkGQD2tNReL6/tmpQlQFwGEdRUKif3Amd89QKfNnK5uWNHpGTLW1t9Sk7
NoWwar28LWYZY49qjumvMK2ucOq5lmcG5DwODRAqeDab4rd4NAZHhcKu8l/DP7Pa59pYD0yjuiqa
Q8gy88Z+hgovj3FtWiT3IHP9fuFHugcRY/k+cgP41SBK/xHauwxWLSrOsOf3HGHJqUqeaAnsuMWk
YkFeMHB25hSRkFWn18rDGvAcBGt+PMLLfj43L628aZFfssIixkoMZBEyY2GSKOMaEs2C1Kk4IEU5
+xOY0BbdPZCxAatDQ0DiWXtmUttTLKy1U5zQft8TvH7Lge+Fko6xGmhoXG0Ewpm8VPP6aE1RalWI
aNpltOjq3NYmtZeOhd0wMny6pHDAR76TnUinOPRUve7R4pmc9jPU0pz/1euPzfA9UBFpu5vz5NCl
3OYUNfX1ib44uaMWoEGfnfhdOdvIYKf+Xsm7lJ2hovGeYG/7mkkblV8m8tDnUeFjPqh5USesHUX6
RsYbGEa2GrZfFAR6yFCBkVT67jaMI3s1ihr5p2e4eXXzRj2ucLVMmvleGW9YuvfbNGgGqXyYoTi7
khxJ/cF2/jdKhwrrfKYYo6BgzXCQ68UF8hYCiAk0pLLl+MbXsqTEEHERUpDeYCfhoM+TDa34POIR
wgbR1FFl1borRYDHnqvsHeQNSYEczANeSmVmilnctSoDXNIMCdUJjKw5hEZQLa5alTbXoHLoikaf
NtykHgTS1iatdyGEak+WrMzwDoz4sSn/EPumbKssBri9rOeqF7Z2hvJ7CSg1uJmdlZj6HlrUw8Fp
kx9FPOTmjJ2mwOLuGH3nTELgvdHDguwSWugpjTDFcL+VStzHBZ/Ntvfpaa8UVefom5VqfEAJzZyB
rd66ikudbpE1jGTO/nfSiOt4xYMIVt+XM/lqMpvUB+K+pPEHUaHthjgc/GkYeMgOPMl+I8Dfp2t0
97PuF3HDWpLAJfntjdVZTZPMqv7prwhXei56k3JhB6rZkD661IiNA3X3cdIwIoSvOxiAlE/OSwbT
j0hQPD7o4YVpZgLqDScnYfIOtZmUfrqoYNXYBjKh1Z9qUCeX1ix8JUrKHZged6GzcRJnev1iA1UK
hGPFTlYhFRLOgyULwEEoLzWwApTe2TUYIThBIugXWyH+BS8fqjyu9kitFKtLF2NiJSGwhxvN7cCa
btNsxpBxbUWjFFbN48aQFpKZlNlJvzzve/L2d3iNeMh0s9kV6uvLooBMHs+41V7n6Xfk1qg1akNR
noF9RGudz03PDbee3oLw+halew2c7ghhhoFhV+MSruHGegWQDnBhhhzP9Y312QgJ8GAFuAa1COni
7k9k+IOr9vlrFzd5fOCgoLSjCSlY2KwVj157SKkLvXiuhPKqp7f1Ypro5mZZAa8KSXKitqbNvLvb
ou3WNZrjvNP8q04xyaVoc9ZEK5GChF3L/403hjcg5VkVhaZra7gNstrSECB9NCy8IjvhJXyKLEcP
K0NmakKFpqFb02Zjqs5ZFopP27WJtY1GpLQXq3mz4wdznGoUustLRbmJ18qeF82sVCBpKMYQyvk7
zCF2rZzMNCZPLnPCFz/7GHQK0LcXOxTBNWMzAeOD1/BIywJ/3xrYClga+iK5naeDmDwX2fR9awKd
2688C0D/ccW3ZPLkndT8h67TuYD2l+7gv6ozDiIHKudE1nAuo2ytcXJKFBgad3QN9GokEWhYnUc8
IBbpR30+bSRK311G2jiJOnuU5hfAlswlR2n2RrdisWgFzFane26b71RJzImxuxdmDd7eUiGxZ1t9
GtBwlTOZUZol4j4A0ooph44YBfc+w2fOZjLP05RhsM4yTUgYBFf4pngYU9lAgTNZovb1FEB7X3Zb
qzGAB9txzHQD7s21tyZZKL/FxqTl8KTvv+HlQjH1ENjpMtz96iF8CP2+F931I/ekN32LJ73XF32e
60f6UVZ0Nr4WD3rgpNXRIJj/Oqfj9zNKnZZqEpGWa2o6ODyE0EKVQZCNypajhM+MSIX/ib1wOEH+
EZ+xuD+K5kulclxA7eFBWY6C0c3B+GGHAHwxJMrJN7wQQQnGRctIC46mgEzi4DNZ4CLO2tJlNw9Q
7C4KWI1MmcDwQB6wXtUP/tkUyhYS5ECkFocSacFv/yOZQ7zPkhahyHaM4qPY/JFbhGu7DA+1hbG5
mF+WQEZ5S9OQgr04xW4cBdEZ7NNcXOYv3PdDLUtZ5LaroIggS7dTRGdMdN/PBFLdNxPW5ycUEHjI
rM2zGTJt+OONQYwbxqNGKdFKW9J0AkpoWLf1C566DkliY3vkD9tll8jDcZlZGsJljGcnSmn2s6fe
p0K+D7mtsdldiqY+GONF0iBvUuy2RODYSJE2Bv6iBNZ4kAT3EDCvG38so99ccei8hUDrsvd42vI9
Bn5v2DuAcTtRQ27jsR9xk2B72bsqldFv74l5AKWxm9bhoRTZ6irVy/oQIZtcV2L7Irj7/woZfuMb
umjmn0/8Z1pObvK6bI4nkOEoSuGDZD5q3PzIUl8uzRGRq7yVTNxwkCqaQS2NGa42W+VMzSc/xODZ
bB7N5yurq3dhkxfJ5VUcPtrGL5ozR1tKOetqfIS8AvSgq38NMQdTvbLLQ34KaFmoCJgODEvtNKYb
ihTVdqB25UwCgWXGXF7FehVRIglJZRGaXy0TyS6SmNQLrYC9z7Hrvo1yjcIMf+Ga2TpKjDPS0k/9
CYvanm978Edr0j3PtVQR0vZAikWi8B8X7Uh20WIR7mHmUqoW+Awao/x85aakJhMS4g6vZeiskJrM
lBb3ZuSvK67KE++DlxzATbFkkeLTZw9FST8MHZoTS2yxxXknVYmmCYZ4WKO+dzFwIvNHOrbkW7UA
powP/Kg9fMvEmVHIGpIgTnoemnzFv59znQBptUuNseP6rHUoc+OejSTAcKeEhUy57o8uNDKguSEC
WCFZ1Vk2z+LV13rv4qrRvruGAp2qb9E38r2OLD0lXXYzJ7YEpooesJ+km90d1mqz+fK569Hnu0uC
xhzGRYCg3YNF6W7NhB0lVls4vBZ0JuB2rAB2PYSSTGuwL4fROGxxcibRzgA/vVtXefA/l0PnJcRQ
npiIpmcSuCHJw6MlKlo0RaXuhQszGcSxLz2luV5qAU3srr257vNcTjcttFEDVAWuRZvNaz/1gw4Q
yerMEdsUCR2hAHSUwt0WHdpsQ2iPCKIBmj9MSqB3vyJTpM+dYmM29b1Wg6QTm5PRpt2iq/j5OmnX
yDh+LbrcY6Zb+28lB2eekFeb10Kw5c05HvpVeJxdoJwe/+IOjMirjX893Qgj+3oK2yYfNk6VZB/y
lk74o4EPPYtejNpqw8Hf++d6i3qRo/zwib1PS0Jkz3Sqh8FQcJm2ZKeTEgcaDeZSNAvb1wGmorgu
hIZ5swbgfFrCRqgPjLthFrBlpasYosxefiyrnDPiPdbP3PsLCnBcgkEFabkD+/13Rwo2wsv0H9oT
terBI84UAWctfo6+3WSULVojcoqhMtP3fHnfg+5JqaPAjtheO23EIMRtVylYkXDR6YkV+UCQejFv
+TIgGSuPzbGGYEWnwXkEFY0GLmyWgKj1RdXEXlLftuoD92C5TLfxiJSN704Wsd1V6LmTRbWQoN/F
kvRe4cpN7rbwJpDEbTfvNhh8qO7bUBut7KETtOywhL7rt6Oh5zJgVPdxLUZCMh3UWDbdQOCMvZ67
7hHasAXjkjTn8kEo21Yj3DyHLs6OummW/j+M2QkEoYM/xJnpGHMT1+ZbI1eRpMcHKhkBzTm5K9I4
QHhoW7RmRCnodK0ZcbeMYxKCwxDIW2WJvBptyZROUWqPAMTJNf4khD1vKtxmnK35VAXH5bE5MdV4
leEx8FfQUsaVeknUWEeK47HHYKdKetNl5aK7aH6IDO7X27IlUwqnIK7o0pcMGO5vZe9owpl5gjpI
7XQyNkXlLtKwIQCm+uDcB1sIFolPCtBG/vVd1+FvxpCaufgOarVxKdKE/SpnKhus36IXrsGKK0h0
qLoldxip8TzFM+21xa7X8WhT/YFILIxKjtQ4ejvD14/fXFpf/04Wt62aW5eC5cffKdQm8Q/M5sCm
y7HCxOaKKEAkPXFtCZO+SkGaYcAIx+WgnI5l8bLGsBEDf9lXKulzUpMQyecnDQ1FzuNI+NQIhYOU
cMtkwhVKIlmiISCX4PITRtaVIdWkecL6l0r56MauOc+UFX54Feg7e7/u/IFIA8enjVZ0kQQoNFwv
R7SN5kOagolLloOLsAhoWyFnV0ComOOC0ac5pftWFyWrREgYyVS8wLZEdzLLtg8+ozi/8GmI/eCm
9OZ30olBHKwYeZv0xKrWrlcqH9jrILkzR2WLG7rkeYRIE7li04yqiIdfdN+ZamxTeJsfRr6nklLI
qvfZvL6IcVeglOGJ9z1faRsLj1UpdoaPB3nyyZqHpcPeTAqFWRsgZh81y5OvOhcSSOohWixi6Znr
ODPBi3SbOWaAlqYzIg/Elxo0FYSArz30uX3zAQd3/xpQCmS5IO7BtRMkrpPZVH+WeEYXgkyk97Jk
22fjFYYt5FLDVQ5Oz4X3ZHp298DfBecEmLZY4+oYTAsmnAsGUGOUmvRV4qx7bikw/QmG7ftNPPDB
bPQrYMnv1PLHsi+67jZRm9zh7+yTSj3fRcmBL9O8PUoJaeP1QbN6ka24QM21eV0kNrZpiPUYLLxP
C2JMi6igF6vzzF9rbserax5osYbLvHy3H0LD9a9a/4QzOArWCuY6yMnsgmhI2wMFjhpsd0gaf5R4
edPnuAFyOYBKK51Wud5MelEEba2rJ4HkiVNrBhnh3T3BXBSVWzhpU8agviqa98f8uMXhCKeU+IRL
gEUKQKnmdCFtiCr4fovAac+32dLpVQ0XlJp0AxUvz9+EPJuPEdMIscFlowwD7iAynFxLrgV7kLX7
UHclI7NmGPBr/5YcwwhiL3rI/tZQ/57UL/ZYUVmFCVFSuOx4kG/pacyzUmLJE85KGEbglRRWcPtJ
10jBGmtRp166JiufZzjBImlhg7mWFrbhwoqTWslip9RoR3yeRX7MEKKY/NJyNe7+5aAwGypsqzVQ
nks59x9IJ4POM89ZQaM3M/yzikN6CWZcO8rYEzD1fKp9NvcmzZTzOzp+OyISfesByW6NPBvT4g1D
2B1SrRFsyg1RwNSFfDKlXYNyKaqN1nvwWbfdBdyY93XMzglmada2XjMyoK+UHXhQ6IiMZdLSR2J9
mfQcVMG4MOlYZrEUSURt8mrYC2bDiyprivuDPc5l5uXp2qRChJ91poPA70UD/TEfWMdoZQgU9uIe
zjFfcK6tTLZh1NR2//ppDMndEtuDHgnejdg5HvtjFHT5dR07i8bu5ksPDG/sXIgPopHXxZNTqPHM
vWC18KtiyjNDT5dhFoNxSprpOvPL1ODsAW3lzranjTrgvmpdpvmwobQWuD6JtuNtgHZbnaGm2MwW
3S0O1S8NGgGCIDvZBj45JFWolwk6gAFaChShpslPi76JvTnh5tl8ZVDvnFf5as723FBBcEPYctHO
ZZi7T/C/zUEBWaYIIAZCc7sRqXLtp9KnSx+mKXLHDkSYWj6lTxeDTqjP4fAPu2QYj5UktA3hHjKB
OpjbpCdGQKJiEC8a1eSdGh4N4ns/5xxBvZtF+d4nont4Xd553tV+KwHyAOc5J35YwggddKPXSTyv
tydyrdSm1e2pdDFDpbFYAcdztFW7MqKhtMq/qlJdkCWQRAG3AsifNmBjza/PZGHyJO12O3REKbAp
Y1tvEMa2f/2UVsxG/XQxqaY7q/SGMQveiTQKaDRWnnMcIuYkWegv/tthBAwBnio9hLmymBO3De6K
SVsorkjsmPBPERz/Zi5zRnRBY9EXm4gUppSFJ+eXTcFDe/QyVSo0HCM095X6xJru6FUCQRE8wQvU
KU81pOwSOomblbOr/w58a7Df1ahHIl9/FLOf1r3rKwsoioSNAgiiSJUZJ9yeht2751B7BerjRxMS
AUHnTBZZQVghLf42L/DSol9xMBnGPYnjnz7vERnvvrqkSTIvUR3t6szSGDVVtI/p0g7l3bjDQ9Qv
wynSKxChHGysoA6T2E/DYO+xC6P1s71hqambtt0m9WiiRT0a9Ugel8DZg2SRvl706bVfrT/CBN6A
b0MGNd+uVNQRgtcgRuLL5fJx1QN0/8Z5GEdDCXOSsC38hRCfmeOcG06rp51kKiMjF2tnSt/biaRc
ulnt3A7VFoULFew+T76lzkM9GEvdDLc3cIY8HvU3i1E5j3nOhHZFpfP4UAaT+ME9enoCtY2jL9YF
EOUFqlRkMe2IAHC3681jvPCJ9YITTK5HQgfqIhxHG71CD3InzRGyTbRKz7Ykv7ILSQHb6AHWuVRV
MjaMnsUrjbx49PTZ7hH+KAjaPJ8lcw935PSRqTevKfd8TGb67iRs333S4YKGtr1cN1g5HsoU1vV8
m18ZFHZOxBa7/uOO904Sweo+2vL5vN98IrKh07pG8LC8rzt96B9Jpe4UnOiYtzaNhMDSsVT4+ldd
39yqvlMVsivo9w+0z+VD9XnKUTy+Z2WwG9/YdN5MNzvJj8Ds+iylXKKGzevM776EQTKEa4/pGQRJ
6XwgW9eEEC1pFmYNUwUCXcUy75OGXZR8uvS78hMIcxtOdfzKQSzvhlpYGTotFDI+GtrbOSJrFJn/
u8NaG1i9bROgoouNh0lE8PhTngqm9u0Cp/IvrHUNDkeyjWAVE6qtnaos/Q4c1Il1DgD5ml5WmJiu
M8QyUat9OF2ftj/N+tzTzH0X1mySxxMnKuD6HY7k3UtAGM4YzFjscZjXd0vvr0d70roKVHaYdJAM
HoZgr7crPNGFRYRaRJ4zJ6eQIfG9n+nCKadTJ0YLNbcS0I5SQvtujjxHaQmvgqS5OACavh/69pwu
UO4MQe+l1XZRdBeLaItar+bEv4uPyQx2R3VeJbBHmdzRgeojWMSSt6q4Ttu5MNC/b+ddA8exJ6CG
iE96XvM9rtI/274uHLSfKv92wc0Zo0OKiLm8Mhavjut35Zagxi7RX47ThZVHJxcChNiosHMXgfYg
kyuMg7ihK/bAUB1XBYDQUehemgCEfmORLEGONMFjfLWpe7XOznPUbOjHOYKjIZDRnFCg0t97SFpv
oCa8WxZV2cPH9vpNSOVrgKpS2gBnX4yL8YnfKuLjXdV6Gr/2loMHaDFXwtcG85gphBQzi1BhwenT
KORzAk7VgKbRSXa7qQ8DGonitw+G393h1seHAyUk/gPXbQ0rrevVfh6EYr20RvoK/7qpgx8SUNci
Kb8qKaAOjmpK1AR5YAAKYsXDG1DCKHG29igP0GTNf/zKthJPT2f2+0tYQSbsMPhMxqbX99Ch2fBZ
JPk2Kz/PAy4Be0NpnDlzaaunIjjf3WtzQ+gEoHAIraH5tKEvWwZZPHZfqnAVE9R8AXmyhnrg73mq
Je7UlLRkmmJdBUyQHeuYuD3ZiSyIk3GyULge+EkIivz0r3ewIwVMKRQ6DxQKlf2L6GWBXGyTPnwU
rLfXbiwCCBT1dALH7l24Fdbr49skxM4ZD+7h89i48HXjUcakNusOb4GIvY2hnavjSBTyJDF0Sm/F
+NQz6ct8EFmVPj1c5ho/y+WbObca61TrClaBFvMWwz0FrkDolIOarH/68LTHefy042xGtIowmKVc
vtzCeyogr6LN68GcMPr+1novHUsPYzcIVSr6QUF8lNpStjtdLBVHTQE8/4XRu0PwXRVS+vaeD7Fd
x4XX6N3vxhsTfhGgGIdzqrkdFRGnMFY1dpT6KR8jdzIFe5t9Od4xGKILFoShnNO7dvkLcKOwEaEr
MU0jTmjRMEyUSQPynGjcrBHC1pIJ3HYRz76rECkhKSICukvsbzQa2J8l8Aw3HffT61tyMZrCncMd
+iL9CB/TtXBKNGE8Y/qyzG6ZbMvCazE1trC+fDi1L0wk3uSE49Wl/IkuAI6FCcMDyCWBwIjGfgaU
8KSfR77LT2PqS1JM7i0XP10HYbSIgZiaRCKGiTkjRJZL5htQdOb++/f+grBd2Se1clmN6gUPfWoq
S02dCMGubiL3SNpnPBCDwzLXV5GARTGGjQZlKBXJ1r2YLxp0uUVh7fHZizhsUaPqrQA8GYbjqzxt
RTEIpC8jh9KBGmSMXwvc6FXpTYLV8dVT4JZov8ErbtelD5sDzy69GO2v7Lgi+nN1G6Yj8vFxKcoc
vVJrZWdJRJKybS0KC4SqD/qj2KzQAZBK+nNPY8AxgMHOus0WPbvGppwyZcXbkILugPNd0ZVKsfdJ
1Ax9Uo3/JEiBEnXTcs45D9r8RoaYOUextXPIjFwttVL0PDmv2inV/BOkanBDHralEOj3ntK29nBX
yq7AL4VQJhAslaZANG/ilwyjY259LKmZmmXJVko7fy9bUWECfKgKiYAyh08lgnoGLLZLOdu+pXjq
1RsKQTwLXbbCsrsYHJPcPjKxm748yy8veQRrkbd4lulMlzzUMkFtLFvJlWSoUyfVxbXDnlLyk/ww
nphYJm+AqPylKDlHGpuW87v+xc92/MK/7FmkfWvYr2UP1vDTWniGIEta2+0nlFz4iU1XKLgMAFY1
Y9M6VHjjoc5v+O1BlXBQ0cFKdF8aaondlLEzYL5kGjnaJHVQDTonU4oCzlvEV1crMdfZQiHpS3DG
AgNA09qBA6PPdrWaGhPj4Q373htpJLVs0upYN+exRWZuyxWugJQJ0ivh6bmX6XG/sORPG0oeEeaF
sOTevDCH9Nm0umrW9y7OZnlEPikkKQY1XRwbD0j8ZdJlS0IMhSgNtTAiRstvd330xW5EkuUylsph
JQPQaihjseobvRrdyraTvVcDf+RXY+PyW7Ao7ZLyFD0CDzcaeqG5PGmisCmv6/szJPZq+vk2DXpA
v2+jNrMTcC6lXj0V0NGyBpaE7K2XXoLhSd5AztIMx9eFok2spnxVRepJTdUqPE+gN9fmg3FjvvyI
8aefqXfWTGd5IMXNmvTpvZ1MhjHJ/gaNtLKObg8iathajdj3dBwzXgu92SUEPhWL3F+IwxFPotjt
bx50LyjkRErXCZ7KywVPPHjdqZSydADF0JrEGxaz6rQUVP+sp9qg8+wwb23TthchhGjXtbQeRhV8
mHPFXEGXnlZzaL4DjdKlLqzcZMDO5Jn51XyT0rfdeJyuqfE8XOe1eFjyskpq1FgNe8LLz5YEPG/M
4sY+QtD5MouGa2ELED9xCf9q9MLuLmVPxxlrkixKr8HYjOebWQGN1Z6KblYv/OUy0Q5x0R9FuquX
CJf0pxVlZpK8yudo6DczN2JMZ+1o0jwRiHQefQhQvck+53HZgrUQGeNGmmM7Np1ZebzYAKp99oZ/
3sX5Hwi3U3o7sJode5v0X5HUwfqBKfxOh6nFBRP4WNoF44kNgk6XHhEi5mTA5Nf9G/Fa0iuJeJ2J
3/IzHhvHSegTGmDaIYfFDlcKF/wBRnyaqInK6S4bvevUwOwPq0ig2y07XOcP5XrwEhqyA13Zh02Y
wqorq08OTfDNbZ3P2bf+aGaMeK1cxqShcoz8uEa1A8Om2DQ8kPlnwJb1DkSW8nXi9V3vharz23+W
31nwYeuX60zqUuRVoRGnDsw44VU9yTC+Ey/gRXFQ23EmRJHdD8nZyTGN6T94gAAv4RiXbYoI023u
/T11hRoX3K5zGnHjv2q9SpmK2iRGj/I2Fnh1f7fMF0PwnvwqqbEouGHtnK2Q2xJ11r/ugKZu4DQS
+6l6oWMCvaSMr7q4n01EA5bcp8x4c3S3aEOBvd1eIxMWlxAjGQEbanPC2Ts0Ds0ln0VxhXVXLv6p
Qlp9k5SqnQ7x8aJ0Sa/AxeJWH4jcfaTAiAb0hVuJK6I8FgLQUWPRFbUGpJmuT9QRAAAjE23YQc2U
Zx8h96qw2eBRABO1SGr1HyeYlhg7I9eQo0LQ5o3qtYKSzUFFJkXy+xsCcpodl7ao9Ri8IsdE35Vz
gG45gb6++D9nPpa6HkoYA3qxMoXgMCRcYZIZP4yLu1FKZPJ4Xb+RROHxYp15Tq/M0cNmbXiBB8Ze
nHsSWgDvlsELRjcZiULVGFkEBP1zVxb1y3/4yp/1ALNmohQL2zk0GpClRrVOjCbTthP9SDQWppLT
qHUsojjjdUtfKzKJb8AWKf6v5/pt7JrstZFoGjqFm/msSSRcVVdR99pXpyJ4OweRPcEizq2ZRYu4
JSWWlPtSSzNj/vq8wdr5E/Z+Bsut3i2+cLHlCsFCGA8WfqBy8E5BdPXmLnU/EiEhLA52xm9CYFM8
Oy1Tm10EPo0b2DrgCu6wEmBSaNrAEce82bKeown5nGCKbmhr/Leo5rCnBqRno1gIvO/DezLoBqn0
m0pVxDRt0AdD6x5k5aPpJeV45z5Vc2khBvHioUdiaZM7mneEYopwRwGGzHtxHzVwRBr/GU0RjTdJ
vnh1cKfoXRvA7zzNp86EWX889gPkMQJDuBQRLXFOjCLS8udqfmfb9t+wdSA4hhITxj2yxM+xLzJ2
NlLF815O2+mHinH1wruhw/K+sDe2WX/xnBXzFYg7CN10a33EIOj0PCSX6Xv8r96kNNHUeazjMDXo
tHVDusAirqFWU/UsdbLSHgyxoff7V4uV/SdaHN4LlXApswz3PAN6+YVdb0wHsF05Q6f9pFKnsBHM
B7vkXCWeCJQFnhvoFrXZEfouFkTOEOtys5LvnhtMXwod0h86M+5ZSaxEpEkqpUgfIN5ijd2LVx9K
sqZPG1AHZxv0/bXnrnEyBl+tYGWZO4EsAIriKuwppNh48HSJHvZB8PkmMO74dcJ92RIyY8keOHcN
WOePy6NIlYvbAttxRSOXf8Y8ojVgu2JVgrScO7E0rhO9rNbusmTFpc0vL08Gq5Hl41kt52nMdRkO
R9M0Xd8/2TVzkJY9YxhYo176l9wPOdMeXAzaNqupRYZJGxvS1uFh1zVM8j4BkPtTLE7JTklUE4PM
Sc0ptS1gogroUuHnxYOMY6Wb75Oa/DlnBwJn1qA2OQMfOYZ+4P15HbOHwE9Vg3im6HxBpyc4XZ7o
aQgisPPwxJCeke0dyFAGg2V3cctEVHc4ptcn31in78peRHaILB6FT/QXWtNPNcg4Ae0TPdnPpT6Q
mwWRowHMcWHkueBK9PG4TEcVcHdQr65pnwrZz54LcgQMtknr6rfzfZ08ubrlDFSrce8+ADostJF9
BHfGwaF3TBiPnrc7tu+KW3zQ7wKcGI5oHDKra1dTaQm6plIzu0bB7rA+vOpngAF9D2R00IdHJsWR
JvzBPi35iVlmfobLHLmyehTPWi7t7Pewq6PgZn7mk01GKLUlyWYs1IK0LdxwHBpIK8QVztcJIqFl
jNEOg9ddvVk5zVXQUVhaYvkAYKlaLtA61oE5UOaDtrsox3IT/EkzQELaf4/ACt+O2PU3kcP21yV0
VYCeyd2HKKv5T2WUQielmQUEcckIMj1oo+OB9ChiL035g3epy5tsfXKWunEPqm1WK2/snDCSEYgf
0VxOUBw36gaQMjOi5XUGPzhChj/u+l69RU2MoYqiCX+eBohn1yD1nUvoHQ5+g/uvjW9+2PK0FTmP
AgQPHI8vjKtSM9DEOmLuGJ4poYTBXEpzdUHp1mikaHBpAZf0hiDl/fxta2GYtMxgredabEWPhy03
9EpV3L5Rkp5z+oyIYABtAUemTPdz9e0N6P6PlYabN8tF79wtUOCo1iQzJuTqb9Jdxw+COC1Wqarx
KIIUC21cOhvgPbIlU1LqOuP0lZvIgOpJErVz2kKNvbv7a1gx5SturazYV1SqHz9MSgOJIPxyRazh
k1HQmQB2X2YYCOjy+7a160EQoxSs4JignU6zoGRk0t+2XeAieyjdjp+66GVcRoza48t2l2uuK2K8
r1RN7r1Eqzb19qmfF/+RfbF075FO0+SvouTnUfRPQivq1VWji7tjHmldm6zZrwLYvEELA4Dviqo8
qTLc3sXaL3v3oSgCMOpjMZSp1eE+kiJ1OSDx3YeB6CSZZZPj7H9tmZw4NT7m0enbhJxC14CcGeLI
lZIyFSdbSKZB7nIAwJqA6QwgJeCYIhLOIw82o+Km2/DNe0di2OmDmyROTIBQlIyR1oXD3brCfxQ5
YcHtLXA/Qj0UA0SNrPRbff1lVAXPGvCqZTh4vXgdslKxEsatSIpMG/++n5RCo6se/cznhcrlyXHm
N0RYnwl+kJn67lt+qdVJb43z5FDQdyLSRml6P4YAVCo7+UYh4keTlmzOLLklAsF/o/BETJpGcTD3
y4YIBO5VGDKuSnMdZpDxq3d6cD3KkXc5sZE0JWLkMtS4MiS3fPKG+9EAVgSsc40jQgVwZyP7S0/D
OiGqMaOj2XYpTreCl/Fe4Bwi1QvuSk5GeWfdyIAaTTacJS4rQqrekOPJ35tAumzTO4ghbphu991H
MhvJ1Z+C/qYVqAUYoNJENYRQabl3lP/SbrKT3JHpdAhsoBRHcTLZninJFJbgXLx7tAS1d5XDxJkg
YehlZpPsTstgoU0ddg9g201V1TrnrU2+gfwXA2m7V+SKW6SL2HRZXUUiBdMZwFRPh75FMvzm5On/
lMR5r4JV2v75u8sJ0cS9Rc9cuF7BDqekccbh3h7722r+kp5K4CHdmSZkJDQ+T5avmagEAT++BI6l
w6ERT9sAEAfWq1bJUZ3PyQ+0LGKrE1pXO4kAalGiEad5pi+4tiI99niJeMN/r59UzsNoHIj+eDRl
kRfSdBTPq3o3KiGNLdudOUfkzixO7mH4UrklKcrvqzEfRk+/arkyJVG8jYDfMUHyFNal6e6jfmSI
MoveWmrJv1S1w/GAXBAMv6cn1zjCzUyGrHliI+kdQmziD4BP0nrYAqwxHyjCMkkVx211+P921dpE
/7VwPIYGedQ1+0dAKLDJ/4JmG7ZroWGx0P7R1PtHokQ12Ya3DpulSvI0XK6hWEoZ3hyCmdrOI2qx
h15G0NorlXhoTP+1pMdPmZCoIw5WDC50r4uE1Ir0D3G1WmWF/gyY/1ZwyWu8LRJ1kjTQD1j9GVzy
vwY4AxMfV09uXfAxFkMR2KdMCqhnv0KbjdHoO5zbnb137hcbg9iPdFb4OezbtxYjkjsBuoZB+fH0
0OcG2kJdmwUPm2GYjV5BNj/4y1FOmaeF6NvFghjWXocaKLDPAeJxN4n+EoQYLX/zXd2c99Nn4P5a
277TYc7Z3YsUoJT5ugOm5uSZNz7FOYGjEGKLfF+GfXbmmLXZteAcxVdxAwIN1IZAFTiRnu+eiEt7
3TsxlQnXzH8lzFMOJd3kwAGHj9PsiQl9I/64gHA+p6vcrsAEMLme5nNQKUgJC2t3ZeMGAFChTWkS
oAszxm/TRezLRbHQE31fW0y61vzWPfJcJ41xOTeX+yEDNZmGdYBbn4riNTdZu3Ce8oCXOtSp7Hq0
mZ1Yf/rAA9bmUwnU66ijZIlMmr1X++GxO2POhMmWolFQjOp0nvt6yR4crjqprIq5IDxLtphs5ZJg
Qwxc8O2AYq0s6f3O7e/3qFOO2lkmApxdmBxdqIcrbBrLHcCI6nN/pyWWX4+3WMDHlRzWMvP0nWfN
fNS+TbZ+v8P7Eewl5yKhNGwQzJ4fno2Xd3sQqpYJV2ejszFMUKWcUHfEDEnezXp2kAkmKVbr+0nk
2HSwi7SRi/N+GabLzW8Zv+eAqX/mRfA1jvo7NsCTD8VLKu/j4Na0cHInuyhM/y5Od8xGntcb+Xob
9ofnMFhmmqNX3D9feh3GNKFW9WK/tF3m0KdXSU2lu2r6ykuGKpkF8U1gpe0DlGNK70F7dchZVy9r
rj5wCt2vm3gFQzuyZn0jD/YNCk18GEbIScjuv64mDJlOSohmFMbb3dZLlEqiibOhrxUjIfopyBJz
UE4pwMS5cWobZcq68cf8SjIJw8REZI1e1ihis6rTNGp1vLFhr1JhWLIIvbE4cuW54FyHO7kUoeG0
93VsP3mrpeahAOE50ctsc/dG99+ivcFDi9Qx8/wqSywzGAKXVvu4hHRAn8swteJ0FBwLs8zeLE7o
1D5bvGtOvSGq34OgcRkwtC3HKVV44XcTc/UyxyRj++IyJQ0DGpYdg9ECw9FjdsylNJ9YmFBXA/Xw
zIfRQR8uj194jyhzOA5KT7mSxQT5SJncLY9fkEOHhDJWoY2NApnyZ1G7qQERlccwDyIm4SrZ720W
egN5HabZsiZeeEpLitgZsSTZ6SF4XoaqYBXsTr1pTYK+jeQZVN+04gzBXr6cgd5zrRO1WkuUfX4Q
46IBNHqIE7mtLzGustF/uWJp5SOgyHZ9TqXZRdVB+4CeifjRw4J8QBj36nmexxr7geq/dEzpX6t0
ZWdMcgTCz3N2NdfXdXdYKwrwa40BloVrCPQVDA9K9hDyBDJ0M5aST1sK+mvAfTjC3QBXSRbPpnVZ
rRH839/hBXZNt+03NYFgkRY1FhaL7WwoJlzVXjZcjNDBHpJPXhcigtYV3m4CEX6t0Hff4YOBaq8T
2cZAskYQf3ui8na0F/qD6KxLBzi5b9JSXQ1Lg3CfHGkm9ninqPGMZTU3UDoEptQteaUK+39oA0rC
r/gImPKfa+BR5QCOlvTbHGzAKfu7+tFSsW7LCb+Tdwmv2LiWvTFIHIWn8Yzvn9MvxDZxujbMufbF
ArEM0yD6Ol2CT5GechO1i+b/GvL+BuQGMcKIK6UAa307GCLtt8t3Bt/S+EN9TV3SkSIJuvNP8rgI
yzWHClGvxZrbG838jY20eBe0tcs8zrg/WTuAky/i7qvda8FvnV0MdT5cN3MH2Dart8w23Zzb4oo9
Zu501FrAsvPHz+fYbpeQ07UduXRK1MaId7JLFTz7YBbBv+6HhiSVmwSptPuQIkBDbaGyeVdvgmSz
TZgi+bw4z84NOoRqENILcNjO5zpNyxSFFLThwikIQIL5o3/ioxwfIT6hbfcVFLnFkAx6dLXkVfMH
dOqI95piwom65fTZCaibh//9jSGvPDe8avPo+0y+k56ijO1GL5vh/ByvqpWqeCSSDhri1X5YLtoD
8PtVw0GJJeuZkV6Wy0qdR3sPEvtCBCFZzwTIl2hHrdrDToh3JQmOkGKAKwVtgo3sgG1NMxtkqiKX
95u04mFMTWcNAR0r84RoYQWntdBazFcazUIGBibZeXZNJ0Zt/yH3siry9uEEi9d5A+2C4lmZ4LPN
XRE8LRdhgnSIsXVqa5gw/l9QfA9Xz6orq3PjdqZx5jWOgnuGrRef5bcto3bF3q5nwI5t4xgH9Zje
RUOwf+twN263eZSH/R/6gSWnTQvtO8SGY1N9QyjaZHOMrRRlc9RRjTcswxOMF4AmMEPw9kjcfqZe
c2HfWlW+oILfMozH6rVvhTbfx7LkshJfGAjPvLeZbzo1FgdxvxKh6FH9q0IaKVkHsc4aO2CLw1MT
p+D2z60laC2nD+3+/ANeceKqv5KnxmW4TDwc/TYlh76GqvyG7lbSnnOxNgcNajK4bTKXqhWN+h8z
LgBP31I/hXH0jWpX1ug10HdCi1FOUSkztU6BpQBRtlaXbCSb3xSTtN1HQkw7XW3QI7WCaFHK5ABv
Ft7Wol0Dx9AyGQcvcHT/v0MUpRJp+mWL7SjEVxC5v0ssdZrqz/YmbClyUyXDyNPuGSJn1quDvEI8
XS/T/NXUXyPinRhd0UpmT623nRMX355g/ncV4mc5FRuuENr+M0a+0V1UFLdPTBwAEhwYk/0hTHMj
blwEfp0f2OEz9xwdRlkvdFvDlnF/bvWtWd8qL031drAFEWZZCfKg3NofZCO90ntAZmjo5zoNlGlQ
xQKy9GXalVAz5SBvwA+GVoWq3hTRFhJHG/l1SObsCcdG5L5p9Lz7/ulaxz0sDXV0z5K0Hole3Qj+
zrItec6tz/57ecxlLmCwMYzCx2MtAHIn0nio31NmYfqottjElGqbAc+KZ9VqP8KuS3OZ4v4zf7Jf
xuGIYUq3WNxke+2TH+adg2AjHy/9LmV2tKxo1n99UtOILRu9cYuwGC6Qo2SKANL84s1MhDm/BghC
Oc7BdU/o9N12yMVbP2TdiPLImFgQzEwDOk2cqZDVXsJK9qC3jZrAnZtjyQzrourUErk0zJK5FwBo
OOi89JbxRISL7g43rvgTlXi4Kanqa7dZVFGab9shmncoqb7PF0eCdsQkgqdNl9vaOouvRuiAyTIL
BDHjb21ROeqv0prVuQQ+XMqFhRhYf/7rB/Y42da+eYNnYPvsQFXTxEP2+Ce2qzyPivFyGsxmTD52
253TaM1SG5LTWZaYcFDQaE1j4QQeMs8sHOBHo8k8wqJQJcKTciWvQRe/uJ6El0a/z18OE09MAgoY
oFon0GxqJgr51kDFuOGEkM6KDA5qSTr605q0id2i43wWAI3iYt3pLDJeibGIu1hgRhj04DnyyjFW
h7L/9Q7FyYbxTPTapvqT1Ex/R3lc54AkFTG+yhUANOSknwibN7AcBzkMRL91Fk//jkpaFvwLibJJ
hDsrHiuEbokB90+T+wsFogsino0CQZ8sD6KE/n+bhI34SKWPpjM47Q0/fLSFi5Od28lcxoZI42NO
xvK5UQF19sNI+wcjK1pU6aWwBUC0Gfgc6Jw/XFxy7foGR0y9MRjvP3s53GhKYGAlRrSR2JeWu8hB
CYas66wY01MIuSW7TrzMraCVhYveRbBUcvGZhHXjp4EAp0xiyjVUM55QlASYQGgcTniK+iiiaA6t
8cmo0d6amFKZRyDaHu1vWl7azAuEEdfaZ3pjZTBHz+P3EdyV0biFpP80cRXvc9iWShvH6NtNlfXp
a6CYOqJdQwT9nOFUnN7RWzipd/yzTweT6TDT9NgZt5x4cnUjyxmvB414RKejYocNzJ456v+Uyhb9
+g3OObAolxW/xu67v8ZDIVpGLGEb1QBtH0QEd7xwtYPxbCUGM0PMNbc9ZtzHBnoh722u1kDluYaK
r/xNXZyte/pXMHJmRARycm6GJx8S+T5lXfVzMYuXBTbYwwyDpPoKbyeuVFW5v16ARMulHzEN4mm+
+mvfjnKmm4rqxpy+An0PQm2HDfNaXbZsF733UAgP1ZfssFB2UiYK8NnZWz/oybrNyfIg2FLwERrn
unSpLkcyBV2RP32MEZ1ZigD4sg+XhnlKVXAdSSnPJfp+Mq65mrt2VdD1CG0UzfU4Utgu5Obwv5jE
KgZKy4Ro2NXArgPy+cx7h5ufxpFGBsuDtu4T+M3g7kLxbPS1XZ0IRQfnEm+QyLF9DBFY0ViFhDXt
JMUiBV0/EfWaC/hQ/Et7ATL2/1XppPtXXqNAnSpdcsAHpq74XIzUZn29p1iZJBMUm+JR4llYI1qN
VBHNWH8LxB7M5qWFfDMGFnqfjiJf3ROw+6hk0Ge9Zwmr1V9p3lzcCNRqLPMaK74ryP06rLeCzwoj
Cm5Jbl/FLPXQWvgiu7/7Ccyz3hDEae5l4bi90rVLSEme14RJMYhV/IEbBgmSh1Zj4lZHqTceNUtL
gc6rYm5Egh4Td9jRutSD9b7PlH/gOT3JF1sUuy3pa0nUaYvqnYlPy3MsHgudpZBD+EMjJPcX9q9f
S0g6nuIeJQtuEBqwMBOAHw16pjj7bQ7bNRdo1e7sHvsXpo+TkrT8fe6BJ/wzCxqtST7c0E007pb0
ODOfIerQC026m4ZijfzcwXlEfdVgH8Wl0dUBmHwQw6ML6uSrGUAteV56qJGvVTllLiaLW0uAo1h/
g2Z7EUaqKxIOIbekiq1wggeP08dJM1sEaEMwuCTiXwu3WUBbcPmo7ks/VmX8yopDnDXVJ8S2adhT
8XEMCQmyqpx/0KeRUMCCTRgJkX8OiNefrQWWBNCscFyGEl7qdl44L16NDN6NOdXOiNDC88OiQOFD
Ta+nseOoX5XfeNF5Jd2XE1ca9c9ZJlT2QY+ZQ5GcxrTd9/3rcGKSwlYHGL6lxt130kUYbgRjRfCn
S2mpobz6X/dvI06IbBDGRVXoSr/iMUj++O2ZD+yeHmH60pYTxbycOTzjFjhQ2/L7cqkI3YdaGHCj
XP7EPgP5w6aCjtzLAqiLu/FvCsxjO+AZPAL4S5pGj6yRq2f24d0Bi5SLDza7eAOj1NWS0+M49dTw
+glN3ylCy8scm9a/RF4SRjMUC8nvMPsvWxQ2EA8fo8p79IAhsilEZWbrqtL4ajVeDqOGvWvloJKa
7puQ5m9z06W3EKrs2kN3S94oJXAhC+DGjTdo8YN3i/MofHthctQGBsOQtNAIL8867dXgdOF502YK
WYup4CJk0QXPTKRT+Lh7kjpx38TVLzSFq65ybW404enLF2mgZQ5S779EdutTg53Q4lLz5yM+qNVZ
LTd7cGkBWmfK3Immxku3en9Y9SVraJvWRSlyx7suKNu9XS/msKBmDUAmzkO5CyMW6hZ+mGZ3Gv4b
6oZ+3KX8tCF0bMr2j8CEXNf2VxSjBd0O+TLBpbxLPL4Ku1sar4aDNAd+i/bY1q086FqRJwhfnS8A
zd7MKL2/Tn7DKQWob6RExUHZqrr/9VfQUAlm1IcuAlPMe0DgXT6wg2Gs/12Jaa6XfUA+/oGLaDN7
zZYo6Mn9wyw+6F7kvpsmkkTc2vM1y8rKqq2BSGvoAG5Y0Ijx5rFe2Lv0DrH7cUEypAoOsatbqO/Y
zu4a1DdANkMwKnwhTG0uek83NORDhK6EwliE8wOoEE/kOhIRVNOIVR3g0P52yuWuDcH+1c4HMdM8
HhBSMF9/n14aolegI+upwxwUiNEUwzoBjETgXxsYyIvFDu8sIcxsxyyHAJcPJCB/YeS5rcqPRHJA
5W82awgnNS2vDX2XzfzePNhOyFoMjuNoIT5OLedz8IW8EfGW9Oj0Q5bAu+sEuKjmZsjLIzW6avt4
N9KyIvfu7op1//qlmIgSgVBMao8TK/SjwuuOUpMlKN0dqQYh5evSR9OpLx69xVikqwOToVIW/wgW
4x9OSK2kz/MQLwDDjzZI0QGWxcrUQ8yXb4oRwK5BBpz3pxoWvuDVzMa3rUR8M1pgiWgBFUEYaDPE
OvBRdDTF4A30ofjui644t+ZST6V0CJtCRFrf3cEPkJn9ArEGRvYNjl2xIM7xeFluZdLiFaYt+TfQ
NRqVJU7+CuMsog9/S+ZIM37dxfCRa2+B6D+qFvV7rtSg3WAsEzhFbw/thlBjKO/yCw7qVYgItYqR
MkzLUS9q97by5xVn+z4uCYarREiMjueKVpbPPDAyxTE30/2wPR9axUpksixu0K4x4mqOfKaiCopo
fWsd9/PsLUY9nVUZTGxBoAprQZqv5wFX2tpflFRkL0gMbVsjBwgJR2FCjiW1ahsldMVj9p6+yRLm
9cq28rpnEy9/rt/ClDgRpF8rH/D73B+ZH7C28M2W6p2TRfyH05+H1i3wgelgaBUoBSmBgru4lNB7
P1ToThLVTiHWQVksVjlBLEm4WH05Bqihr7YKHpPBMEq6jhTw6VZ7OLdId6eKGsoULSGwij6rK4Zg
4teGxxmdYS9SvCF/wL1BV/W/aAude2cW1NeCrnCF5lQEcyIlMBTF1YhRdqsl3yUYF+NO58b/HYaF
uz+8R3j5hIK1sWLzZ8qIFY7U6z8ts/dF5PjBSpQ2cv/FNEpGj25eOxIU58mqLLmt691UQBmwxFDn
+1jjTlzakRISIegvTwCgi6sB6RW/r2PC9h5r3ZWsWms+XJPa6N2fUUHQbLLznsy7CZtmsoWsC1/L
NYppt8AHu2YdYllDcyShfcfeUdh5c2wYxfnMiRpqi1ioAQYl7rM/Wmd2/BTg/5yW9aXiuLmaTzZ4
L3qSzv37TBxexcfHp74Fh26EjoCUFMqeX1BylUJJo7gtQQeGjBeI1EjSVrWD+CxSFPWEHybnJi8C
yPHHfkDVWUopILSXuXPLv10PjLsMeCBABmyjsXjlYkUILoyT6Vwck28TAh04tue2OZMsKa/HP2XB
Z66PSn/9U6P63ZvwrGoROBkvnMZfGWgOb+nkuIxXSjW9Pa38ps1s+pdeXeqRvGQA2okPRgmXYTv5
7TVdGCMydhqZTfFTh3uuTs53XqunKSOfaK4uxZKEfv4lcbsVqvI2fuemFQFp/K5zRoxr8qhgi62V
4HUdBPNyEjdul/X+xKk+ivbHDUzwg673TrLODB7Z4dadBF3fR661wTt+GYjn8CscFcK+j6E0teRp
l/miHL25xOMRAJVpKQonRvZcQur0CTdt8SYrj5FrmGzuPkvCOPWqxrrTJmW3mZIeR51r+8UExoTa
nhIMbKJgAhv2KyI8tvEF3ZL39UMGnfqyzcI1geTyvZPRNhiO0EQFHDUXUpvDAnvzwvOOGDb3Aafn
VJ1qcuT4Xcy8mQ+a7pu2ziWxulPNfPCdVVnsjpJkNWvyLMdhNllPtOszyQ83f1WwKniybqvKaRQA
IKtpqpVRRiVBsgHcV46vcwG8sfW5ecdD8jbGbQ6uB7J/+HdBOToFn3PoZxKrsD5uiDlZ8yOjPOYK
qX59YorDw8gsBrp9zfNZo6LePSE1CU9O41nf7UZNBk3xFKmLTLIkvkP0SCw2IOwUQS7NUpSydlYe
pDfU1U7xxrzP5WRdwq9SrvQruOnRRRXyYOm1iMQBJd0oks9Zs5N7n69z9RNg2hl0xLRVLOtjo3ER
jWVFDiFwQpWu0zKT4sdELZF9WRUI2Z14J8RMA86fEJH1VOlm4t/v7PFFwXggXdXEyOU1TlKQPMSH
A3oac0B21cSxsU2LvMjYWN6tQ//T1h7r6Lh5WwcZKjTj27F75AvRuzP4mlkI5AGRrlkvZRwyEwDk
ZPWtsQ3nmiBlwM0+gmZU0k+BzQikWNrw1JeKYAq6b6PmneZxGRFaZV3tbwXNwBzKZwLj9/OgdF3H
/fNpSrky+shnYRXJseNQmQjbUUJsc+m25lL6ZsgYKdd9yCJgdB2Pd4u68Ar3XA0bRNUaszzJsp2F
esh912nVcGVEgniUWn0a9kmVrCfPQ99ZM1j30d7L5J6Eh0lLydeWY5Vp1ZVFCS30bT2s/lsB677g
JjenXjFBO/o9ARVAWfGF/NERMOh5g5KUAaArFKK2K6JAHzU+aGcn4+9APnYzBa/qSUQmpn8DSFPh
N+LWWuEYJ8z6TwIFq3p7uutKjqYKSWFKT4hjiBUQc/CTIrhvPRQU8WpcCPhkQNn11AX2W5zfv/eK
mG/39fRTVG+svtyi0vGA9gqt4YgbAn+FVKRVkVG6AwMNdh1Y8dW3oajxX83Flsm2lYgnA4KjG1e6
AMDVpoolhRRFu/ySFiIkPf8+akBuVjren+8QGSBsQquk9nOMYOZ4DNCOwCzHux43WQJmxsbsa8Kb
ohTqhysqqV9wW0q45ufFxmv1gMUpRI00SWo/Kqnsfq2Lda2FellM7ijMjjuoLfBZHPOA4Cli+H9t
0+ZDsRsaq0+JPmCUySOKw19+3dEnCSQOiAhKSVlXRgvOpxUbr3eyI2CUNfXjZRCr9oF2c5NoWvFt
5Q5JaxEK302ahaHb8a5UFcYvc9z2Vzp9yIMENBERGPadqnyxGDopWM9Mvu7Wat0aDQVXsYDWk3LU
jk4Vd4emaBSQGl+zC7xyVeflpMpK8S5tpwy6yTLqUNzWHRjSqWaR2p5jdDHqC4Z4qQDiRAUdBwd0
udKxzPZYaj8GBbbWvAhmJK6YzADObvODme6bMxYz+FEpKXFugMAqHNeYE2kLZZtHCgskUIbQQOSU
4A6F6ZQxRbRicCdHeN7OtPdnPoOVqIT6aCxtLv4ykUIVTAaXvbR8IwfmYaw4QmHEtO3iFydEtemS
drhpj4jBw9NUfjcE7oL5CfbtkXATljBbjHWQYU6DCEgRfSNXabFmwCO/JQO6GrlwaSx5S4+p3ZTs
Q77fZG9rnJ8hibQN3ZAz/R4C/C4M5XniIcKX14XUzx6h3YRXk+f39iabP9wpYmcV+1eYpgHzdugo
hWo+uGFMlCM/aeuwV2FnSEJmQ47i7wSwt28vj4cWQdGKrqCGKdKHLovOOeChmGXlLSrWYh6KOKPb
i9WYGWTLWzRWG5Mqf8LJq/zPmdx1mNcJQ8vlHmuYnGKsDa8BYmejudFCTkzCbFtcho0AWPgiUjBc
M8l5QM1+mmxB0ogf1iKZhccn1SAW9a1kAR69awt+ldWcbpllqp1vdVjPd1jfV4uDsVSFoKG5hZ4S
TQNoBfBIWeXyOxnQ0JZAdXhgOT/BBN4fghTTAaoKuLys7QoT3zy66VU9FEd0mRI9i+9W6wt4Y6j/
2okkFIxqSRzuBsmsX3ochtd3Oo1eMPcZbsCpvGqff/1eNbby4t/tViTtOFvhoqOzN//K4H8j8sKK
aba7hGVK+e+ohF3A6sr5bebFmUfIYaHEyjDFFhvp4YXJMQ3/5ODHtAfX4xyYIabCDAxRrlYNhI4r
4PW31p1gxAVI5gbkbju9jkVY5Ozapq3ufHbvhxvHjI2nrWIb4L9uw325Hwie4I0s9CXiblfgAm4p
Fm53V8oxCvponBl6hapfCdi+S23sMKsoKjvS7Ovx1nA9fAc9IUkMW9KtWIXBGo64ZFPWgMas7ziA
U9pIpECsWghlZnULGiKXVZGUwt8fYTJ94UpLQPFRwiefIfHVDZrUDj+VpJvStNlJtjqJ845kpJ1x
PEBFUZxW1SFD6leBSgLWXLSg4FZc5Jlm8FNuwTYBKBK+amlnh+DH5Y9c0dHEhMksFRgf1oHrCl3p
dnS9vbAMNRs2uAYlc7fTMd9QO4/ZqlISYrzJAttx71BWoiaPlmXu4WZePEk7dxq9z4Y9pX7USwbg
WM7yFWuhEMk9QscfiQFGutGA094AXf7yTijugOFQJGBIdkd75Mi4nYFyHDqxcViSu5Obt4SHljs2
d8f0ujNoU7FS2oz/13LB8T4dvne+YYlVsUgMrbPfHfvSAenGj5arWAidaiM0Aw4GzMv/wAUXLt6N
AhxpugbgfPI8GExkPCH88dciERWts4xsVgbZPl/7lifsYbKxlQg4u70nU7gNR7LaWtC7nDBNoaqP
ScFUkQW/Iwf3PZbvVPD9y7nhwPpggUZTOYWawaWxmdcf2B+8sXaOOK7mjY30nlHUKIXjQdksT9/z
hJ9pJcksHzyCeDlucVRBWZx7Rk0Ofnxhc4yxGN/xODu0mdSr3/RzFpb918vqzzjzKZk+wa9HS6sG
xF90D993rAYfARwStfMxxAwOwoP4EM4gurVklUzCNVES/zzpPQmnpuSGHnOFRqC2/YyQQO8StWgM
2tPtJXAIclRCwMRzuP9BysnNep4zi0/V8VH9ptGbzz/X1IjOMv/Cs1U5w7SOQOcaDThCHOUXt39b
ngLFepluZPJueAN/M8agXvYd/2LoEZdS/+Qsq/B1u6730oTe1cej4vyd9uvyo3mMzioBjVRqWkp8
W9zy5KM+4BR1D6kLg4cQnoenPCisX7jeRecxYJpRNdXo+6x0bFpc4LJm7Yf7MGV8H0ojol6tX4Fx
A0Ja+2NdXFDv6+5bTnzTrRLZCoaJiDzOW7oDwqm52yFVkqJpH+pJdVA32EPnlEvHDIL+VKxezVkd
IedNXbxrrnHhG6aBfzC2tcQHdSZMr/v7EqYgwqgk6rMQiIqOQyD/478SKaEDpmnOok78R4T+Ba4/
S2oSC5V4/tEE7KABGQvhJyxGM26SwIsXZzeHLniq1vJXvtP1gKn1cO0Kk7PL9XNhnTyPMS6og8qj
LfHH5fQf2FKStfIygKCajp4P7PEbeLVrVk/QbSmNDN66UL82y5EUbGeQU36qR3Sr/22URcoe7KqM
BuVBfhZbhVlEntyp8wbUGY5zFKK3wjhlzKTmrCaMbo1mgXQaUvjlzv1n4GmFbbE3UEodHmWYUKZV
7kJhX8XDirq0Tbje06LoGh6hoZj4r4Pp7e+Sv72sipQ1lhPw0ZLzPcEqVlM8LWNbxVzhS7JfeR6D
k4LyHl7/y6/wS3E07qTmubmnAVxaOd1bZzU4fU4nwyafBqMJZiwYjtx3YfUyAhKQRrNwL3cxd9kJ
kjDNorPb50Rg/3Kodb0o5sxXizXi700nCcsC4IKgVGlbkSgUonkMM6dZCIBzg4ICzLQHnTnlzAKF
bvtpVnUukX/UTYdZzvxLwDxW2MUK4nd5y4AaLivyKve1Du3hDvCdQjewd50dA+y2vXSou4q4ERZj
OPwJEfWe9hzoLMdPRDAm2Tl6TeM0QcbOZUgCwZbpHHAGPVVclFkdp0aRtu2A1OA2XvzfhgEQY4nW
LkkV+t+T9RbVCr9M8qrtk3LR4TKfcqs8lOpoBtz8ooFGYc5tpIVBExyWQxSq2qsWZBxftd1jAFHP
BhgNnXgFLHCsBUpHNtlME3Ieo+mbn06V7fumarEtjF3JJ30a/UFwnLvcqp6FJMapDLc4DeKZglNj
dq0B48jVOovtn6TAJrkAGQzGo2ZszwHqQHZg2rXRnYVWksfO/cmyQgiVE1+AS+tp9bWnyARKJIMA
dRKb43fpsauURFJmY3iBE3H1iE/L8Ucdw00IMLMvNfuV0uMHD5kx+DrO/t+XQjsT5qBuxAxbRerU
Cq8/gKlhf/e9wvVqvYBM2xt6S7fypM5rCTt5VB3qyzm37jEh6ztEm91EMy55HW+6mRuOj5kvG/NG
6CqmXsjTEeyI2SgLvdKhts02RNxJqJpVkR8yYsmZjOeZrIMSiF5IkX4upPD7Cdn+qCywMTA0Qvex
7K4WGH+xbVMSp4H6uzjBKii0N3dRkKT/Q/A/Aa5RhYGQC/qJrR/FTlxAi/P1Zg+8YQhqGsryNDGC
M3Lr5VCniJpHMsailUCMIbBZ4FqYiS2MlRzSWbgGNI/h/3uU8uNNUeYQwwtsFSXicUgV8lldIk25
1dDfrtYNRJGZOHnSws/EhPvqEHjvm4DMYSSPoz+HZHAoY/Hlh/h5d2UhDUQxm41Z49Cq9O/cmYyo
8thxL72CepWkifdoQdS91G2+7iUMBd7Xru6Wlga9d+VoYgve74YsCS7G5lU5bxHximmrIMAX/HAr
ws/OE3l3QD8Iz3H79lBYUk1mQrX9K063vCiWfFutterPyapBw9dHE2doZYQpwt+lNADZwU0AmqTI
eDXSuSQMhhiGVCBRSHAd8/tnW5vueXQ6lYhxEDAQSxqsoIE/aL4CVXvy5fYthsrwVsGDaUBBnX/2
ZRkygjsvQuwHlvEfGHOl1o/JVKMfwNTeP6khr7uTJ/0RAQKRY2atptRlSXcStQVlY8pnFQXGqUOU
aNg8dgOs6T1AA7bNFYFM0jSJsm61SAR5qideOjjRGEE+miS/EI491IyFd4iA43eUxpxiBFdO6NuE
5KfZfq/cvPkcDYu2x28flWu1O0mkwVy5swqoGnvl8TbwDd2Prm+I6lcTY8uQU/IN3cx3AFhSJFq6
BwwA/ftknkro4HL7cj50yPztTsMGTAoEhf6MPAeRRLgBxRcI3prRMkem5ouVn1cDgAg25UkI/Xrp
0y+g9XrlL5jiOq89rTp9bry/GqxpWbhZ3/hjqcvR902vpqhV2d6hx2oXPCj9GDOKi2ibgaIDCNhY
9MhHh8kqGQQfH0ROxNU2s7YykWuu1618x/Z3f/GBwWRFuOCR/i8junvWGcPRUjWPVHGfkkDquIuB
Ya2FORey4t5p/AOxtHigTXocDMIbOl7vPkHgtnRkgigSbktU7vkM3IVcirjV919FSotfTkhflgqu
s0nZ2d4YgLfVndO7TnDltV00cU3OOwTwSdAwAxYdBhmJ4hBu68uuDq9AufFf3hEMdjLva8X3f4uX
woqAtwyQnOdIZLVvS5w37xczGLNDTCxSoBClUIo3V7dKUpIF46MzvQ3kNV9sHk6y3gDRR9526Ld4
4UZyLk2Y9Xv9g4zCqOW5OTQUKG+cRNK1dE0fCMi1j0KjEM/JHxV+DocjbqIqhtkd8dZ4Cp0imvvc
vRwAepdtAuMZu41fSw0ICZG+kfn5P3pNMvLUbTMGklKI97b+S3fXRi5yq26x9KSMZn7N169Zd0zt
E/gPYZaHL7rWt+oXQzBYXb+v0fiamQrrp/4wxhaIvBiLQO7GZw3s0Ofennb3zOXKjTe4v+cLubjb
kMm9TmCKlPou4zq7OxGcm8GTUxNgMUvWuZJZjffrPBX9CK+EQaMje+oL7C53GCK+WMS9b+ubQEkd
1C8h+gjxbJxxERyCb6Fr5uEJ+CaYbxtVk8V1+VpKcdiKlA+ocwi3i0N7/xMUdokUxTaAKBslJz0l
f7TqJYg4S/NYE8Imy9CkztoS7XAHQ9TYuIaA5fSBQ6HNUBoWH4wJioXi49kBqAsJI6jmy/zywh1J
QDykWDxL1Z8sExzVNXQoBsHPTUcn+csStcxbstGKfe/7cZyzsif0CkhZxG+whbDLDNSw8ZjtvBPp
NSPeSDPXsKHXTexiqLmuAPiA8pI6kLgOpJ+FsZQ0SGrNL9GKqolGb0TfcQv09KzrTyc+G2/xLoMp
acpVGN4kShBIu8l1KORlVuZ3pv6vH2FTyO7GYN2xIqJitM4Ch5MMvmvlPVJpHqEEfql99+l1K+nk
yHMGSXuLs7V1ge02a06O5MoCANiV1+yHlzdzbcHyYC/QdpT1t196ifQyMXkXTwMB0lv5BGITi5qH
PgH/c7RszFSpP3+TJ8q6Eh4RXRh4nOl9U7tE4dQVGNb8QXoSPwrCyLDJF3pP8ioFevO19M5NRiPv
Y/nlWsELVoUCLVamtF7EvElTyvl9pzAYsPdtsJNbsvmTj9U8WtbvJsKiS+E2Jy0JpbKvirwcV86h
ha3qWtXSfRy5JeL6/AvUQ40eyFblcX+5XGQwVGFBBYigmu2vI9EQwqVZLJno8NBXexbmJlw4J95B
3hgllGb4NEcr6ySyYz6PkqlDryQkQLEGMVkyHsPinyf9fkewdhtHCWi9m1CpMk6fr2IbzQA/MOuM
V5jxtDeSqGpv6rouIyy9JO+LDlf3kPVgCkxq09FofPwL2xp6DbDnF57NYNZsHWzswVIhiwTA8Xhd
I0R1X7NYvtsDKv1OLU+TzMYWJQUhbVnrpYyDKXKcFANIjLzPNcx8nWOkSC1ANZkHK6MEP0F9b+Ty
GenICUEmzM0pwvLQrvMNiKqrRMiFa3fNfSNahUy9tYKCSmKjIxo8zlgIqhzv9ku4WBKBCrdohdPI
khHmZQng/nqH3IZ7eoLKW/YfwzWbuPbLYq2IwymO/lvaWQ+VsMVwbmrZJRNjYedhHNfcMiBm4i8O
eNkk7uMwpvmWAPGUS5M6/qf9sBJ14yks59+xh7sRcRsdzDEmO/SQj2Q+ycPclJqxxRk/wjs/gODj
ebkMh/FdKRa9mrRK5qyaY6MZPLso+oYesaUuLBMjnTg7oAQMzuFyxib6YEwaY+7W5v8iPRhK3+7z
8IDFMqwOh7NqvS2Lq548Wwku4+YowvBNXZmn8oZA068amOnhlqlgCFb0Nk9DYnTran9pEd3HFXp7
Hmg2MMwv5kUm48CKCY7sjL0uc2pn1NR5hMov077DvXJE5qizf46hpkgLj356TuRs80UErCE5ALQq
cDFOX042ckHenzeIEmY/q6kCpYbRDsFXGoC3nf9F5xiUekXSZsClb15oekv19QeAFyHutJhewg0/
psvewCFxwAUgMTj8KRrwa/zI7kT0MdvZobqQrsRmLnkA42bZsliGU3C66zcgkdpbo+5niBsDq7hH
KJUXiiG0KDxEBPF197miSSupReWhBiIxBeoy9zgX4iH6e0bZzxt3QadFSvuHmX6rMCuOaCyXDqkp
UcQq8BlVW4TlCvcgX66+DXzTxjcU2tio6rfqGuj/RV8OMaDveAdmrHNABEEAjDxXgAG5eSA7XOp1
eMZdUR1PPw+PAW5ZqMrOR2Wj8FvDoAnfLKa/j8ZA4WZkwN1CtEOGBsqGToGEpA08PwVflxTrgr69
Q21SCTwDah/ttf4ov3MChlhWnl1C66Bq0P4BcXNWII8hd+bQuLrXy/sBVWzPHwi/jOJkt76GI2Bj
DpmqFvmvJt93qMQ0pRt6qokw4LMFPVt66x6Eyzrmroi6O3rBIMaCYW1rpsPfJtcGwWSOPcqObifE
scYJX8q8GqIwOFfWJWP9OFOPItjf8/iRPEJOmNKKtQDGqbakas+prGK+LEJdKqqbrD9N6IWnPCq+
aq/XSWaBtpBBP5OgCoJ7RQaijtLDWYc00PwA2tx4GHrI00oO9uw4aqfQXWgMxIt8BwZw1PxU1KSj
SSx7KXmNayONQTfCzZcwZ/XVMUEmD+7bkhVOJttu6CO2ygcWzT2+sEMEwvpHWKoOdZIFJgKI1sj5
dCePrY+4vowgspqihbjtMzZlCFjJB7O8hf/ZxD5e6XojR++jhehq6eNBky22eUeYxwHkkaVV53ml
3VJoWEOMA6JNqkpuR534K/8Yy1TDSb3yvLVWYrzDLJvhdR4UF3qCIqOzQQtqbCWKfQF5yV4ukR5R
1BPIWH2VPYQqtAoK0JjVdiomhlEn5alhJnLCYejpjUQO6K941lI+u9VPEMqOlIqRAHPAkMuDi9tj
VvlUa4scEB+9DVfV8YOC6twQLNQZYZCJAgndW4s1ysHLDBFhUH9hMskFLnaKlwj5z/9mzU8JLfEQ
3WF4KUd0ZAYIKIn6CmnwX9ogdcrFML1+hIc0Cb8tUUFcnHneEAzNDkgSH7bj+axgveY8nhs8yI5H
yDOL24bD6RgqF0bLLeJfZQ/lGqOw17Cp5ldpg2ctTTuNrNtM07AS+aa1I+CMqWolvpw3fi7gSj4K
VAbXb4sIGnv+A6eFc88KhDhngbK3orDEZmUoATCPZiWJZmg8DKIjVTGA9eQFUpPnBAYSS+jfA5/r
lYdQyXuCq0DSRu7LbsyUxb0lPzUpZ8q+ManrBSkwixvI2xOzL/aPOnWdcAmMTVuHQkpgCdkwFObd
0EcCMs3+KLct/w5n3JbrEFIbxqRcT++0rSvctgJZ5ZzMtWYx3S0zaAIwN0UN7F6yvZ1QnpZzGtMx
w/eWRdYZnZoK6RVIyVi3w5tBW64Nh9aEEE2Bo5Q1FpeXyaisL7G4xBu+mMCPwjXrwSb4Dw0XMMfU
EZCGY0XdwM+GsNsN345hemBlzG8E6M33RgbyNeqs0LITkO4SN5hwKuT84QxFmu9UyNtOXGcWDt5W
XEBmfafMAkS6YdDUz0U6zaznkMTSsrjk3Oz1LRWselHoo6jQdij+jHmdw43X4nWsGn21+HE4qMtx
jD17Tuxm+lmriq01JAl/1wX8shv5oKwgbsKncn6hC1Ya8FTI2OehJ2+Pr4JjkRMLZaQg58v/4Guk
wj5lwijlNVtdRyEQGWtIJQ3gD/JAfKWT1sVnCoB+lKOg5hdRJqWfyiTt/DXwHhFFzrkvJh9sfjGr
mKWKHikwfsg5jxvSWNEygEhtE8IRp/m2uMMDlvfM8yvny/DhrC5/CO8eKztGpeQcvxjam9P5IGff
EF0h0hX00seHgWFCRHorNrQ57vp8QYAv72f3Xj1BeXG0nlWwCO7wkiYjb3CkcTTSBGVm6sWTzzNo
EslqbvujGCpPRCuZhDs4Xi/LznytWJLXCPZsgLuM9gqld7NELwqQRvoPcr+S5ZontY97Vl1AHWor
Aiy4PEPvoTVoBGzouPs5lTTrgWFvz8Ad7qnKRveqIom3AlwVW9og2/DKSAactj5aZ9dcTabiuurS
mlzyb8OBzJEIV9kGJc9cWLZ3xwCEVL0ZZUpJPrscI9eCtgfXARSK4SqwKayC7AdFHegGuNbSt7fz
inWoNuJUyeQDgYYkSlkJqLAIJ6CIz4/VkVRZ2eAbw33Ld523jB2Q7EA0fYGlwfG5LRCKpYaEd7hw
JVEr3u48ajQ0rpjf9BtQJn2BB7450qAHdcANTCGZoyzH7flryFsp9CPnvOCILd9AksSzuu9ox4P4
Ogiy5yldwsZv8PGmNlcWqOehcgLz3SmNjo2kv5+yXoqHtHN1tMSkSiUNyVQncxZfmfjfXVBi/Bvi
/6qwe20zyx5bD+4+G0kkUvIibskG8kEIQd+n/Oxd/2LClptQOsx9PsD8UtbSY0TylpinD8bka22I
ViN2jnM4R1wnWLu2MJdIS8rylB+EIYlaJTp8NbJHalYf+UMo+ILf8II2CJHASUDBAWYXvrSGXBSC
6LIyR+JN7FClkULOaiK4Mx9MbGeRgQ8g9vcG15Qvgzxj7Vz2NY7i719vu/uxw4PTjX6EqdwTHSTU
hAQBvzloEyCST61ys3ZjhCExv8uijuNUkRHk9r7aAevzkXHO7FjH28VmJ+ywxXXh6TW3YAupI7C8
FLH3oHcV+qdrn8QGwOaDm26S56RxNkFK086FmQ1q+hJJUlQ6oeh5eyMF93QKJnrpECqSf3X8B+SK
0YyR304eIq8kkj1/CVXGC3vQ/+Z6vya/pxjDdhGOrm3FSvfuN7jquVAFw7ryPG9oXb7mV3zoH2FK
PQKd/Y5T5F8LhySImej/PzD8Ge5T1thdfqqKkw1IRKv6BcTTHkAQ9rdvFs8F8pHj14b1BAcpDows
MKbHdmYYP1bIyPS81zFnCbg6IUSdZoJj1xPopdvVO4W0Ve0C4bj7oLr4d6DeDz/ra2/tpfn05poa
/l8pGF2C1JF69nTLqa6la4IgeNC4jfkSqtLFohc9Vv1BIT7FtKEx05ExPaXN2wwdscC652VN1aLq
tX2FzubHoIQsnQPmOOlvB5/BNf9kpVQZZBYOVM09v7/IzmAXaGbBMsQ5IzLKLRGwcXzJ1jGINwA+
jrI4qU3Ww6zvV0ILnCKco4ZGtPfCexTt3fMz02MMRcntGfkIkn7CvyNZXVh4jz/VaNixkEIvSKoH
taxwJyCjcwQ1bEqE4oqVBgVMR+klnI0xlRCuw3jsKOI17xrDBRLBzAzFWjszS5eeqSApROsSrwUr
sD/BsTpfnACOlt4+TqSgOIhawYY2MST+3wrvjc32catbkFSCBzwyk77QaUqti82tHf/Baw9cKuwt
Ip6Pzk8aVnOGn8Q19470jqe96HaDKg7DKqzghwO7LXgtw/N+tkk+VzmtNj8WRdMLf4Eww+5IL+1B
ePSJk7dVQMc3K0vWpg4mkBrwubKJoIJH7SH6Nuu9n1hFj8Ne58150XOTHgBA/G8DwTE/FRdQ84TW
P2MEa3oHW4niX0VD4onIbp4YG8fDRNfExr88+7OmzLCfdx9OdH1Hh6kGapVoNQkIcGa5olAGDorH
1EbxpfAPCZvk7zEmThy6fdybrfqxRZfBwJT+ldCcEBoAD0ML/eJxBFBrhCzp2X35Ah+VTsYd1h6+
D+eqzJ8lRo4LByR1Tv4HSRAcZyvxlDgYywT8LaPoEQSzqb0CgUZLtgOZjyQKJbpdg6S46kXeBpGa
G6Wu2YsxsYdn4P6ma8oXAV8I0/WyVSUh+qQHTsxBZRAqFaQZHCpYS4arW7ra9M1N6IrhsdID6UXS
hATzAbylNxgG2a55MlsTXe2qruiK5ZM5QwVSu5Q+bIOjyJKa0hdFde2edIXr25wenfSSjbwMFSkO
OP+34or9fiibLGCQfB2xrAVliC/jwGawinodLxzEm3QMmGbZOmY7pDMWvLso4QZSVM0YjeGsDPRq
u2kqfnZwwEc8uvwPkRaXdbbtpPvIwx6CL5DFpuGQMRUaecLkERa78vo0lB3PDYP2qiERkYyZ66aa
A7CdGuvmkcrfpBcyTVrAkpkipEIcI1WgG5RYxs8kuFiEpvvY2R6ls4Syt3JcR9X6aRvaEGvk90Fd
bxApqSk4rp6EXIApQ3asLsI1VXMGP1WSJmoOb+YWfguwOR79kaklBTDFJVO0WtY4JLfHtFOL0ug0
IFfFBToQpDmyklPjtMRGuo27jDDN9bPdYWl+JlNfjVL8T2kIyI7wXi1URj0jPQO7knY26PYxmcw+
cm7iMHEGLrQ86xn90M/wAecNk7Strxium3f60bvhL9KHt1e9VdqQBZXTG4KqiAmYSZYzfX7iLtSC
PolZ0sZZ6/PQziKMFPzSyxCNWzbAWnGzNonmLBZJZpKHZufqbPfVXDcYKyRS2hrSGbH86l6sk0nu
EzcuET6jgwQwSW/XeDhoZ54G6jjWoKQUncpX6lnJ/8h8SKrSFhlKejPOcJl7LhqZU3JWSCSRm3gW
QYkDiY94wKNvbe3ofuL5LVpajDc8oy57tu+v2GzGF3Phvaxi2SqnHZ7r1OuPMb+qTIJhvNL7xbXr
iZzOEdiDqwPBhLrqz/KN0/Umklt8uF4MIg3VZEPg3+UiPTjrlsw2hcLiD3Y37aHDCUZNd6UrjjNB
M91AG7JuzUmCihoV83y9cihKmIAXV2QSo4M5RZ9x3EcGnJKtAq8h+qPkyb0egTP0IDNlPiAgxpsg
iQLBP7OVLdo1wJMa5fftX+/Jxt+JiPSZTYhm6o+vW/387j1QI4qNRnZ1cJTJlZPRqOJVstW9VHP3
8B8NyQysiQC78Sz03vI2nwDIPH2GXlbZsRn0yeR/EetP/1LE4SMw+DXEnzE/+N46jCxlJ5R1widb
JYrBMgLy6/oGF2dmpyW9mBqLw/kJ6FkWySLbcLGRE9jMP3beI09k3oePAQF4lW2vARe/5HiPg4N0
4aFiF34jlYjIIpJVOyeR047ZRmlyRBAWR725m8MtHo4GkcdPU5axsmEl/BrE/JzttsRu/teBRTE2
UWcfrAiElVPL/DUUxpytCjDq1MQP0zo7AZ6alilz0pVKyb2fjJc/gqRlhsyXJAvu64ipSOYcacYm
shUdccdWD9KshCyDtejMluIbmimJweA9UEWG2t8X3J/8kMNDt+KNvhmCzBJ/ROQU2ZBjAYJP1vH/
+rVz9DgfBwMjHbH/MMxkX8WwJNhdcYQ2lihbeodqtgMHhuVQ9JZWEBxeeRqRHPhn1F/uXdHv9Mha
COBI2eQBhRgUnB/27EoZLaBEroStst3KBfkVhy8ry2VgoOLZkrJAaNu++ix6ag4rY4VsciDEh9FT
iLzMAdhH/uk8KSVmQ1T4p1ekxxoSe2H2Ym9k6GZ2TOu24uJXPMu/YWMka6szTF6Nl+O/BkvGV+I6
OhdQcTcXE1vXN6gUAmY6UtKEBwh2Qed8YMHBBIsidcT2zz/0zNct9ukaP6IIybzwlxkmD0AGkFRI
BMHfEISicinO0bpZKSBiUGf5PtFxeQOxdFHa4bTDsG3RgxDB37LteMHAuRQXCBPph+vyK2juSw3s
p/x48RcJM++aI4unxbGvtI6y5zexkL9rlbfqmF+n8fbIO5FA78fBRTaDYhuJ4VHB5g6nhugrlHVi
sxZFZLM50b5VGa6CUCNp2B0tIhbgZ/Kb6KZj82yL5XGjzrRo8Djkz457p6XPTz7mkEQwmIUHJAQG
+Se57GBwD9aUjAI2aOzoTwT2DG3EsGkCKdS3SWbNKfZse/MjLg3mHvT3ZRqCW9PyX6zHpcz5ft4T
ralSkiKYOs5zDoASdyTN8DEDsvtoNJ+YxQY/H1YOWnq/sq0JX417fwrQo10QONVja/iIRlraq3TT
+KtrZtPNpZkonk/LwcPhYSWcPUozBQGMGW8pyysb/SE8LkikW6cx5RxdbN9LtwRrlPD7v1Me27wW
z+S7h+ObmqliJIGdx6g0cT0sMhKALYszkMCRdMn1VtUtHwIbsXRGDVIHnpyX1BxsboVoFfQ2snM5
pfLpi6A8MgBz1/SnKLMdjd50t7gjqiinjYc7KtKDa6zFSVr97xT0LRRh0s26x4dD9xEc5ADcP547
xjopElGOONAvU7kf2uL0bZPtptSfGvZqR6y/WfNiwx6WeVotVYbf0LwJVwlUE/+V+luhz6CIkIXW
jJHk6NYde5D2vvTrOX3nsKXsRE7R2gvMlO6kskp1LswKtnq7i1VXy+5fWC9KprBM0sRhEV30gN3t
BKXOhDBOOpfIhZ9i2cd+DFw+ZYW3IuD83oNw8IDrhft4MwgCXRiJdI9a+qv+kTYz6fuWQgLDi64f
mvk6AIqijI2PVp/POLKm01JHoTODDuTKSC0WQB6x0HWxBv/bFBabxUzy9udIvqWImw1NPxw8aMSR
mu6DRwua9PMADC1j5JxrNkp9Pijvkvn/rg1fnkNQRYDhLE/AxjLcv9PMcNC9mR7riKzdlEDAAqEz
bZ4aVzKb5XdKcowNC9p8fHo6Tus8eZgrvSXTStmxmyLniy4Cr7kZe+aEpBO7KNlfhro9h4+sJzUn
lnKUAvVzQhjTnRvPEpVn6weUEmmuWojCJRIU58aEJ868cfPIbPruE9L59b8Wu7d9ypENUu6f3H/u
zCtfgN/c5tOK3d/Lj+sEJt/8ru0rELczBa+K8DijNZMz1xgESsckdeth+Gf1hxSDitSkEB/7zuGd
cMDamIiVV5DfrpaGxJchtyF0iM7XKnQOhJ3DLlnuN3F6mOwoREE2vgPGrRQqyINRCbF0yFXyPb2K
F8vCHi2Bi1KYGVBFcNDBXedlA4rq9VvchtkoZG0ifF7ReMu7h2odlkPfGKGW6z9hJ6H7YKxODs5H
QuIRTXuIKnVi1upwrbXSOwgGTj4+gt2r002Q9AjGtApqLvPhl7ca15BPx2pc+6G2ON2QaGiAtaKT
Tu+7oTmmfIOtuD3g/oIH9TnIS0CsSaLGLaw4FyLruSuptuwNhElml6bY7GieYqLm2J5hY76LO9dx
B/opzsMjuEf597TvDAIcDSH9DiqlWRoBBcTD70AuIzhU8Dr/Fj2ofku8PqMRasHPT2d4QjrQbTLd
qxqotgoHG2Dmbgm3G85EgGsHVOu/dl/Y2tWUocyNnZw/aUCtE3KZsNV6GTdNFMaVc6oS6uTdizNT
NHa3lsYUqwHa0YjOWmkO38TWnsRMJQICAhB/fCCwwdVkhK4gWHDePhMewIvASw+fMVwz3uXQmpD5
j446/uklZcTbzSAswRgUHspUsfJhQHrPi5WcZkWJhpEfWOffyrpX4zM9631KNBBssf7tdNWICr5d
Cunezlgve4e7snTC/asX5PcG98TYOmiyUtYJ6Jdk1/SyrngMSo94six9oUqHUKgNsRxgOpsLeEC/
a8R3HWvcFoQrqihzbHIwsSyqT5GwvDc3CawB44IVX5yaY1q731F/BNX/JaMh4mAjKqrl9Ove8ZSx
9g7TjsnweMXmTIEzPZkDiXkGJygX+PugVYnE7hQvIBzbtngsWx7NCmkuFS5fb8hxiYrV6rXdWlw+
Nx4M3IQo+6bQoyywYaLcutL5n5tGbppILP3FinLtqjPAc5VybIdmjECV2e8ZrWaQWDf5ATS/cwVZ
rHHW8zZM45mklWxXUYrlC/69kq4HyLp0QUuJ+l31FiHkppoTVpgJ9AgV+5v3sQ4Js2Lwr8CkJZXV
fj5BJDnDwKv01QUxwDfaygySf9Nh3gBeLXzg1QoWzl1RaWSgq6Xzp7/buZMB8Rv0jUM8EY5PqKRI
BHglQNZUavcH55uSyzrF5gacqPMAE5Ylcgff/hQj0vjqsITcDO2aHFxjseeIvU0NRGB5ew7br2WL
U2QXLqfos4f1QdFapZmG/y//CMDewgxTbexjmIPXGJtTNlUCq7QiWisvvmCZeMMeuAOns34fVloM
jw0owJf2uynmzeqN07LkKMWtQIgI/c5aT16PhMFSnVAcRkX+s8CWFEBSf7BeSpJJgHTMri8jiFz5
nyodjf2YrnemW/5t7JgX6HGOQIQVmTrhnPF/XipeAEGiDYYgI88MfPO0LEF+03giu17KH+xcwSM2
25UqcMNZ7qURDmtnNSECDENYgVgBAOGEeUzg49Y1DBR84CKLrP/zuv87vIkwlQetHrJIOwWdcTBC
4FI9OzgwE+eYeJTVXUUXoohtqXWNOf9QVdbOpDMdvrgFEbbjfH71rXZgrKof43hRiJq5/+3L1cRh
rMEu7b2ZAp7TuWog2HvwhZON4tiUMT2a8cQujRRVjn/6MgK2olw2rpJEkaHmkckdGGaSNArGCZvN
k7nlcI/6GX12g/FPkT0DN+rzA76c460UnVwHvAAypf/eCoxoTZwpH3q/fGBJ4GRm8HApO7L7v/Jz
KNUVfRg9XDn2fWlA67O1KP7Clnw0o2LXURc7vr6Y23k3fD3n1lvJY58jyz+ttcyy8Ov75eSt06Fe
WOPiHSceC/wTlCgLHg9BFe4xQFBEfk/jSOHyV+QAiIJGX29SjfuPuPPbkOwXTcgN6mXP1xl8+DcP
NiAQDBd+PjgIdzA5OJNeijuOQCm0ZG6/xUWw/w73FuV5Rr2yOmVY0B57B4f68mXE91xMhvaz9Uf7
iXBh4Th/XfDV8XbmC61OoVCsI9BOv5n/vSEloC2aigMgTKHQ7AWkEsRXJ8RzCOtjxXUddkfL76z0
o4icQG/T7CChutk364MmVBoykua2LkbV0WyWp41ElCzPVxHZdNEGG5eSpPJX9GhFrL0qrcXIPtsN
xmCpOdMGRhznYYGtuEvipCsI9s/1TBgdqETURxMu30RdyUsT91qt49jhCAaeU+sys/K4fm4g+/CU
3DkmGPwUH+/W0A1m3bhAwyBtf+00+ZZd5+wqrvXQwfBXJUPSSmqOiftJgi32fwff3VZe4AISZTUg
Cr+cYjv6jN6I5tSI+cKcKOxnodShx+KHZuScgdwVwMc/Ky8gg8wNYiTDgnHh
`protect end_protected
