`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZaIDYQkL9fQwO8milqwdrsg67fOLp0uG3CcXzB7xhmynauRDFpSMeLwaF9WeOUy+2qHOJLta8q3L
TJs/uACyxQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
khCdPx434gR6tFZjkXzNmrh8TB3aJmQPGJ+zVQtZHaHP2R8J0ou47DB/UGjvEstd/qN2LDHSA8UV
XTtxj49dwmEOEbaMF1MXG12CYEFhAj4DgnCMsgt4FfvSIo5tLz0ZDCfWjOPiSrDd1LW/Aej0T9LL
r6chvTfQNPW11inAWBw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nn/n2JRoMmNkmcFKurddLbjLiBKxSjzDogDR40dxSYkyBJooWa9HcvIVzGpGjl1jg1ljaMtgwWX4
YqBQtyh2J8PuMMLcWo9gQLA+G1sHG1CpmSw4rnftZe+Rzf7oiFKmY+M66HtAPjnFQOXwKdKpTPLH
k/HvxW8/je/E2wsyA0F2teSxCXxYit6hG97MPiKK6GJH8Jb1BW6sSE6kLGhWfvIwFEIGyAWtthoI
U4n8fU8trc6o4H0SM/9MJWIVe6CYrORU0CnrksEtNrGRzkKHpyIjVpUBAx3rX8qiR1IIjaXjqZBf
6QKq8LdXksO/bdDyPS7y4vPv97m0HV7uK4Xsxw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
w0dmpTAQPjjFEWkh4Rl8NC7hd+oKdx4bvdiu1z2Gg7BpVI8EKoQRKkrUmRIzt9amptZVctxhK+tF
DqQUqifkL2nvGEXf0TgHmp5E/xqOExSsY+nBHVcN45mrldHoRScIT8+Q+Qwag+TWRb2iAOA4wrZX
ulCFaafDTf0bpWPyucg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
muVlZmArXgh6BRq/5ITO7/Sb1rGC8i2InoA0XD0Cb/wRK9mQAYpwiqaK5zDnG378rpKyl3UndlwT
8iiLiWnm+jTGZnIUrQwD/dZ0FUL5Ew2JB/tfF7ZLbe/g65DWUmrnAqjiVCkpIn9wbzFwj/2pkGIP
F7vE20Q8jl5wAKvZKx87ao3HS7WeNI6Ga+BSug8+djHwg3DfU6B6vIxWAl2wc3fr648766U68Cld
+gNgbTL0FQWc+1KqEnBK/EDESLGM+ouJBmIjXv26cTHxb4VckTvjurzS+H6CKeJ2Np83Sunjm7ur
t3fzWfNYnphpwchLmOyZtPCVKiMWqSptRpL+SA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20896)
`protect data_block
pdiviNaT2vLBDRtmj+ZGskb/s+ZuGCApajqdGKdufWDyUCzSgn9wpogG82CKLWx2m80NVpJ2RzwR
CGc0EegMSA717WiJzv6pHvzKUJIp14GiboH6N0foOoDZXcYZxZLdX3PAZD8VHhOXWGrHRuqBnEOJ
E4m+lE4qlr12PiDWPQYz0Yg6x30xLALdu2zaKoJ3jkjuIZl9LLO1Dk8p1alX2wn9gHkUm5vm2+lo
vPPBtJCCuUKyU4nAaxEGsT+7o6iXsxun8dYumrPhICNpRkJMvGbJj5Biz+gW5JSXJoOHKkcgdXdb
Yjaj1QoimjQU3msHng5x9D5OIIp7HVb0Taw/EwzKsAIVYNuK2OA/IMFvIEccON+nCKaqmMzVpS7m
/oDOS4xd1ZHqe1OAViuCal4heBeD61vySaahhW8VT+06xi7Xl7YWE5xyOGmAQ9WBta6w6VmiG4m+
UzYHU61MZMhBbvvANWVRnsRLv9tq3+ZpJTuow6pBbITR3LrIpH6UmSyMQV/e9ZxWsK9h4Rxw/EQV
hrA7C1k3k/ZZQ8orlmZUK1frqOmloFwqA0ZDvNPGli2ex5FTjp8psLB1zg2p1YGvHP/CBu5wiGO8
fGpw9Ug6SwmSDW0EMbMPiw1vE2r+BvUtJZTBzc551sJ+EvhPQCukAgw0dJTGvILpDg+4a0E9IRfN
9mNZBfT3Uj56rYblPLXBg7siicgS8sKoZnd95vEQdDPQ95z3Al8yEwoaOWNYELT0Va1mRsK5z/US
jNSGhgyxvcGpLGxBO0E5J1bU65q+S1TGymCZUkX0nWEQ24t64XJ1AaTUU1OahGYqJaX7Qn25jVz2
2S+WyYRs4iQpd9DVaWIbeRoQYngaFYHVZGJZKm3xg7mNoZSsSVPpXofVaj3iOUAHuT3N2eDpJbh2
hz56d43ZsPoUgChrF9yPpCnwGflzLsgoV7eOi1ploCeQ+qP/BHSuS1Zq7vYDnxEpIyl3M9VfHT1w
R8YRb3cSolNkrqfNCSbjCl9X4Wrp199snNcsNwbAwz/OSqOdr5PioPfnF1pV3i1iZxT7VOwAsDOE
VOi7C4ZkrfZR0U5id2b8lBWMk18/PZmRXXDvaFaD1bpkDRL+HT6TZXyyH2EwMmwTu4jF0m6GjAHz
6Cds+IrYWEPJQ83eoRwL+kefbUIvlBV1HvSiHlkkkOQh/4PYLynLfn4bEWV7bln/3Zv/H/DHXOG/
Pi8suAVRhUl/gug1QQnUH1kacAZq8E8nZjM+cMBqMpb0innH7QgPqKRBRhaIP6zP9M+4UA11Gj/8
n1ZycTD6lgPC9MJVuPT7BhqvLp+UePPGUikS8n3zoHIKnNlae/bmjR622Yd7xu1N8Zp1UoIb/+hq
Qg11LL12WCF9NzcFFns3mvHlYDJKTVrnTEsdsG/Ue67iRs+zaG4mDw34OvNL3HnIhtwl/GqxoWrL
z1Nj45eiVKBStv5SZIWbGa0gXctjm3bTbAEKe+JUDZMQCr012QUTrTq3254V8a9ESkMARuLptzpZ
7jbQ96e95Xc+/aL9z8uT6jGFNX4FeFha/9EVyY5NsbDbNj38begLK++iDQUVjY155AkQw+z0WlL/
lpLGGufhAqsSYM9I8S7A0taHwblle6AXoHbIjm9ykeEsfNipAcXM+3yKgu/B/xJS3wvjbADwV2AS
E0KMznAh8nqNCG1X6ay/2KxAD0v7tOTcLxDLYr9Z2Mc0O84GcqP2iB0V3C0LzK8Rs9KBMc/YZGLl
0l6jbLnklA5UVh9FEMxmlyLIPAwL8kC32JM9v5GWK+eu5VEh+vUXauVv0oj9aBQAz0nblif64tFl
sTZT/0Y6zsGqdrAJI/EWYPu5ted4QF0sFrBtby7pkObsbj7NDAr0zHYJr0fxgs7zzUss5FZhO9Cp
g//E2Ry/c7xHZbYfYyUdqp2LbbYeFAJiA31WC9an4lexHpXh13Xs1VfVi6pYvplq7TwrnCDWFjV/
05SyGpmrKkg5MjLZ/JNeqqGdqjunn47oupfR1XFMWmyjzf8fix6ZfO/9M00VD4JBQEwwrRAffNoZ
KgAtXJVEnSfNbYf/04HURP7I10oN0Imiq3vaSF5ZKZJIebbMPejEugFQR6UoM2H15+rVuU7qUnI8
YgZZNSZZjRFAHq7QX+6D+pCnk36V3QVC/O1wONMrdCeLdr0IrW/qIFutQnO+2Mxw4Sd601xPIhUv
FyMxF2IFTc1K5WCEEUlQoG6Wusj0K4VYIn1BxzSSRS/8MikTDGYto2mRluJJ1jazx/QfO82gyhT3
51wFD6jJ0AUK0+I8vItVl3QxGfNP7CnTbBvWib5fvzM8LRS8AnaT7M7ToyhZHG//9h0l/M+d5Qo2
a4/tf422QCo2k4iBzGTQ0T3JhRhrppNFSw+ADTiUihrbLgoV2rfIqdmDNIGzDPVr1/QuTuHkRjvz
A0x6S5Cs6vRFAXjMh+BiwPvj1ia88Tj0GeaV9qaMgD+RYy1O07hxJhrvvSvXPkM8KPf3ERJWaX8v
qeUVvibTgIHN/u1nUh5VsH2Mu114zjBgc301Ci5LbEBTUNlE2/MlPK9Fg2crF3UbblOJUxAonM+g
giCkspoJQwU7OZEgh6EYRRhnvJnbHNPnMSr8/Wl36zV9isTQC42u7LOEx2UsLsZ66kPHjSynbb5y
o6xDNftumZ/WdHW/7sH6gA0ZojYwPkLv4vC5+bDx4I0rp/RSl8xOXeS4l3hIwOByVVlixNQmik3D
6V2alPxc8RYcICtgZJuz15rwo79eWn3VyeHou8h5ezFGU0q2Ih7VLOzZT0miRRxEcFQu93xErrmr
3XQH3qEVZSv0yUBZxbjQNUWulioiOm315p2obeUoXht1mrPe/xOS3rq/VmLkKEj3gy+j2zoU+wBK
TkqSO+nTKCsko5++hRAWXI/scZ+RIgCCJHjuG9xLLM2cN4W9ayZDfKgM3plSFB2xXanqKsMcx4Aw
vU3Hkwf6TIPYUDmsU5hCs6wirLqba3jFBrJ+R3CyaTvZm1Kl0fBmnPMdYHuJpUGrFty4NwiNkqbm
IEhd+nfqGwlJtEmP3I+UZLtcp4OE0F2IqrknMrgcZQ5y9sALL7TkrtnVs7gs3/vvRzMNLLEOtJuJ
lRk+fQL2VZRTsh1t9Qat7GpIVWMJqvswGcYTz7omnLM7I/fwQTbFc/7JYBYiSZt2CNYlUAdPtLAH
Ui6FO7tu5XipkxaddJyOdfk8Y3L54+MtGsxqMYbqu8BzbcbfK1J3++J2TH/9FnRdaBFSjv8GmFoy
cS20l4y57iisJbo0DMBa3RO0LBCNyv+tJe02SaE4YqlgA+EawCKSZrnN/ZrFCsL8AY3khXLAwtmw
OLqsPyaXK+cSl2JcarbNgzge1H3Y4YxuBMiEzmnxv3aHKVtRVnbnzaTRgetFDxC0jyO6at7vSaOX
BjBa0q6TKdJWSOJ+h+JFJ0HD8cNVU6qasPzQ+qd4BJREkB5CBLq0GixcnZCLE39gP0me9B09ZA+V
bFuYI1FhmMuzg8OUUXsGDqH7UFfAQhBS1bZ2dVH1x3RFrypwV+cNCdWg4D47cAxfErKULSglhUwZ
tFXIHDnWDqGxXbya25YpIil0S7jaLL4GQgk1k3hGERAqDz/XOH2yeQ2RpO8Mc9kcdr8SyJ1+IN1m
LCE72Zj5+Xdo+OnldQxcfgt+MvqamBxKJEU+fJfiWf9dYXz+SKXx47hY6/JQRsJblnGEFsIkgKa3
Ka0ByF1PU5jvCDB/euGQWMqwEgWjnRPTM6cr3PXyiweqfFaIhTZLxVQeCTjOm2njEP68V0TSSl0C
SRLhn2IhyvYeO7D6Q8nNAWdSHW1HjrcN78+Yw9itNj004ZUJPOc3LI4Qagg+EH6B9kACdjVBUaJT
gQYcj4w1fJp3StCgCZoZnsJIkYt6L2k/6WB6I4MghAbd6GTe2w8xmC4tA5Hy40CDdnlt5JT828rf
Mflkp2QJ1PKJM21s9jqaF0TTIyjKhIAqI0O9Wv9gH/miqzF3FilvInrDJb97mEbq5AIZ3iLz7OOE
UnJMjRhR9IWkTPUaKGC9UCKKob1vAn78gdXPUjz9GGIKwwAmm9EWv76zT02JiFUry1VdYgHootI5
efdPfOYE/0Z2Bp3+YQX7Zb68g75W6eSYPPEiuBGHHoItQHubTt6rPiK1K0cBPOYVB5ax9P9XheLK
i22TPG7TMrBJuGSaXqC/73WHziUTfQ7idnuUqDswT3kf8dHJj1CFHqGNjBWel+vSiTDk0412sOhJ
RtSql0d8OS66DUoOlhP57E9Pq8nOjq4gUCEjMts4cwm4686nhVZu4JFOKu/WFxi4XZI0oRhaedDL
YyMcZqZHrnZFizreDE2MMxv5gkxsmopn8QnlIgBY0EFC1SpbAib3tfTBYRwQqsf+vZkYNVVKk7lE
lgHJuOfyk26u8iyF2vt126wYjgu0jsqCdQ3RzVbYug57btwKRsWtj1PwniezpJxGbJLRroQFjtty
LWzTsaPYvVNBbivZUv9KBCN1qGd+a6HY8r36v6YRX60uCSwFzQlupCT0YEj2gz4vTsl0Kyl36c86
9s7o+JsaWkdNt2kMaqfljgjCN/+nMzS++ywIvBt8qTE+xwb1VJLqiVtRBuIq8JTlb9RPpcmM+GW3
44KX8kPzJ7k+ogfiO0JyRwQIjunhbn8s0O7qD6nx3XqnET0mJ0srytvVk6O2voTKheD3OxkXlHBk
gqheoUP/psFPQhoXcy5JKyxxk19jLiZR6OF4lDD5qwdvOfKbM/G56kv9fRa/N7YmWbCAIlWNG+Db
vTUuBl4WeXqbPOCF6ZY3Y2CR11qLFUyHpU0B9nt/EYHl1xLXYlGZcbeN7oTmbmgbvuzeMhG3Pwk2
QjhinJRkBdS+NnYg6zhQCOxVkAsWZPGRf1sBvb5aJBrA5IzrKmMTeBg1MDIKQPqsjQRIXelJcGKl
RHG145dU9Hnxl96iQfHrs8N07tC/9X5Iw6JSyb/gLUws0eOzE3ycv3AABTeMdpdq9HeKTXEexohE
fE4Dkrak/4SDQ8+EJo6H9AEu9PWfJltiPJzBaT1HOcgfbTzBuMZTLf/3iwN0sxaxAbRFdADJ2hj3
w/bLil5+5iAnbF2lo2rNWoDZlKVIJpvpnoxRxElU2T8bxGc+z7iumOVIbRw3vnivB8i3NAlKWZRT
WYMM/RwdVrfvWVZGO90AJhbb8WKVWSmKoAk0ngOchzPzb3EBO93sZ6msUJBjku1atOAUJ/KRKxOo
2QIjcVvjHcrTmw4eH1tL6f3t6XFO/Gn7Qp6hCSUz6MY3icPlYrac5bPsKby0qdPc5ZtlAbz1rTIk
8UjuK+zg2382KlvsjiDcclLlNgo2FVdqRxhX7j7nptk3mSuwOyoaTnJL2kELkPY4viWxgjGkwiig
ECx+azb1ikrmm6DNfjETxBuelgawKBB2YH6Sj4NW8+s0Ds9bGxAKVOdw3JvN5B/j9M946DGQusvv
HnMBt9ySnzQIo2IlFaSfYb6i8q6V91xME+/8SyITlmV9jxjN/vCu/cMh2jhISqd7yidVtdNRWxLh
KnarUOLr/n4k1D139WMWOsQd84SxbokfGPCB/hr+TkEsNddIrErMjxK9TCceBleAAbE4xumTJ+zd
j5dfRstGmAPmLXDL93RPgnxbbNd3HZbZyGC6aTJzWywTP0WHsXOhpw1xrQYiRlNjjdoezIU1Jn9x
uXUZ7naZH/RY8Y3JWjjaHjCz5AjXxEE23n7391aXVsKqQY47U912Yh7x2Bwz7WybupKs56r44d/Q
nbanSFIO+QVi9DPCS/1UIDasmjvN6Eygkp50P6GO9KAmrz0J45sccuPz/PAGXjtgtQhADP8e/cl3
SPNxdBvGCKPA+gibsM8ey8cmXmsQbEfAVW8hJh4Ng9mDc67VElLa22OPy5amU2hq5+/y+FY5vBaQ
84QHymErNCRALTYG+rpvlRT7bQ4XAYq4g7YcGeAmf/LGEgl+A1w+HvGjohZClArSbajBLgZALG8n
AYDVohKXs6868OqMWhbtjQwSxAF5M3RtNn6qioPwDWrOAB4cg1Lwv4zg64mfIN3M1bsiIfKzd7AM
2B73+HbHKks8DgBtfDpCCC66SULPfuiJsuym+14Ni2PnjmgqduKwviYGD4ouwn+QZjmeh6Zoj0UR
pNzxzI+f4KMW4yyuWkzVCEFlSRBMB7gi4ZWPQFrElV2ekIMfqUg0zitewjRyuv+r3pO2I9Oh2rxx
PjvDtf+01+9jXQa6YJ0fmgEOyLYOazo7udtGXTbARjrNnKLewpi7r1Rzt43wt1abULzeSgctKaM9
DdHjBRqimDoJ+pr8wpOu29HKtE5zvzdxd6ZdQjcrin9anbDV5U/qhtdg2socy0SpSvE/ld+InUjp
TiEtMxRprlwtf/rrrZTcoQumXOF/r820hdDgixs+kkiFBrhcwJHsc9onERPhnXdGPiuE3mZqnD1H
YUcF4MrBTasEY0tWuj8q52qGl6uYIXfYA2b+EVoMpjzpP1P1BAGzqCkwj+V26mHXKxaMLX8I5i2x
G6tWqepe9pchP5eyjxnCF3Fj35f5FSif434Je1q3UnQdnxqLXf3I2GuV8lKkvUk3ms4Q3127eA62
e9VaiZ7Weg/Syl1Bhh60Zd2D0huX8M1xr5VXS3ZbFk5i8HC1P554DVNeVrZCmKlRQmfsY/Liai0j
7SDJiy/ttiLK8xm0mZbfVJJkwq80gncwi2LH/WEH03YDH40LzF0md2THryEDQXasSWOht3iS3VzQ
Tt0R4IbvmVW8teGYabXsNbeZMvrRuYhWa9rZ3Q/lzHipseRHQi0ibXGPMAjnRqSwwHmfajR8hBFO
JU3UgwoKFmUVq9mo6r1XTlFgIhKF6Io+Bk/bzMxHzpu4koPfeRiMRJYWhv8r66tKI1IRKZ9GRPHo
LeJ9eYKObVBtDytCeyB9YKxY9yugcQiQcGWMpnLS5zwpRyYvNlX+DAfEeCnO1vcjJM4yNzJbPoyM
FpBVQ4tjLZiQA3bMfxYMmh1xYmUzjuwCorDK/4WrFBchJ4858Uh+NSlaEJF0M+kB4wU9trV57/yJ
Q8/Hg5IWYVMl9ikaUd2hOFNsSpcWwcEw15ibfRGM4EOwxL+Myc73kB6pNKuMUvAgZADBJDUa1w2w
t8L+8fvewHFajsQH5MqwEYv0PVjHEhiFCLmATWB72BzIOOyVMGlXVR9hXDCrX5Pq03ieSCU2g5Uv
4akurrDh9WAvkmwjUrkvC7QB4Ls5ITuGvFNcghUTvT9abKIxd9NVcb2EoCw3Sh2oAOuPGjmVdq8j
IyZQ5L0hOGykISi+kAmhBYrDGqf6EGctoeJVZafPAl63q5yM0nEoZU6uiAoBJlvZaicBad8ZRPJ2
qqAVS34fMXyUR297Sn3IEjDFlG+4MVrs3whoobmf0Nf1MSNROBiCPK+hQsEr0hmhOG3qyu7BlJBP
OyWAOpSZDTblmviq4PURUHNARYpT3wmQ4jHJfEygUj5jch2J58Lta5mRLYdMrxphygT+pPXNe0Fr
VwTse6oVwiHCa33KWXPXtekz4rG7Hsno13+QXTbSpzbq57bSDG/p44YLOwF8Jfzwa9CftffeDFcd
TkYKXXP4OV/edWeGXLm0YZkMYf7Ie20m0mPn18e/0z1wrCoNrVxAYEO8EExXDIo6EgdVqrguOHuV
KErujXZUe644Cxmel2elKW1GqXPWlTSB00TWopE8ditocUZBBR0V6pLDaBp3Ty0Utz4rv5sWvYlh
FKPZcQ0KSnBy0Rp1SawLs+cEA7hF8V3r7POaY0bfG07HoDjR49XHuedKINpgKdQUakKj4jtH/jmd
awEr20CKSRW2oBDjt2+MYUWEV4wkyywKcPmOhIT0tESCGICQa1ZWL7abZInwSWvARuJa/gCW5I1W
QVc/P3YWrrCfp3sVBlcCZEBUUa//7HL6ljrGe2WSoX3tgd+j3WrLGQIp4oyZIbXgGMlYrew+Om7l
z8InHrn3n9i6gk1b4GmtWHgWxq9G5nWq5hVpVSd/CtHwS7Il4stlLGu/GEZRTtNFPDzhmXuVoyJt
5MMmW/Gx0AbdmxRYY6etERurkzzANZvIsmFjFVtTbn/o/i9dQZtiwMzSheHwy5gK7k4GqfzX0qeN
ma+BArOt8X/9kxh262CxxY+HnEgmnLCh2TDtY8gC5zn7wRgnHSb6JLJ4P5UxwaCS1BKipvKfnXgZ
vtum62G+VeJ1ezYdZu//1cTOQqbkALjQLpqkXcraghxfJeWAR27PDllJ+y30lnKMIMP4We3D62lM
Qbph34cV1cApEMAzz1a9Uft2g0e8rt6jJyrvob52Jr0foFZDX3TwFJWOEVyUBAqJcfXbrsILUmGX
JhtMMAzUq3qk+1eIt9Ct+avAp/h11pH3AxlJgC3BIOz59vz5P5uo4m2eBEqn6Vs1/89dNbo/ekAl
ZTzPhewhYry+wOJsnyYQvFrzgVLlahGQAhipBrpH26c4uPGqNR9Uf9vRH09bPzQcp8XPDikFWu4k
rwChihWc5ST82kwO4rIOOglsOCulkaxM2FKk16qguCR439ELANvmTlPK7LBS1vbAUqtRhCYgFha1
Z+fkiAPM4SwuPSWrmIpa+D5Y83CSLMrZfbSrNDMNVB4a9mDrVL0lyNZ6ClPZPA2C+p9Cv+TNT6rF
1JZSt/GmlynJ8lAThRaXJgeCxFbyCdj3+9EFEy5RKwOhCgqLTiFC0ye/CxmUf2qWyk8Yo5tpkmDf
CW2h+QP+b+afAJimS/A5ry6ra4fOKlPQxiLQE2Qq6AlycvX0aMyRT9zf0Hmac5hG2+qOPxumKbdm
QNgMmKAc05tLJT+oecbwDAkx8j3JSQtRG6q+N2sKTGWxETDoAoLbb5OQPo8MAKPT/9u3UnUFejUv
jIXkhn2EGArlw1lsRdnfK7uRtSf51QZmMyVFcf/+MJWWeplrZjbv2SA6BFs7H7Exr+v0Q/hjo9eU
cfm+hDOZS4ekE4IyDzzL3D3vH8U4dPfyfJbGTVhfFm15EO4r5bQ4Su2rXzMKj0CDeXXseB36yA61
/AbYdzh/tpFpgVndAH3YGgPVQMhy80W2r0k8UmIhIEkKrjaPQhtVRMNvYbnJbo5qTuNrTjBpEzyt
5IZUvedD/KklnnsYd3FEDh6CttJZAG0il7K5f2MfO3aKvZQL+GCaOyVv3lPxf0WyEfJO4zqOjW0g
YbBeSW5caySxjoRr5jUi7Pbf9SUKIsBPjVzsJNBtoLBlxA/97B6mlS17GX81Y8dDiX+up214EHN0
Zjpbo65hqmfZDb/vzAYSI0Y60NiGPjyzo/23O6pfj1StSUoI2VuWriOsOFODM+9NHeB+pYdomE9q
ajviqOB6ptq/W8VhlJ2InwV1ci+06kZQ78l6U+2fsxD7bWWK2DZTi2bPUkOsOMjmcM5b8AUpEB0b
aOAHWtkM2RktTu3YeY3nZiANAD7jfDsmRoFx0+gblq2jqJ+ak1QrfioAVOjr4XO39a1NYE2CXRBS
28R72cI8of62WJ1KgzC1JpRJqaRNqLXvN3EsvNu7s3i77dGfgXDEgxaXmEj3DyOF7HdZAYGLixJx
gL61FgzmKDVs7pX//oaF3qjXbuTb7F6vl6EZeSl6qmhAvczNN5FIqLNhXqzhrpkWjqsH3vqbXIvJ
2hPZn5vDgrDwqGY32aj4o19H320TShs84xps/AaqzLx80vznOk85CvWmaOc6boW0i6l/gL+6zGbQ
k5owo0pfBlncIc8CQrP8ZocMPeEaFf5XDnsfBdU3v8RtK7uIPY0KDUjOFKJJQ2RXDpBL0OrNaiMX
S331zn/dwGj1AiSgNyF9E2WswPQ6+W/qUNdVCDsUPHmQiz4SQv6NfOBPvoApZie44RQ1lPvwkR6m
68rvnq3e3vFBi+r7aUPQG+FgDU0ypXwWqVzHRf3gsIY5iRLkSgIbxBEwhQgVkDz7C8gP2TpM86jK
0flwq4TMrNMihe96wYgvSFKBT0C1eKqKMBF//0LQoNwBSNw+SSOIzGoSqiSx6RyWZTfmZKZjVt8i
8uyIe6Rh8VUcAS6Q4tu2QKUtwII1cPXYSGvSiqhjyJ2y/U/yJHTl5MiCMIOZICF3hpM660L/wTD9
RK1Eek0DnNgUa7rleHVCtUIGdEYzS076atGvvKl6yVz7X7LKIinfVTHD8fQHxO0HOhH+i6HBc49k
RuCZ0r6FuNzTqq35ow7CgUJkB3CfvQfz+IjGoTBRRIu8Kb8Ys8+YogS1qAGDJA6IRHdBZ9s4LKIP
5M6KDwXUyzd7r3pmApdYb9EQBZAy8FJ8xVXuZX0puGJY0My6rL3jEe3uhL8bYn0igDtSFFNB2qTd
T5njEAvh3mY4g+Su3Lja0Nr1XLoNU729Ze62p3r7DFiAm0rWoObo443rYm9jvHAc/nfKXgZqcGKH
AgT0i4rOzqIBTEIypWleJVXW9XlXvUYxWAd90A9MWS/XpAMPaX9kOmMseXwARET8RofmTLSIGNTD
4sXuLOa/Fysbek/0y5n9jiXZDQvL3vQzvAVKn6u4D0+6X0WKA5rHoC00E+VftNDXLMUpcm6sCv9M
fTquxfCL48y5sIRwNxZxSuqNEgCS8cooEfXBuwv7RvqInJ4tKZioIfFRZ19lTSWhaIr55HNkrlvy
qSgWI7/phau0p8c6CzC3Xremt7IUSB5E8fOrB3MUBdI4+SCQdvKZBsLIOiqyNdC+G8iWzOXVf7eo
ks9VQ1yxWbdS6DlT6k3sDoEyNhnd3nlupV9GxhB0OsYUYAk6FlJTYYLGDSIRvDriftGx2g4FLoU+
z6Snv3td0lfxUnrYsh1+edl5i9ZfvO8oQwq0trp3HzTZB+aT0mnnn6fk3cJI4dBT1ciH9Pw6pHVr
j2Ek473uJzdaiaoJEjxkNQcg8013bzKN+aJADJEWOg9Ktyyjg8j5mFZ9S7OZv3/4ebK+DKx1N+5P
JvswU7+erMdp65I5wUOINCKbBAgATx2c2M6G7HPGPfPHY3yyvJ6m5/Vv1qs33xgHA4XoYjWjfpK4
vS0NYohMsODzKg6sMSa7E5dH7gqP2W1MR86kOP+4ry5NZJ2VhlRxw6HgcPHDcXV8ZRvRidu+X+D7
I97W/7nfcRZFTuYx7y9907RHyyo3fmhJKai/TNzn90lpv9525qMiJzKXaV/D3yvRTvPoyQRReJHF
wEKbsGULxO57IAb2GOCsBQXiHiMcbfOyHgALB/IVmYpPHorvYiPFDcKElqooiEl8asbYS1Sbvr5A
hD3cpTqoqPNHhSPYDZ0Asj8S4HRTtZG9B/PmhFhtlxiQdam9WmOtDuhpXV/M2RR6MTMFBbQ3+r01
ChhckimKrgi3Ksiz/aoc5QPsbIOTL4G3FqiA/Vrn99ZVHkjhsRMHzj0WuYazEZuicX4Q/QTzY1Ei
ci/MSVsGsYyr+M7MCZARQnxwwKgKwAwKx2Q66p0ImwIDrTqd7wJdbBjvrUflDmvVWEtmdyaqJjCe
RtyZHXKXntkPpBGY7rKdrTvQGlYATIVLxuzK5WPm/eOc6mr+mC1uS4fMJXmIOtamBrj1E8Qxv6vT
126NzrWd+wuvHLZJnm9tlmW9pxLhzjykuTkyYH4FSRctIhPTg8R6EqmE/td/DNaWSwEx98HLVFrW
tlGaBxdsdg1FATDm6v4sRDwuHsRc45epFhjEeA/LfcCIWGBHSqLNBjxDRI9ueFrFviVdJuzu5saj
lJXRNcRIPh57Ff2GYRoUdFrS0lSKqn0B0uNXTtGtFdxSiMOIZdnTGHz3YmTk4hglAUyeMV0F10Gy
RmZH412xj3LnYJc5qgLmN+o0zoTDiCjVxuj7UJBTgJfeWoQ+Z8MY45lZyjklHCQMlvqiVJaLkD7R
DoUtvCGkQ4DEFRH287TAtqKUAas+m9r5kaCeOuGq5tuB1oBQOR3HPOyAFylH9APgd8sLNVT45/eC
eUjJ36iDJdpQJWxXjxf0MG6IWlP2upt4YZzP2fwdKcEQfkmWz39kFPDmXiZ88yX9oDLljiPCKad3
wU2SHiqRGVz6DpVRHOngKh+4H9JQuMuRdINQW20iHlrdOgkP6IuxNSCqLTZBW/bgugzBkUBHc5P3
ArSRnNlUlc6xMXQVuBbYqaMqQ/7fYZisUHMIP1Vs1K47kb2SCtjfX01+wL2p7NJpC3tmaRmGdYNe
sPbpWPFUV4BRCmlS/bxnCOTtL2UsEzDNCkaOs5neBNw9j0OETCTfHQnstGqZQprX6iQc5OxtLFsr
TlG41BGpLfCb5pe1cHCCcYrwcmlvhdDXmuObQG/lzOmQJPzd77h6WV0G85VbKcyyUQwbxgwutHjj
l2uBD37rHly/6VlmLkdlN2RfB+BtZBRCyUKH1dx3hCOzH/QgeABsw/t21qatNdlzuGnA47p4I2rM
UFByjld7NHU4B3jvOJZFGPilcq44GAX6/9iz4zyD5F6xuwoQ+0EGXdTK+EmM9gYEf7aVdGYQvQ1y
8HVYbYPQ3s7nb4zzSmmNt83Qx7KYsTilNWt5R8doAkNzlYZ+jE7mcXY5dQgspz9GL+T0354GKTMu
MzM6sx9hcw5BmlT+p9jFhQKaKPhXbUWAAkV+WPGGgEc3PU+9hpe5J3wSytO94v+grG36fD3rVQIV
vItJ2iwto5kOkqnSaLXbTVCj+pDf4ssF5Ws5jVars9nb6CeZ8EVHN1eo36Nw0moT3FySMCNIyfVm
S5O7gjnuHqOeZmIFbKwiJqH6El0UrIvSJG4ZqxE+6YbNtWDM7LfOXE3eFsnS1wPlA8dv+QhbRS3o
ukfzM/fWlr2Eefv6C+CS36Gc2lPFZyObREt2I2uj4wETa/2SbOmGb/+3Ujct9391YXi5ISb9FVK7
Wy7PPrjXC/YSLUgxck5tMN8a0o8TwaNrAJzTzK20cAtA3E4FndhNInHyBQSCX/OFax3W0jGx/BeX
v4szbz81/ZQql9TP83bShXyrWxQPWqOJgT4Lhe5WZVysQr6U3DwbDXm5mXXGD3eTL/UwqJLpa0Ws
rylFjf+MguTUQfdKNpzCXs8KOBQgQXwk952zG/ml8XeDCXYFkxfiZUo7gsY6yAt9A5gd9TvR1z+l
7PrvLB3sUkRjUKIDoOypPT8Vp+RHvHStJ36iTfXJ40lMsGyhIiIz6IeIkwelh0FU8GSHUI8ILgMH
jpA71Vcdad0H7T2O1TE+nXRmHPa7syqUhuoWwBcFhTg0QFI9tpI1lAku8+6ausABQkIkg26gmAPX
hYIGjpNVS08G79JWKQqdw0hC6W4Fkb7KkOK5WkRdWj85EnbNdSRFUJjIi8b7F2VwnqW2VuGcYWO5
XDe1KsEHpHmS8utFFhNOcAibQtjgmeDnubJpy8YBg44MWfgsc5KW6j8J7ihZwR+Ns2ar2Eh7gbzh
8nHFhKyerZDyiBUNmoBekZmc9Ze2OGChDA0EpGui3pbOA/05gl5a+uDzzoGKbOvPwUZluK8+rPH5
gtK50QGSHhBvSifEabC1weLXqxRcwmSkKcRRA0Jcb0e1KnBAc+5WlzqXKxL2hadVQ3yiGR2rRjBc
TO6wmE+zEua5I0aMCjc7GtjwdAG8l0jpqoVnX7FEB8luhEXvEkIZMuWl3afxmbW+uL8mdgAWK+9S
Rp+KJKaz8AiMGmy7skpLvP0PMeUTSO3WKzz6UBIfyjJ39U/7mvgNyLJwJRhH/mU2LN9U/S12ITa+
ZGh+dWSA+1l0DRF1SxBybvYvLOJ+vi4acIqsH5SEp6FWfHLCGCD35AROOkJgEPagM63hDCF2M810
b8NzI+LyQiWaWszw0CXpw9gIfjqYNwV1ZWppkcEGEH5YsZggWEhkoLP7D0e8TKrxmm/RAO/YEVoF
soRWajSupIj0YXpHBHY560sGY9DNtoQIt15i2C2x8P5F11+hMwYTJgZSY8EnIveMj72R9e2uj8/X
//k9FDH5dr0jqgs6NLyTUKLO4q34ls/MXSkK3itqIkeLZVli3oWq+Lr+ZfxoJ7Il5LJeWudFF3QH
NjHgPaLNlZyeB77gtMmPYZgXcYbhvy5wz+5hV1ywkMBvCbpSWYfZIZjezmftSZsDJUGxdUKbTsRc
Yk/BIzQaHMITTBw8q6xjzu6Sx3+JuaPZBM82+hVB0vdzs5/jBMjFud9w3lnyi84tRr8mfCHjUlSs
KEgcyWqm6WDbezthJELPMJfIA55Vlfcl2jzmcBRvt/nQ/vGVOvEPe5014TnoMIf5/Ga0jENlqINp
3PihOm5GeFhoNPWxUYAH3dYEZzQcOvP8ZXc+7l9zDR8UYaSFkSys35eLle5wRU6VlUBdEh5rsg1f
v6LYikbPpiTzh5GGELQu0kMjIYz/ixiRF8hszaWcsyYCSs3lSYVGhqXzjbhqGi+DOC0EKdcs5qAL
vooh0sT/vRfce/1/VGraJHXjpWaZPwhVjW4N1QY7oFjuZgZgWaIOt43mhWLZixMmmi9wSBfLN6MC
AzwHvwDShapSzx+yqaoeYazMNdloUQwe3N6LLbYP+So+IOIdkQnfBSKdEm3xPC1PeElS2m2t2oKi
b72ltbQEL9/IMxsIUUcj7oPqNzhDOzguBzGNX6evK6pCBFYNMqYtZZqGakOYx+eW9bQHJk7Gq33T
ca6OLEe+O7exsqBRCq9Aq7RaoJgQ4iY5V21ys47Qa/dpjAhRVt6b2SwcwggoAM2NFU1HZAabN7OM
7DFSwPXdMFHeVD/NeHg3OxGim3Nb2p7VTMiqGDjmFva5VKNFoqqO5tdxZeRerUNwMDSL2dYWD0Ou
zaZAH75MJycv65KiOIsz1Ka9Poldn3KRTpSEMN24R5XpcOEOJKO06/66U5VKPPVHUe5C/7wl+tz9
1iddlvg9EEDGVmZLZ4cAybZHfLVF06Bo+kmqD+LD1LPSdDWoiLScAvn30o1tWTrEB6LJitaowCAy
3srrr9cr03uD/ZpKro8hQpb/mFG2ClbwwWo7hX2WJCrCKOHk+EtUvMo0kDB1lrEt96RB9iCYYeh4
0PaC7CIE2ns0aoeLQCgrc+v0aGH87ObRMiNxWGofXRbmGxqAxlof7IE50eq/3RntsLRXbX1Mej4y
Iif1zhkH5XLzAx2thG6tXshFrH0UoRKuShdnS8l/MSS+1v76j2GnqgL/KPwoQJ1vmsWvYCPt/hIV
CApKQ90ZChMo/pEpabwgItpzi+zgfw62E+L0Z2Qiq5ScVU/FfFYtF2kVGBQrbmnDJYKuIfNsUdux
43byPycc+dc1cGMv6VTlQn2E6dJ5A4rPFlvolzJXtKmvYjF5H7q56MNVsYsDaFjME5qpU3QRJE2J
rI5EDbxQXlm2SE8Mz8e2bj8KHWEGXnSMYd0TNvg6rJdwR4cOdrcE5qzg/1SrH4HGVV6QMjbrtuTT
Fa9GpDQuALsaL30615UeSIrJEN3h+oPphrvCC+y8We15KlScwaS7Q+WCUUp7+Pxbv+xq/0TY940t
0z8rib3ianZ/LyDlN1eLqOFYWvB1dBDAN/Xe4zhM6tyAyzOyvYr2I1p5gd4pSjzfctvI5/wpc1SA
Wt3h9r1onA78WZSHuSG2KhIIlMGbOqNVPyMCVh7+AY9yoRNhjS6YzhgZf7x0km+5UOBoVHmEKg8b
v1yoWqvyys2Diu7+UoLUV9BYo066f8tpyYWhEDilZaMOterDyvHIuVpqkQlNTTYZg9+kkSL+XUgH
M6KznXXy1ggggyZAdmqs4tiUle5+qYHDxefDimXMe8VnSyVpLuiMNpg80YWZ9kcTKIXrHdEwjog0
CgQORWyQ8IZnrYxcHgloB3ZH9+lqbJ40wTIJ8Zkd36ZNygO4GUE1YZjXCXNv9/LRWcfpRqVAVpWm
gCArKyE0nE/W88t8WtWwr33nxmaWNK0jX1No2wKZK5JCtRhT7PBq14farvYnfMrBB2sh5D1JoBKX
eETpwNlWWhhWUvZVb6MTGucn20GE9fG26e+Yx4maX2a950Z4lJvzdLBSgqKoLm+5gd1n/G3BPehg
R7bx8NoRp9+SedftHpy6GiRbPDZ4xHREVZgTxGDKnbDFKfbvyww9SuPq9oVx5K7HtL6moVLvXlRr
1J8CEyaUdZvQqdPao+3bGZlI25VNYIRn6o/gM4e4vR0GKPK45u/FkrKNmfDByOhRo2BrN1qK0Bbj
sZx/FL4vVR0avBm5am8RS4NnJPhAOSdx+WfxQZe1oPg8bJT3mUPrha36bOHUdvCR6+I83+n0FUub
6ZzUAEAGQHroq+QFkEUT6EJ3nWnEzHEnbA2yQ01FAPfsaux+8a9yeSCoPvpGbWes3Z0tyDkzjaIL
VdlN26wOqWvbPe5hQ8foV8m5K/C9zUVFAR03cyJKR6Cg6qw8scP8tLhvEF3CoeBG5sQxUGloVEkl
J2OQ1AUajF7dNNTSYn0iHt0BXNRGDHwWGwRTGKzgOgxHXoiTcIaX6bPSzfEKjy6K0cWo0jpQWU+2
XZhiOzUwYaTE5oZiaQ1Xv/L9APryl+wztJD3WS4gWaOLU/e+9XAqq3olTbTeg45a4XHE3uaCUfQ2
p/qbAvIUtenSitnMmjACCJjZD3rAppu5NHhqE18KtnsB6Ni5bDqCus8Un4wUhHg5GYAHbotpE8mf
D7maOr2OPRLgBYNXn08eZ+SCYvT+aCsdzx1CSTGocwI5rVJRO08rX+rYe03HcUyxJvgEvtWKCeb2
UN5JOBWzmO7sDLBTNJhiZv1KTWVpZt/f35NVOFMenCgXFkc8UX8XyUwwx5MOBaXErR16U4psngl5
ffdNjEzt2mj32yqIf3FZzW8X3IatLaBFuFXL+Vql86uOE07Ftx4IkcRQsHBPMLV7FuZioiS/cwaB
xPiXmPMKp/vPJpj9ryfRIOatCH6NDQo7kMQP8euRT2ZTZPlxUZi5XBs522TYAuaAxQ/+PhKKc+4K
dAXD2Mxt4A8j14N9mB9Ntn23ZsNNj3THO7J+8geTz3/7oFoN5CTYGEPY2T8kaXqUznddbQ5u71+l
vn4n3Xm8DGZGn92rkoOyDZ3GWdjR8fpUiAdFKBFvZyseWf8EvtkmOs+3L+PdkRxFZ5cOiQ+kjRRp
uGje/ThEFiQy8azxKNMUa53LjwjVRA5RW6h6a9VBWc7bXojsv31L5u8ejU07W8sp45wmLscEu9J+
e57bHGjosIyJmVA+p+X/x79gFpIZLJnYy2uvQst+XIEM99mCRlM9WXu3ahJW+L8y51GPPFbCMk83
DOW/cmtSOIsOh3f5prx5pDcjR/5+EjLh6qUcsUA6/hPbbFARumxtIj/zfn1aE9auy5QGby56xL+j
22eXHxKQKIDFBRoQRD2zshj2GMvWjQgo33AZKdRdZZjRFvG/Nsoc6fUTkUkuHX7DRcfVrvDP4Fgi
JEPp3rlza+ULUYF4x19E79fCVwZgnqGO0fiv6EIWIeudmAGConvq5RYyqfDgHHqPkyvFIE94NuLb
32P1d/WFSGPNd/zPnIF5wcMu2TgBF+7qLMrCVM7xZEJZDdntfXTxlo0PGFqoQQCVmwIhXlnHuRz9
9klhCa/3UQIT3k5gslB4x6mfAF0EH/qBxRfaniG6J1DvkPKRIr1nW9hN+Bb2WGh/d4P0NYofQZtl
d+VgQEc1wcYYyePlJyge4Q4AjTfatv+Gc2jKqrE2w/mSy7mjuA7jJ9W81KOAMgVhs2ZsrLzMzdA3
o5hVwwCC0aKsGMjR9Zmu19R/q+IM21eAp+S1Mtw0ef3TBC0VKM+GQsJosKHAWR33cZy5uAN7sXfM
QwiUm3aRCJBpNO7E8jOJXhcj1ypByRK35HMuOkdjCXBXhdpv871OuOcJCLmznkrpxv74eCxD2jzJ
UPvT05a9v2nhpUR1VCy8JHREEbPMYj2mBNCtbpdhOcmCfYZehzKETI27dejPMHH4kLlVVM1MT0HX
5SXfXiqlF2vM8eNLotWFGEoY4JENKfb+GfVW5GJe9JlISm+EbTBB8fZfySZXUIx9FrNAbBTFyND+
eQDzMC+Ljra3OOf7bLoTrfvJD2joGFDRXgvk+fnVsNAwdSlRZMztT/TR/Xj/HV7Ie/5zIGV+Q+xY
c8ZIORdU80XFPDSDVfQSnit+hiFgXC3bB0uooi/RB04AYs+FsnrajGdH+AWdUiGXkiXFMVyCUO6Y
qWVHO2U0BqYt3pG6T3zqlx0GpDEoOELgj2rxjeisphuhri77UqUZKQG+tz3Ravuq7KlKR03UdyEW
xB5LLlnVxXEz8QnEW1AZU1yGT7enEMKZ7Hoj+rYvRq7clZl62g5u1oNYyZtQLmdEyPgu9ZZnrLzH
8DNaDe1ynH4bq7SQhbs9EEWm0LoOTkjkCI3+xtmbJ2hOggc1lNCS1qXfTVKTtI9AEY8QKMvhI8nu
VvqU+TN+UV85l6PhfLqhb/uh5LW4aOJ8W7WpSvmzggMjfiUdgVNEbNDNY3/ez7aLcH1fPEiyuW4x
RD+garkFbEhST2jjT10ujR/Ozpw6nRMko0YGDh18daArNLfAO5ASYft8n2ocywc3QY69AMPb2EVT
1BcsTlYKAQMO+rWFNHMgl05Nus0Qfa8YMHcEed9wt2TBXkU7mIc1yo6aadR8k0stshQGCFQ2viSm
kSaHIpMmRfqoPA8yWfCqZmR4kDROx64BuiLNFvSVRixqSA+yGtvmuXqbZEnzcPJ3hVGWsXO7HTSv
VVVHyzbsAvsdIlE4yfv1ekgCXf27XGSy4IqnOCC0fPKZXAd+u3rwmfoJIahehroCL/3fNPOblsWa
CZQo4RfkkgHIlIvX5yrXcQk2kZnTqbOV9ORURDaVKUCQzTt0fzpUHTDTQ475Jr44z+VxUAqZ9HT+
BSP62iv9kPU3WY6TUsFvxg0SKgospoLynOlD5BZR4pi1ytKsG/tsAxoeA2YhxksldBdiDmFPh1Yn
9eD+YKwjmEltgqkdksTtf2bKKahzhI2x7hHNbciieEpyvqRcqsE9/zj1N/eagS168uwr6IVsAMfL
r4S2SKExzXuPSXiKJFqh+O3O+w8vIhEcMNB93sicK3CDNpeqbQxtyWXMDRL+0QWTiHB8Ji2koGzu
smkCN67hpoFgrJN9ZdK2gGi5ZGZjGLeQdZLzVsJZThlwhbwyYcGEBM3ckv9zq0SAKV3AAWxzupqv
UDEnEnxaJYOc5WgVz4ntqglJryZ32+NyuQStW1ebZwRGMoP96WPiWomfnorwNy7Y4x58IVtWzYUS
wxrDFZBXmqOicFAd4FxKMKIRPaCRIXnl1R0DGxmg8Ud0S4kRNsH5ZUl3X2x0XsHW1l/cTZkbqVXa
Q1yIxvfcKeALH7neOVIUVZrWLmC33X2N2rqyknAhwuvnwvRwDPVlLNkTIg1NSA+xj7o4+V6Gd3ac
ni0RjEMzCiRXgrjtJtyuCTesqlu2RxdJQNCbXnkP/5yZAkE+agKmrHTq4Ob5WlRh2WY8OdwNU/i3
54mPwW0hzMYxlcTzqrMKzWQW/qX/ofPmLi0U2jjHXU65xLrdkedGzBK7aF2sCQOmlV1a4xOd4deK
TTPZXEVoGHMkomQYo2CH/r+Eo8Tz8b3qKhaj8i+U6NpUgBZoboGm+oghtmPuUlGj4VhKmSAKVGF0
sAEusCBfxNWSIrE+ZV4DlCywl4eKzP785QbDpTbvm/sQPSbu6kn0y02tffkFSW2diErHHEKFf68z
kZTJ01Luk0edQdgznKy9M7/+oN6Pc1QugBRnU2kF0FASgJ2dYOKNdepmHRUVZav/8S2DX2CN6+/d
i0VtosnT88o9h7loLNXHuj/drIen6l8Can8FvxdHRBGy6P2GSGhKLkEfkqa51d3a/FEqq0St2tyf
ncaoTkUMu4HeUtkKtaruwUQhFotN6bBa+h2RzSxGGWBsSdYQrhFybgq5Ux3YMimPvTUxqwL9V0wY
mEG+lLEFrC1lNQDvlMYnw6Tr+uDDY3ZnyDyVXyFt6ItjhzRRU7n/vY2KZeHnDVv20vmTWmk+egzZ
uEsb3ufMIVJS6QJ0bn3kzlyoqg0uVs2HGu8LQdXcDjSxnU6auf/d0wHKgqermnUv3jJ7fPvh6b6W
LtswW48yebYQlnmPP9HmkjRGZP/dLML3Oxoq9+WcSz4Rbpfbtt9rM6M1APMFKQe9/sqaJsjqUzXl
8yR/eqLSP0psQQFI6vEeiLRxNCTMnjwnm+ENfNUVmXL9ZjMhPx6fg7lFW9Zk9Ic+jwZBUHcSY8hZ
+HP9QYBs1N2uC9hzAxjiQ45/11Q5NI+pyvPIKHIqyF6tr0dqgGRayQFMSYysG6/kSek4+Mn1Fzbb
ZVKfmPf9QzJuGLap5xT9Dv80RnL21kAaDEx3dIh7fUSaMjpwYA5Pwc84G+LL7pWLKfu/eNlAgQIz
JNU/avBdvasuAH5je9AUHhiSuDt09HWr3rBsvvS+TAj82HrVvXJQobFnWUfjjaLsRDij4WdBC34z
2B6higK+T/LIlgN9iBbaKwihTNzPugDUGi2iEUBnmBXcBBEiprEpwv21+1JgdoizgEAWwUyw+Hxa
cUJdKfDFzw9qvZOqRZebK08f1PZFWuFugLepygsyOfr4z8Uqd/SFxV9ObNFCDSxlqlDzvRxM5snL
uuFWw5vNd0vO/w+AqJnnl8zdBQLbPfVBsp2/5EotEwhGRVfHeSFOWbSYeAEyxntS6Dhn583yIRtt
rN/KxAzVEiJamGnjgLAzEGskBI31z1JfBb32X+uoc7j5aoLQuUL/P1GElnYzTKiyf/X6XUggKNaX
MCEw+m37V2wJfWDSQiQEKLL7UtwhlRMaisyU0oorbM4eEa29/JY4PZeLmDPeB0dK5JnnheoVz/or
5MQrlge4GdjrJqqlIkcLKQ2WsM2ObPC+7jyh8ZS5T0gdjdh6OjuhM1y7KY9BNt51ybqx7xbLqvGK
fQuS+86OjIawwmV0M/F6aYkskuzaal4xZjCso5SsMWOGyDdWT8cMpzK4YbYN7mzkZjVQUcHJ6u11
c2cvXVDvOYajuyUKExUYQnhrfyswrcqrLGIr0juVq2OI7WIbdRm6bnW+DGX1JJbKASXRcFfcRgp8
5jjNMEtzn9KLe9yajgZRERWLDUKmhF6QhGRkQlc5v8RDhDvVjilvZuHTcrqAAKHR17OFEW8FC0IF
OpYMiENLbVomjq1gsGn0qNzyg/rSdMnggIDMe9i0d8Tnup0OInVNwx1LD37kbidDS7Ma6a8QhfUo
rGd6IAlgWaaRE9IHTgHiAJ7dLMRARAih6dZc6ngQeI/W4AzOcmAxYowM92sfy36Z5tRlKLZeKENH
j6L7Yv18LALnGy5bvE0lWYLbwX7sW3PL2Uzy0QMNAnqSEJ5VfSsedCu7a3F+gndc6X7vQTft2wcJ
M/p3IA6sN1htbhpD2lct1KS6bwNa3+Tbp1rBWxzClW7aZ7yoB6dyCE0nx8gXZaxC70HtUUEEpZN6
Z24gwf5Vw9KwD6uKdVMTYUHsnH5SJfEwEiekIeWkSJWIcrP9cDvktsE0JF8RAaoaY6Q3zdGy+0hs
9x5I5IoRC9RS8nPPkKB4a7m6ZqcbLbrUYJGTervc79O7LXmrAJUGluywl7bTGY4XQUd9X9UuLU91
2dn0oZUxxBYZ5BQ+dO50S4zoJoG4a328FmihAETEwnpouzLJBgdSc+Z1tMAKVjAmsKdEKMabP0Dh
TGdX0akUPxVqlGihh7BZkFHx7lwAyXPJizsPKIEze2ya2ohFbs+DnyrmIpFzESAK1NYGwfAIIxyl
1KmInaRpH/tJZKGdKiFopJhhBTfd/LqSnbXNPHb/wuOVFcbbctgSc7YDjkd2zt9HiEf4izPNvew+
HwVDf6JXCMw5CJxhTpIfve2P9htWp1H21+eeJI1AnaVxw/hd7nZ0ztAx5Egeca6Qklo+M1smI6lM
ASgmpoBpLrOGG0phRJpRS6G5hYxNchPqegva29xkz8tnw6xLVmZWet7i6yp92qh3izFglp+E1nfU
AgteRwHRUUsEjrfE5u6klkPLaO3cIRYed5+m3YfpmaaQe8Ep8yGls6ToStaM1ZxqYmID1TWvV/vA
vAPqa/g4K1VJGlZ33JqNBT46S+kv8gKMB0aUuGTAIEGhpVC+RBSB8iADi9jCQXV48vva51+4njPs
RRCVn4c3ysSbgTdugbmPUqLqN2PESUSrDcmjUYV0cpNP7Aw3r1C7C+/qheSRQex4/xw25Rb/ikLX
6ggK36OPV9q66IIAM27+Nig6epvBpNxcqCGEvK2os75eWpkWlUPQv8yGlPHZpT0DSlTgbZUm/g0/
o4fd7KY3+NMIkVK4xuy68LIH1Wb5+9HbKaX50VDH+01SR7dPn0cJSxp03LPGJk/dpCuVxlDAc3NU
REWI4jg2DRV3qMMUo9+xoGysla1KQVvwDUYzUJmnge4nsq35O1YSor41vy8vPk7ND9dpgOa1+Bgf
sW3prXhksCrrM7NgCQR+wLMV/ykMVvsRJ+niKK8tjbHjvLUq8BmAoQ+X2RX8rI2AqqRDWqN1oyJn
gRKUe7WTmec+3INF2R6z6zTrUJo9BbebfvoLKhPrl/zC6tUA8tw/UYi4ycxEdhFU5w7Bprtnx+Gr
NVfwa2cRtdgNFGCveAXPXdWmEv9+oe/oEXMRpcf8oM+yTXX/nCHWtsuZoG5hU8BygRfWzlk4Y6qK
jkkKVdBVgGHe0PnE5B9oHGMRGzMMxRx12FLhcSivhIo+KyCFM9uIzgMMyUfzDT6q8oZ1nV0WXYTc
kl1X6Y+za4j1Q18Cew8mdy1uAaeLdmmI+qe65mXpXUoOFpUxrozae+H2Rd5Tt2P28KZi1wkfc1/+
XB3NupVcjGqfxMQppyVJVwIWIL0CFw+4bxa2b8ooKAgXWcXrgG1iAWlUZH4gltl/IQAP3VDQgF5o
B8WPCgAsqh5TRHz4nDYz0JrV1KPLVVhs7IzwpHyQlZjCDbb3XE5RnXov72HJkj4QQr/1vqCYbyBb
Xcp4Ev2H31cUqXR4B5ZnsyuwHO/wzhp9q7LuR17IpBrna2XLgmwtyKHvGt3R/1B4BV5QZmoN/NwJ
JR7sUa5jljTYCcIJn5I7KeMFwTFLllt1x9TbSzwnWWCUrGBUiKN8kzJOxuVlp+6002z+F+fR6p38
dNWRUu7UiEbAlNOEI2p4pUUBtYzqMXS3ln8ct1hdFUZvazBpoRh6qDaL3ybCrhQaUNSeb0gsQtIQ
LjoeH2cNUHTP4XbzF4GMeWWy6RRryLLUftTf+mxkTKEyn/BctepTndxJ8QUjLQKi6KoT6sq0JGUd
J0DRhCG75JUd/ePeOwxqQJYrg08S3NMbeOQOdejleTaHgkOsuGDWnJpjdpzHcgrqC12wevP5sHEI
UJwBOzES7w0WStfmvArwOrPte7sWXZbuw25ZVnWdwMj0oaioHh6pWakIMI3fcCi5OBxSNDeb5z1M
UoIZgS0kbLOHqJNfAqUVWPGIbOTaVQdy56uq3Us67Uz6tjdqaBgWftTH/RMHtBzFVB3uLXpzTP0A
Vv0d4g/NaAY2jJXfswInQh4CYV+qExdMrbjp0vstP0eV77t1+VVi9qRXX7mUehncyUTxKYcrPE4A
7rMgOuGB5BP416HQJgtpAju+1EBFXhXCNRBafulPmBdqKjXZqKzWyjYntEEm9T6sB0VBJlGhqjyP
o3E+O0Is3VpMs8QeODyU1b4gjI+b5yUTHjiKCsm4AcNPnesdgWvz/ychS5ImgLl99Zo7V0F/BQaJ
/mhi/fWz5TnZvQKRJcNE9LF07JpouERxkUW9lYG6rMFsgItLeLdYEL02G4vxfd9zrfBi6j3i9SCj
N602xoGqFAQ5IxPzqLklh71jw+nDi4zH4YRIw/vdyuvuNRsuVYTAUiKAnMB+2Nb5rfi4kPonIMPB
N8klL9CoIxDsHJv5G4d+3xNiSqiaGbeQXgs8bVjDVPzrFzRIXd5HqBf+XBpT9g0tjcYIe6AcQSO0
/zThgC2BuH4/1FFazY56BKN/oKtIM5ZsXdoVM04cjMlSCe1ZjA/1F81hb2xR1ZlVeksGWGue3bkM
M/r0m2Hu+UaN8y7RRAoaHvrHUubgLGXIU98nGwoaiJZ22tH9VJ0XQ37kJIZoxxKPMAJmm0/S+qBR
crUijQrtiFliiDiX/hhYel3mEjd/+AdMyd02DVgToypvUGX5Y8W9asqbn5HAaqmW6LPOSRcBb6vy
OJ9YmaZk6sfO2t9VGVy0bikOyBvkIDJdwQvJXk/XCGz+CAb5iWfCcCeNxa7ASEhp3lNxG9O20cIb
r/Xma8VQOmVaSidPTRjAvJ9rrPzMrFAGDmRHKHqcC43bNVVxDrVpJAnmvv1fSZwMFh5hx+FwuFAW
1vyEwv+/sQCmXP8xNDEVlb9Z6vJlgGF3RZJAT88ucLdS92gV3Wu2f7uQ8orj9qdMYZQcJvq72diT
QnASMmURieZtEkfxKAq+dB6xZKsQvsDzfr1CL7a1MELoUxT6GU6GU4XYR72pOQymX6rzPzYKXkfV
IVuGTYugBk496VdooeXaTy3VtL1WJuZpwpdWRbi4zuRDTO1xTzpqnXm0HXSJ/PWlWLyBb9FBr9Tp
YbjJR88hMqGUff/yPOS3HjRbTEakChcn2UxEiMQLhUk18UrEzQa8pEFtZuUNrNjtp7mGPD66+Tlh
idKBd/b3E3RMU2aFvDbV+nsI5d9t/Hj9BDHeS5+lU3GAxSWoiP1mOhOB2YInqpylJVsnYcVomtzF
PvUQFvARkkLe6heRtpaytYIMdtSGMnh7QHyNWP0tHx4I5No/QjkXD3NQGbBzLX31rjykgDzfaIUZ
qRjJWPvBa8fjlGtCA1OxxDh/RgxNb4Hw/CVqUwlWArsVbmB2Z+ereuDxCzKT0dOWJVWYsYtVgsko
Q1vKc7MxtdJVXLHIr48k3dQ5K1+8IDfRfyF47CbHedwfx6LxcQnkqt/C/YDoreBXTiJLXUUIzYVu
6Y941Jcia+DsmB1o2MLKg1BIbKAuAYUpHYioPCT0ie5Zqh1hXGNIWN3ajVDr/oCndZh1kyOPYyBi
YYCyDj40VciDdg3Cz2EM7y6frLpoFPZiS96Gqy4WckZeaLekbWsuole9j/SOYngRduD/G+ovz+Cs
g+ERxajRzRFwfMxR/5m1qJkkcglRSalFfVYcB25IuNWppxKHkh92AiAwYeTAKZC/Ydbnjm1p/YGT
BSd4A/ZLDANdGv2+hH211I6VDNqII9VYMQitNm2qxYCT0papm3p3wfegs+Xa2qyxuBQoKD9thlxD
rOjf9kbFac3inueekE9W85X42Hp32HDjadJpDpzd7UgoDQFwKRpcUxmbJyZjBMBq9YZpfpxl0oPh
i8lQ+omb7Y5hxvx5JEQRiatLg4UWLELyH2kIbMl8yvXO2s4yZy+0tzHMy4nBm8gyZUrtMz5QkjMr
1Dp4J5jle3k5AO6nTSr4AzWO3oTwi7g1fUsdt7qmztFQDyNqITVzt3uh9DkGs4GuHWKsTOfnhcvh
wuLucl0W3n5mR/Zjdpgp5xhqbtGyT6AG1QdVPOPmY1P2yk6nCHSeE9gt/Djkg7gK81wAjB8NYRJC
4MrXye2VF72A7d6fQCulCe2rd4SmhszjWXP3Sitct4uWQbbiXoI2+LQdInamVpO+k62tbKjZuUE7
nVki+KenXS4UvcxCrHi6OyIidMmdP/lM1alQgBVckG5wB+BquCEXo1BqtFkKY7Myra9ZPYpLtjFF
n83oWXAc6Wt4n0YDlMHrSqEZb8XLOdMWDFMs4mttTMj6w3kksZo81rZ9eXox8EbtqZRLkYCdpR1n
E+4Gl90THOC8F+27aQgKtT7eih09WFdB8rxHloGDun90MOk16Qwf9b4zdtTG70tQ/X1r7jjI1vEs
iG33TtXbgrWSxeYq3U9uCZDi6IoPdqEb3RytEpeh/kBt8t5ZnT72DnZHGwplzI8rxafIzg2u9pM3
PucfGYiFgQCZv3PyBd/+7ZGkTCd1vOiuXvmIGfqMckah+Z4OoL5a8zi8wZTanU0UfIlCtyPmQQ0B
KIdvR41RGeb9ZpMNiTfDvF/ADOsTsmOSiuvqK9I/iJz0rR/5jadN8cTNHweNScAMF/oC+CBb0J7z
PHEtMLhug/cUfyLcx8tOjejutk9QBom4H8nz0ygoIFQgFiauyIrd+qM68zXkx1XBEKlTkBXkBnan
YbalQ8TvcqQubCt3h5XIdf61DUz/uWbZ9H/w5ohnXgluI7v6RxYMA0W8sulUqA6PXKRMyMXNR7y5
xgjy0eT+j+PxJ5YeC65cnMIicJof7fcGId7d+QtOVkmJgZJzDSMJV+YOA6p4B1U8laZc1bR+1K8G
AuxWM9mUHc+ydhw7M7wur43ovPUG0vSTE8f6xTOjwzPLDw/CvIcx6sTl0+ZHCKNWEeE+0gp/Tgw6
xus6hmPETVAygEPTUIyTFRoJ8g/iyWJF3znmFWQPVEah3JF+TmZCVexEh9wizDuYQe2D0MW1b+2t
O8eqSqglkjSkYoxKmendJYHe1MgbnOLC1Y950brICajIgUVhd33nhf8tyCpKFBwNSk+A/n1Lr5LA
aNka30c9Tl+zPbiZqfNT/lI0NZwpu4RBfoutB/nYkurA17MxRZytY+0mDyUcNuQ4q3YxQlBnAxVq
pA2rWcu2uaAXdiKA2xhhfKriKOzLcUGvnTwQxj+3DJ/X/zzyejQULG0xUIqx/QBD41UcgufPkZQk
TmahpJ1RkxF1FesohFihW241TlOYYnsyb59Nej13l+oCc6shT0bk0xHH8zDrI0sNNwddTjj+95BY
DIvKrx5F4Lp2ETr0t5HXdu6ffvHlYbY0I6Sd2Ln/yEggvJ21nEQPriEHRmcmOWElHxZyyxYE2POm
FNJho1LBHKHjp+tS5k5wZuWwmqXcNkDNaWBMxEtRbbzwB2H5RpYK86R6rwesWjk5wTVE2GvEvpR3
xIZqGncJ9fFvuLaGzO5iIQQ2fYVwVEvbRXyV7aCI6r9TrFn/t4/jiK3IadoXcVLm2lCmYlVki0EH
4X9xDsY3wClN62AEy00uCyenI48N1REFcP/19CLcW4QBJlRJnI4FKjHhRdXra1LGiSUSV+zGjiR8
/aRA2iBgUlGUgmO3l8kqiXuYZiPi/qPzxE/FX71Se2B8KVFDxZ7O/hwUdIXhFFCNDK2w34iBWwiR
0wS2Vjomes9xpOXKpIziw6RZv1dc29OQW3Vu80FFdkGO0ZF8SFpTN2926r223sZQIUoxseG5IAhZ
i4W5QtfFnCZ0Nu8G4m28O9S4xE40hdZ3hcF7cuN8ZyvHXIGGl4HfMmKpNSwdoXBBIrc1Xl4fP+tP
rPsErqKaBjGHLOE8rBbPW6XIrUNZsU+QxpusCqejJCKNakXZLsvZMQpO9Rwh0FZVCBeCc6Q0no67
rP6oNzmFNqRTfp/yJK6jKXiJXM5Sv5U7y5O6wpu3+yvj5VFMGDEeK/dPzIMEteqpyuGiBweZVBcE
R6g296wfSkIkQ6elOCIo/DWnXhZfO57+0Ajnx13vxM/lAydXPxuzqdZ1R6lplALEhNPE6PXl5iOk
uaZ4yzoT82UOkNt4y390XRqa42oKWC4+olrYUFrx3leyc6nyPEhnXBXZqLvAcrweDQXKKkqhkI9Y
ujWekv+q6/P7lpJNC58Cy3NtWEQhXBSqawvJ/CVf+cLB7/k3lbfgvEcB9vdFW+kOW6DbLdNVCeR2
8lwcVl0HNE9OLsCDpzN/ps2wuSrU+68vZzpyANV4E+83E3JNbD+QIfDBLEf2m8crA7UNqZRJucmt
GPQuzhs9Ob4VhqJCdABTIpXTb7qY7YIZr06ET8dOzHiR5HVibVrX0u1xTwvP7vb8Lj2BZUAp8G/k
ES05aT7TjNbqcS2DTKbAPo+7P/EhCqA5zX7sO9XaUexZn3sNtdhRNDKFET5e1CHkRXUSMFPmH54x
4btT+2EeVpWQG4Gul7ZfwhBKKQaKwqiPdYeIzWXyfEk0pw==
`protect end_protected
