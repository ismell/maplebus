`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dx4v6c9vYvnygASNEz8Wt9YQDwnEzFYVIAcFDiKIl6IJHPQhwIfrhThphA7cw0XGZCiW3Ti+sHaH
g7gcATmSFQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jQUaZcrD4lrreCa/AI+vVRPjsaj8XGL+l0O3lQjviya17HBpMdVHt87HDt/2g4V6uw0mR2Tj74Tf
F6Ad/nOtd+o/vFSACZ+A5+r1AB/0fClmu/2Fzt3kOUX80dg214rrWDmxSc8/eXiZzo6FSOckGlzd
KIQOe45QmBQw6t5uWY0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H1WIk0GYOBW3hj8vq7cNJi2se0CigSbj9zDeE5/bvzzSDq/r5nY7ZOJGMTOOWXaavQKPdpWSXTsG
jTY8ATtNvY/EqGnQ8Hid8EAUXPZRWSWNQl+3r+1l57f/J3P03BH2ZYzcB5HTxd8umm+eVf+n+lwJ
+KsilER30PDLwBIUCeujtE/Ul6S1aUFI2QhngbEFeRGceALTb/CFiOTqcGFC22YOCOBYNMnIRmFq
1qgJeeCv/Xz71bfhEWD2RmYWA3TFru8NKofca03HRHaxWyjMPbA6/s16ZpER58CpeMd5mXaMTBLi
JzjtDS9hOHRwAO1Di9/qjHT0DFG0auA4xI9ZNw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EKj79D+0KVH/6ULSwK5yivwOJ/tIwb3kcjRk4TjrYUGSjCVc54FLjdAEd7KfBgL2TBPz7nBj1hHi
TDQiYFXmrOR+2zUiSCwO7kU4ToSKXckj3tfqtrpXZplZIgc7LKaVD56u2q0Dnm0h911vSou1lQqS
OTA8qJ/wAOLQ8/HE+yo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V1vgE5dAU3bFLw+cOfYP9905c4uMPNnOA1LzPC5I923eSOcE6YtRhf2p3os0BybYkU57rhzkXYSX
+TM758npt7m9mXIefQATfe4w3Ih6C/vGXgt+s/7xP0D8aLU0sAX4Buxyx6EbvBr6KrCp6h/l/PmM
zFS9uwgUh1NumTwqvvB3Q8Nab1NooYuz+0K650gJKjbQpKvp9iI9xSNBG8phF7sW2UT+oklxTuu8
K37kaKdnLVfhoYNWvQhXnUYU+Ni4pmmKzPXHfm/Km5pauCNog/Xf4bNKHDaynxRweVCDub9aYVDq
MdQ67fEKSvy+g9Z1bQKqPfmzTSqi+3GGLQ+fwQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
CejqOhuB2eRTvExa17JH1CufcrBuHV37NqMPpeReb7RNIPYRU5x4ky0++THIgV4P5742/zqTM18K
3sY/g/27goUjfKXtLIRru76Ku7fv0h+wLvjnOXrCWIzLJqY35uZYp7Wzm5enuVxBxEx6buQy5Tr2
C5ErFQj2Vx3oKA6JnPwO5eSenoFsddS173QAbGUYj9/u90eIZFAecaFMgUXX95hpInlfD8lGDRjo
R/06rGa3Zm6lxgfibSFuHKke8egKEVFu/hIkHYv8cMnoeB9YsAB5l6XLc6jM84xxv8eN6gbWijN8
cf26aIfhjqAF7Z14146m1bGebNoLnbbw4+I1P3M4c/jwLZTMSfzfQP17SVUcv0us9ZiKYoTUQsoU
mW+bcO1mH97Gx4VMSG1OtaYRHd4/zF1jNcQdbi3jD35kabZNADgrbYH8wc3R7MvKDJm7rfmdfT8X
aOzJWycLRq9GYE6kUzN+DXHKNqRlXgT8u+oyIiY7p121MXYEniKtQH2SkDsUQ88QMgbMVw0y8flk
sS3hjZ+Y1+v4leVgiTxQkic7uEb0c6LLl6dR31z5Dw8iF3pCsbv/aCIMBxspoKyWD6McbjgiQGO7
rLDBja32IT+AlkYt3vNE+cXqirGe4pwbLF6NQB5qV8KJWmQjvx1CxXf5J/RypKWQVi3v8T+61V48
smu+T3YIa3v9cB93M/U31tVH26eILtBYEd4szvleDtYbWNgEnA8+0uchu0dAMMZ5yK5B9BQCeeJI
/I4BsZZD06uloRQPJjEvHGU5DhKhawtNOpZzS8hhan4XA4fxU2dBTpwlNUIqV3B0k7KyCvVBn7mj
BSn8VtEUCQiPlKyoduQGQY6lQYlbeH/AfgG7YiTdi1TxMyActvbKQJNPFlhv8jEjZFVhbmLeNvgI
N1vjZp9doRiQc0XJEqxgoA+VPIpUZB/ODYGyzbiMJBIP3o0wM5JJShbbhUeCIu02fP/an49WOlU4
9ox+K0pCLC9IGI1fYjwu3dXG+RvBubhd0RFB4sjXyche9Z0qHDai1KKKWylE2BEdSLSnSDO46lC/
U4PcUX45SPrDlOQ+dpwhHMYSc7Rwsv6hgQfY8iQ5zeqWsDszmLL42Fwug0mMgZJ+zWlihLP7QTxy
W6i23LiXEVJTPhRGkVAtv4GsS4DzNPRGnC9QDeaZjWv29Or9slgN8QS+TWI52N8n49U2jTwMFleB
LT+EBeClW6HxkF+WkKwrnxa3Vyb9Be1fRMdZwr7EhclM8E/QpUXRIc8LmbpK+ldnOJSa/M8w9OtJ
lQX2e83sfBpEDlfgkEKiqjyuPQR2n5TfAvbh4EIhjACkDgj3xhXH/oH7BTwvzVxaD0V/vpS+xoZF
PIVtbC0Zc454rDCDkRjn2Ryj/7xekNlhFliFUq952W2BEg/yh6kxxHM6Ur5AJL2qlYjjrHSKN3FK
IE/LkcswsSJpkIF1f/hF7LF8orTscFGfWFBrVTb+gAJCqEmH5FUJ1e6elIltBs1ifokEv6eVOzjN
Z6KgSF17aMv3hRqWvZFcsjOw7d9yP29A4yd0UdNrkzFfrBAsCmVaNbMJcD478NKjo9bWMuOIBqBZ
xhYozTrd6TNRtb62M5WAEHuvbvr6o9OE+QZEOpgT5U2lJEjZBsrPx4llSKVJiwQV+4ATcuQyqY1M
7anUcqF+KLq+LxTXUA4RAElHA8vTauwiRxU2IXMbUdmQC53up7sXrXKOr7jijVD/EIIsTUU3Fa4b
DBUfcK/ZFAMnFe6x65yShUjzmAaqYflY+B3TozR36ERC75ZvWS0Q7juOaaOBoqP7C7hF2apaeBfj
uNe8f01wBvkM00H0P1JhbYk3qxIwYVK5hyB8hPhKj4BZ2pCprgavVgtJ/8Nyi3cHaPjms5LbFcFz
dGFWwkao84AX2jYKMsXw+A1LbeEHaGMLPe6oriG6anpWnjTkOffdO139q+H/NKjPZ4GDaWk/J6pL
HSEQ8HAhG0aIKrcKZeF0NZWsI/d4DsIlagWk7MyROQJqkI2CQHzxBs77Q96Gll7+3NNnx3/LpPEe
Njxf76S8uYe1+s1Q/dIyhCHBY02QtB4AuCOP3MISR0X7HtAcYDm2ubAjskezpOr6XB/eP2x/icwB
kPdINDOWxTJRG5T94mbxujn0yVkXaMn/ycmlRKTtVulve0YBTm9XLcyTM1899SrJ7VH9/ugt8GGe
u8kzWkhHapTv8vtz115zvtSq8vnXvzq53j6XJ4th7Z6YEGNBUo836XmjAeq1v/O3YUCK64d52cLD
BXKvKtSZogWT9j9X7O9VWizMP8StahwgrrlxQChcHSiQXmhBElQS4Y2ZVMD21zq4VSmbSVrEHIJZ
qqtoU3BaEZekM5zi5vM09SnIUSIOdYvux94EE2aSDf8z90xfnirC7Qs5ZZTkgbm1k05rHjJX/KVr
Fxlipou3o4kXRElWl8XdX49QVfXeMRYgCQAtPt05dbhYSgWTS9daeJRzTMW4lflfvtUrpkLbVMK+
VjhX2E7xwBC9LsO1oAL5Cb0hpWqZ/AWi0UYWJf68w5yp9s6sGNHYrSPQSTfBUo5FGqiZPsMVb6fr
Y8imIokm48Cbw+4pJ4owu3m4rRrkyqgmdm5XfSP4F838CyBWNdM5qxwiwsyTcx0h/Ra4ByuP6qtC
P/EtC/PJI5HlXOGHExRUhjkXV+xwNiizvx5neRirBu/2SqvTKpfNgL/k8rcnCGfQTFlJD9it6m3f
OEX+qfOlieR8l8vN7T3PIFULxS5Gq7P0LcnMT908b3fZhGFYJoi55ZEcw5hvpvEzvBAVou++5Ftx
LQ97XxMmX/mOU+16+Cw4G2g1ZDzIdyU/n4HrYGShLgoPPZNgJoqUfddiGDyP0aSXD7pKog1VgWDn
BN2o1YMwdHxeTEXbvC1591e75RypiL9oxV/fNW8RP96QgCqJkZLXrN0fkSCdj9jn3YzjCtDVVCk9
0mrvJaaRDTHFiXFunHXgoaWss2XpIDlIjUgFbvVfYHRaxNloWtBYtjch1D4Rk0Qb4JjLUc9OYtXS
MOmtldT9XicY+j20l9jrz87sjKNu8fKDF/GCGo7+Zq+/JC4j7mc5zCjEAmMWo+hBzWktv0nLA8+T
+h9dLFh62/jYH/PaTLWP8g2o+sI8Potmaa09F7uCJVskegWsVoi6Wte5NMCGM+WV2rvUjKcNHFZU
0VIfqqR8H633NVN0g7KxKg4sHUKb9w/LkkW9Ot/A7JJoKhlZscHF+3Q8VftGGu4wnBTq+pSPYi9R
t2ZGAye/AsxljsvGZ7SterQWbkJwzsehc4q2LGTt8xr9NpSPVrzYS368YAOPKupGqbsjz8p6ACyr
o31AFPA8/YyXYKrjwZLXKSiyftFXhuK1SNkNcLPK9+PhtW3iqCKo40Uqj1qTylTVYejJU5MUuv9Y
OowZ/udR7MqGXK/RPl+Gaygr4FMNUxCCAsi+/DUX9e0JCoeDIxV1jQEoQFBNCxqzSiMWrQi0LuKN
y+VZ9MUovcD4QWpunF7beHO22lwOJNkj/dRb/7xTEwP8DjtEWS5O8ukGrGXwiO4YoIwxzp6ZLTvf
MMQ+vDzetTBz1Juv2awoJ8QoZisTvuQT/w2xXS/NJGOXzlSeM0Jb05byRnX08xi89XRNM/Pb7Zwe
jRkXUZmObRu2cnf/p8JpVBzmiCfd9jLg86DzS6dlxKr/j/ibQCQXfMp7Dx2yvNIcJLj+wJdO5GCm
oPLZ9XEW0O9ZLEFqEUPjn/OCktnxWAYnQCh9ctXbysv02rM+5yRF+Mk/Uxqh8DELmuObrzrYl5+s
Xrfgh2SpD1G6vX8g6Jem2++XMCTM3btMfxAoU8QTE9zqHTs7hghdqX+wrYUWHDKrRrXvJOzUTDaf
mUadWdxWhhVcpMqlnOBz8iHBO7USzMdCCd0/nyPGQSXTvftOp46ED5Y4TxBXuwVFaSW5x2LYDobi
CgnJ36NXrlcH6S8qy+jCA0cvZBh1Y6mjnIG9ChihZZR1lpz2YEJKx5xyNndDQ6c5P6ucwmK/gWio
beyWqM/g06cwNtN7ZzGxG8dECuerhouVkbmEqYfVM3MFjjk1bUYK7fDDAC34rr+0nqf5FWmZT6rR
KkSzekp32ioiprv0PeUZOxYJgLdqqKbQN4Xqs/aQ5/53mi9oz3zrxwJG0lQmUonNYRUAWWVeVGYM
yRXYeWlNg/kkLTI7kJHaRQAKpPPInEIIaUtGLF+tQg4IDSbxxmomuBTeg1pJExyA1JcgQy3oK3JI
go+L4/R9POu6EyMMQM5unPhYDfqrUibrh6JUphrzYSHNT2+I5/J7UAe9mZIkgfmtno53R4/Ix8oM
4vwxrk2F9PuTHAyYd6pP0VfP7QdNsFhCwlbcz3TlRsVpYZz/dshIILWQdyvoDxshPfUx4vlxqWT0
wmo/UpZoFbuTFrL8uMxVdhYcHKbgFTikoG51zqEkNSdAUAREr15ZSMhsaVFnrFth5ySszcom9xqP
iwwdUHVPjxaJPPGZpPy3mIqYOLG1clnb/vJrJZGeKYFIyZ9AEpNL8BY1PAEMWQ6md87e/p7Yo/wi
1xLHxKgiQSSaYrvg6qJm2H0OkG/NI7qOgSck20pFgwhPqSqS1ccjF4nkbtuvTj9dvIj5roYHjWSt
UeItWUWcSedFDEECe6HRPmoqdMWGlMfPZYkPINH01+MmiXrycuIUNgYbcmvgVV29Pef/MWZUBENd
9m/qNZfRbsppvhWwSrajbWvK3Auo3nLkNEG/kj0H5yeYSjNkPzwV+b11oxycrgaH/OASplubDLxS
io6Hj68CUVN7+WC9w4rRQIlq0M787GkGbsVLQEZpxDCH1f17YKcpe2Kl1Sy+6Vq+Zt645G4yIiZT
7yu5fTGvhX5bXfCr0J7i/P4i3v/eZsUdA6jXHhGUpf6aQ8IMRCJZgVRE19v+Z686Gm1oppTKkaJJ
HaR6TH3UBxdUWyyoaNG2bFoTbwsyNf/vqnUMORCguW7mhDlNltGF0W2zxKJCr/JpC7c3Kbo00W22
yJu2nGW2DApk0gI4/OyYyCo2wuNpFxfQUTEd7GUCxvL+a/BpU+rdmP9DaFgx2McfYGLIZxJRlGkE
gCW2brmqK7OT8s4N+5AHOIUt3IXlzO+SjU+r2v7clhOSCHJOSMHJfjhfyK+mo2uHEj9X14KhE3Fp
zrXkOKo3xQKISTC2NVDQslBhwyI6Q24gR3M/y+Y45t7Rt4R3omzkAKWjIgAWoIxVUaC4Mjy22Ogr
0QmMKy1KadnGY4Qc3lRI1iiYbfGScnVcP30zBAjRYRoW6KdZUfYVJqpMemZd1NGvS7XJVfbGwaYR
c8qnnzD1JZqnbaNlWmYjbWweRuhOILiilfNvOl+XTKdTPhRO7qc5OVYm3Qje2N6IKENpV5Johe9A
/uc/ZBW5pjXwvgfE2bGzS1djHW/6b+KkRHKFKz9fZfJe0CwHCRbF25SHgV3OBf+uJfRV8Qq41Q1W
ojpb6kQKhBeqcegImNWqklIwN9cVat2qSIbCPNgxtFrYwapayd9YOvrX7jI/h5+047yTHVZxFprr
7wNScY4wKA/gy4GgAQW+ElGnbbng1/NI/tcGU1vMaOQs3ZKJkaqagDyhcVO+qhsd6Wx1jWJxEe3x
z/RAQ3Q60Y0NmyzgU0TNY86ejhYkJeVaOryZ0sB44dNu0dDnKxEIxf1SgnFtFDNh0jyvNi6y8t8s
5clPJRfSF/+4fPxPc3iJotcqKtSnauY+k7GZH2Mawhb+/fsV+6yvLd9mk+fznwiHcxMw1m2i98YI
b+I3iBYd6fkE8rUs9r6dqZKfcwyV9ZOb/T7OijLHOpQS9Sn2c7hvOaJfFmhiMuJRnX2M60aBl238
r7vG2AfuUuMZiWWGi20XIYeWRjrTnE6wwfqdw8CrW4hriCeJIin8ag5aqFgZcNLVEZTszecLS3Vw
JepbJ2FliSbZNfwz5Uhh7psYFs4U2vF87k/8UucTjVcH2kw8qE4Hs+bYuAYpjAmNStWg0hiHSCVV
3ohX8E5zQ7J5wMea26yX6nyT+X2PZw0nJMxplujbqDIp4L9cPSaXFfv04CtjiESWz1b+6pVPHxqo
1ZAo7DZ3xlsaKtd75NnsOkyrYNRHzC9huXkSHiJ+tklPnD3XoiOFq/6KfA3oiwIzOipVTnAQ2V6e
2+ODjeSbNK6Cf6QuDOuorh15ScdApkCOWJ+4BDzlqKPqJqFTQJ8SJybp4WgvicLixevVS4U1MJnh
Q4/ghWvArGpnIis1z5zwhYMDP7C+NgE6TFB57FSE4w/TZG88cZB853PyeLtT/fiwY82P53G0N8QY
ttS36NkYuX2GXVe3YFwWAfG3BBFadYCY5bWqCtBxnFmogBzNKlECPf4aSBY+yh2vcEdCTlg2HKAX
ZjHCQY+quboCN4MSabiYRt7E8DNCSUgTbe5JTk5V6PoHt8QAFIoiJJ487s5ESQYSZteUPBiwdXJH
jClr+ELa0NV6hWpxAmBqgyX8T3LUNSt+Rn2qRtvLIfhe6ZEr3HdgwNP+kERloevNHaIGZaJBqvFe
oiOa8U7u3ra7LTUd11/fWHqYU75BkNbn/xeprLaBkIxwAvz/WacyOFir76TSw1dejOQAfH0Ku+nI
GPCm6foRzYl2qZ3kQD4YvI7wj6td7/Fij8pG4hEmd4/AHVJkRkNKTcY+PSLSheA+jvrPYx1KL0Zg
bd0qSEnMuDjvpL36nrFqySdjbcw3bBYnyjVzY/jI7LdVmmbadIbw1N1ulRlt35djb/7sGOUVaOF4
s3V2RxSnm7v2ndjTdlKxPh2e7mIb28NICfUF2hXeA/j1bpH3hTDxtlVTNDJ4AJSrkOBY3J8v+hNR
RsiMijdfxVDTx0m4zYyKinc0SvW6s15vLkrRxQRyFq6Ani1Ushd04yfSyfNuHduLx7GMklQwj++S
fEeh3G7kGpSLOeQxg/3+jG+93MLZrHAeqqninl2/aIt00EuXPbjnm1PGYznEdZVS/r2CpC1kQSpB
ikwFABzDspkt0QPlv4gnMbhB6Zo9DrD1EkLBsqyD93hmMTLII9XdzG47Zi03tuzEHr+Gd1pSrvRF
HHRheqKEoDcrcM6yIwiUW9bINFXsD0GI8ATi/HvWz2XpRLw/DgqPMa9JRAREGsJsZqCk7982Bxxq
Q4GXLs/OMhDH248WHm2KOLL9cmiuzD06xNpLtNgv0s1DqoWfU39NAWZ4/4GMYWyl6jJtT3ToB5z2
XNjpXSlTUsHYxYZGovuAI+FDngpTeQ1r2pwNE/zf2C/IxbSKDrRNuE1l2jkmv2P610PnQTI40SK+
VoCVJTmrzFCyZr8WZZcAX3wociw9vGaDBbGjTfAu3aBao33sK+eHShv7ieF76Yeq+OzS20u/Cufi
VT5Rfd7kS3sZ1A4iB4FewuScq+Jk1+PlyjYwAVXKqrDPHPLyATX/zcpZy8PEvFN40duALNpPB7+u
gC0lsnHgVhLE2yiZVMogKo4Mq6Q3HPGxoQ5hZnIQnHeE/sLex5QOy2TpX3kCQEZ9ygQsvuaCF1Bi
T0QEU6ua8SM0LzrRnt7taVPQvvd3BpMMb/paUrmO3yB0L/OHS5fDjDXLNXfTbWTumaulsCXz1ALI
qUs4UqZan4L9pMfRalNVs3Qfg+lLSSEAjgZAxULHM0My3UUfMLiz+prLvvr1FKZfSXpNpLsqtM3C
5Sp2CI9YoL9UBnr4pxnxmmxDamooYRu+BrUOYECFjbA7g7T0R6aTfyP9Yf4mpe/ktEmcwx92Rltn
cC7Lic4hyP/XoUjdPye9m9o1dZCZnhmADEXOTiQ/egq8yEeSTS5YNVWMPwUITQB+5HlRMfmYcGEn
OcIrkJCUYtgSUz7CsKF5xdd+EwIEESkVEIeK050ylNp9i/nBDrIAZKH0wVytdAM17mHLxZtJa8l6
RGirZcJ388iZXhRUJxhOx0HvaeVbNBHrjPp6lJzGCRujiViInuijdCKXMM36S+ExYq3iKCZ3trjx
srqCYlj8c9K4S2Wkdaq1DGHolgV5g09XJEIn+faeNBMItZzXe+vPODlXr4MHu9tUAtKZ+DeGErWy
YMx0tKrgOcTToQDI140Xi5NXbyjF8cRMrx3C3GoLMqO3IQ+WxbHulpzHtgbSrQAAX7xPJb3/1xkf
+1y8x/DgaosP7OlOkOjomjffn3S9/RZyKfKIaLBY8gqIG7xx3941IdnuZWnNAlQaFEU8/SfOTWP+
OlH3BAodXUOATgwtCzx7BzNGpKsYGDGsV6RDIfZQsOLu417NeGZNLPp/46Nh3Il6tVxOmVGC1TBk
G3qa9SWW0OKxSbVedeyCDcTaG4N2kpo2x2LdnAy0FGRqlvfvChZfckfEHOPmIQacKCjRpD7liDgO
gez1UnbTm7TebM3WnDagbVFvinnnbLABkFNjcct4uVtE6lsUR4do1EphDBD5Njca5jGB4WtJhIoP
Lxm9/zUvgp93AGxPob7vbIApDR0S/qGb/JnNQh5Zw4e/oWZ6KvR+TL82VeP3pnMQgFam+mSG1Zgw
qGMPz48Ijrs/wOt10U3oXtv2k7PInwK/LAbK/khzSFJB6GvkMHyoazvSPf+SSif4whsyc6vM2QHn
IsZxDobp/2q8OXdiu7EfB4NIw8WA2LvAa8zy/+IWuZjPEduZy3I+Y/Cdf8rll7F6L9pLaa4q7Uf1
GOqsX9KPbX/ngFwvHY6RdT+goNm+RPFkXEqo37Nb+9F5LL96RMHUt9JVjLWvBuv2r6f0jYllXHLc
2eW+bpgcVI/UMl2oclEUfacj4QYiNlhS0+DPCSiNg1749clAw7jQ7LXeYnY74+Gbx2ZbA11RTBUn
eb39dgKKNKCzIKj8AUyuRujP1t194CLz6rOIC5u8tqyEC9/azOYtLHX1GB7/aPKVn7XTK9tXZmT/
9DMqgzRrFmxHOeC6QK83Z7+ftiTMvqjgj3P4MQyR53piymlr+SzTrk7nT/b7tkkE8VFZlMZPOKIl
gRCr3LxG3asw4ytI9tL/oXfauDC+gbkt9Mgcie7fE9hDjmaSUdFKsKTrF78yqj32CYdG5vXl8x5u
q0pQReXCt80GuBVzmvKWUSMcT0nOZhLWbLNd40xeDAZiCOXmpfqUuLSnJ0kn21vk/57JmwguRAXt
pZ99j/wLyTbRNC3wihixILKnrtUEg/lUKth8GLfeRbG513J3WLhQrstmqWlqFsebV1fVrUb5C9XK
Khru3zhQTWoaJEHDM2SLSGDzQxrs5mTSeuHgjW71NcMx7LCXuAQnqbif/ppy5MjYSR50gQYfA89M
9GNqWerlCqa/1qNbUM5LrqHLIp9nj5fnpOAQLuMTBPpFQLPrBqa55YA+WaEoa4xcxaHJGI6LcnOo
E9H9ZbQaQ3KMNoli6YZ1bLGCWxe1AbaAj31ivyW684L2/oClUEru3KHy8yvUkkphE/en8/0vinBm
Wm7BG+xM+YHQAAAak9KF4o841ZlNyPyq6O7dwBWElyjFNxFdTGVPsF+GN9a7ZpFYFr0DF3fJf8Wa
e7bh4khCP5P3KcQXtvrHknI3Z6XsCPSiX8eZwEwJXQtKREyjktLeT9/IGMiVNpmzJ+1ubklbH5LQ
tDTphwtliywKXU+VqwQMBNIPyr7XKKmZ/ohgUW58WtcKFOWFuZtdG4JC7flzhYVGD1juQ+PndLC1
xJhxGOx448H1hMgOZzq6Jsk8Tnun12kY69o9a7fXQzCw512oVCRpL4BGaEmrqaflox98o4h/Ted6
GkjivZb/0Tv5Bs3p5WaN0+WC/BOujNu/8vC8aDXPmu7LRWFfCo/PTLEwPLMUEs9YqXontX911w0g
W8+02b4ZWMkmeIoRMXpZvr/UmNmV1pInXLNFeYhiN1FHcNyMHMg4IJsqsclPfddGKuyEJ5hbwzze
UvIbhtwdkYB+OCn95r0TMqetD+u9+xRx6OHVW0v6865DftxZymnDkLUQTmbPjzIU3DgBRC3oANI5
BSpnU+z3x/kYkRkKfHLmbaIaPluUI4XC/iLLJsqV4VSFHIAxyGBSJSFarwgFttYgJxXwmFQPFXej
NimNOa5b4Pv3/z0fygxxVTyrqUYBd0lpB8FfzdTvXLL4wEhsWs8HP2CZhGIck8DLAnubGlx1EKb3
ZXBBifiDx4TYmuijvEA7UzugFM22MYG7AkQw3mnJhDEuRNAEzuMVL9/0eTqylL7klW8Sf1jHBQAW
Ky4niy5xtgbjL3O4KBckVhAiSGi/+wrXFwwdGDEWkI+H8SLHp1WjJuB+v63XPA8YJu3yvU+HshTI
5vHP86n19m9U9RIkgvxz4MDiFStvNbk68pOQtZ6FIQuH9ScgWWWJHCPIV6Bnb0cZ9kdEp1z6Zt0e
eH2i+7u+7bs10t1m8VXdb3ddxG93pxjyt/BafA2DQfFm/4h9zSBsZBtyuToEyURwFuNqAybTaUQ5
UDWwuXJiNFsUZ80D7xMjGqfEAfgBM+W6e9jRZ7HnGfyCz+aR3GcdwzbyPjaXXivmwax2SE2i5enB
F3V4VzmX1lfcs27PQp7AjkJ6UuBk2GCJ/zBDULw/YhW16agviL4tN8EkHY5F5nEibIpMCKCCTf3O
uPiq8ThjdYP3GoXCB3eiB1qntWPQgOXgnEtH3deQ/wgGg4NJEhp5l5o9WMVSO1wmkAruGu7u4iN7
mr0ua+T9fo4Q6Sphs1BMZEMrtHpkiuII6iTYaR0yFA9ivu/j9XohYc+fA0AzYbKgbl5y4yiS/zPN
Jzeh00GzaJ/OGPmHFXEw8W5vURsZt015I9vAHW855DAOsDazXBXkeUz7YI9VNQ9KXrr1YA4C9r5N
2wuT15Is3rdhsPKi10SOj0YuBvQXfSDQvhctM64ziRH4gK5Tn5POzTfY2MC9simWSz7gYHD5KXAo
YmJj/9fUStZSKDAiu8NmHvg14iRSegPqv4uycy1vIA2U4JwJM/pmpw/GD2YFiCEbQy0pVSpHfo3l
RBwjYEGdixGtE7Ty31qVNPhea0VEB0fm7/IzGIhebKINiuzwFjqwvR/F3F5HQyAunt+8VKiF35/r
RGfw1ug94d3QQqaiKMrOr0XJglC1gDNw3lsy60C16sXhxuw4WYgf024Sz3LOtcx/ZQKO3WcOEQyr
9aMRxD7DTYyeKYpYbINyNvbptwmn+rj+p9bVyUTP++zBT+5D5gIay+kBUCYtfr068sO3369iWV/7
HZCsLRSKB/Nuwa/6Dn3rjbxizx0UIqnMgubmxisq9xVt1KPElWugKtRaULU1rYvd6fUjcJ5egq1n
vF142OivZ9LUpKhp95f1SM8tstFr4I9+R2ItZan4BgAUcznCDJtNYtmz7FUoXy+WgtLv+2YbUvYA
Idjmm25fFJFryTiq/man9wT/h1nV7uN8dLY5X5Qko2fAZxN9B2lxhSb0hucFZdiY79z5zevLOqKI
8UX45YDMZFMRmjaz9zrMwRNLigtI7Ap9lY7XRxRMnkjmFDiLMUipOYS39ukiAuaVEM2dLNVTByDx
coZbZDeaPPbb0FWMkTmC3qEonxCMVZNKF3MMqPEuIb5BTe+kLQHhLSvMoRqcUhpFFx8qNS3ZLpTU
2zAnT2NB8hwqKdaCSNSWtLQZepUYQcz0dqy2y9dX5H4JmE2InCWG0PK4B0K/ucirlG8yKXRqn4Bj
w5etH4fU6rNQOR0lVmsX4VCwHMhZilzzhxXux6yPlBfl3Z4o7Jn7+mqDRZtBO+iybnFgQ8K0JOKN
d4zZBxpsk1VEDunDbNWON4ESH7SGaPWbAJpiAx/P5keHbGzOXpKvcOF+hiV7RVrhmxMbiIH4NWJo
bN+yoYKQv4Bwuu802VwmxKuBfCwJdklVMdLzDskVnHUNYWeTSyvriQB/MSZUtPrF3G8w3UMFeUQL
SJgPKOE+OgGJHi9l8wZqRR+c68AnU2qkl7IJq1kSxw9uTK6ezJWNFFPC1XOzPEbdT9Oxr/pPnZPW
juuA6GlGk/fIxShhJk6wh+bVGarA9a3x/7+Re1XIXI3BvgkBz9dbDxgNpZMBO4vJd/YYSF5//4jH
z4L/0qz8nTWCzOKvMZyWJehAMBf/mRxKkil7ooqBeIeMYzwIsFmQqE8IDuKaADCfaIZcTfAvxL9/
z6CHQkKJ2mhQzMK5IZ5bxhh0wGNdU2WwQui4lBg08NzuljbkhTf9CTCeTXbQ2ajgAHpoHyB4YYQe
jrpGgU+6jrdZBQrxpWYp5mgkwgb/7H87eTL0QDmqLBeLZUCztyhiUY/xblE/b4K4Tt8/ANoRoOux
fvCWQypJq4WHOEXXSFR45lkVLR0vFcxEglmKj+dhF/3KoyAtYuyjsHuRXyOfV8BdLCnPtL8P1E7o
inKIFrMZa405qCTiFyo5Ol02RR0u0dYV1UIVI+9a8cNoIPanuvX9dY/2L6DcI3E++PMv/l4q9DRf
pwQiFk2b630Pt3SkWtmkwG2peNrJkP7TqQY8UqClx3o6/SkB8FvCFx3TmGSSq6pwN+z5m/tFxD56
9CTEzq/KYvYI3sZ0nsBfte21SBo/vMUM0DPeNpJWnwqQfdfdPaZ7ro+uVfO86ehsjdDC7M4CNbXn
Ezmy0so5zAWvxiUJFUJU7GLymSg7fwZwnlsndVSxy7vWDfUL2UMeYCnIRUkHvt992t45L/q5fIEt
uUexmXPYwLj1wMiz/IrUXJreb+paaPlv1m2IwWBIjTOy7cVZ9m8k40V9b/AE1jUcq2IFIetqsu35
zDkKzdj7bBzGo6yRVQaCEO/AXy2zqJRH4yxaBIhXHzaBRTzwpTiXPvas34NxPypLA2cD+Gv6+LN3
UH/8RBzuj8+cCR3pBkNyYx3+axTXgCS+s0ouyyAxNcaBmvnwfS3FUCBjVlnS+gIxIVTpVdoSYBfZ
y5siSRnIf+Iq19L2/YwqzfxfwWFuqmnq6SB0FeZH6T9fr1r7Mr7zAVT2fIu09B7wjvtc/fdnKTX3
5p0sTP177BnYDKEkT8hlqBPBNqebAVS3Rede8BHvsFgBC2w4rjikMvgiP5WZra4crkWWoaJU0qph
nX6NL9icDwEj0TBCEsyo5PM1nxDnQSm8ZTN5q/W+cjCj5IEpABdvywhp/RY4Ehd7nzGrRRvQkV4U
r7gTXD0P6/lXsAIuboannK2PM6DNl0NK50q2Fkj6y/7/u9qdF1isTiOnYZXgSf4I6WrdpDq82gIA
Ie40pJzSY7VhpgnEYiIhTCs4UygJP+bbrez0fFHTWcGibbGHTYlMbDDYBGskRdd0+akYwiQ5M2M5
zXUEKKkBYKAO+V9F5GNXT+tQxitNW5eDxCVt2MYqnte3hb8gxqDMR1Ylygs57kSD8x4vTp+xXrif
br6rZFyIdyvoNcn+QH1de8nP6BQhuvCiRkVAuuOeOzkZuHxblpiXBNf2EwC9FpfKh9L6t0G2Gms1
VFMEbKHOjnATZDny5/1zN7sNHdSKfogpwu+U9N5RHF6tgAz5iRCM2kY7hgToQQsvPSceZIAY8XfU
Jb4X2GPhswXkqB92Z6DM6HMlX4BUM/EJQQfqmkKUsa1UXLOWNIXGKguysiGzNQDn7JQ+PidWfTei
gJZ6o0yz7d2ypgSnRqYXK9XbRbgDzyRr8O/3j0tng/Olojr5vgdZluHBFIEJ49a6RsImV1t7RQKX
ui42six9LiaMZ+fOVopnvY042uPKzwh4CTVotdAwYHfrIk095aqii4xvEhkbMZ0lm0FkR6UfRjDv
0EwOG9TwpGlaKsHj1DNT6NIHFfKi944UbsM7DbLQFapYAL5KZ8OfXhPJAMK4GMaXZPDVYyhi816j
J1hNDIl60DSeToECD9NHKZurORbeUv0A1M9aOD4YrcTr7NxGAMQwi4+Zs9b+P99BNM23axf60rXx
CJALwZpyPG6dOBb/Du/UaBF5VBomkQhczZMxckXkmcRP1tLZ1jpkdI7qhnOj4H1qSOWyWTrB0Ke0
xIgsCg4lv7mPzSp7Gqa7HqXxAH1OHpq282AS1FfMes2cNekUsMsjr+X8bNcZagKDbm93YfqnXpBQ
M3oj4wAnZGK2xuT0Lk25E2llN0b8aKDjD1IuVdSSJPn5ADtrS34rv/MTUWnrBj03kxggg/KvkDio
qYNfN6iRT/JyIy4LdIUpt6G4GPZfR5c4zxePOhHQAtc3Xh0jAfcLz9ZjeAzvsyQJ/LCDBAIzaLxT
LC7dQ5GpsyO4G9cn9ZGeB26VQDpf3KnuhbVALOYlIrhyaf1/FteA+pM9nPAA8G66c5cQB3aHtO61
+iYfNC3ZpnuuY0rjHOKZsZnmHOBQhh7t1b5wqFgVK+u7A2lPu/KjXx9AObihKw+/ZuqRq9/ci8SV
kHHyHI0rzTxafONLMD6TDJeydfrT6hB9A3VJfD7p6PgjSoxbj1DKhV0cA5dsij5Acb9MctdM8h2g
ER3p1DoTGFTakZROyvPUnj+oeKcbhcisCwyTIikLlumOHwx2t95F/bWWmfyUszqr7MGH612bjenf
ObjShtPI1FDyqsORl+ktECkaI5B7EbeRMSufzP8Cotz80YKkOEuvoLt8nW0K2ElQVxnX5YAqcwlo
/KuQ3XgYNHnfvR2LkzLQpxv0F8H/yqB/xitl3X/VtgAvAjKzjN5PsSd7077uSreHJ9HxXSU+Bmfb
z9MtlxCxCSJc7AQ2xUZy2Z5egiRXEPB5vYcdj+/BU3JnhssS+4rcIePVp9vAuJeMy1UuTJZEbuaW
aghzjf8wbPwYK+DO7psyYoIZ59KTMH9eyFcHHgSaL3YEfNSeitlrCjRGdP6IKsLiQlKlE81lvDY8
mOABOjDOesoIHIjSExpMlT5H5uu8NHo9lk6g5Wiba9Y7M04lEta03p+52JAD2f6deh5LSsQ+9lkK
sRJVCNHs0VcQQ2gOY1OhzZZuFn2XY6apJA9ADsDBb0oCiyQ656N6PYitMlSL7fBrmeK7psVBP2Lo
GeyLi4tDZeloX1rrthT8mJNbmdwmQjvLFwKpr+uQUNQDD35R8NdZ/iFOU175rIZEEdyPa1kF7yE5
zPH+KDtAAsCqXsJLjgVROSD7athWCF8uKd2KBqPF9pkNEQIfa2EWhyBEB+mfFfGvRvqeoy1yYIL6
y3r9u15WL9iec4+HsRoB5Uorjwl3emXzJvHjhx3iKTv7ShLMs3QMo8jIZBEUP7YRxZolZY2zxsZE
bl0XiMg0CzpZiVBhRvgvr8nDKjBHbC/+8htqstjB1RxpuukrDpPGhMGR1CM3JMTreH77Gl82M8fL
1bwX4BbYq8QC/phYOLKBzyRiwowzNculQbr6aH5BvFiUd22lI8Kg5Iv13gSRU5zkOf0tnAoU+sSc
wUuQQEbS4achiSce7yO5ihnAUzLxvK//Y8cdGChAuZll1rAuO6aC1Y7nABv6orRDf+9SwTz70kkg
BeKBBGyh4dudZXKtm7n9+8ZO1gug7jqW/qm3ydWPVXNZWj28h7AvidMwBtUGTyuyD5k1EK0M1SEw
RlPathFM9wdHwBNX+XxnDu6N+qONi2kfaEmmGzJusI5RKVXOWKLsMfUslGNmEfqJXKKJ7FRacxJe
4lQ3coaVs74umZjhPNDtbty+bZ+hrlD/GIPPPUlUa/3yfnZhLE8n/wOi1+9DNP2SrajXLdDvxIeW
Vb1BxDmM0o+PciIv03SjJ1enfbpvPYjcYxLwTVEnrOBvFOJ7KOSfjvjZcp51yCUEOT00DjwK0Iv0
BjRK2b/hxrq7b8xaZgtav59nqhQnZIS2asOfHHfZyR4bJImDS/lhNTgUkdsl6GWnCDlFbO9tds7P
sx/3+I62ccVRTJHWdDaLsQaAjDzeHY5KIH/QGOze9KaepWAuQ39A5S3r1AneML8hpuDTecfu0ldH
qpPKBKT4CUUefssCF/Y2wT5TrU3AS5bREnbaovXBieCmjQMHbTPBAZ0+VgUpae3qf9eh5uA8xYAW
YmIWbFn38dMNhj4ljweJ8INUMnjpyFv6tD852cN7QCSlo0vkiPwys87kYj6jwmlFUP/C7gB2o3CV
Tyq+tg0JWUfn+3oeWE7fZvR4q23XYKfzckjLPmDb53sjjnT69+qARTixgPTkTUYxnBYpdfzAj3Hm
b6AW2dLtTqw7tbb30IM0g6L5v2PiMVHgeP3rADsTwStcg1SZ0syCay9UCpWsrefEqsjVxxqTFU7h
05+v/frQvehUZfYnryOhXApw7Vz4wo4iRyI39Cw0ykHOgQZ/OoFmx6jPC/YO9rarWGy8cWMyB4Ld
FbHbC+SpTZu3sFKR+xo/TNKZLBpkFdAvygo8Kfm0bns1WGqFHhYgC71CPLFDYkt0ceEnOhJyeP/0
9N46qiXpD/3HvOKKuEsgplCAD4cXn98naxyHBhuBKjOVP7oiu/5arJlX8SE5ayQl6FTnPk6TtUXP
r96JhCT3NWRXUTPsBFbU0AIjRg4j80bf38iXzX9IzMry9floX3v7cko83xc2uprKyu2XKlY5vj+f
W7iFKgNkBjInHlncJbkJZIQ5O/V9zPF2KA6xA81UMqSxe9FbrthJWfFTliV8IWG8mD6JecwXTCUm
EZs5YgPPDr822XCHsdJm0FNAweTiFi+6k5Q8qD1S9e9unXGgsnCwwkVaTXX3c5RGsgclP8n3Kepo
CIO/RP1WoLIA3ZpoA7tNlctVfYLcGLGMfjGiJI8Q7x/8g3o7RqXXJBu1ZqdAevl4DdDf4XsZIzXU
SNfalGbjy10VcELkNinvmq+aIGyiVJ8l42QhLKV455sjHqHLh//gZaZ5fl2e71ZWowb99ddb3n97
t4oNcuR/wz8NOho8HooW4sgR13wsM3Ts86ZUU6J56c1f4qJl1ro82bOZgJeuWW23hFmEZUg1ozDA
Z9e18SWmueXfo63208ISpuIzJfD/uVHsOjqKw6I/EBKmlrLh632xEVFELjNC3p2lrN/oheBDb42e
UTPb1f1UiokDmdj/JD7vLTD920b0oB9N7hX/Rh3rhMopbb2xlg6Czusx0d9ajfjpaW++dXjHYNaS
haw6QlDkshrcdf7jArDS80i3l9tj6ScJ+f6nu0V2Ou/CD7v+f0d2HwfDVCfdYKDatMFcBIB5Radv
XCOaUoLYgAolc+HNG15KI82TUL9ZIv4pZwbGqiX2TMgVCRksVhE4oHZWNcFqyfsq11lgHrpGPBaB
UoFgOGkRcoP/lOJnVpgGV1BAHNy61RqgDtzhBL9T4FznP5oXzOGo6WxM9unVWtZmeI3wNduZyEDA
CaSxzU/+tKIfxZDR/WGhY0hunk16zOcr02UUdi6fA2PBCRHRke5EcmR73BpbECxP5wnZqDJZVioA
P3ul3ZYih2dFkbktIRilR2y7da4MDRmH1bFvWx/EIiPAP8gpEhC4rxKmqj214EQ1WOy+xiCSys3I
OYkJi0YYmF7k4Mkuq0sz3hu8BC5ajoiWhDpXh+UTkwZzYNEpgUXb5kzjaCPH+Ml/VFks/0Ciuihu
IDrvBzy8TrWm7fTrblWBI6/K1nw+/EsSZoUvfkdlB3bv0ac7F7OwcXZtzkhEULi6stOWXrTLWs8c
2KvWZgESuMaZ5oXKb1ca7+Qye1PUyEZlDijmwyLkTUpG6nLeNRkmSASE0WTluIPHyfhlJhloQlCR
P7gGlwWWMIHgHKUniMIvmarPVK4euGViC7AgHl2aQzoQIfSYztAs6p+i5Bxw8KoZSEckdIdv89MI
rrj0HPy2ewc8RnldCpjmyaIRUEVBtEXh9IEk1KKY5TIo/y2w+wUeWVTINAF5RT4J7xHOXBvRuDFm
Yn5jA0HX7dWc7NIo8WJVG2PCPjBd1+yBXp5PiBG+0NDcyaBPVGdqh6DsToD9iuhKbHlQJr9CF5c6
b/ctTg1wtsAgUI8N1iHagxjnQ/H8qJGnU2h1atdDe2s5SwFshY4rRh2ziN5Bu+KoLp6tBHkAfnhF
UsfoO9fu7Nze0Y/RBn5d2W3zUtLmeJJLVBkdA8J+r7EGjzCubtlP1m8FI3YnQ6FSyTKL6Us8Bdud
TdSACmkHW6whBKRh8nzOsIUFN6V+ubjPAqG45FOB/vxk5/sKSwmKhGJPKYWH1AnevIKiZmxGk4BP
W9qITjhACIwukM2tyv/GvqKojRbsyoYY6j+SPnbW4Mdmg9UzDKXepYV5+fXNvVFd3fY0TUA3FS3x
XDHBq/UX73L1XhaaecBTqiamVC2QWzGpP1KI1BzlXdYZ5cpeiHd5LJqq+K1wmYkHh49xfwCXbvGm
H3oIzd2U2A7NuYWMo2tKDmwmS3GyPeZ+rkJ2jT6UhptHvSGXZEmJDEsqKBsuSMkNI41yQCzLbhFV
TeopWHigePwDpkc8PA28zN2eTos9WbBJaWnKHMVBqZ/lvjQ0gwGZBjrStSmHZUdNoArqEZ2xrcPD
XWpthwtoRB5N1BBcj4TGCz6bV5nh4KG43ey0gMOLeZl/qcFxPFCI8qqLXQoD62BVDlD5Aa+tseWN
8V8w+zebHSWXQ7hal5T4a/tQJ3hkxDtbOL4c5SoOMigUt+Ne/tvqGIfpGsfvj6ADXF5ypUerZyVT
1AhjT+zb/bJpnGweuNPkucR0ftmutiU6N7a0rMKSJC4Han5Dg4Nktr5WvM0yze3mPCtxoD1MDd+m
kCGTzblaUINeS6rwFtVPegamtQfKddIWCeU9JVpMdmJNyLouMsCipGG/6qsVbVODv7RMNxt1NZCu
zDtnVT2fZv6nk992d8WLlXO+VQnfK6TdCOG7+Gw4VzxgxANfpl4MmppTicykA63Zoc3m4huIUWFF
ZGQfkXH2Wa/LOTNxhpiSzoHGQ/VLypys4s/iXFB7EE8TOP7TeFZKzD3D08ZSOCc5uYlWqgXfBUCi
l6w6Tf8VC3ICGj8vqAqozQCq88/zMbvQOw4JOWfj5RX6WSyNJgapelm9AU1FpMhI1NGPtbjaEYb7
fYDMwIRS88LOfa8ey0bsO6EzIgh8eR5zb+vWhygbZlJ6xzsuz+Zcp7ih9YaCkznPgL9D/U7LkAzz
0OlTvTm28ese8Hwxd4VgMM1MaIJmdeuJbx4Z1DtDNqkmvQbSrOoXgR5CGKjGI2+GG+o7hG2zqTC8
LcA/JLe3u0Z3GaDky6SrY8oGB8wkuFdGuVVykazjBaXwTqP/utwnyZnbjXlzTWwkRMMAoTx+2OYB
Tt3u1i854EBz1m91gk3xu40djWtat1y1Kxnhhn4Q44GcfLm1P9kGe6/n3YD6qYyv7X5E6/My79tv
P0h4Ibk5WU8+wT23B56OsQwPOGxu/fyb+thPEZCnCsd4n6SxJL2kQ66NSX6kgrkv8Y+qofhSTe2i
6IqvL+2MreUFKhNgu6nj5qvAEdK/HcKEX+MzhU1LaU09UMH2HfBQzLzAkjciGD/RAKw/dCOrTY5I
QSKDdr0EhLdZzDMFbi57/cIeoOr85x8K4wwDNQfQpEclG2EW4HaXL1uuzbH5VjNcxNDL5+sWvf/p
JQ/+Hn1FgKqeDs95A/YGon9evYmq03hmjnKBqs9XckStEgPFVjjjo9YlbaDpF5L+g4vS2ZnB09vI
Wm2RFm91bIfRCjjs2/Q0uXyrTQp7vhWqFBrJcY2xxyy54UVBIbDJxPl9SIwqEjaqZ8oauDG5DoYO
50Ueu5fZxjpDd2n0loMYlZ4xvIH57giRkrA5JElixfndSRD8n1EJdKUB/jU6JqV0MXCK225WXeEL
SSD7K1GsWZ5yhdQAfmhs0e/kV59Yf+6Ye0dBTvJstZrg7hISG8A/etpvD83eH7+V4V2xWGDwDV1L
reWjJlkdz6uHO7JbRjYXu2LsHfphC5dmngTDkvljJKBRQWfQRP0vs7lX4GHtBbJSKpjNjYPMXuZo
NpE5APy6a4FgIjPGw9NkX/Jnye+CTl3GLJIyMSDDHr0Z8Fb5vCcxU2KCVg+3tiMCAX3vtZ6anTD3
nz0llXFZP16kFFPQEfkNxxIe3bxx4YAI4zx1MBekJkLYNnd0O9lhZjmnweWTQ0/3QxJxh34meGfh
XUiI4RAf+iGDCp0DSZ938wgHQcVr0PYol5wl/erDoBgXkpvb5ab3zieEHleW75dwR3H38YKay5N+
cLXHxZzcMgbQX6Da82b7GmtZIIm2ilDDkBJTBuS9XAcq1CVK9gnylI82IKLrPZoWXeHu1UIrpUtd
1Ny3eDBu2IWLCoWJtPQNHOhydMEl1BMFgIPwhRWqPbdtgUlpW9XGrZMgYl427Xo5S9MFjuV4KUbr
OCHyhyeE3fE5rwBRwCF4+Zt/rI9RoT5G+XfulVRFHlaMh1wfwGeOUJpDfiipgfNuEbS2YM37TTFp
0zvTRS3Bz4jhRF5gBDDR+6Cfp8w9nA7r+0BU9HLojhtrqz5C/QICbg1b8Y/n4PQHINy7uAwN/qLa
G3t1EfK5rJeFfW9EfGRuR1svT/yPCsBwIhhylPzvIcofFCuVIm8XGRKV4c+Zmo/2ljnh5oRn3bpv
7/Un/MuZ26ZxauBELWNiDvuK2VegBzNz0c2fIsMHjSsADVrG9KFqZJZ0hA+1LDOF8uiB4iGQLJS/
Ag27rDhHVUPZ58WOm6GiSmxh3qwkurHa3xUN1knDUZJRghzoX3yg8F9Udq7OzCufp9ryWc6odD6S
HLbEa0aUieczdgh/9Be109JJDuq+pJClZzKy2N2v8h50MaFjfyRuRSAuRJxQN4GXmFtTA6iauyjo
4gQXyI2Wqh9gqq8063XERRQj6xtryX56tQQ9z8xNEcXZ9eCNwMk/LwQlZPcsy0aPfYObrvA8AWBt
ylMp3Q9NVeZiwp2eMLvnXjxnB20i9/9XlFQOLYLlBWkxe1Vq0g4fH72edeOak9fe49D64iRrOhjx
/csiAstDBeinbGaxtPaHySPw9ywqWjKs15jtuvDrznF7mB2HXOsUVd4iC7PVbQRBjGwNQhHXw186
9BgA+vJLAMwH0EpJKswKl8vJVr+l4eno9f5L1hrq5DovEhzIE4QJnmGG9VzrOWsR7qlB3JVHT1Gx
dUusTM0Og8BLMYm/Aata1QUWELoNZyjgrGivEkeAROeNQrzJ3uZde+K/3uVmGb/6AUFPGhOjQme5
iunRlOngXI1aHsfM3LxayQE3dAy2/rWh+EJzxlJR+foIWAS4hlHWNKYW0WULoGvyAU3cjmUjBxSO
8IMyEcXt1SOx07kGamvR09Uz3bdF0otGGq8Cp8dzklZQ6sUEJQeSRVKchZYJhhAXqZyrtC1F28w1
U0Hy81plqeI+SP67qekWrYMJlpQthYHK5zx69K9QDsvBX9/wDxmRSv4vmcfoFSLntZGK9j+eraJN
Ujx76Qo36KXSjGLoRsfJWvWXC6mQWWhxJDxWdTtGpneXZ+5UaWRk94gpZ/31qgsxBsQp0PNjCg2n
8ljqCtqW/JzvZKnGJfpHmwF+GhTbqsfpsFQlkYxtKJUDQN5Hze3mI702ideaYySAo3MRj92tfe57
dYrjdJSt8mHGNU8HI0bX9jWdiFQL5wceR9jnCkMuf8xQVvxlXUonY8DzYiYzFh1onoH3gMbil/SE
lA4/hE85AutOsBuA+7D3k5/oVKUEtxCif5BoafRbQhKdX5LW708kgL7hnsM88xzk03yyN6fbuOxE
j932VObSlNUEeII/ecUb1QLjjyAiS5MeUAoQGgpQhy01pOuPRu7C17ElFi+HUfgtcSemnNbPFZZ9
IH2YLn6tOHgjOeT7h8/20Rldok+vfmYt2hBtrsxHYffKhvTHpa4TCyt1RiHhLAIsCB2zXzSQx3Wh
dBEQ5G64b4XSCzmnLn4WLKQ2d1MCmVKhR6mz5sqtn6B52hEhQQjdnZXUlNF4Sm3qnSlmH+NmwHDc
TlFa4RMzjlrs0J4WalLxgxVVkT6vtGBZXEDMrGA4h16elRrlPnPqvMqXfO9dwmKQfcGRpOnEOvE6
M20yGCAHksdGce0vFFKq5JcPJI3fc7yay0tLH1Rl4nJdrnGm/42Hqcg4Q8tTXZ6gjlANgwQKQ7g3
kGyU7tu1LhoFdyMyjnJk9PDi5Z/AAAAhVhI7tjfcd3RmRstLI0aBfK8GIZ0ZWFbp4UGDNiO7bTqA
dv95yNcwwEDzyoZGiYfSPbZXdOeApcehYC4G8ctRAGISSJnndpk1uj0bPNUE/SuEdKpiqGjQqvw8
CIB6mDijoq1b0Y2Q5JqzDdUDXv7WuptK6fzqZg3NkeQTykSowmUZLLRFzQi/Qo37t2PHiPl4nNZo
W20V9W1E2Cy922QwEs1lUn82u+IWSm4yxOPFfCBaD89HHduaLos9tSYy41PwixAEKg3azsCo1inY
OWCc2ee2qxr6X3xcN8zgu3nuSE3dg6r5YDQ8S8ONX34pwLF8lUzZsLPzoPAxCC3QGA9oaD3I2yP0
Yy8MCYnIuV2EsJguQNUqc9Ngj+Xq21OblXkkmW0GfPfc8UZcIz/wruoqLfAzeC7bgcfLc7jFjFL1
nFSMrZVJuRrkYfgBSFUKN1f8DNI7dZ0G1d9RtllBz+ZwQguyH5o8z2F50BtVl+il2oC4hGfV1KO+
3BG96vOn4Nl/+njLcW3JbTxcDhhfi9h0sc19Pe3TEr/b//7on7pLghJdpc3juA2EEUQbaTCTvDcs
GLv1P/fxSOm5+ivglfaeRSg5PLnDm7ETBjARP/KslebJywS6ZuE+A4ckFZHdyXX7hbkZjMzn2hz8
bDbyOiOKdSt+qdQ64n8lKAwMkJn0sdcPBhAwWnwG2sKQPY2cOhI68yF5xZOPWntlGTa8NsN2lWsA
aJT3nOeluGCqqzr7tHadDRgys13ed1s4jguH0Oj/RQJJ/aH5g5otFsXGMUw9GNEh5fJkeAmaBY3a
TOCmvKQelSrAKG4l5oeDJxReauM6gLpcdxj1EtmxAlgzQYjO6ToRMmUlXJFygBAdKHxckzf2qXN5
75MvTDbW/nibLwKPMgio3JkMdT0PQjR/PfDqsd0WoJ3TAXMV6EyDQfSWV/WFD9YjPUwLoNFyd2nE
ySyizpY/egD8QkOJIiTyBA1ebFb8agmhvXF7qDj+Qob8KsTdeqoIQTYnxPevAFK0QyUCcAhuSvfV
+ldJ24IIN6Y0pBzkAjttQmNJu3XoYHhTk+QnnNGHyV/I4DY9bNMjMxmrWwVIz0cqq0DrPamXaOXU
M1Mth+NtdA0snCTmCQcls8SQQSm9MGTkXS+XzQonatSVpVc/Yjck+tnVoYVSTH1a2eZA55khI56k
k/T0mdYaJ9jlu1vpsvAUPL91utJoJqmPbD2TrnbTCb4rQkUfweywFUUrjziypCpMSoMuyaRW5+Pc
URmGg6tdikPKhVcKpGwFKiDn5MGDUMyxH964nYRbEEIBGkMecE5vgzlF2X1SFo7EHIXiehU2sARQ
pS+mp1ZhIxquDL/8Bhg+YJLcaBzPXHCEUCqInm5WBfe7ORwA3K4Vf/669TYbzv54+U27BpHMBxNs
YA5opl5DNebH8MU6zbLrENvex120ho1H99zkkH+1zFF9drn3krUqp/sDzbcwZixFNoVyhd8wRZzb
a7NUddJg0Lc29okMUe8Yl7SN1vEHTj/LdpB6GlNH1hGZDJX8QmsbHqHNSwUF6L5FiNjs158Te0V+
/EK81G38nycmPLgcLzOKOOxJuikds4J1g66MEdDmsf8V+8s7njH+3IJKCmIwRyeddxGNDdxPmD/T
7W9ui19/OlDz13+hHvZ/aXSAqFch+TbZLnvbl1VjDEFpoB2KyDvW6ry4K64DznzkbkmpOvB9RM57
mAnYNmwQZt8mCIT8uJsHcPLkjqo0PogNHcQVE6Xcmyo9mXnaoZstl6/iAO4fpdk3vl97yViMHXZv
1eVD3YCglGtm/SRzvlVbXsNKM8HlKK15dEhFQhWEHeMunXsu4IDqX5q5n5Ez4hGYDf7B3+PsuVUp
cLX0kf4olxtLquVea/Q6Yex/x4HeIukfbDAM69FzchdRCeyOZQZPbVxPWoBJIUKL38WjWfVu2ELp
T0cjRPF5mg2DZhivgsdrnVot50MREGLBcNCyutjDNn6cpf/gZc6DCblbGIX8dpQOePa9HVQ0XGS3
TsJgwMkHiqTZxtrqeILzj4ZInc4OM+Z+GLmwV0E6j9YXe0UyST7nqF2GqYGrFzcfYSyhhuRUo0vS
5x6NlLEVlsI9eTEK1am64zLuPjdLIkTclksUyHbXsADghJIaU4IPeQMIIQgDNZIj7x3i/cmipaDN
QGnqip0eEc3+ZYYzo3wQtZRbbKlFuigcG2U0aXiu87nEyAoHIRfcBlNZqPh6prSPXZ712Xs4Vega
/YZFwDpBPy/nLNDoJJwcgvwxGI77XHzBgiXj7zECE2lDQ3SZacwM6EjMmxNu33Z/kAjgyXonm7vH
u9UN/CtzS+CutjvBUiqQw++EwWsiy1r1o5IYCYGWLhs3K0xDfeC8shGqcKiN8deFRgK1Mo4vRKwB
/5gcd2JaEZMbhrIyRAG8aAm4yNSl3uMGDRdpmCszwbTcD4Ia/AXYwI++pgQ6SVjtSvxzv7MiAgSo
giYq9G4489msjNyfVs4zEpWChtIpJnucgVm6K6XKj/4gbzJy+2BJ3VpMQwSUAwDAANK/e6od4t3y
gtY47RVjTRQSfsrPF/aLtF4A4YkTi3bJLa77qSbPxN+9FBxfJrpdS9eQ9qcmGU3UPqcgYdqLhD5g
0nvhGW9lQjbW1f/Haa9aOhNgv2G9+QVZf0IHE0l8o1SmSTROBOLuyUzPHSLvsQcAsV3wJGDlXG62
CS9I3LZfFU+7m0lAhdBdugFXjrr64gRFcJ1g5hbSxQEFEGWWyWnKvsixfpououWRh3m+KA8UFTYC
c+x3cVzosYWGWqMEXUN8JJZL8YprHrM5/2RF2b+Tfyqx5a077xMiab/IijGj27rF3Qbb7IIhGZen
eOM3Xo/TnyULfP8ilw3PFoSp+0dZeYjPhlfHHGCLDfUbyADsarmJndYiqM4MB+6FH1Lbpjp3k3df
u/ZShTX+lRycd6omKGQaqkXLkAs8817k55BihNyZ3WxQA/FOzJoZcD/q4L0TaSUH11CUXrd1QhTi
tPoxsIE3Zt/kndwCnSpDsCikBGVodmXz/XQi3O6lKsVjx4UKRFqMUfz6U+SE6L123sGjo+kjrcK0
HlABL5wyHBCNhGxGOfG+NCLS9qXN1W1I9JBa1EucoiQP1BEz1llaJhNC4tPd4cgjzo2zfHUSG4bP
3LIlb+o9rDgqf6L+bKbCwlrtY6Gb+UFokSRgk/El0giJY2oz5QoJ3lWXDQEMkFLsRhw//kktqnHU
R/VR8NxM3PyWcznqrgYNdQ4CGTizN960kbNk6mdLuTuCtoZqWHsDvlUznret9IFdEbdXqH/qQRnf
cSoUwFgUQjpYcqaTIPs3CW6Nf+X6bqSiHZA0BVsd5i/jIqWF/ZpOdKNYKEoIzon/7x3NHYPZI7Kj
SS500fOpMSgwLAGTSuMweMlJ9yCGrsxqXibazqVqRJRuij8y+jprBRE6hTM5B1G7nDxUfdEppTex
FfzdR7Xc/O3KQF6BEW9GgSVdZnjd51EHtAwP9B7zIb6dPejE9k3nvWzF5XZvd1p/CF+31HW0kuOk
q/ErnzV48KJo5ngBNctpkJRtKhNa8fasTS2FdRnEgHMC+kSlBTZWcOrkyAWoUO8w5lTP7B0PdID5
P8ZwvBI13riD1jEzvquDhn3iyat6DuUIdYY3n0Wl7tfQ7mMkSkK98B2sHWcU8Yz/EEnAajQ0wW9d
Hgynt9k3N5ggp6mRC67L7GP00IwNuCPFCO5BSJkhBZsIxCaacZpPa3icY1wOBRYxhjFp+EB4IyG7
i2jGOVxLMcXmUOJvv3gchSaoUhidLSNG20/jbvQfKz8YOJk8CRcxj2x+n5JE6wGLd+y8E/r7qiyv
S95hRxbOppl6op3cLA6puijSfb60wQmJwtbusq/UhJFLy2c7e+3UUYVZD8QD8rOc3Et1L2coauCI
Ksxc/EMeNHReL6JAR6qHxocwswuNDFTDITwMYnNtSkD4i5Crrcwqlyk6kWlbGE4PZn8aJBh7xa3I
eqwh/3Ye45u9dT5TL/9CDD7EQ45ZDYhCae0SyCGqYQWHey+KNmoUXM50Ansir9LeqIqN6ki7aldM
/l3C6VmPOtF+YGxkebOr4hfVuaQYaJDNJx5bTjuROrqJGfvjgIOih3JEaPZWyCsNbWzbN2Q7gUxG
WiQDFC7qckbapQJ5Bb3V6JSUh73a8gdb7wkwpCdym71R09qEmWADl4VojiDzLrt9a56ijuMyHGvN
NbWUlaxmaYLWtxHH136bviscyuWi3VWho6YcVmuOrnfhWM7Z4vi/e+PNG1LL3K/z+S3ILX3dmjHa
2jw+kwVyYS7/dIXoPSj/EjFZRktnHWSj3v+XFAPkO12PnK1hwZ1kgqI5fnJY/qpjkDQNi9Xcxs8w
InD14KrzzOpbjUqYO8aRAjqxfi+usfACdg4HjJGBdAXRVIm6kWIo77UW0FY4lsUqnumredGQFGn7
oDupLfOgNZT8lRbE+gj7C1bh54AOPZWD44ilYdzTqvoXINDFBDCjKdkUA2e52uU+csmcdLuMqSel
B1koy1F/5r0fPYAlqPq7FChoslhbwMOpBXNERJxtBgBabuv6HlIsQHWfrQUJ8KZg6rxzlDWZQxl3
2+arOG/J7QVc05W7SuGZ3KTIsxZWezPHfVFoPDxnnwFZbIFpGR9HJVCzUE9bPnFmfduEapX2M9uR
HQ/iq6sfHV/Ndx5I+BQ016DanWY0iRh7v1goroDduAPFRUDsAFrnLtl6ZHVZfaV80ldQbWQXRRv/
YieG/5SDgQ5R+pGLCk/ESycKtTngc8qrHRxpHmYdZn7XeKDzsKEiy/wKTFdicbvv5X4xxW9LRtv4
WYrWROeKU6HumEAi3h3uyi3QzUER7tfDdZSmWiKaLWgkBSsduExM/TnLto97Tlz1PRWGfF5Coq4y
6xhLaYzEl4MWBhFJ+1WWfA1y3IiGmjNxptGRV1IvBARYNyam4NoHHmTfk4xaJmdWYGHqNraS9z1l
QcQTakjeIbg830JkduXjvIjXy4AwEc9t5uclRGiAXs7h/YSnaeMb6ChmBzZyhCQT62F8MF6bxFbg
g+UMuu99U/1VpU2iSpHfxe8VH9FmNSqU5WOpp2h7X5x2hKtzP0SsXCuNza7Zaz+g8uRx3BhISObZ
BIHt+Dblj9GJOuoxElJksUksP7Acmsj4UgRKF3l5i4YMmzh6RTJqhNxNjbNSUSs8b6IVXLxgTG+h
S7FjK5gcKf0iZlKAOkquXrTErt7/+2eB2SY5TwsbA8xoXJ/pnqF7gNhrXNupE6Sx5I9AO4ugKEhK
Czez9yMVdgv2b83EXwntzKRBR3sWcumWe5hshPBv+38bBEdleTh10SgMHhLax3P8tOl94nRWG/Jb
GN/OVyhNlJMeO/Y6Wcb0bGSeH7q1EXbUpnRxAkXEIr70pYY3hGI35mz2fZS5LWe0B9m4erk4me/c
VDvPG9dNMenp7Cfo1m9L+HRztxiDHjV6DL9i8QTrJUxRNT/qVOaQpP8VdgqP1yqCUJJuJvIRA7wL
x4wvSq54pJ2owz5v5ICxMw+BDlIf7bIP5GHjDXjnLoMLoO9A/3PT2CwD0upiUOg3rLRuCzXY3dCH
BwW40h8FwYpKeUfEZemWSRt2JV+GswOunsJ48RnXPGkli8UMxKbywQ+6RUtYAOcfV/6A/86Rql6k
kFXc15NwoyvbgmBfwwvyrNoH4yd0zlvGTK0qNUCQ7ILhLSC9dasXNLwUGa44165xZzbRmVwWjQmM
OKpn6M99yiEfXM4KfvS0jtt8/tE+T1WdL7Bloctk4X3q1/KIbyFUtLHeSwYYFyKt+0X01Y8/51Ao
2SW2WyqMOwhK1zRtnOj0RvYe4wNFF7GJiyUkxkIhJs11ofKU1A7hkhNWuJbeT/mSYBOw/c2NSbVq
phgZW9LFgTLV5shGG6zdY900ZoJC6oa7qzU4t+9717g0YNqWa5p+v5dAVw8bxv/nNXLgwDnoCkdr
/73iI0zv5mFl2qFnQZcfUHmHcC0eZhACQNcmAncXLyka68pgYMwTBbORZFXIFlfi+2rdPWkzqLta
Lu0TuPD9JcSNp9XJ86/ERkV1zWchDpIiLIq8VRptn9jGRfwCTbuRss9pqAjGgrM6JDf/8LqnqYoC
I3k+CBKJ8+uyB/wfTL3sjb78b708dfqnOt66sD30dnGmg+mB9+7Oq9R3exbcAYLC8SOlByQleUE+
ZmDJ6lawu01QFoLfA3BWDW+m++OFbbeCj01mpugq/huceBFfVyvu5dtfFzcxObRsQqLG3Z3CKhyQ
2DOQlczGFaz6B095JDfeI39rirQetnJCeH09RoJjLTsIeJLobjZlM0D6Q77SCy0mu2X2w9KhYdBF
PBWouxtx4kxbb0hgxpEYgAqEl7ZbdyXLG4YpHUy41XYaw0rrNHp44+Ho8dqnPLVeJ6kEDE98qyWX
5JmbuOu0iHdDXMDtqFMpQn6LjElDeoKyVnqnjvD7P6PJgoYhvvkKpC3n4e+B/B6l556HvEwDQUwg
f5n6C+n2+hp2dx1A1pxMfElZsbO03InlydtNVzzhy+Kk2WN0bVOStu5JvDYmkwK12Lkj+xG/mwEY
0npdsFqiZtJOwqTAtYTTG+jKEVWCi3VSPjgHegCBnW751+ux3AOPJcsC5DLZK1c7PU9+MlFPwCiw
dtH6FgUxz5KczK6aUpUgRJHkM+128QAdyWbNk0ek9FYqRp8wHsZWEldf00md+GCY63F9sdKfIzfi
zvrCN3Tm/0YHbZyqGlwXiblNsSNyP/qDdcVKnrkIaPPKUOfe5bQDA3t09PRosjGXDjpByutqJChf
hJQR0dzWa4zeY3mCguSgz2Bb2OTART2KVywsZ9GubHe2fyoREZiy6/i1Gp/5JGvpRLFQRQKXZcJt
4gh6TX2m/qfoVM3qM38NzwXiwIHAUdCoJma4mS7HXVC+conaU6gME2tQLdL9KsmX+Ar/gj4LwCCp
qlnjF8CvzfW/jEFs1V0K8UEjiKLDF3ejX2ZMtnvx3wHEIc5GgkCn6yIDENc9bzxqUiPlbr+SK7EM
YPwmYSH0yhDwNha8jgwA72H7p7Boin18Za+RK68TUQMz/5mQz6P24XkWY5sKiP/T9v0ro6o7PK1L
nkqczi0roPwhZAhbL2464plS2It2IXDQDslAhT1BzoWajd4/RujUGWQE/kr18tkTwjM52WiY1nF4
EXEjeyxBroaZLAxooYNKFcJwD5wgccExw5NDIoYfZjE+vensmDWMTenlaomkgAF9ipAVH0ohPoJX
buWeLOarU+JETFE1RdZY8F4CS39Kh3ctqu1u1DJF52KDbzaYEKtGnIxE1xIc7Nnd01pSxejnnZkc
kcSpZJX+hYPIduPKqOPM5dAz4fekRsBnsqOreyqrmiv0Gh0iJqWxxSmYcE/N5t62ePsRoKsMaQpK
miQvdgqE5hTaDHVXYgrOQlCQEpD0UDPDxKk4e2vNhXLMtsS8AYKXu3jEyXnnznZgMMmXf81RLz0F
twNT3E0wLzwCCBUnwTSm7STI1NQSAthkKbeWhxtQE3r6neKbeC52teFGxbtEOL7OdK3OXS2c71VH
UA2KWiWOiFtRJFDZIGO1tq5zkn5wOYFm9luR/vr6WovZRun7G23Eo4NSCpXNHOdgEIkvd9edaFTL
zhJzLl3hTghq905AEesLTPKB4OazOedJ+ZoMhNuMTUfeGKVCUAZ/02Fyz39usZWyJgsj1ojeu7cU
LWEs87neL6OvkMPMWtx1s54wC3sbWdj/twne2V2hkaY92HiP35SUCd6j97hrjeCy132r9e9iZXS/
fqdG5FvfQQpZZRyE1etBndFew0iMgnzRnxOJ9sGaSiFWYPCagtKqCVVBmBQd1rW3CXaXzqlLfP67
DFCoLKFqV3oMikj2SjDMkcKxkQemrzBoMjPxw8YeRVhG0M2lqGurGRRn0FV2xaCinEpbTUa8gdaM
gVS5ohXr8IfNyUA3nKLerascFDh8wsL+MQR6cYebE0ty+OGGcGR0HBy3t+gB0e5krB+Io7jbKynZ
ocYr/Tj09Vj/rjkrdOTPyrYCax00nKu8CGY3PjKIYTUkY0HUaERRFKPbrgTJIqNYZaV8FNLtk6Ww
98GBgICyisbDRu68yUvRnyNEIcN0NeU8XegXH8Vk+o80DJi1SCeGXt9Q3EhiPFs5J6v1b2ZKrVKH
JctisAZdb1fWnpj8S5KomGs+vpXWC3PnJR/Wi1zK0dkqEOmxQadHo9i1kwnM2kHqbXBGWiiLPBB/
VAZ4oA4XRR732dgpriFXkdBBH7oEZnUvtYqor0lZYOWxcA3FzBpX0JSNX8GjjQEbUw9q5gJ+WlW4
vZoTKr1vIC572YGD/JdEvn1CFAcMbIXis6uDDsfHDrpIMDerH8OOw9RnNf74pvS/tGcEjIDb6Fgw
NMF4N79mW5qwVC8nFv+f4KnYux2VbBiY8DxIuohYV3iGTE0T2WG9RSLRhC7XzE09GXbEK7ViVtaB
/954mMbzC49P5pluYXBM0uPaVc/bTOhE47L8b82YqNjbSxy7qMkbOGOwhzuKsxM+e5trDqMLnR9+
aIA1Wvhg6CKBUFxiBh480zk8+qZyeLOCkESiJQy8o8XzdJ0qp7FdmVa3ReXl1zibq4Z6sGugjJoI
pbBds1E35qPRk0DHdx8kN12nxXYl4fi5zN5H2rhRmPCQWqS74/dO0BW+ZL8mde+OT0b6ppOTR3/U
yEqBuO3j1GQZkqU4HmLu38UDWa4MyPyDriEpJaYUCbCq0TibKP5romB4vApHbDkOfo+SQFS3ewRM
uLc/jLgQLrcKliZVWlqk3rLaelR5LkRseqDrNS2j8wvhtvPHWiFRSlo1wM3oKb2iPnYA3at8oorg
c28rnQ22NQVT+ZPOWH3a4siw3f0+ZwIcQmhckBgxb+GsF2Q606eerSZbaqltuTS0ecBwfskNqoQB
h9QH3LNIdIOnuEpxQxQB0Ii2xCccp1uRokfrQQ8goMXQ8W/gGpRm2/1WT6LfBa6rRiZ/WNjQ3olZ
RiQjnGqsR3jV2hqPIKsJkFEcscbsmgaztrLwmEMmsBnSgppnqPt6OxLBy2cyGfKYNMR/OnCb2jQw
n11qnjhe5KlpYsi/I9zISoCx6omn3uyKbIUhF29VPbe7QFkshhrl28ilwgYQjFu0jjNlnU4/lXUO
kfE2cgWwRQ3sAm0qHbvG4CWjRYSp5Lc4VV9ZuSIkJgbmMK6EWBfuoPE/V9GGHkNlHQu8ZcUYooFZ
XUpWOANlhwsM3p13ax4wOnWW/29RNEtrddyxyeSX2vqdGD4jcAupkXagswEq1e7i445juGgeMb7U
c/cCHZkWAheKOX6BCyq4JpOFiPcYt67PFw4XsYcWpwuq/zCOZ02isUPSUDL4JCFvnu2DMJh0npIB
n6hHg/VQ1IqPissXjcdQnPGPJb+fZGtLfKjft6TEtpnZYyg/9xTvjT+ObkSrDpgCFi8+NZu+uwz/
HLWRqBrj1+b8BWOJ+LPdjPcC1tsi+CTUALFSzcoyfeKCfE1sX8x2C0Wp8QLuiy4l9fcQ9SmwoJ4i
7GyvBDu3b5UOniRmrfzfTTblMZk+o+SaJeQHH3nAWJvaxS/U4i2l9h5LktnLiD6HAd1bknWzF1V+
CWaHIYQDXBeHPz8oXR+mxZY871UfJ747JOZxr/IG4oOD20HXQizjoFhf7LJNCDXYDGW1KbTMSAQg
eSPuCRGzVwPRfO7fM1ix/5zLtxhAYmtQs9Uv15C4hnfvkHnavYzQs3RckVpnZxJKQV9Q/2ZuGeUl
CRq8k8z0HHV8YYxdYJDs5lTH3QM+qJoojC/HD/kQScXJgIYhHBr7A0f9qKmGzQALJrLHwx6XG+VY
gIw4yOduD8tT/NkIJG1jODeqXCBZZwhSNlskUdKfYf/9ErcaXgcJOWRQlA8pFrNJvBSOXEn6AKPy
srtkCKARuhJSyih2b7JSYIjC8ZqZv2SYg86eqgM6A19pl9PzLcyOycduQ/4sLZv1qZp2tGn4iUHY
r4Guf+sf3hbt+jKLilOFOQlSaVLom/yGG5ys4WfqnyGFz+RdxGhKe8etXvDn4GhyQ5EUhNcb0YaY
xRq1ieHJyDgG1aUD1stzQ66RL0Vz4pfc0vEz0lVGcpJlOHq9MxMUmUGM+2M7rQfmBt24eVSIoY9G
wtg15YaoOeSuTsPnCoxQ56dKH12sTy9gdKCon4kJRL0hKjntTNHSHNSS9tspz9R8NzzgbS0mN1Zr
HnmA+5nakFTMVU+rgNaCK62261ON5RwtIA5LQt/RXX+W77DtEvWTVlRIjmMHzTmgfJz0xn4FpCwX
giupbaXLK6cizIHWx5ctjZ5NsEvnZ6u+/3B2PmSl/KNhT00XHfVp+y7DaldpyhqB0yiQC1vhRZyI
voTTvQFpcfyaI3R5U+9UYEpDjDR10oTuZrWc6yjGrhPt5C0RlYVTE45fOsYD5rNUON345Ytz1zRR
ijDU1VqfnzxkoFKWfcMetqbjNegvdJTKtW1zq3QgyD8XyS4PfadsRGN6a5h6kG5fvqEM5PvJ55Dh
qKvrMOhMgt8BzWgutA7BJmuiS6xmae8IbqVAdbW7ZpOa5BU4eH0ieoynPLRKuegXmYWROB3Tx55v
aaX9BLoDuyby5i1jdUPAr4O3C5+HfroYdQZSpaBS6R9bI3sbXzwOx4BO2dBLM51ljVfKHXzAr80v
eat6t5UM6oR1zpNLte/2rBZYrc+mCDVwR/nqIS7+/ryOJBr2ABj+F40xZdoGlC1kJfvqLTOoH1Ur
I1mM9vEIPqP9qGx39SKMfIQoNJBmPpwE1vItUMWe91KwWtNBO/G+A1Gd03e/RlYtABGNUZ5fGppf
YHoXmY12xKCwEFMxSc5fSJ7dFcAi6iNoty/p32Aoxm+wjZUyGW/zp8YsxxxkplslcqxhcUEwkRLW
lZM+dEgAr5gt65rv0AwbJY+NoKY+BtJq76jOW8SX4YqRaeH/H+9WHRQC7zYZQWxL+KvO0qOz+eeT
d6eyGH4YsQUUcMZDreenDBTzdJEE8834AKEFzJH30BOhF1/7OMad/0JhFadjGe52toCH68/oBbK4
HG3tTV1yYAsFnf0LnNkYzmFSfuE4t5F1sD8ISIgdmImMY9WZS6NJizLzJ8uJbp5jITQAegwNo3x8
amVcGUvehtSYf1ZhlZ6HCj4MY3w3ce+jBNIm7sHylQcMl7QXnzfTZw2zYIY8Ids5FJUueZnQEGuk
+99o0r36VRYXrwmNp6cR3wGvccEo2FHOTU+T+uNCdK1sMA9vekPAAhsh/rgJ3qkWp4XoyktUaCIu
JVTd+1/qtbSo45xgy0iMYMGtUmdG0G+IYp3P5lY5HJ5Hxtkr9UMjGW/7AYxDuy4TzWiCYtC+uZPy
spj7YtLZ3NfeQwHFrT7GfjQOroYPT6SmAaz0N10CDfZnHW+irFC49CqzA9Md9odGPHqyymc5fYdZ
i6SI+u1dSQ3Jdu1wMgnHFBJLoZEUahMYeRj4xG7iINZB09g5ReY/Y4BrGaRaHZcS7Wa/Riz50xeW
weAKhGZ00qwzxn5PKA/vWtJEihZIgtu2fXModVXHEd7SiyfgC7AsZQxpA34ldNjD49hNebYN2bUO
x9sE8+cdKsfFZBKv8KGTmQvVmlhAHzlQLf4ixxzVG2bhmUt53GjDGVAWoPbsFZXahQXEP9jc1BX2
ye9WPshkN1oSf/G3N7l/w0GaBDRkBRWPKXr3AOa35SDrEtMHozpZsn9GBBAUamTTExhIi88fjW6w
pWejdyC4vifUgvN1V+/bKLEx1O79Fpojl5+bIO0wPrGHF8SXRozq1/01cq3Ih2EOhdmar1k7FoEQ
D3e+zYd/ZnnDhSU50zXmghmXkluFHjpR2l99j4ZDeC4Q7RaKhOng3+1YPy3+Z1lFtljsM+NJv8wU
CxM5soew+9BC2loSmwi9FhFNfSIGFaeuITS+aQtUwmDq8M94vsZa7DSUJkuM5BsqnFHmwCDb40K4
lFft9VJruABlHerieBkMTxaB4FB+BNWo4oj73qp3wfvb9YO6EqyOfRmY/Ic5apcN/xSZzEv4/8Ho
2p1+7c6v5p52kZu+lXpfFSydkru6jdZvgbPeGdcTz8Qxq9vwUrft02QEazYfRskcx3gvuFNb5TXr
9jKwmfeC0deH6P9Av/+dnLaswR8/rYSK5AEiNEgJkh7rPtIwJp0Qopjc3+/4Ff8nCkiIMQ8QA3mh
CIwRNQTxpDlnhbKVX7TeZR5+aJrfaRicoiAr5FPbv7cLEucJVl8AJ1mKIAmYBBIsJeDpoltkWSzL
ufsT7AOeu1GfFlZ3Oc2ogulTWv2cieefXYXGTt3xQuVrJ+fyaH6jUSGZNz1xSGArLz8cDRKUanU2
IZugPXtmEoXWXUkEIXfI6Fdkl69y0tz/4CI2ZSLgnoSpiJROouxtxcyRKLXRoevEHlIDuZzttxTi
cW+1HHmMrrl7qzAeDUcmw/mJuELjnE+nuQqPzY49L7ohPoSLlAVz3iSEGLF4FrPPzd9AOu5hBVnI
oGpfqe2Njxwo+NOd0XygZ46/VY1C2s25/lfatYck0bLw6SrT7FVHkGCc4sVrBCphu2L+TSIaWNCp
ts+v15yqa3jNf8F0dlqewqwypRirWjznxMazy5L9cyGmhfPC1HTrQkaisCbJOIvbfDLcSjfgnqzV
qol2toip1mS7M08+t/qv+Z6fzQEVaScY+fYDJ8aprej/QJzrTE8MGOPezromc+QCsEmT7sNJ4m4k
rD2S6VTraojNm7NrxIcAto7UEt+w82PDAhY2Q4HzH+gw5UGLj3t0wCbRK3cX7LaWqcIpNIjcnVub
aRLmNx/1yLqSI2bPVt2igX8GZyZJuVvC5O9ZORdnnc7CHMjo4BxhllKQCjZ5miGjinQOpTYV+RAG
ERn2AtDKHcBn2vRz/1AnO3RaE+QF6XmM/ozNqtncxTA5ppb3dV60FPXcliTumYN/ueYFWeT22C5q
3qcYuIvKDVxprtYkS6BoI+kAytIymYRiCvlHXq9Df3me4DMr+pejacFlDOx+8zN0IhQbjakgrkD6
WO/DnqoJ/bPN6bWeMqFUdgVAZYBhHJ0FjXVk9NdSzOPmtGyHEonfdrmFYYn+cG1Ly+nPRb5it7R/
BFoXgXKvNzPpKSMpbAqQDIyqCfi7QPFazm9MYM1fmceCODhgcjFn9nmDg+Tic40I6TPPML1/8wAu
Lr7oRpGS1BJsnGtKtoLxs6Oq6Qsnml5RT5CzBgHu5PZmnqGPNmM87XK7PUNTqYmNmMdWhPlDAsjv
tNK33Tx2sKGQWxnt0sHgJY/AoEDXNuoQYnwwgqbZ+rlX6PNJeWMjcaLd2hopysEYe1HzVIClNPjL
HR0xL9dv1dtlrMC99scFQxbr31yh34uMp7D7b7lbhbhwV2vjA9u/6ElYehGpF8enW4UMJJGJ5zla
4JKTZJYfzP7J1Klzj6/xbeMHAJH01qCBtonZDGk9pavKG4cqRM+Qg0M8NwuFhX/q14PxuM31Kq2y
MhypaK0cfRt3a/4T30bPqP9A4y1dyiDb08RJ5rQ/gL+Kvwok5zXiJxGSazX7yLf5SZrUZ09dK9WL
n5VSiPFTFizfSDZMYioZfk2enelaOMbW/hD1VWI539MNRUMFmirG43/dCYVfaxx7V3sbVZoO481L
C7/IKuoBR9DZA/jxMFKB0SSWyEC7kPtOkRwlUdIn/xnN2Uj7U2F7e8pquKhW/ZetVzMpb2Ev4OBh
84zS0BrCc0EqMYTBC3umc3VzDgLp9Z38CbysLzfArgjHezvD7F3CMctWzRodY2VYeo5AaE5Qyu8T
nRpzDY3qZ5i69E1XQLVdsiAJvTj6vDHlzF5ex4h0pUYP5zfoC4gLqfUzOi5gWqbU69N+IG2Rhtvp
1LvPYENwHza5rTOIB43I7FE41PGvkgdEooKHc+eZe+hlzjbBCZQzaPIEWwvwRDYKEKjxzPbQ6aQD
nal2M+M8sBdIYSzcG4RuImZBLwaXpy54u61qt8Q/GVWS25qsm9APuS4NbEIgJH4kiA+iLqkpxse8
HZX3a9+NKbUbASant6bkdSBjPDGIR18ZYzQxcIIQa+9RkVXdcSu27XbvGtI86HM2ZU2tifx3Z8Bt
IwN6zDMSA4+u0PEBtXcGt4Lkn4ztnAT32+0tqDe3j0kqeCy7xv4PDhKlK+37BZBtLVbgdgltQmQ6
BsSti4wLcnR3aQa1LbfDeNK8bmpTIJY3MgGqZc6MTbwGoOQ1bjp8qM9I4uAuz6pBKR0DK3qgUntx
kahnGvm5xrDbgX1l2hjlCWhiBK3kZ05Ju5y3ZgYM6jr0XPh98xXXzOPDOoeISX53gWOcwdo94o/k
k1+Ri1tJ7aQ7b9iwinz2ZtPuVkb+R1ogF5pG3FwGPC3o3K/kks3hh5Bna52cVmSRP688HK4u8jIQ
WGOR7KLTYx0Kpd7+j1wBqIeuSeHNdn52XpG9d/yKNMEMy7FH81WIlj5bZqDg7i2QSyG+k28SiMjm
JGwtLo5bHlfPpt3w2jYNqCJJTvnVvCUjDREdVvKtWkgW3pU+jUBRuWo4xwLb2BnKlDdg0UxATgrB
GMTFKYl67bP7XrLnEFmbGg+J8MOJ/Yoy3ZBy7Y/ebHOsIbEM8jwdW53dewwmTUf7FaXanr7/Kl3x
o26rDhBBqny0Hv8qL01icSAS/H4MzNjaStI3ZDJh66x5XB612686CuT7PBzoY6a8FFDS44lWgw8K
caH4NfWRQ4KUdM+KTkE6x6+G0pCbmIwwH1nf5L0gAgir6Imi2NGjBs/W4Kz54Nsj+176fnkcx8/c
DUMH3yXm8MUs60gvFCPi1VMFaio3X33zhgSLt5fYHLGMwlrXGaC3A19OdqWZb8FKihXG4d4lUdEv
9Cv/AF0mT8W0MgdjOsitXMSUg86GiXSurkid+3KzRw31IJUJayJpR94Azn6U9fpheRMLND7AzrEe
bYGhQKbXQob11a6XhdhFPtoWT8zy6F7gzJDEuWmfUgccapD2/W/PrFjsGCr4l75c52b8GgzBWXgU
EbHCo9R1bBJrk3T856Px7bOguQGPC+6R+JF1MIC8iP+119lwH2njCAjQ7ruh32kloA8gtxWtLAjb
AO9ThEOiqxh11HwXEalCNXXtwBFO/CBf1L5s8JIatvHuVvpmPmy7zniQA3Tjd3FcPY7DHgMYZi4k
FNOaCIrWTb6xNGqO0VB6KeeD4uCkalQQxOHLyWmZQLPtBQeNSP+BFVmwn6QMUOHqwnyRKuL5dpp6
jV4yhbU/LFHUc/LbhwUaOJ4qt2n7NgZauRiQjGV8PtL+lai77biZFiXe9LckytG3FjqLBhIKBMqO
CFmIHh3ixklN+EUMUF0Rnab4V8eWuGOvOReKS+GSQqoa4QGSv8Vic8EqR5wo6rNYLjwqqAI63+m5
9MXH+7P7qYDsItxo7XWcOeL0z7d57yj8e+S0EXzyLcgOHwB/awxLJ8abBTxZ79+aNwe4lCuL/Kt4
t2uxY0kG/ymE97w4LME7BiJ9k8r6Z3gKZ8ZTb9Y0u015ItCAwFm7ZNVQ0htU0xbM3Zk0w3iqdGXj
DcTcPwEhRDMEyuRWWF72EqVj4cU/yFdTeZHpXS4rPo00DSe6Z8Aw3qFgLXiab86EkVFCBPL2W9NA
m6sRSQT37u1mz3IOU8btF4cfL61gU9oAAm9Y7/Xa+/Y4+oPlu278mdhaKiUBJzVJDrfxwpOEOgBo
P8oOOn98SX3z+6pP9kfkAUlRqMQMSbNdx8CXrt/ouMxrnNhwfM3ALlVhpyiMn2qt+4SVvEmZwrDr
J6Y7vzOEWHFXMKu1GYzjzhIqqmrbWqeHHhGiFx4XpJdU888BuRoa+a/cgh6B20N9MQMhZJ8c7wVG
HJpjnwOEhyXMFv6oNREenUJ5wqur/wMLPRxAFz1L3Wp+29yT9Bco2oOliIC6V1FNlhyr5zT+G6Bq
itdUYar3lZdVTePgY76PugsB2hqlj1A8RVkdgtZZ9736YX0DDjw3Uk1eyUXo8EmgUsNtKtZIoA5Q
c9wv8I9KvG7+N7MJPVheGtp+1S1QU3CZdV0LjWpEoK0pL1IXzzCYlD800iaBYYBYjlMT+FK+oDyz
YhReKYWm+2whaBjEsZ+lqyow1sXfqz7TceDdLJGI9f9RlXJwul43RBca73NuPBp857jtGhL8gmGw
JbevpRzFXsh+HO32CWKUdBRegGRhEQg0VgDag0iIjWyQKaxw2joKWvTnHnLvhalqbSjT0ZCU45d8
Bf5nVZ3jISwoR/4R3cJNARAVROAO4CZFGZ0zQAbB+hvXjRAlLGkS/wRaE49BMl232o3N/WzlhGi9
zY9c1W0GecXfCwt1B37o+MiNPfO+cmgYId50dlhQJPMQe8gjQ5AxaB1lhtBUA3jm3ZK2t/1Xf5Fg
7oe2dQkM6GLgeBI5shxwD1WqftLp4UBTyUptqnX2pgsj12wUQYzQrSPO405/xGtOcVJ+YMh1Y9Zg
AvnOHIHNbL2Nd+FAnejMsBe0Q80mb33/ELGQ/+2q/ztGWPS4ARojBldOFoG5ATD7QGy31Eu6XE2v
QQAEwkEEGdkEBo6TzZNREtCpWUJURhTneHsNk1mde4K8gls82XhkRgfBXz8iPSqhc/ipQGU4/NwC
D31vteIxmqCqAbfkNIFWKXqmp/YDiYOZwp7fYVbHnm4Jn8OfsLWCbZc5TOO99BUlIrLMZzKTSxR5
iTC0kv8VOlpYobrt5VqGETJhjs4KQaXzGr6oCCZN1eBtpG42MNqH1Tfw2z1K1YALdk3lH0OPGHsM
BVY2a49JFZ3pevNAhqQxRMUtDPdVhI/KzRRVG/RVEqA7dYUuMsvQjrD8m7UGE2iGuw80Km987NbR
WCZ5MgvhPNJIlpqYtWpK541adWZDGlJxBsD7Jwdh5xtEpGZRZFdhEEv4L/fBImaMzCnq0aizHxfb
BbNOamZml3L0b/f7PKFNcF8GtYkILqrDIBs2IID9KmXJ/UiAQnVmqlWVYSNUj4Jn2uRGHGUR3Og9
OddhDVsCl1dpaDHakjXgFQtORZdPYsKKXW7R840MRwEqu6LtWGgp7/Fg8+zyvKP+53Um5gy+BlWL
gaYYyj8OLpMxX/vrBllIeF+dq8o4pL1vNBDcWmOUGC9UALm9lqbB/wfzGPaDN3i4UTcUeZnMIibJ
zIeLSNY3gT8AxKkOywqw7na8Mv2HgRuouHM8A6aYtRv4pJeLHDPffLh+QYercvG1DgiIioE5NLdk
yfZxAssFeTjp8EK13wHp06e4bm5zywCQ+esdjSkohNrN1RfFmw6A7UqC16wFnmTnUY+3Rki3mkw5
EqGzxLOlPUFQalrFhmVcw8TTbHDE/+XZScftlUH4eq7VsP2WnjFhSWVdjtBu3SF9fKtKWEH6sDoa
mcJCn/uZJOLzMMnoeM6zttZHqTH5e432o6srvqkoDyaGDrRj1DBNOJF7Rm0Kqs2IDGDd3Y6ewfkk
XdJC81HSCGXKuZYT2U8LbernreRqB9BgaA2/e/moIwngLY9MYbZkGBedsCVBmqDRwuhR8IPo7COn
QCz4NoWIKbG2jxt7mkYZfhNO3bUC5biRRpSyRhIoRQPrsbueP+9XtnBmfEjzTH3pcD/6lDQA0fJb
hbKRFY7APyX6rbi5TwlJrcf1lmXp2qTqGaMT1PxK815atAgd23mR5b8OXcVBTwMqNbkz0KGboucl
7ihQc7E7NK72HwAmowkDZHrbGMoDtQmjZbWPKmEwj2JJz8HTPjllZJvDTAtVEbnfFW20WFLnjxEP
GZQhh8JAi/WyC9yAjbSGFKrzVZGNc9w91tKyKfhKonsDDdm8mGqbYc9BPumc7f99BL8SqbfCABqJ
y57asNaH9HSOSC7gYmlhPw46QYgMhYFrYT7ByfgM/X57iS7Rz908CSW/mR06xIV9Oh4HXubA992R
sXGfJT/RHT/Zf5Py0SZWoi27HsoLNoK/KRqD2DWERwMrYi9U3SU0fQbLrs1fZqxuIABVHktr0MN5
k9WMkuysYmBXOonMtuQgocIf9BIN1Tc8leJGx+2uwqqjAUPAAdmS1LXaA5mclBdorf8iWZfYPBGX
+mf0LNTC0bmXjWGKZ+g0TJGqlygZzhIppv16Itc9VwqSr39+yjX5FNCOFoYi1oeWAlrAOQU8oCW6
Lj6sd0RHClgyDSqhVCstn7R7xlv2SAyikTIzG/qf0Qs8CeZn4O+1SMRtgBxmYYMwTim+zLzbDhrw
mHb7zimvPAR6B7acORR8ffRePmbAqXxqj+0JC3qeGZMP0d3p18lKF/izTSATTa1xw/GD6jmtqKZX
SQUk0Iic5qrZGjOGo5Degg5yUD4zIg2mu29ZPX3TbZkd9Z8VLgVdG1epzwMu8SLSBXvEmezEtPyp
HMXBHy9BlxVnEmO/4W5XfMZGAd6AgjLpAagRigfKGAamdjj441uKg9BCqjRrPfI3nALAsOjF/0Za
mruWe1In6LU4RrHFbx1OoUE3DHFJmDzAQBZAGpV2Oa2nY4MZ1Cr1ih84Sf/BRWSMT87MGrQtuMVs
iFfF0Uo+LENzjvJUBMNjPNV+XXZffcKFRxaHpJwSiUgO2vjdNM52xqDfYLoIOuQL/0z4QBkIT5Z6
4HjnzdY7xV/BjoH9vtEwOie3khTTG5wk5Rk2CRd1wEcA5TCp9GwX53hygJXg3Vq29DCyBRkUPIP/
QxrOhhCA1AxoCymtRMJHyYC3Z9yNw6OfvxXUzqLuUZ/Xcym9gFk+1k1B7xMBiOEi/9gYrtg1sFlD
blKoSOeD32ThmoKlawYyiADViFnQfHY7foUZNIeOooTcj3tQRgucEact4tOYM3GMMFXo2SrOO8Wd
j5gDWlx28UXw0XxzNxtQz4/W/sKNgJEY+F4FKcO5lRhodoQH5tuanA0yQ7FsHQYNTzUO4C0aCFNq
W3gISmq16XL9i6ItUXTKORCVDC5PwcI0gGJewPCSWD7/7R+g49HMofDLL8bB0/esM2EejTotYfvJ
C4uLVwAWgVApf3e90ch8DosUvu0CDDmPNeq2Tjj0phj8JmB/dqfk1XXwPrElIjPlA63KT2R9eYlQ
MlXLTgbTfc2D1ZsdDHX/zuh3wMtUKwmyuADJ6BIA9mAqFXt+axJM7aX3koj0ICxxIXQSDESRSzRh
W/J07UY/35PsXRJ5HV7K97D4qnUeMShMQJw+aaz4RhLWXFCrAtS0/SOZkIKK//OOxMqB0pzfi/Rw
Kfh1ZW4QWMwoerhXBXpr6TcwTREsB5wjSH6rYLYEBas9Gdmy0BmfBTI5Dc7HbQ0BeYVlYCYJ3qPq
Qi2Q9b9wHsGjm+fEabMa2iayKpd3A79/MzKAcJ2+d8P9iIpboLYnqNffCN5YyEUvP6rHzwpfPSSR
dSjw2p18vRj1saAMt9DhmiqqvUPiz8zuqTTeAFWbsnOpmlRhyadcgiFhMQYJ/651zj+aEQcQ999v
5IYlnS9RB4tGtJzl/3T5v3O6rLD55AEBku/1jYLJtrbqSe19RDTL1QQ4PI6NJ+l7MGz+xz9Y72qv
UArgMX92IQ4RgTFkFeh01CS5eRUbjqs8Ck/ywd2mLWslwcaPD1BmkAnUOtvVIYbZFFeiryS1PuZL
mkIWxVtOz5eTsOqMV/bh1Qa1wDwz7akxo+BDK2HwaSrjPj3JBGy0Du+dGGukBfiV3z7sj3+sfJMc
/4omcRKGUVIAS6MeUTTTQ8WBuiI20gxmnZVrUyb66f11diI1Kmua7aMQauCvq1u40kXHPvCVocGT
sFqNT7tUqb6RSH38uAumFNAbEGhEVXKSwfjwaBfXnazEpOzOPj+QOeqsZmajCtfZSCxYYruwXNIy
T/X2IjJRwBZhAZ/IOL9jt9iwSvGlxoDLMkXfxHl2Z2nP7MSgiGRhYH+4kFo5fBadrwNmzeveKwWH
uqd/+XnDCCg8JYtB6mY97OjGBAZUiJ/ZM+w32w63qdWqzJHVWG6KmXHnW7P2CpBb3tor0EtK6I+d
q2iHJZ7MFQdPIy7+zMDrQhhrxeb/sl1MRLqkrNdVNmNbTkYwhpuH8AV/ScfKTbIUT8gjqfipFfLh
e0kB2J8cRPKNCm4sFzOkL4dmf8jOPbA4fxFIwaLOcBIXFAVuyyjsGkwb9HLtO1b/McQG87HdLNi8
g8KN0Ay1CTwWj4oF5TDwC2n+e5KEBOA+VaF/R/3m7msMfQnNOJzc0+vubG4Ah/VVq7KSY+bQ2B10
t03KmpkmwDJedIkSHftY+3Y5H4jAin21bZ/OSL/1dlLH23GuqcpUlp1mNx9avckpGMVyKPXa10A+
R+wKcKIld1UMgYLt/JJlFJz5YhhUUAlpat7bGF7O0One4e4Y7yJJ4133hbPgXzmQ/27PGRaIVwa+
zfHZVfmRcCJOwMCTZrzjescpZrZiLMinyrC01UEcy+YL0UulPxjPWEpb6In5g/fM3QnHt5djFMS8
ih3TvbOmWkY6xLbr70fOzabaNoASXVPxBvuLu0ZdcSAw8ONVTkRmlcqbrqcYJ4+UI64br/2rViRj
UPowHWzgEnWB9AmdoQjzL/ZlVgwkaGMiuAuCTt3XMfNInqd18nn6TDhSFCKCCeqN/AQR5MQXQanO
/vGNE2tq0Zfi
`protect end_protected
