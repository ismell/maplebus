`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mG9+IxTgHDfgTriVTq5VvyapY4jw2nANbER8aQiMAAHPjhZehVoU/LiaYKHhNJBSdW2E1PggKKWU
lWpWRnwQgw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ayi+iJlwwFvprL3+U87AhBxWUgsxuMOzyI2CQLd5jAk9Aomogem8qJw7tDFgIBy1lcFto4tPehdK
pu5j8q6peq1n7vmspin6wr9DMQn6D84DCu9WRRHnNn4TndvUg/GIWEkKV5q2Zqt2rU2bJHbiVeL5
1A1gkI6+LkiPcaxvFkY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lYFjTYFtaKMAyny6h5Yo9NnsT9jGoeCKLiOzx+jrceZDT2RLWhWpMdBl+b0y/r1g9Lx5FkSPy/m8
EoR7nLuiYbccMOVwn4mWrqn2oipMKkcdaQE8WjJ5GvsOJx61XJD7zXga3B9cf4vlQu4JNFzjW++h
Rbw4I85rckXIL0nuNGqXFXV7NXLiChfg/wZ3/8lvQHaKIc1AZsd3tbRlwIy5ayc5Dk4t3BsXq03y
0hg+GehsVkRDslDrtJtDlKvq5EfNhnVsbTUwuxQIupwYlN1y9yya4ZbpB60F2LnilAK1ECXziA2B
sYeW9MzTVcSxJjjyInkF9oRJD+iYlntcELAS0g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ev65y39rOyMBMEtv29o9PUGnQ0CAHNw3Eaxu9WoQQN/+bXJrQNrgbYXihevpLvhldJHjQIrw2yp5
l9E7PAiUAwx9H36V+JxRHVwsJDoMumT66nqDttiQbMz64CkCg8g5rttDm5V3dIMDZ3SCH/Y6lmOo
l64FGbnzPpyT8FCzCgs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7/saSCzH0RXahQ4EGTxwWuki45+SfsQqCGA7IOYqZOv4vsA8SUZ/0IdCjmkhRcJn5dR2eOnjfoA
ZkjoBXhTQ5xkKrQZDG8OnUIvJ1qvcWFo72t9mKp9ovXShmL4uTdmwM+x+Pqlt5wVxOeqUtbWjMj3
6CLC1NuCL4amODhEtg3Cy7hHFg6+9THqA6vR+jhBUjzhH6VqpsSX2tPRa/v0OPbtLQGaloTOAtSk
kweCeDXMB4RvoPyUKg4Q1C3siE/NtDcYDZ4oljtLfw2LDFG3X+CBzFk1j2AefpMPuDTJQTwrwnM4
JGPdS9C6X2iA0Fp/83bCHjDz7m+rfTKCIcVr1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
GYLcFJ4SfNMPvFeZJB3Kw49MPkugrxmYdlJZv0xlQSzQ/Da2wXlZB8uLsWAHLsXX3jIq41Sf/sMF
AQF0bP2nYXXG4DVqNoa7y4YeYXU3IOC339HbQWFf0ONp75Vbr9mDh3vBf8hQpH3pjBxPAi6NPC9q
4NPtf45e/WFHUpsGpu3jtCtV9Br7/zYpamI/bpNaadsVhtsDS1q7qvnH5DZYBh2sahbijIy5+OBL
l/bQpPrXb+/bSnuC69xP9o4oOYliUMAbYWXDII/z5yqglG+nVatUGJsK5gFkb/n9y9g31moI2SFI
rJ0ELnxm0JWKHiqPDYl4RNNAsMR1uZSZoIpCNbB0TQ+adVXpvWZtYKr+wh5YwuB98Pecvc3hzV9P
61CH+z3LdYD2kwWwBkru+L/aSpjy96+gh87eZDyTrVEQSmPxy47S+onyI8068pN5lKy8uCKVa731
QLNNNQXrNJQqoX/gJB4HTTIik440we4pE/79JYgg2nKoWQjAdPbr1WR74hAStov9lWe02JhRm8mP
aQ+sgHGey1ngCmQBjdhAAOFTt3BFLXhx3pZB4M9NXhkTK/vQAhCnrTbb7ep8+NQjq/Bb4Zlw6/Os
mZ2PojDIv5PwTsVGukFAJPP7trPUP0fy596rPAGWmwip5N1kH53ZAqEOmqBKkOMA69V1mNtxFhwQ
vusEzOWV/FFGTSkJkaC7LRSsPe7tRYFbZuY6V+XObkdQRlHTVq4YgM+CnXXW+R9SgkzD+mplnWtt
2rC6G8p4G8MBvXco9GvB30i2WqL7GQJBWtCIMpnE6C5hbA3qs8qiwZv+IQccgKLZ76bPv3xX6zp+
/FzBBM32DPbtT81jqvmWObvYQnWN6Y4i4XegSvBcf3qpINKzTqQJQvajeVflve5wAFsgwyAwH6Qq
qdF5kGqhxYfTWYXjLR167MV6iVHgbUp91N5txNynCrgn4rcJvvHfpKC91b0m7g4F5QXw+5qGC5BR
pGfm985X+HkWRPhSUjVFRUPyhX9b9K6JNmPGE5uFZYdeJnWsTHC7skuTHr1kfgKsJn2ovbMpiQNF
2Wwif1CS6daiKP2dl75ymIM1XPiiGdBeJqmuHAERiaNqidvBtFyoX7DS3Zryi0bjtlX7/4qfhDmO
0UDZMKhiApJwC4xeZqKFed6ApvZXuw0Yc4p6PCCHBXwzoXvwuS+4EL+V5jDCDGrVqVxtR1znJkPM
E1tXpPjIu4MfGLdGTjnIaYELWNS3OZh3jVpNHub22sHzb0K6BnW+VzdROK3QmO5Au/Nk4lCbbMAj
3p77KrAXxN9MpfdUtv3hiFabi9ByAWvkepoTCsMDjHgupveB3/mwWHdF4PggPvAeC2i1kA0Ke1Oi
5bxz/25s2Guuwy+FqrKeWwPNw1dNWI0Dh8wq6AgvpXppr3ergBgniipxhmxX5gLXjpy7HiPVdjya
YzXx5iIlrMIYlpCQZsuyqBlDaXRLfjWVxHphBdQSLES/s7BbUeVBtfi0ws0BxpmrBsXKd9LPpL5v
mqjfGdNtwMXzRzVHqOyqhrh+pZVz074xQlMT2R9ueZCtgjKM3qtRmIw/bXKxsZtvpzJFjFiIHdhG
PG80+yKORzOojY8P6l+a8GvZ6QIwSK6JJZWRHf4DYx1ur/3B8MLvI1a+L4b5Ii0Gnp0JX3toX9MR
IY/93zfKOWrTPmlLlGlpYqZX3U5UJQ37P61Sbsw1m6jziiXnyE7sHQ9d0ufQ914Lz2O5MgTccPsE
14kBWisJIjdLUqAYBcrcDmbq+uynozAdHJYpsj5goWbw0YJSC+EbsGXoHTgl6t6qrXP0mpjmKc5C
8B1Bnh14LP3Qzk10JiFbaWSApt2kBvfh5W7aNHlKRaeWUg8V4dTlcwRDXL+rugHUQFe3PowsqWzA
MGMLvX00BsctSPnLZjIdsUPnuOqQnfcnXIMwtMMsvEO9OMOUO57OVLTUx3TciGxKsB0OpHLcVc2E
ArjvA0NHg/gAkSm0AB7feTmVs8G6xUx5sXJxaeCq0inrm4Z/wa4YyS/JC2lQSdQiVno5zfhlbntx
hM8tdpRyyUXZ3acmcqmSlNAb1jtwcThC2zVxmLywBc6lKDlg3Hb13iicFiCdKHrOF62MgyheAJfK
wdYhYpNmsSB2Z7iTy+pVCdxM5QDhOU2xEwfISJ7NHVY7FUW3ui5aN9Fq2XKcfk1k2Ck5vd6zyZhv
k+avZCiJVbOzpqI2S5vhI6ZdTlcVo3fIfLBA3kbGuWUrdjpzbZowymMvBSW8BMO36udE7SeYuq61
BV3v+JHlRdswU6vP72RmuGVf6bVLAhu8RBNFqezgoaIn7/zyRw62CWgp0EVjtV0H+pYq+nfH80xH
OAIholFYFrl0KT+loCczcLhKUnrNnxGRaxMWUlk3qIXpfPRGyDLv0WdHjFLcAUX7pVPrA+sx8RnW
eLJiGvaWMRPXF0Zqe1yvqw599Lk2fbUQ+gXV2qyoD4Xb45SMF9uUB8k4aWNZmGFXjmKVwIBLfsvP
QT6jXH+7eE6L9OUD3cwot3TFjmnFgZkaTCAliyWY+O2I/eZxpCFUembrqH7eV/MRYzAXIwC7COr5
Ud9Az1lE9HN4EEsSSWhOd+Uo6q+nu6z/Gaa7qHnNLw1N3wihy3lbGGg8AwmBqZyvEa5awK34vjWD
qUTNAFFYVVR77KMWnwDCobcmFQVg0Yzs6o+gfi6JEdh1cnmUzdtVrBjER6+voKWcL+OASkvKU2Rn
fnSVaphkCQApNyXb89kTqARuaRAA93EI0Ro1N5EwT+4+WMkgQBGjkLJ2MlCG7PNy7QUsJlOAAbPS
kHc48FKRyLr4JtUmPv0xN03UskZ1F/Mr9SHaHgUbN1XjHrPMZ+Cll2oLE/A78dtlqHlPSn1wvpd3
2aRJdxIy4vgGmK9YbWEsiujADoQSZC36VfdfwwSFgis/AmUjW8p6y3QnFeBjpOSMlrVXZzBoG0ms
m83OWV+agBSKTtRHIwPRJz3/pgceXvi7lVrGEAmN2AkdmxSTfh0/LBP/UniUR8cT/HKbH97bRFCZ
qRKjsyQqtulH65Af1mKTSo0U/l5dnTliw7KcSmxRO80KL4PF967nHNvMiY9YfbtWVYWXTP4EGgd+
3BdPFRWAIHjx2BMlziW2axMUkjgaTRbeAxFbcvyTgTKqpHJarxCC7OKPzVlaEBhsbTRQCUQzwSz5
+MjiCYfcZMHyK+BYlFrRsDlqMksFY2vI+HjvZETNE9cOpvLKPSaBl6PaBOkKY1u1I1B6So/JEsC9
8cOSEPrg4vgdt+bHJOTmCaDkG35Fije0WAdU3y1bVf+xpbEUfhru94PFYnOJqozqWcv00KilIdOU
8SR51IGebtzDOzvWWoVBl4qA0xLc49HYxcde/dksp1c3DceJjsCbYo1URqEsCb0FfcWFQ7GtJHYn
jo5QTRGwGdJm1k7IDI7xTjTT0ehyOhp9YU4Zmbdqxc6KBBMMO/vZo3QOE9XBQFa/FSCEFM2vVFBT
NyjRc9LCUhfzs/OwvSs/bEuqQ3HMUFAbipNaugk/sJnoL+WI0RaoIzXolXScYUqe5uKYu4cTbAb8
6knQn/ZnKxzCpOWkNSbzgeIQULSTWKRmiYA+yuziYRZpZf90tCvW2Skpp9fmuiw2W5Ms6TFDOHJC
RaaMts8o8juxBHoIIc9oSuAUiYPbLmbcn0pH84qANHhah1QYh3nf/bDcLYiIu83pWHFEF9feCeRp
CK0lQiTjW/Zo1QtR3Qs0Evpfd2/XmxEbXA+qF67G0+dp+BCWV+cEXDqGuFGo6goecgRFVJyIVYjN
rKW1qXbJU2CdSbS1dwSUKC6M9UIHpyJcVrPH8eVlh4buUdFUq+s7SrXiK41oj5zWJXM5klpkD//N
N+9ZM4rtSCcndvpW7BrgKdWFAJ1u55gG7R8U+oVpYVm3DWf3xK1HCGyTV8UtiDVUeMFye3TvgC/z
ioqQgCMHx3lw+bRyNigBQiNgXv6ReRjMuvtbKANxDfQ3OSDF8AJYmgXoxcksxegJwV+iiOpEXuvI
guxQc+qdGkLiRZXGtrjpbQO54zo7F877Ma30ZO19fbFRI+fk7jSdm1Fwy7k8Jnm96mF4dpcvAUrL
hhk5j2pSSSgXoIzdSlHdz8JjmUAXH1eP98VGGnzGRgTIxcVolfYUaJ/iClLP/N+wEvwr0Af3YCtT
yX3yWy34OxXTdUKC1QouXqUwLNOq5IjLP6f0Sd2UIAqTwZyf5xFoQAzPx5xuxL7nPv3FiEoRcipi
2HZBmSbtjJtXhmKXeItoOL7NxyEsgAr4lvc8rv0LmMwFzFVMlj/W0M3IMMu+I243BfqiWcegXk2Y
Eqs0xwBFG/pKYS/a5JxTkOYT93fjq3dvAV+iEPe5v+FbbUAtn+VdKtqop9etvD5Rnuq+ty/VmA+8
dkgOTh3edHhIaOMj8pP5T+jWlW4e1lFDX98odXEKKcMgkTJTLKEz/FcSzVDrIA0suFBHBpSMmoiQ
m7/jAs9zlUAUvUS6yLU0h2JbbZkMiklJiKKXZ+t3smO6eu/QVk8Wq2h78LHZAjMJuh2lubFfKYQ/
4fEsXFLB6WPiiAJ58IVpMmeqCqCMdD1zlrAeAKpkBgFFPt7UmPA2+MCuahyv4GD85s67wZS+js4a
OEeIPxj59QCDpeiZLhNgZDxs2KYTHJbj77gS6EW/N7S6SxRV8Nhp3WZw/QXXgjCvasznvp7PQ0Ee
B7YFP+0WEQ76jD/k5JF8qPaJZm/MQ3nz8/6uwQAFySXvXFP5lTZzHTS6xyM5yn7Ai1KzcBcImx4Z
6thzvMRa2fqdGLUThlLqRrLNMAPFVvIjlr9ZvPlf83qz4OU1vdO8Eb95DOnRz+E8kIThxi7xli5l
GHAdXB+GT8UkwrfEFmRDKmDtaocOyUXM2fXoVltlT9N3gXLN6NtG2HtqV7bTShR6mYykHiaJhae9
oYYZUxogIIH7Cl/LCCpZ27wKQY9MkxY6476/axC0j0CXv4qZ/S17SyZ9wuXsBK+gbybcfuVmDMXC
PvbyiZMwf4Mrgs6+BVnAd4FVbOKZnHnRwlI0RBUXL4WmxsqtbRP/vC9aVhwqZM0a1nQ24UGibI4A
3JYr7PXpMZ5gu2dR8BF+qZt0vApGPBngm2SYR97SFSaQFzg0WBJBre/Llnm5ENv8UJ+eLd1Z+EsN
8ky4fr+uzoT4+vzScaYdaTPrEAr6bhmZLAmPvjqaWA2p0surdgvSwI0y7WM1T0u3Rlct5SiTMnB4
pRb1uOrUUq3Qw01jDfdTxdOcZwrpdz2LKUvc+dC6toHJzaoqSDoNESmzMXHlk3TavVltJfsq8Oas
fy3tZyNs85gOj82l3YbpUnP2faNBY2VOVxIAD5m3tWQkHEaqbbnUYSovmBeAYRNX18c2LFTwEJc2
jQoQY8HYPehnFI4RWGIPmzpYZsqgneVFddo6zUMcRUvaOl5bgXkF+vkr/8x8WBRGCvtIa3NIMOB2
KVWaQlDB8TKuIq6JJjaqeyFjFdM7u8sVRdFpPvHPQBFKiP0GcMTkWhp2QyTEe3M754OntduQD+UJ
GWyrv3apwdBF/ezin3j0oewpPLEwJQfr9SdIOYUfyMgOiT2rS3I2/93c/d91FdeK/sF1OEFzVTu5
n4a6zZMLwGmnfoUmY3HxtXHlBK8BP9kSPjztyGkgySXwYG2BDTq5U7PDPPBPX4Eh6FowjsazI0Hw
C9ULMFI5zVnu/+pJCsNczOXIFnbd0AE0Z7YMZYUqe5ib9pdvf1ia6g8WXNYvPcl7g2ioGDRo72v6
w1W6OmOxGMBMdnZQyi1+3+M7eJGcsiEUGPEF33iIcceybAyDC/3rA8NRsu9LcWWFnVenh+7USSxL
Rr61QQxfXN3ycY9tsAsjDZhd4rQkiT/8TcQFEg2+k3yvJeAZMFFgj0CE61uVr7yGm+d5COwarTDi
oRkqyD/odZOWUTQYZB+VIoP3o6+eZ6J5/q0f50TMuVPZDSulQIY8wHNZXLm+zaaKTqLsWKN/fOBz
pgy37DshS9MA8A97amNGlzi6m7omlG+lKZv+zc0xi9KIFbr1xxE4xj2mx+FmW64AUlATFixekCSl
S4yrmClk3wfv35wEWcRhZusWaLSfvPSK7+9mECy1MXmESFvlJEuaWqguNxrAimNcfd6BQHeDDIBY
v9P+NhLLdKzMJ2i3KsvuesfFwdmDJ158eH9R0BUgJB6rfK4XxBAvgNZ34TSNPWa3K6/jM8CywMpy
HRP6v/q3hSathAnjwSqaMgdePABBVNpqBK8ka+DEgl1yH+OD5p2fSu7AMIbjirA0Yhxmf8O0Lzpf
V803iLKvg+GWYYvPLKtiKRmoh7+xWE9GLYuVjmRMhWg6n3eQp+6MgPpZSbLP/i8uwKKaZEADB/Ff
Zk2pf63Du/BiOQdhW1/Qa37TBtiONmUu0hh/CHu4ugEZd30Ky4V6Zgh/uavPP4m4jUDhqovneHf1
gXQn4Tmgf7M3pqDFd+GuVGL+Eelv6DU4dJc2B0wDoOiPEjhM736XZ7xAq1cCYgl/X5t4TQcry1Nk
SwT9E2GAuUMNnqhBVEx8dIRnn+GqbS6/d2gsd9lnNsbbI7h5F6boF9Y6sbCm2Gw2f/1oV0YqiKcn
lrgeVbRu0Bb3Bnw9DmQCNMsGwicwRFmPY6/P0hVUWp4CkZsak/BocJwc1Snf6wLl1AboPBJY7M7A
bz9JUe2z41smYkh0bDh/iOtL173mOK5DDiX+9oWk/+mKnbWKBEAcJtpumHCwakYq5tMYmj5rvBhu
g02TB7o/9zaIjvQ+4JqkfE8fPoVGOquTYx6GFqIkXLoc3che8XrXGOJnPiJqHMVsianGDXTUVwKo
Mnc+XeAC+yWxi6X+n9UKu69HVAb1i7giaTa1h2VOnUzqvL+o+SMcCn4Uo5HiN3FKXBJaW2VAKYIc
9UqyJbaH+VrBPT/aVcAi1oGvS9NeDIFmDG3gMdfrY7MTgBuZZb1Knpgp64XMMMsgSmrHdim2rtCW
i+XkmuSeKqRLRnEzjXo63z308ucTbTxHgvJNfIvBkCY8LkSKG6Tgiy43sOoKPg5/+/qbUIxoMZL6
sqYym9aVAQkCV1zKuQzLMLdK/DO7vow46avLt6GbY5PzcD1+UxwtXKYvAew06p6QuND1lnndm2JO
yMG9pnRBJ096T4YHZZbGpluTOFdqaZz4uzc2n0hV8LsN0SmM+PkjJAz2VgsZJd0ibwx91VrJyIZA
NmDR5DnxWlHrkIQJRxiHJBv1sSxn9jX/zVhhA3AALXGFYgN555pIGU+LmrIdpQ5VO4dZLyP80J5v
Lox4PIJ4MssC6A9nhLWtPXDxL3VcBHSHU1EsNfra8v9w60rPRbKytuHYKTC3JPsHizhaZ5qqddj6
OEgzVirbv91ApacyzPQECMt6o2s1Mg+5hZCS/TXJZb8Jg8Qp/WEolR6TJKQNlGYhUF5u1yNoVA1e
AXww01artsm/7sH8MjHMvkcXX1y/VtKrRIcF8B1SY7vP0glC2mW2949FZRwvXk4or+Q3hmzMu6Tn
VUQJfLGoyV6/6byn+4A5QJbxDks84oVjFXiaXouOl58LtaFifQI0phrZ+pQJQoS3a4rtvaVK5jsY
EBfYSeApnl82vI4ZwPxHzZ1C0ak2eioGcgfNw5cFTsDElCJ7uhflmjpS+S2QLyHh7rRBHIOo8c94
SPl1/J5b1h5EZcdHwc2tRjWWfcKrxJ0PqDQbWtbuRl1g8s14ZJKHYd9nJd7T3QJZJf48uTaMOUEW
O/0GUCIuTKWwBoh/pf4RRIcL4cHGUtQc5y2HmoBFQ8VlEqQa1cV5iHtSMaW8mjqMfKGPN/1NVtWS
RJBkj4qdAv/A0EpUlI+jccPNmKTkAxHNaSZSttka9EYlyxiYh6ttuGZP8InUbpmx98XF2fD+YNzp
e/Et1Rdd8BJPyC0o9H709p6XOE2BCBBeO0puRBkMPXPUzHl0v+Npz2boQsNZbnxlhk051fS6LQM7
X8pP1hWvyJuuz/uu5hR4g261rAnKG5l5QtQ9aFAsNLZOqvurAxNAgmYLER8CfKQ7iRgpUnTjl6Ae
gaNR22naJJkyAa0a4oQaCcf/6cAgB6baLFYtGk6H/p561C5Zcdc0G5YiGy8zXcJWfNu7zN1m0FU7
MwJZvrYg2UieltbGOcc85/yy717XEMqfGSQY+f8mZAJLBA/A7pMZ+uiPywHFVCG7UC+gK0Sid0Wp
z+iGyvh26I8hXhFyRIgdO3zBPK0/fzsdN8IYuGn5cmdXyRll2k52LmOC7jSRm1JdJXcaUI4cpavK
2KUXh87SJzxjb8Sqi1MjcLiQmevlkMciUvyVJjk1QCRumIOeAmF8f6D1Aq+siro76IkHc5DQKtDD
TXTQlaM3CbVl/rAdQaMxMTH5C4oo9jqRyVQ7PHi7n2RRVBMmywnJvt+hdabF/olgp6Zh+M6gbe0S
QGu85GhxFJ8DUmg7rousB4dx8W/o0BrtRpn4FIhk0JLVedZ8OzF6c9F3+gmWKlDyXkbS1Lz9oyDe
4Fv//LA8aZ50lUcaFelCmCXvtj3390iOdcOJKu/5oRvFh3u25SuzxIPGOqNYETn93dlRGDoGJ4dK
H628kkq4T2eOBj4JrtDhNlOGUg5ZpjY24c97VoJX2B0WYmn8y8hGxtMTrspW/8ffXgOuTQjOcENg
3gWBOHYxqmiPAKfqa20FiJ1vCj9ssUxYOmjTwY5YgzsI+W1n93Zj+gSKULStl+zvEcdA/SRQHv/b
gtBWiOhnMYAj+BNjQ8WvOiTTIwI0bNqHEkV3SVkCvoDUDLvfuItA6kk3BsRbv2RX68tluvQycy0+
V2wXja7hQnt1b35hJQ/3CtSPjt6kuMddz1JMkwkaBcQ2gziqehRydRc6zCQY/nEoQoh/87RC3eUo
3/p7rqHGyP0UjW2Sp4XQMd6qpm9FILoDnICM4H4+EMHGUp/lEeM6htwfi3KcMhivpdYRiJQUTpvl
Am/EcU1EoxWN06KA4iUBmLRQfMqJ6VKn0f02lXhvdOOHYYl44TxjuDHV+0omlo1/B/63PgU7YR36
3T7CXUEqI9bAMx4ErwBEK++QOqV5OoA8dDLEzpk8/y4GT6z4VNuy4AaHZi/Ih/BS9ahNX/qEaXBv
VjND7OgzFm6LgKw9Rcfog2BF1EdYUDcf4cW+ltjdcXKzi3OhoczLGu8FekDLWpZuKjTh3v/YLD0w
OkW02W1p6B+OXArHsStrL8Gl8y/FZpvlMIt2qexJ1VtEDddN50OmdtMVLT0INYSkMDzwU2jnPlUg
w8WudVgWVR5CDX9glSlvERonSnxZ5+L4043kYMRuKFkvJ0zou/ylFG0OhF8CiWpnkUShhfVShYqc
YKxIAYhk+/sAY1btOcuF+Y7DrZVz0tVR0gm81zH7r7H4Y/DUAjiTTsi4nzIQ5RmW/8YdB56j45e6
UG164J50hHgTm8Uz5SHzgf3yY3K4pJnqG6DwvNZM3n9SyLc43CKJDquOpY2HXGE/fvOMsef4j+82
wNgYqrAgDWFSxvbRTgghug/Qc67rcfCdPE8IcsZM1QMn0hfJdVqZU5oZX3pVMWOVb0gV8E4vOvAm
QGa1+2zS709PdJv0Xe/A97jn+oo87WoFAW1Zelnq8C1eCbys8UzPKF4KkbxU6eT/radxdRdUHMb/
2gBHddU2Et6TH4poIm4U91TtGjgSjebqiht7LJq7NrFFsE+F9ISTJFM4VRG62zn6rsSdO7Ct/EbH
iwJGflpYa63Y1GngyfUTWhFqvAcctCvJ3wWx9mo2J0kzmE1qbgXi9PdFcqZesTys1HKMS6lRnMaB
Q9Uge8PQte3vH2q61bA+NdN6Z63RODFPWelx9/Q98DKvO16ZfEimopVzWONPl9L0vN9sYwnwiXAe
KFSA0HkCAALlmmlKG5805ip5OkwDhdQt0+Gu0+Wu1slrGNbs2/kE/k+i+GpbrS5SMDmmgcn+BZgC
j+TlhNipXohwNNeB79fI1bcBWFWl9K149p02JZuSyxQ6Ys/zQxWAqPLThORVf3DA7QabJM9hGuur
fvGye2IjudldvASq7tsaSsuo0ZPLCtXZIdAf0I1sfJSWgJ/TruzICYzCo6ekHbLsr3jtmh8sP3Hd
Oy4c2HjGFIObh9GOIc/0TNzuT5kc7NGCF16sdTAPWfTy15bCl+D/Mv5mlAbyjLufa0MHhsFnw4M6
Te/+/S/8Tc8f63iQ2ge50nU3wcm2NdAbWzM+ggpk7LbJBcUELzXq/Cd7/2RS0GU0Ryjd2PPaQKFQ
H3wb6y7ohzPy1I4RrVYCGIHKVpxBXQCTlk+8B5LNWWKEVj2PBNnumVVxC+EsWj7z5ub+zz3G/Sln
bg3diMmTJS02YPMUWVxtzl1pW49D3z8+fH+e0mLnxzGH3ShvngvY8+6NyA9azJ4JoqMmmI8hi4vc
iZl/uqdhCy+j0aJCxDqWAN7WGKuuy+hr/jzIUBm0KLJ214iEWHwng2BFeze8keAigYNi1YLHLt66
hxXH25ix9WbpUNLeSzPYzYhqgEt6EBaZFn1gwzJQingwcdSyJGpdWj4ZyB3FgM7ugxYy+z2yBP8V
xbMt6ZmDfkEU4ab63ZL5BUEUYUNKuga1mvQ7YuNpPY+gt+FBed/BmpfJ2nP5DOXcRIaBIlICihOY
ZohoqpjngNZZdPhr/K5mf2omZ1i8jztanbd4hdRDw1w6KXAJOL0LgqEr2K/awtOmjl79ArLMW021
T8Arn2NFKQYnDEuFRsjY0fe8CzdLnepzXKT7hmLuQyD0MjtvyzXveKz5PqImmeND9kYoetPjOvMW
Vmew+9toiPvpC9u6uMBPgJQUqYx82XcOCS7BvIpUgKiDtIvnZA0uI23J1uaKMywSMvj1uhaEj1CV
rgnuhMkSb1bGdReaM+RGkOpb0CmU6K20x4gfQcHOqI6ThQPMmjl/u85i9YIVou5YIQwNRfBz4JTl
S4Yvn/8FBbIwK35/EiNfRHRrlU5ov5duqOWfMPP+v3/5q92xgdhnl2jT+3ifpSnKWNjBhYQVvLtn
pwVsoLXW85fHzgSmu8QRaPlYrWahO1QEeVKpDOpb5Aq4TmKffcebTJc35Xqwxw9/tn4olXJVB9g/
Y8OerZuSEIrExT7KOvTA9/ktXrG1uBoL8hySENApYqX4VQvCyKEPvekYelvT2nZjm3C+M9byXila
erRw1dKljy2+qHJ+TDVU7G3Ox/wme08XwUOqoGM/ZaVus33pyq7AkDCxMgW/ETxTakdtlmQA9R5O
qYWUVlXeb8Ee7G6L188I44xo6/KZ6VBiL1vbbaLv7k0r3CAzr4t+P2KjMND7UA0eqGjIaHyFN1/T
bt+2uwcp3O67sghTvZomIdhz+mLoeDC2xustitthvnoT1NyO9C7Fkdi3NVTQAzhIhmJITEgfEXCX
3FbY++ks7qwiInxOrDhzbV5JIJiq3EE3AjmO/6NrAWz86fDAZNc1ZhgXGnDuna/HX+xbz5ZXLT74
3EO4CSJ2L/mtLVp18mteChb9cnHD37HyXGFFpiYlLr0jRswKebSg0CHmUdwSY3+YnktkL+oNqvoD
CGjRsbd21vlmtD7Te2ozBdkCqrDSnfJWtva1ut4XG/K4cq8PTqYLsDbqu/G+Ci4dlJVs29M9AJ4X
uCdaQnzVRMsYiBiJ27rv9OtL/ykRfVENeH49IfMEBoFrNzDwGQc0ZBgJlyoJW968oVg6OhVmL3F6
M1zfWAcgFxZJjZ0xwBfwwxihz1NQ3rxplOYK5LgO5eMkqWCTpBuzydjg0DPfOzYwy+leDPsAbmo2
XSQEftScjBAJzaLT2Dmg6IBPvzOtAZHzrHc337VtnPNtfbWq+VjRBVaV/A131TQSu8pZ25mw+8N8
XAnR97ginf6fj1rb6COEl7u7L/ZnSc/FNxEBQvhDRYvyKeIzENovpVWYMDelzcWcZ/98HlvKk7OU
PWCRDQnZgvisEepuNhzh9ealEAtPs6Xc6MoHLLt6DmlvjS6xrKpGJ65YzycAHbBxXEgVlCnp54fk
VoNw+4hFtMbH4Yq/GmGYu9BdZVWg9eDkCCMQ/JwOCM/DX8Y7EBzVbsU1q8sbMbskEXoHd7rtXzzI
w0aMaZDr2raQFFR9TfC7HYl+zMNCZX+bvMFtm5pffA2AZ+33ah0m/N/4e1sqS5s4cpobGdBQfE6Q
NGz2PlmE2B7rcJrIQB4hqx/eH75oBm07whZQi865fAsve59AviJA/uBR4qj4J2RWnv1poLME9cSR
8L8V8heKCF3ynikB5x15xDGbGdoJK6wcgg02wwynaZgsyekxPuj+xp7Dhwbr+WTFOPDIxbnO6an/
RDlpP3aiSu1G2dIzOLqSL3XLkZ9/YS/lBT8hme4QeKUb2pa3d7f/m1lIN6d2YfGSObcAjX5un37a
keKpl+wAt25Hhu2G64engQRf1KLTF1czEEcLfx/fr0tmX3VJcGhn4jHRDhg/A6Zjj3czZDSKeYb0
P9E07XzICDQevFJkwyAVyi6/JtHbtHZ8Qf0i2C66cU2USShumbcILBzqgTECA2aMA46ci0bTdcNE
3tdzpHuZIc3tx65HYv4f9nLPdw9YwWgB+oubrrqwT2k+yixPL7BdS+kZzkgkUtk8/tMVuldTtnbm
vFJRf+FYRBf3PHXrnMHTWFTHS0GfRIrFnTQn+/uFrUETxvySUadZFyK9EEtBhdV+Sk51/PdLMsPj
ZkcqjZfPzjIZ1ePzIJMVAK1C/IaAwXvqwwPQEB49SOPYDkYh11QEcdGRhlpjwatpxuUmjVsEG5Pa
4DurznTUPOlG5kNCo81d5418XleUNB3vjgyswU4JIMvOkiW/rJWhWWTTJSVTo62PR/DPMVLq43ry
BjAKXMKRiF2T0mIHSosMm/tXH07oPl9WGLOnBkLcSq6O3N/S6bNsUPdHG9vtU7pZ4IxDLbdt+45Y
dIf6tbPqxJ09swUXxXQePPFAbbM9H/WuOAg9dW3x5IvlrsBS3KXjLGYc89U9h6EVdwGMHrXkj6Pc
c7ifeV8SlBT24jOBMZj1Wb48CQPdvL7c1UxnUinSZJDVK+XhZrvSK7YzRACoC20YfWEwocuIzLfp
uNrXRkuIFT1MzwcRFSYxEavEHIiZQhmMF/sJZaVC1DqCIOqUYAUWN3m6sJ1vdl4pkXo8RfO1yII3
MKLKbp6Ht0ZBLX5RMWmFrDrLt0BiZtFrlUg2Gc4jAULK0tr0V/9V9UZOzENi+xXGZibgezUr/9EL
ho4E43aQkCEVRcdIS41iCCxJ6rxQSDuauvMFgz15tPkgfU7+5ux2azP2CiAac3Sj3xMclQ58AroS
lC4jvjTjmJ65l/KJuZZPFqcvpYi8RaPECGhycF3F1AJpNaU+v1b0BFEw5QLl2CFvpR/pzUYrOIAY
94kiXB5IjEFXg42sEPtZ4s78X2qkVIpa3AvolQlgL4aCM3G0NaV23YWWio2JzPgwMdxr1zsW/W10
PfzheFA9Ml1+uddDr8iFqVzLPVmXbtC0apA8k+i/IxrBo25blidQEBmHBZFTwGavYksh5wuYyttS
rHGaFleVnn2K4iPo+qfqO0liak8QW91pLTPQN4Vk2v+66it7CXbf+iWKhZV/zfn34JpvYp+s0m5H
y4pCA1FFKSuO/mi568ncUlYDlqVJ7qPHv4YR2xA0X2CM4TR3t8s7Obc7/FKreDJO1aCLWjM4kU7Z
o43+gCgmgSG/KqDSESHmZbdnlTFfbw+dHo2ReaAwa3j9DwijXS9QMTWOhLWmbzij89M9Gko36dnp
+9FXKhFc6w3ysQJsawwHoNZ2Vp5vUfbY1nGEh4X58ep3RADgGcWRBiBeMcucPW7vFCW3snBq0T6J
ZohdTM2gOkk4gUnPQcdb4sHO757QMYAAJeQbnfgooTXdNw14+wQJlPj+JUg/GEKI5l/2mWW0hWtO
HQ5BoJi5N97unR4YeLwmufipQgwVoT8ja6DbisAT1Yvq3tjNOZm4YODeTfVODwHMd0J6CWl4D81x
cnJTc8iimClEoClUpmX32etsaaXDKTxU0uSBuESuWnzoRqDYD7ZSVFoJkoTILfM9MXl7C4wnEYBC
m/hy2jX963AbKXA9EbMJU0kzPtmDNtETe0VrrcKFiIJJqeEgREbTJnU/zTxQZsGZmSthA96COjYA
/NDfNZmfFHi+SBzoqKPys06QncGg5G1zH/mVF4tupMMb4f33HefaXRl4aMVq5+xtndqO96nZin0C
IY14Uomw7QlQMgDL5F8/ctXIfe9Bs/3KV4ecjmpc0i0gwDFRnviEOz/VbUGUpH2aMxsU0Y0PfEPa
iposHKgCskup6YrgR6O2CNde2FxVidCV7d+kyXT3Dbl9ipQZKDCPTheMbbbd/4Ho0nrwUpen506A
kpc8xejet38rSsrSzjN6lprewnoX4tY8EjCu1gArSQfoBixSYaM0vn2ET+Zof9BX1HQpD1DcYGLF
75ENu4kgR6KNuuTPOh9ofXdt8/vHvuSzzOhdkZFX4z2nmiLuNMP2C4tHFBpl1WJg7vhSkbB95t7t
tbCRk/yq/kX1tj0e5GICiavH82QxcKpAp8kdAOAuuNbiiGqMRDBML8fffFDAaZy5DAJgZGqvrOZ/
ANddNpz+YyVX/ky6KouRhy5uWlSeMi1GKL+mcfWRa90297u4ZDnPCXRqwzEh0aJXBdVsChdmRx7a
NOS2UMo8eYR6ryo+JBvkN7oX5L0FFewfzSScoZdwX8tcbL06mBV2j/Kg92SSEU9KTJudj+39vY5S
NUJQdlosIb/lyJ2/3q5h0HwWAKOC5xqtDOz/oucO9PFzrfY0AFYLs1bhSrxMU53ZQJ8Q9uJ48yqP
wDjzlkiIVRCLmHK5CYd8yYHXxvHXFp8ZSHIgPGZALg199WT6opunYJRkJF1tOe3a30Thn75b2zjH
MtLK89JJ0Hb6nhSYg3GwLXB1ljDgF5v33tqLhv86q75aiVBiGZ3KiirWXsyfSkYN7bGubINoEFAJ
913TneDVMOa/BDDtRyb6Xge+p46vBrqN8fJ72fTPQeb3Amf1P3q2YCgKxjQwmdN2n2JUg6S3I/Yb
vD0JayuPyYtIADW3YqrwsCEAJ853cVUf+aWUJG+FJL789d62X51oPUElCxRtQvhRVB6xdMfMDPKg
5BG5vFnaFlFDoKNqpUlpeT3hk8aIbGjsXnDaIbquF1vLpAMZb+eNIdPUDWV51nk+gTvjCTWnaPRZ
Mg2OX1r3Cf4ye4Cmk5ULcCTUn6MB39OpzBF2iKwTp/f7MVtlL++r4ZnMc6ufXtCbd0ZJYwiiCyEB
8A6/YD0C4gtuS0HX1ct+D5G1WSgv2GC5kgddzrG6dZfUmvUeY1EcXM8oFv/HjtmirQVSCc7zxbnW
CAjRA8vH4AwP3P5UbfIUIjZgv59SoBvEXYnTbt1BsXKszAQ9GUapJhgaGaWwvT2zioamV+ApL21D
A4yYhJVTTyqsn059jBKoNbSWj007Z3FsEiDx738kzRKChJmEfnganQZyEDt/PbjZJMTkKepBe6rt
csuI1rcXOtIqfMqgxFWotWBITjQWZJXkbgsozKO7+ufcOg7XCnAwEGP6q4V4idzN1b+MhsLlwNzf
AUAkzRCfTZN5xfMQ6RPOLTROvgBYQ9jV4j0/yPGpJMv5p/M8uUFEsDI0pyKEBZubGR60qTnTj1mv
o4L2neY9k3uWt7a11GX5XE8YhDH5l220ETqq9jqUvtNF1p4gG6faXCd3j0aVE9joeGffgGtVZK4d
y1tYqLSHiext1s3hffUgw0Wb2mrqUn4KGdc1iKjHecXZ8N5xJSzVJAUaaQg12pimQgUzzOLhRsRx
gwWjnQQxsNSrR6HTSGZLSRjILg6dNJmrSKgVhIUCI72OunAnCFDOz/hhLohR/YOy3z8rKkKwNSW7
K9U9VTNLyfKFcV3q1J9t+NGQKZ5pA+dvXzCrWvzPL92gtrf2Ktg5B4vUb3HdkrYobdFiW1ARATpm
yLVasobNPuRMnY2WJDFm+L1n8MwrDnqtH9DJ51f2uQkELfy5ZQWm1kV8M95rQs/r3LvW4mvCf9D/
yautpKLlQPz368fge0unzsQ7nOz4YRzGibSYKXPvuosPYU067ubQq0XKX+EuPw7TKwTDN0wWbpwU
Q0u0kE8so/UJ5zpo+V2U2LjshA0r/WE3JSkGo4aY8nY7lsL+7wNPpxaSY6akmC2ydZH3APxIhiFw
cX90hZSA7O4bXV0QLtIeAkS9ITF22cNWounDu31YDtbxS+vVupD1Dzxcga0F78NLt55f5tBRhllj
KlKfKNGxigXKhIbi5RZRQW98M05ZUvSx1iuMs7gEGs//DMVFUbxeP/lWNhzexreWtW4dvI9vdO9A
06Cf6PPtFjr49Bqdu/fBGOsmj5JZjSiVUslCo6QTXQzw5K97Z645G4OXamuaOyS3pr7t0wQt8Qqf
eRyodg026JPjIO8LSKjRxNS4rjPh1oxRgFj2lT/aTD8pwBHkKMlHL2L8jYV1l2dNwLZA1U9OH1eO
0nzAppkSF1Jv7Yl1J6Eh8KBz9A1+/V37/xapaIs+WA/DmiNcMSJEWOhEDuntxkLFCx93nRMXbs7A
OgTcIMDJn6kUp2NXIjVy5Oow3M2caNfxS+bvZZXrAkU77tMTsZb6DfBoyc2nvFNFuTZ9A9orOyt3
yJcFK3n8gUV0TdplGg==
`protect end_protected
