`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ro9Uy6Pv0undFi4fHs6c8yhpOwPRZ6Z2m1F1+8SP0JOt1KXqaubbf1mCOZdKYaaSmtQhF5ycT3kA
gEkisnzvww==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IfFFT2r559os9FAUMtgrdhputqUfsl3j6+jBJe99FmkIN/7QgiANUNq2Z3cT9CElrO162qLsucWn
ZIxxBOL/tZ9URaimBvt93fOjqr5B/lURUSbg6kIJHd2/fHb7KjG7hjYN3//m/JkYkMVUnd8qxV+a
RTnd0/DuGlHYHqre47U=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QT9M9Zk3tRRumRkGhXlo4JpDgHjRf/7iQiBMFbiFz18pwf7KBYTyFabrCLexxFmdviLRR+KB+sfg
S1SB+8/3qkpI+pxC6mvL/Nhui4ydEeO4ETkbmFnr07fT8JqlqiD8azCXFZhwaiLYq1ZfE8RVcqBA
774lVlATL7RcuQcMdpds2/1fC/p2ckCPtZZPPBX9Vk//yzgs9arEK8QJESGrh5l0bGxbjHmbk+Ld
nBUmMCky9Q2ON54nTSslEXpDEOvSZvCOISpjOvUVJnAPvFHK8dnrPIiIpWaxFImHY7K857exsj6q
V9DYD4cBhHT9qEIEMpVECyomTSY2SfsE6g8SUQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V1hyvAJS6HBsYEZvVzGZjF2UzwgBpTL6oMWziSiRZ7uQuBDfIvdXP77FPPoCF82Jbcgwu/HlKzzk
gopOBrL5mylaKNAZiIRegEfdehuX8Wj4nacsEB9jFj3vNmuWB+/tLmcS519djJKFm4VcIE+BVjcq
EXxdICjzvVHQIvhi8Tg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m2El048nrbQICF14If5+r9/kPY5L5cnMPZy51iwOZjjE2aeL3EP6yt4piTMyzdSyujWKKskwrzKv
m+j1qQMbL08JgO0FiTPOydO1Ae8xU/IfcCfmWLnH5MOKpBfnnDlmD3H1D3MJq7W3FFkFFt4mTQ7a
z43HMQOct4gVfg78njNNbiR5Gnyu9MELmpB/jMFuOYxfOL2JS4zC/SyHW/ZxKFJw2EZdZTCkLjyo
H0nseCZNMeRJkMs26fUj5ukkQT2S6m65G3v5xwDYG8waHOkS0QpDYbmdM4TDg8EWX9NCJDzSl2Z/
J3orzClpNwF56lfR2etX7uwXACyX1jIYZH9N8A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
4i8V/PWWkhIICmI+bBHVFPZ0aE2toc+lsDu/untaHTq/VMKJ8ZUOtVi92QuHrmNYwDCslQhx0R+h
ECGcD1bO0nPe4i+MpgUiHuwRaQgrSCjjN3+qNLsszKFF54ZO9g1rHbDKMu4o2Gh+f02nOH84Y0Gj
lfT3KSqI1jrxWPxzxtY1dTQnv3YJTkuSBawEaxl4nUBb8X07akLeNDfLIeRwXLDxIx/KHgxYjSMw
biJWPAESSsdcPQUpieOE3fJ7i4ByqUQ6FGMs/RsYWjpk4f5DRHDArPU0n/bvCN0QQr68ufe45k89
mDayaZx32SytWx9qiG8KH6O5ymVou/iT958u/Uqp58S0LT2XnVVVtrWr3ePXgZ4lU2jVDulSTeML
Zbx7/DATUDOneKuwetM8xaGwNMtoCgOLs7kWZelFjOcWulXa88iPsO1yCo+FGUyJ5x/PZYPTC+i2
ABc2o9+0ZFpN3AdJYZA/YJqBey9+kPNQHTmGrrP5UI7N2uKiucp9qUvAUjAGCzM3LYhv2b7Jur9k
CX99Q+pRvsL4Df9ZKz+zgbzYt99mXRLw1LitfnmPRo991VY1hYm5tasXhqaRNlmAQgrp3qZGvuba
qAf+Ehjr9hxHABdzwTrcVLUTdbs723cYLSF5XZJRTSTA3DIK7jrKi+h9KPJjjODjrCIgDHqo/+8j
vRDZYj3KgVBRhesBDbCGKSMFam9pOuZOfYvg7EBOCsJjk7KRAE7FIPESnbqb/My2JdLEt6YxmDPO
gMTi8Df+x9av1B8R4ykRLxfbvXjBqyh7C6l7gT7P1ZHqB0HOVf262sFyhp9VljzMjYCDYnpQRjl7
XEKs6MqvszTyeI+juQqlIyBHdA10wmato+UIxi2GNVChCdl10fbFplR469PlvDtp41T1if6YfySD
WPcrE7aCvPGPrk8eUO7EHN2F31rIrotciqC/A280Mo/E7hB6YS8XyVmPHMS8I1JvHQVUThwWH5A7
OM6ntHmd04vNFxKrEsFYsTO1Rdu1dlwhKKHkpFjSem3noi0gI9lWSh0lsWNz9rIBQyUbXQw1zlgD
poZcCC0AGYnZwhHelPWrgbMiR//K3z1pSGnYDE/BfL3dcvHDBDX2zueCbeX7190NBgJenQ/kepCa
lpbP0qeGE6Vp33aQmCcEY5MTmu8eGFOZadwekStIrnGAX46tu7bFgKvXL6Mrz6SiNvIPLR/I4U7r
GducBm52zkSOrSvbrGYLqtkLPeTan18IN3BwtPUFIiC+eAadUXZ+fqeCyA/tnoQiMPlkNplwoM/R
3BBUJAEfGV7m5jGyUdp5be3SORWtEu4pds8PIQRhmyys6tLoVIZfiCiwMi4+JwTLzPhtIhdjRTk1
0aGYP5DGW1xgXBrWNwmnnZYvKkdHcdBMi56AMi4WRFZ9gIM04PujoK3oBI6mQ46kJ2n0vHIb73qV
MqSENHLjDL0uwlwmgnI73QeRAfq+qneUDBf0L/zccwSpaouhoglqOus7iE+D7v4FImL+/e/1Wf7P
VCdak0Hlg3YkY6pKl4msj5drwXXJL9NhutzB4kOEW0wmYkgEzayJi1JPdUw94KRh01yyFnBn9C3r
lBS/pNf5e7tE5gTN3z0NWj3bSbwvIIyxVRmn4JUyTM09Z9UyC3pgI892Oo3Yscc6GrzeqHxJHOma
jQ9JEELvibMymdBK7vR54MmkWRvHjfuFJOmLg96h4zF2DJW45TDyhTlHULkg8YJy2qsSM3Qgea59
iqfJqHzYZUjWwJIPR51uccCRWzMpE5SkIQx+pJPkJFi3EQPTf06cKWMrdGfJIR1czVxvLow/LxJu
oMMd6lOGpbXvDYMmhmQUErR78GRILPZQE2isJHH5f70sWKhA1WEbgs+vJQx7KEMS9IntJbvqgdeb
norFo0Q2A+7ZH0Cb3YZk6voV5Dh51YAaYek8LQnbipF3PGjM/0IZFfbu8MTN5kJ4u10ODdYN07/1
EKcXFn2Qvb6vuQGLjMRe740OCPL6mLNPypJGBJjV3Gyz2woIYyAlkAlWrzhzlJSVApqPre+ap8t6
inWxBwpx1gsDkpa6B4XQ7GbyHWhZlfwQ7sbecr6tG0jZRJv/lRbobGBZ6UG7wIpGhVTFoZHyaRpD
/mdHbadwEqmjZxKbyILKr/d3rJPqptUWA0N2Bg1GFGXXpMs6UG2inL5SZZ8l8YUlc5MPSLOec+HA
gb1GW9xPDp/TwHxzAMINdk4iWLYE6XHORqarz9pochkySJs0hIJtjuvLXSY0Rq8T6herxBz2yPpi
KtCCnSd9UjW6LjdPpGY3ES1JTZ2srT4VMKAhIOFE/SBPeN+kv6ys7myJgjaX3Vassk/mMBrM6O7m
Obefp7NO52ePKSs2Q7WDxh/jGhrBPNVEN/HkW4bl7tKI2ooTjgdmXcDUlf/mMJY1WNgAUw1O8UfZ
UW6ypmoXciZKrGqH46/WsAVJJGflYEYPWibnU58I/Q8fb+WSlZ+e9Ab+DSHUu/bJFP7JCV7CFiOY
YsdmgMIGaJjtDZ/vKdVZuRSzVBjhLQJyYdkZWlFUn7kMyfY9z12K6ZszsivLIGYakN8HRz2isn1I
oCadesddwUfF4Q9ptLyT1Pube2u6ta89v471h0EVMiQZaSG0LQuXR1ZlAvOLTzw6J3NSEuwNiMQt
CBVFmZgLofFSwLQ7bQrAda7GCnPUc/EKTjmDMma4rWPqSmRKBhCl4GFjpfl24kkStK0MqfiC8P4l
TZN9kRFi/Ccq9FwVbLXPdAnyjVEeEcFftIpu2QAjLo3geR6yfhZLMj+dfH1XWxxnw+D5UISSN/do
YXMDiswLkxCGx32HjfFmAIXyq8TxKgzzmFqGdjt91tDWY/3mlNXSK/KvCV2jh2GJbqv6qjANTckT
5VsNkxlIZFN2Wf1dFGff+Yr6pEXGZ0MVdM1ixPEBg5ZBmFA3aZVDkOvDgwtg2e2pr3mLzQK0gsMD
6HFXi1QRcATlDnaZSCR2Uy78rvvuE+JPd2S/vO2ITP0CIfBCEVKdy/vIk1jtF67w5TMTrEXzjKvV
6h6lSa1LEY11hW6CXq6jRa+p68HjY5eH/C3/omnPNzw7ETcSl22i6kCek5KJDCUNAI0ai3p5zZTj
aAhQSof0gVC5frD5beS0fRvURc/2r9eny+otUHCSImVpIjrcln8ZuAvLLmUfMcwNQ/3RlPcPMskp
i1erRTTF2+hEtEmY0jPux8Y6yYQAOVDL5A4Z2Z9Qn46vWW1sDdkuoxxT6B7fzUeOiD1Op0FW2NZ3
7Fa3Pqrujh/sMI3a/XCv7NjzPAWJRYiJgO5VoxD8BWAKj0mF/LoRNkg1PJbKn1/7/kDi4ewZ0j4v
6loAmNSgZfy5SsAUccVRU4/0Go7lGzkrDGMP2C6TACDZjyZCxlVrGIaEDsNV0fZ3pYiGg7toRvRN
lzgstu9Y36eqNeL3xdPZ3wx4LoDuhGBRM2Q322JCyZQ/rp4/xh4BXcDimkEb+2mRy3ABEDhOcB1G
0v+frqG4P9z1Usky96plBNo3MoA0oJmGTtur4LvxGQpg/OlIp/zMRt1wobDLgSiYOk5TBSP7O5Jo
ysdsqeHc7G1TeI07TcJZR/gDzJ3wOfrOgNan9EK/l2exWmAXf9Vakyw0FTmgNJIhL4ZIU+CKWYSO
RAum3/4YU13t7Z8jd3fSJFDGuNBWmfwpnLv90KUO4iETugsTa9s44rJtJ8I0kXQBWatmd/KdAjIz
2ONBJtdFpIP5Tj4A1T07W5hW6nqboCVbqxQ9u7OUy3IUGU1WXMdQpPHtZDKQ3TdTK+ylfx7jQl7c
btG2c2SlYSQpN1Qzo1drhofqnCYJf7uR567u5Ar6aFSAvSKf3XDuXLyIdRIT7LpMOFX5ivGKdK9+
eF4H7P46c4GTBBCbS7dDNAlInG4fCy8Itk+4vDysmIU3JmlWYZmLa1LB6MnY95CPKxlWxg8S9NHj
yPTuirzkvbt+0DdAA24pp/BAMuS/UY6ht+6Z+OHuJBNXoIbSUiRjq0qONCn8+mrBpC7cNHnY2+Pj
Fy53DL2yGhGb7z2s/dHNOkJMO3boM4V1Op0hMvJt1LcGkXeM9V1+Ac3w3KzKSMiWIaMxb0XmEp12
qO5cTcuRq9VAbZqdD1Kx7XlHT3d0u7Rr31C6QCl/xlVNZeSOlEGuZ+JGHZtJUaqJK0vJLqXiWhRv
XmXMj4dGORrDDJi4fUR+BTxjsJy7nfLuhRLqVSbjspjsHEJBGE2ZuMEnH0vV/Lyp/Fm3lrf/7pv8
DUx/evPLUoMMc40HbxoZdfILt8LddYZvxy3ncEv24oVRu9hJi5xoVjXwTver7WWtGn7rltrkeNJY
yWoCEdTO5MFfBNwDxwMwXOtVgyaOUfHnfHpmYa3ympWApuobtUP6sBrcE1BvT5L87ItDOyoT/+ws
NHPDa/YbFk9S6nQWqCACKCHg91HKhhRAGV1AipIx87vDMOSs49QSgsCWdFzHkG4kCCAc5eJMvH3c
9eN77ASXtQU/Rtw/Bs1lcDJ9DYfCtgY0sAcp1hy5gg5mdKqfiNzHaQGRgMxHYFusHYF5AP5zPDr3
RTHy4uYgIecmmsN4UfBOAeMwoJ4PwvmW0Nx9UZtL/NQYIoRYi+ZHXQh3ZCgn+hBYLXzJ7X7Ox7Um
yvZqD/a1/QgOun7QqZwF90Eb4LXCw3m/ZoPi2xIaElmtKqsM+J7CrPcvgkVAr6OhsyXcbryxg05h
qWqQc0USvPLnY0x/1fD+6LCY1IZuVTd42Cy04Nrsbuth9gX3oSzGaG8j4lHLdgP2pzsQjG4n6Exy
Evf31LCFtOjIjLcul1RT9t1mkRjhtBubWgOehtuvDRB7uD16xGTNbfeP9F+NFeVVOmX+/47rwRJ6
V6L0wS+BZN8bbJzcSn3xvSOaOgqu4ZmqUxoTn7VvWLJfo9lYbX9meQw/IUSnKOW8nRWvDfz8UmPi
tCPCgieE150Xc778TlPpCF+HMjsXaaVdjEH0ED9Xp3ov9Mt7/yft5LdVh+3RIuh/uQLThLKwx85B
nFptVlTRTl3sZQC+MP/6Us/lw1RlTuoliCUYxJjrfrP2hGZ4rfnT5RLjdn4bYgVTbqwCFPKhIfQQ
AvUtyP2qXVcVGzvc5ns10f0c4fRStf+w/6rM8R5YXqAmLDWWZJg355/DcN1axcUJlXNE8Xa9nDlO
Lqjo6FsDzEhrKkXueYaWHPulFHVyk62ElEa/VIFtQ1dhOrkfw0bVt50Ecf0PQPHctQ3+8YL/4sqg
6DdmREGp1Cdwls/d/4Sq0tfnyMs+GdkeXdqLlscaVfNGp1S1ynVeThLah+6ypntaXZoO7WFqvBmO
KHWo4+V59JU8PPTXW4gpXis9iadOsqBcjGDuwjGt/rb2Cu7hpoHKg3MS1GzFsrRzSv+HRWzFxXmI
heQGLy781hkcw+KjTf/Nbp5fVHRNV9wXGaWpeIedzWxjPE2Tb7iB3LXktrEzJA4tZ8bnkz1GCiAe
isCGhCN/6TqVQBiAQ52lHrp/8A26YUq6Raoz1OlaOWe0Zre811X/aTwZAa2QWLmvHuafNdIpbyA0
L4BeC0T7fPjiabmHHSc9a+cMf4wEt54ksr41b3EMzaRIq5D71eCgCUOC3lQK8EM5R+P9rDTFC4sP
jewe8F7ujpHChsDLJbtvjyJo+7rkvCiEfcK8iMoubsvu60yY3pzA0aKjeRYGbrgZ3b0idUCo89H+
vz3hmfHK4IPFuo7ROo1dbiAQSyG38su6+RYaNrxF0MAweEVfAKrtzIpkjLatYSFoa+Dq1W4b7Gne
C4tLICHwRBxL4OC09IYegA68glipFplaGoFNihQWJ22DXfu08X3Bey1w/KvqToSdkOjwDivwye2N
YtaHjMnyTBNRObLwXANWLn5o80vd4jr0LuorNehgtUNp3NreFe1enDmHZ6skgWGnI4ksKXribplB
Sauv1cvUE31QRyhNjYrDLmpId0tdvb0Wrylik52ZyJfk0dFaGbdbZBBsrbwnQleapJ46Z8QWCAAf
ZHFpUZfpx8YdNe5WnqN7Qmzu3mXmbEvH25+wkp9KiIZ2CAVwDyqRCpHonLOPXLZZ240ZWHrKa/lA
EI3bfrdTk+QJhmKwQ+2jIRGHUCOrZEZm7LxVfo4HbDDYxO7EqpyyK86RYviiVDQ0LDiJB9X8zw1Z
tRxUOpETx/k73GHxulN5cP33aj6XCld4XeZ66XbvaJSUYfTZ9mggbRBBXPv/3k/labx2uXnEfPdS
JVOrda31qrnP/RhwmADxR2EnZHYt0bnbeW3ZPxvjo8caYZ2iZQcLRrPuPtKK+nG20CSPOoW9CFBU
04NZGMC8VZvNRAb202N4avtvoQASyF4ITeIgVetM+ugq2UHa5AWHUOMInPXxONokvIMXUtZ9bBTo
Ok9xxeuFvVUXovbPzjrddWL5FLGbNHh8+dCQDHR7iUEJs+9wLZ9Wy6YasNEwbyCMAaL8iVsBZtsA
jumKmQHlUyognDSbBQV60ZO/8BK392OC0nyNACj0P3tpsqV5eFVkhvHOA+oaZEdJ9PLgxmC7+Tua
GL6UiZ0YV7QG6h89uuW9CahPnfBIvBSR+ijP8G/iEUP5ci9g0G1zqEL/5IvZFDsCMJgB8SgEUXm/
ZRvphHRlFi12fTSXOoMaY1RabqRdVSKMEoNeYekUYSBrAgaBx/4bucBPmyBG/5T0pZM+q0agTCwE
E/+CTeepnzq9osTnMx9d5WLMSEAlbOikf/hldhTwi5zkwAKctNTQAi2UCCLzNnlgTTovdjUFFSUx
ME/TOK1P2++mENntZHqWNlmUm4Nda8w6aJfSLW+SV/PNPUAHVsTgVfVXmbu0fxL/f8EGFPoqGuL7
dXcnUDFvqtvZRO103FLuMJJk2f29Hv6JeTnuDQ9irGsa9enVCmzyj+ItlclNLYzEmuHpaYU6Z2YB
52tNwA1KmE1yQwQoMvNhqegbttv1X1hn6zQDtft+uYI+kKw6ArbUjMbLJTi7hoMQww6a+A+ebnnB
BybHNTxTkq/YHihZ9KdHeNFSJN8BXyDetaJCtJMdxm+gmSzxO+DTYljQY/mtu/bBKd6iHFsg0h0/
YmFA1/l9hs9EhDoIocOZPk9U76TyoiQoSEYEwxax09d1SseALNcUd5Q87xhUVswaq6UGwZheMTwS
ke6cOZ7Z235/620rkR5Me3lwcMZz1KPNvFvT7G097501rGfY3L3PHKWnymiWjYFcrft3cz9yf48D
71FVmMg8EFuMr0FW430yboAgx9JG/YVdk9t5qcnBQSl7XgjYxZSs85w8+1ysz66U5ZmaQXY3STRs
f5iui3zKVWT+/5abO2hyPEiF7scvCAegie+x/DtJR0M+F4H+4bCDX8NkgEpDuuG/1nIe9HglM80I
JOJTfmBeaVUiiRx3FbF6PPyALjiA6/7GuryY2w7JatBaAN3NJUm8MTtEMwTEBYcbUo3KdVnM1Xyy
lN+5aICXFRAMKZWy5OP1PBZnx5hnO9/GVdPAOahASJQ3Vim9wGEIlJ+ZJ8VXyFpQASu7riMlcR+q
utlbvsSALQ8hwI1+JZ352BBFlbcx7KEjB9SMHmKo0dYYlGYnkyAs3ToKmWwpmsqmV4Omb0ekF0lX
cpTWPiQhOfv2ypgmKU2r77j6bPcj9NQgr/RPabrKmFOHeDPKWkDoiMI4g1oNmGeIPQqE16QAHtMb
MFO8UA0p1SZPDmo3NoQb4iQJClyRrPE4H4k1y1CKFpn5lfAfJ+Ubpsk5lvL9LdT2dsvLyTRKhRV/
QbAoav9CvN862stjIwxq63lBuZOtzps9my//RU1qpsMVUm/mGStK+NOa1zvsn5HuYFkQ+2KOas1F
R5U37VAUg8chkkFtVPtORJnnYD55vJTXhT2x41ALMYL0mAg6Iw5F57zpwPi3H+LOYzZb4lVy2t4P
+IkEAUnynRjqLQxnlIDKb4nxl3TGoSUmBB1HtGgeTSIzJ6/nHDyBazS/oLOgW7ShUJLnD0dFjZlZ
K9n86+r2mrOhFEyRDcNLmDQk0QbHuyg0DSPhPJeu0jxyIPvt5vtNDx8HwK8TJ+T/cRWNmJLkxcIQ
0oMrF/b6YDQYiBXdj/FgfZMzRam4fU4E//32CAxlNMsdcF2zBi/e8EQccXqrYSX6D58GIeAbddnU
VJ0iLE0vB9aD9F+hiidZilAAg4Rd042NODBzbGBxJZ1FgvDj2BHcSzNjgjxVAbAEYZuzmWwornsp
jMOvU9WdZWcFwEhk2s98a6E3YXycWMJn+3YviyiLm0S6Ovr2+S0Hw84ahIocmu07CRdcyjRDjztP
/nKqXkf8feWcBhgw+2A22YSdM0GGzOEzvIYvhcmxouZguFBQhbQbyVxYtuX8Po0owjHGrn98UwQA
gUMHA3xBHDUX2yRo/MUPAkb5Ef6Eo+9sJA3aJb25dzsJtFhfqVm0J0qy+jCu4w+UALyl1VoluedS
+mDlFu+o/Qq1By0k1gDuJwU/ReojZr+fJ4C53vXwbmk6ZEDR+3cqdTIy0CWxrFFBOwqs4bg4NI+G
rwPytRvz341UXAMQ8Ow34YfTZK4VgYyOaC/LziJH0q6rgvTeVg+HyX/em8lqvS4qptyYg91mpyYJ
9wXO2LRQo0Eq0gr6r06fz48YsEsSqkBGSMThLpCTDujKzKh/8A6q9yOWQstW7Bi7kbANzOUJrK5I
4In7iu70QNzU7gM9FHRtyTLY9Z0VirlBxzDWAgxWOgM+Hk+5qef9gr6H0IraWLk3PluLLAqgXJdN
EKZuP7M5Cp0aYewM1Z2ed9Fy68ffaHregMqUAG/PQmfxMzItGv4mVAMNaCOemFQEBZQRM2CyE96Y
odk/FB0pg6JTx+LINZ9AdR2cFSPWXJ7Mi8MLBTGOqXfykVQnQLsRyW9L7BHw+cCAasxMADJDmTFe
zfNCYQ+d4uG2AcEs4NbAf9eI0sQmzCUb3IC4/R4apfWk5Ofz2AUJ4zi6MbuDQ6VHntpDRLy31qiA
z/vFUN4ku1QVaQCmMGO2A7SbdjtH/ueWqcmCS27G6aOF2ZpgZ+UgIM3m8D9AsvjO/QsdwK/x7a9L
hHYIrlpEWYnIZoD5ngQJAHDcZk2BCS1gX6YGsJfm3IEqEBQW7Rc8PTnmk5RuwktEhcol/fl+Pai7
YEOsjKcmRpB8kOB1nuArkuXOcMu8ZHU84Sphgf8EJYqRwwBBCG28Gp2Xr/4wTb4ZKWHsi4J0DjuF
XycEUSq/KHHlcUx5SEbG/K5JFIfZV8rOy90c4tijNA4dUN3Gcbj0aepYTviCEZivmgVKetaDM1rI
7hvaNzAEqLfhJM6zJXpd76GSSnBwuID6ikOrhurtK3GKeyT1Z4vh75QF/p1XMMcQwN0F1ueZz5As
fp2dxli8rE+D2qNqvB8umCkSd6LU5ig8pw/l2YMoIoJhBsot53QsRVdYmc8HvMmRI/X1B882aJs0
v9VRCGN3urw/9qqDtCCBH3A8E44ia2YOr4QzHOUoM7YI7tzgbQGHkXHOtn4DRIsEVWbnDOw3pdPg
r37OKiDPi9OmWkDCRoZoGK6zxQ0myJPIBJ0cO0I3P5/vZYofX8b5DW8a3pWnmdK5EI/VzJWHG3Wz
F5FbcNUYRrpQFP2UhbBtbNbJJYklj8w7Ku3CxqqdQz6A4obzCPzFzXcnEACTdBJ7/8GiWQI1/2kd
AwncWqHMJ/mq12uGJXp0w0Ht9j2JHF64wxzl6u0kZeKh796FCXM/PregqpAx9/ldMalnYOfbXAl4
Nw5PWBEVYe1wi/2u4ULdriPlJBvWq3kUum+dtJlambxSp2wwTU2bHY+vTebgyc5LhP5uf7jPq6KA
yEiwfbVFqoE8JnQF1NFsVesYDOGk9X2bf0mB4CI1AXcksWJjxLPH8ZHc1a5glr7ahAGB5d3sYqUz
O8ZNPT0a5V0zOzVS7Uxg9bSVMQDOEgRP78UX5xDSPOjmQSwgy4UQ1AaYqbAkSE3aOvjKc2xXNJLB
nodBoR5pohxHvQ4iBWtD5bdy/y2tUvx7sZErMDWxZPIOMWxo/gEn+JyLCkOzwZAlgdwQpm3/rpC0
lYDH+o3K9rwgi/2q8fHRg4LVbDGoKQMdrw/kL1eIcBUtlS4EjKXH9U1kWKhA08EApqqWmzCamb8g
+NvrFJQ77N+IQGOCygCu7nvmVBSOC6flsCVuOtID7Kdi8zbeCUIHQFVbVfK9NJaIbSDXv/JOV+H/
3s6VI9Iqi3b65coKl46Mcdziir5Czja+qBnESNCKpN1AjNpmICE4qm6K6ZDdCc6GFOqj7jxRcwV6
zgKAJ1T/HYc2Sc0YQ4A709ZAzJHgrePcY38EGeD0vEoBoe4/yoT2WaTOMH0uRy6gJE42LfS9vD/3
ZcTzRfL+BAy/dgGH4ZigOti32y2TT6x+7oo7GLIs9g4ev8zZbshUApiDNFYEmQ830UDNcGpRvUmz
i6Y8zfrRuBTfBgxjtwm29raCdMMHtfX2i3b8hSdvIlzTAZycpTTO7iOD3wuzHO1rHdS4c+YAyl8b
3isTMiyYJ+eqy45PcPGSzXrus18cQzyToF9lurXhaSBJYzvLT9p7CnN1QsWiNY73tKUNJ/rh/+Wa
I7FnVWVtGGJqCLmq80EEPDy6uUDEF8YqxaWHBQQHuUPZWLWn5G1iyn3BaUq7rynTpXf8g8rrUmQE
p330TwxSVKjnPp9CKUFf/eSDUK0s1dWUaMuHg0diflwE5gWla5v+gX7xum5LmVMqCi6n/+DQIvLG
F+r+5s2a8UXo4PRfcQO0fp34FJzmzLQe1kJkgYeidfJRu8XtBiI8yk+MesL23R1jHHi/MThcVlvN
tPl0n+ZzuO5YTPfOo8fwfsecnNfQnutL/FIe+mqT8z9IKV+Ph2QMZh8wfM+3SS4seiRyL2odpngv
nWzdr/50ha/ctV+hpcnYEc67PzLyjTEVUXWV9hXxNUJLcKR8cBYF9N6tt5XQ8wTWu3qdXbCSaYV1
isdupsYYn0XtFkHo0WTqE4WjWds6FCpdDmFzpXF4CeXEDr3J8GkTQ6SQaxuHSNAmfo6SFoOt/+r0
XVwVLGYFqG6a2TD4j/Zr/a5/wV0OBfdvnjPfVzuB2tdchq0CN03n59V5oXK5knaA+sdJp02Y2okN
s7ugRVlK+yEhRZCZTHxCC0tSfGHvQglFmdL+Cd7j6pS26dZen8Y2vANYT7P7pLN8WXs1ezyipKop
OXV7xa3pBS+rY+1TnXTfCD+1SRPrTCfiFBBMKSjvuh+fC3ScKGtWlIKrr8eEFuXK7LgSBynX8I1s
0nfTua9izpQuPOSvuNkUCKwsNNDr/PRNsAMGkRV51V60n8C1nOOHMAwJK6kaZwNgEAoFUl7Rk81n
h5v0QQmFODVe+DKACZ3HXHlpIG/KLBoC1snkAeskXUd8YbTr8LYbEXnO7uRkOEFk+KMPIEw7nMI5
wOjcK4OEFU51dCtokc5CUVLKTzm2ba7H2wY+4jcSDq1Gm0c+H+C58lpRcPj7TF7qd5xTIPRhEJI8
XmULlAUQLpEg9/5xlcCdAPkrF/sZOpt9yCUUQFdjrpIqgNz4hGO8kcm4/Hv4yodEPHLwS+1t81ma
DfXHet1JtAbgc1qS7psG9kslYKMayWIUigsPkUyr2gCoYfwXLX+9eeesKW7gT5761A0OwuW9uJZ+
WlYXsiPAPRQiAko0S7I/91WLtWPXWPlQRNGUmBhYM9F3hVI0L0gdIFxHr7RrNY4oahl4OLl9TNwg
vphQ8BOygIVyn6OFoIy7RUdpjhiDRzHhmOWhDM/VhJdJOvkWJqcUOQK70mdfWrXVeBhFdgf34D1Z
TmIBQv7FHkRbtEvnW7SflRNhQ31t4zWm0+FKSXP9zgzdHm6i+Rw/1nR8aqgMNC5IK1uUwlpl1TrU
P/HQ+Q4Z6A40N9ECTDFO3oNRvoto/rlg8CZfz9tFnVUJR56cGoy2PZn02yHMP2I2cn0UBIndQIWf
mw72rzCEiZKfbb6z2ZhnanghnxCLCyPGLuDiZ8Xje+j84P9VNgN3fKeXW5AuynhF/L3CqJK8I3UA
mPaW7x2JEIhmAFf63g2HF1ptB2eCaiH7SOXmQsIOVIROJqP3qVbeT45ana5+pU1V7H4omyeLGM93
RkSr1nhEgyt7dZC+iMlYLjRn1D50FiR+/YaSjvMogJmrooh8gx6bhIYljJvhFd45TiqFzepIwSh+
rSCU7VGOH+B9ryAeVnjCiMv/1eXLBfdD9/UZLc7eeOWKWhMt1R35EhtoPL+aiv6fO5R6rj+bEXWJ
I6b55J6XU59QwfWFUw/UX8ER5uUtZxoB1ilH8zBvA4URKm7WsFQE3fiV850K5WEiQvqhm9May43g
Mk8NtORT+08Rdw/9SbXayJG+j4XCcBCzV0Gav7fk9WqFR2p8CUbeI7SqjBaUt4oW4ax8ywmTo2Z7
Km2JlbTAGOgoffnNg7+Lp3B5UbnGfC9pubkeVBmGUEmLx6umxn9M8H3XtBfxp8gZQUAlCeBUMXM1
2w6i9j/48awL5E/xr0T/PjLN1o5s22NRKxYOpGzvtj4Qj9zwOPLfBehAoO9ujvik2KnvPqaDOaB9
zt5jmHAmito/jANsGctfuMas8fXw9e+zl13qWmQ3yS0/uH9s+hp1tITIgU2FD+OoegRo34DkDmSm
gqZXTaUuc+58tu8AxQ70lO9Usbc4odnh+GlgiOjbO9psR0RX/psBOsIdt4FsDKnJKPk9BqDu0yyR
r0rEB4LTuCeNAecoe+1UNe3/7EFaTaSttuU1t0WxGsUnyKYK3PYqGPzfIprEzE8rIMWNygIVKtrj
V50QEHP798y0NXW3sVS0qt/940YtOptnmRcyYPOvbPxr1VfXTFRl26MkyIXNsBAQWoOskDxk3Fud
fWQElVWEqvhBzrHhKmhloC1ldTbw3iIFXnAxkq9SbWUGhX4v4c+YBfOXZHTxscjD24kT6Es5wWdr
vKEFd+kg8V7MfpcL704zKGPfpar3PZ6kE8KSKaj82QM3v8WS4grqcOv/VG4CHTkfChdP8i6JjVo5
dcotAXbCZTWAl6uk0WFJ3q69qKCF4fyy80C3YmGqx8XkJUEtkdYF+k2ZBjW5EIidOEuePKZxkQv6
ElRQwc2I+PC4bXBXGKXpCodDiMSYHr+iyLSotYgdhAyYeWhCb2WqzhlJstG5PkTsVk4vsshKdIBq
ylWAv/udY3A4M8GGqSuvUcPPZNftpc1ILs/bJ53kqJKnncMS2IlvuZupQEPlQIyAkT1T76tTkHBX
wn/iNUgY63vapVv+HiiTqTOQwd+jZYW+QCravQywYVg97WJzg2eV/iw1/q5GU6Kmgg2wLtvGGDmp
9ZxcpK3sZC0zNXYTTcLo309PTcqGYN3qdZG7eaR8CGWxl5PhZMglhuJG3hcVYu6AH1l+ABfoHXSs
XABNc/q0unYRasArJqv9yiLDqTZrYuy+sYNLxjOIUKbuJ9WLXGl+kE3l9OGYLXn3omTmDv9g+G8H
Pq9/XGtT8c9k/S5kMiN9fQBAg9AFWDS4/uLqjHUpkG8pl+erMOwzwYBZs/kTnUikMhBOgM5LOpgC
k7eUfj3f7XGW4URr3ab45A7SiKPuRNdrmF6w1V/wbhOnAv2IHtdHrubc24NQKuW85Sb/8N7MuyPW
/ZH5NDSH8gpF8S5HbBdEPBYe8Mit/aXrzNzPAlsVcGP8YlwOG4WKhCVnJg4a5JBMmySaaXEJ0zZ1
kS0aAtLevQtIhorIf6dcAAJ30b234Mv6QE21Ej4oluibSlHJDPBQa3iFDli5VFXol5QUQ2ruwY7S
27U+x0v1mRc37FgkwKCzm0D3YEjjHdjrJ8yHpKooKn1/1WioVamr33iSGk6ERipXymvx6emsf5dX
FwzwjVbNLk3q27Xu9B1cPfS6jqKLVcZgkXWxc7hZwXaBMosJzb2DpXldKDt6UMfBg5xJHkafA/+f
0bJf0VUXHXXcBGC/9Bw1Gq3sw9ljI0W1atlI5NXnG3RVgKxK8zHdxSu2kyt2iMgs2P8DIQs/XLXa
ekCEHsvt4YI+8wGTRcDMMFtbAHSN9UEAqrZDDxoZYqKvlpSWYJPAP6/TzZtgoq5Wm8Dj1Wl2V5xB
og87JMKb6IZs5/YB2K8YWnT5E6fA3/otVGqJ0S+2s3OJBQ00UTaQyajusgkot/RpD3vzlBKU2Gye
9OVs51NznhdVA+mTa12YjHwFCVPe8jmLg0y3f8vokBKEJEmXniDnP7zva9KhBErPt0s/WXQpc7jD
7aUp/uAdzqurNJ63Abb79b9MMS2vpOPYN1zNNfAIBEHCcpjg41mwN7EZsIrR2Minu7jltZyliA00
uApSrbrvyXVvbkJBFYYNkCyrNWQs9NkZJtAQyUpG6DdhPJ6z0XE1xqSYpEcXgmw5KuoQ3WgA0jdv
Q/1m1644NczqfxkVhYyLKvleDoJ30y+hIOlvzEC6hwT/VOTgw+KM7CeOJGETTIYgsUDpArZvg0s9
UsV0K80MXABiTPmIOOPH52M3Fnqn7iPV7Yk5b94NDzjwOpO9hZ+t8lbzIJnjIZ1DbIlrnHmFnPZ9
UuyCFVrH95C0bBJxHCRgoRgqN5UdDp248y2lrJPb0rrKQ6/7CO2FUZQdz5A87x1PAchGsANQc37j
JgLIIbYgT+Lnr3h+hiVcZ021bpPZROQppK2PU0jTDTkgESHLk0lh0Vq5z+XzHg66yhld+fddwvmF
OPwj406vkeye3+tnk8eA8gfLvbQGQvnxwyC0xEzRUqkucJ1kIGAPt0aj5C7vvShwz9AZIJErD/L6
ChgZjCLQck9eBVIua+EkiGfMgBLBbzVCFFMWWECb+csogn1H61w9VOWicqGHoU0N4wELyej4Po8A
C82hHQmfS31CeRwWeKng1gVrQ6QyOnc8oLwjBu3VUtJ62mTULLvI/oonufRlQgrwPGrzLZ/u87sN
s2in12UF/POylp+v+0bYOIz4SZSupNXO4YN7+fmykwqY+vsdv8NNrbybVwZxMpFqWxqD0wJ1x9MU
OKf6JGtiGVNpW4ban1aFxq39PxbMqisq+gD1z+oQz/AC6K1Aq2Db5x2uW2MhPCCc2aSu3WFzVwO+
D3nv7Tk3sEnb9Aso6uR+bWJog1Pm0uvVIk8dvg4LD6M83nN8RXtfPRPyFW4ESpejKLQiGI9lVl0b
2CIRnXSGLTcf/VtbTiIgMvYPz5zJu/fSXbDtixQ101xpGi6VJFKUrOzb3vM3chAlXQoygurSiXCE
bDjqa+KBmZKclOjeYozWx6bVl8+nj6W4pDPiVraL1tveelkpIFPW4K7Jf0+qkW+yNlCvRH2Rd77j
93aRv9yd6zgTh+QTEqTo1jS/LP5D3QPgRi1GRz+7ig548/jqC6cCgR5P24YooQDwXoMRra/wser5
sAf998RyxFQ6bDkIaRxu8RjIkHyQnYog4zItTYoC44Dy+vbMYMOBiTb5LqfvAU383mPCaqr41gI+
90iFfi3pG3k5wsHxKPELRYrs1Jaz78n+4GMEstHotg/2Gwx4UqH8Wi0+HXxmeLd9KejwptA6BAZg
VM76vq3r7MssP/pHOTf5yHowWdt/HqtjCoovDM/I+uNPh/TH0wlC6+dJ1Bc5suy1eemhtpKCZjbC
2O8daUpGBYh/PnPVX+pfBcbzVS27s3I8PZXAkLgdDoW4FOKDzVoJn5/MTfEDzIV6dlufSKDoIY1q
W4wuAYK2Cifr+aB4RvCVMG0hOW1oKyrbkz7CBpC9RJLKvO78plP9ebo8RyGsRknTAr+CyUfr5J44
bfdKVoRfnNCWxlLlq2MV5MqkkJyaXH0o10QKtm4pNfugX4mus4XIJzk0PpedkiXQ39wS05XhJBQ9
uk3ENUpHe6y5CyXdOGPvNCP1L4isABrKPlha+C1NE5mg+ZBQTyQcEKAvYDpe6B4+HskLW4DeEyxi
qjy+hCYMY9cl0yyJrEOsgvbZ6aLHdJhTO8Uu2SMQUB7D8AF9qxxsIe5dnLkL25rRPAPlrOUb1Ud4
Z0+u4rLJIhDvjOP96cWguBG/vLlIJWa8WvkL0YJKvH05HdObflWEkerwTcle5VwG1fUIF4GRFb5a
34bywiryZ0zogphWAmM3aekru1Pyc822XaJ4ey2dkadSUSVX21GEci68ped3OjiBsAe/KYJtavxq
mOePUlQeclN0JmdCocvrHAmn+SRVuVfrdGDBGcWqK2rsijzwr0uByulsk56wIcaYfsI/H3hZejJ5
a9Yj/9yFQYxAE09ZXMM4jKkaD5bZWRCrkOTl+D2SlqyyYK9i2QX6yi13iB7KKUkwvzOetxVfMKta
MdpWmVW4Pvn++mkl2XiESJAqWPPMTBKE8H3b/e392gg5zcAgiv+00xe1+4YCcNrYL/yqAO+aV16r
og0cmzMQS0S/z7nTGnvPJxz3M2wIoWQ9hMDl2EwlCJ/Rsk2muj4AvhS9iNsOM4RoEvfTRbZBVSaJ
wkwLPBrEHUmEjm4IwtwGwicZhHzcyWUqOGmp5mbWZUitiCLJfEhnwhe992RFQR7iLT/yiWaGI+N3
eBfVqpxsUGzHqn1wRml7raPv89Y7JXPjRLzf/BHeY/xpxdd475Y/clOOL3em3IccPGPcyJ3o2Ejf
BsX3k+93M9TwvwOYfjePCaJbs5xmyf2RUU/bL2qQbcHcj5gktXLBN5aubMdkHQhce6GO5liCeQoF
umwolsKCi4l19MB88VsUdmnUGrWIQYT9r5M+mCgISILmbVvio0kN4Ff8vNU1OE9oIdH6swd/XdHH
NUsPpxetnW8XfEloTdSx1NWtjcMCrmsdq6+yme2X+yTn3Mx1vmgFqLE2qrO5B8BDx4IJVCipiZOi
nn6BwpmEunZnUKFjD83QAWNtVUYfTTEonmwLGDg+hOoj8lV6s6wswpl8x6c1wJUk8ue3fZ3p7m99
yJVxU/O9iow8UkBc92eSep9uA2OSnpi+PMXnKM38E9y9vjyrHDcMIxXudMqVpv4r/nehIJlJcYyX
oKylnTk3JzllShS3wxY6PRpiy9akMYyb4SEEHEg2mFZcPJdvgq9iXvGcjRDX+ipU3CcTASVU0LDI
HfDNCvbr9VBuuW5U0ePfNDh5HQlyPDKfmnIXgilG70YD64XrYi7nmtaV1kplr+2eMMxuKMEXPXQN
FUFiD3sB3od8g1MrlczOlRmyOYFvdPFkcTWKEIRftpaMbCHzdeGGMouwjEbBSYWk/IXuobBRKkAG
LlNOXj39tHS/GJ6Tgv5BgnG7vm5s9jsQtOcVcxlg1HpgN//o+XEV1tcTuDTY4Q4iRdB0Nx+IZOEu
E+WClUWCkDvMi5j6AIMDqKSlCQHSLcZe0+TKI5jVMPRsH+hLlOTbTiYf+T21bOXXIb1GGagROtCB
CHmh5dCTJ+ye0Y+qTOFnHDyPzOVMxIrBwnd+q6yb+ZGCs6mGy+jHwsX1TfNY204EfZD9Gap7C1Sw
ZSZgIH1rj1rxvkVCrQVJDwpKq1jedXF7J5rDl6SWVsqVwwilrg9XOyOVe9EOpMBdj1tjc6nLF8dO
Lcls/NusmyKfdikht2Iq6PO6iMnj4gWRgNcRj08SksU5exS7I7eBVTc5MH8y8EIqxrA7GjEsDRe7
E6R9cObHYSNCVRVBjO9qvsxjaEtVcbBTxLN3/+1HWIum2actgEUxaEHxq5ZCdfhTvqSN/mrUFk1t
Y5auBCgrCH9lSM7TShyHbTJBK9bWNZ6ch0GaLX4QyLgo/LEHcId+6oqCetduAEDebj/lanmwSPvN
wgil0a0ifjEKxbFIhg/IdOi/GoEVlqukg3s/fOwTzuyQKhb9L0cQ32yt7QLMB9vGg5+XxC+Ztg2/
DnrDWzx64DwhZEmrBTfLGXkthwmvvaZgoSMlhrKEE5mZLN/t2QE0Uo04i2CEriKEgfohLYE61urD
lUjAysNWTtA4/a9muEyeQibGYaE1IZ6YDnTuSsnmPxIdaqKmRygGXPvdsuddQyuBwGALnGwzbJJr
jWh2XTM5Es4DQsNpN0UwqfO4Cs+fgRrKopONvNlnlsMqnxqOztD8+1LF19QTxo72pdz6GauSKEpI
3AmkryZPkkzG/bY7tHZFWZY/wx3i/GFyjiWZgrL2oN7q90cfd5DP5TY0pSL2cq9Opm34F92PJ39Z
nVBY9jAfLq0ixAakZ/RO28wGrfygxD/1Lgzb+tUT8UPQXNI3P6kDjDyGqruTNOIGQDJ4ZOdr8YM9
ibw54j7xryWD4xUnkdUAme3cZEKyIIPX7TmkhPIUnVixn1skS7UT3oNyppoDa+x0rIBxBGhRjZrm
vG/qgjcQy6KqQM0z6Ca3Lhjk9ZDaIHUp90O8afIsSDmKyfzwGWrQhUfHMou1DyMTtVBr382YNhIE
Mop9pM2kjhtcQyuTkCCAWCdmkpXIMAn+qz+YneYH7nMyuFCdgO4HOLF7jRYa/+ZSbl+KLsEuVTZ8
gQeOG1zlG3pEZkUKSOzvc2OqMBNxXFA1IQPb2EnOHLifbKHnPZWSng4Giw4/2kTSL5fZoKLlDivL
/YoesSXmDljq+0gRSeRXjW3aa2A+GiW+o/SMjqgl4Xs7qL2AdCQZ0zLbzceq7cn8LxoggdFR4tAu
Dp8/S+z8Bw4b7rz8tWtKSVNRJ2liIvD0ddk6mUFf1D+0Y4EvhIKSBnUR5U3zRjXqGCBmh20x3VhW
MXrv/dbbg2gUsFKKBJoMaiLij6Y1oeynkVCiw3IBOGaoYnTjs25HGi+24ZpHMe6EGR9dz/r/Fi7o
MeC8d4GYm5ahqnOQvsSDB/rxwLwi5hVk49ME7SBUU+9FSkUGxXcH8v5RG5ehaUIDg/hsObN7fc1v
Fo4Tuk5qhrRQQRcnbQIUXTA7ghzTCsUBTTFtxeZkwDIGTDaiO7us2lPbvYoY6qHV3qh0g7sSVZF8
4IGr/3sxB6B2bdAIn2wb052NLN0UVbNtPrPxv0TLGEnJsLBmvCgKUFOOl5+Ct1JOv6c5bA9bTNwL
PeCoTjGzNbz2p99d8b37cn43P83Fnn15+7f1s+BVp8MezAiQzn0M9IiQU8Yqlj5JqkhjilkAhLBR
GPIZZH7l1RogshwuEQmPspaAV9IJeVhSbipWA4VMpA+0FTyy5GhkSXlvhcaQBMsbSglCMjVFevfJ
HdSRaApGJnwAOV7yYkhlvVCLYW9DsK5bO7ZxZZjXX8U4MD2s60R8H0bReKtL9ltyojOk3BPxNKVb
o3P/cph0wQ9OftfkLr1BAkWnIBI51tjTaFVWMoIw+uN9n/WJrnoodvC2LDq3oa3VCCGYw2Nb4k6Z
YwmRDNPUD/6qRjAC08rEyzyBSWZJyHTV8whBn1T3r/hO09yTwJdEih81rjHb5IlFYyNOrFXsxR2o
+w+ujvlJrJP4RlIRBOFZ5oZPiFCna+5yeGdK8W9g0c23eB0jim8NsekS5mDaABGinB9BeyHkJl3r
5uNttYwyqt2+9cB1idDggnxyiA+iRKrIIYONkFDnzhqOMlJdvNQOtw1/iQjpNPyjdasDqrCTRxFE
K/Ox6JaXxwH1amWNtSMZfhUMUUjiIg+yB1WYseQxZrtSWgu0aCjrmM4JTiGvkTr0dEoxKUtySnSm
GGQokK/cvxXsj2gcjZ2ECWWczUog8uULLJld/XW22s2Qv3jlDGQq4qhOGNhgr4Wt/GHECcdzfJ1I
3UyE1nxcvo5MtOIT4aPm9xn3S5VOfVlZV1dXWcX99EIh/MhR4DGMahmzcNYC2blE39FCRTe2X19D
2IYIcnm0+vdGepG5wWY/XJFu0SLRJGpLlS1IOMv/PXwpH645hCmNa56N+N+L6P7c6Bqnv/pJap2r
Q3XszzgKyEUHpYx1gUoLko8fkY3PWQB4c7JsTY/et+ZZ4lntr11Uwif2yvV0wgCS1PviwHW974NE
F7g3EfZPxycXp6cwZHe+Lhe5hwHrBMf+NVJhs/RlfNmU4aCX1jL91xFrMKbJY0k5Tv9rAkJPMjsM
izArvbLc2rwZs32Esvnt+r4Ng7ibpneKSC9RKaNYfbgovLK/+R/cELgHKheOZe8+cSWlQvlLRAtZ
TqbgQAZKnT0e40I2HA9NPx9T9pX4tkAROtgUsejmEfv6H0oZTfJ1N85Cd/GitvqKRLd+jVGYysWo
/zb/Lwdk6wjAhG3n/+84Vi1meQKyVBEvZG0zUeuEC5v7qYK/bEjOhX5INt4zbGBlnLqxqBcEuIUs
bqp+1QMKnxoEXE9yrsXltbaqBTpLJEYiOqeuPW/MLNYqpnXn1c+2MishCN25EgJn6hU+CG8guOMH
dN6i6jOEnjsRHnNKfSA6NtQLmeJyA0GBHYHRgrF2f4pucPKAEfDvINFfR3SAcqySHdsSQ01yBkXU
JQbNROn6WfECDUSZmVPHYIyiodrStfsBaXgewWE6RO23DsHYQ9QN8433l9y0LFW1u8BuCyMGAwho
fc9VZij8CyDmvEZNOnRTzFVhB5QvbVwKvO7oTr8zL9GnqY6MYJM3lUHEIfA87VlY9G8g9gsfHM1i
xw1zeIunKXoTgimhjD6bQiedITmhRH+STMDIx1gbpo/XMme6kguCwzng3M/Vq68+LLdnmiIgnn1r
s8+mglROpx3K08mS8iysv8Q7ZtemYtfcGZhw8ncpQkzCAEshpzvdrGN5OyztGifjqqMgxW72YCHA
+rim2LP/hbwlFLXfNOU43MNQtrpJV5LxyieTcF0RrGy9qegnWXviR23w6B2YDxy9AknVIY0PKReB
7LlCH6Tdyt59X7MO5hC1PZu7mYNtfpH0X79NE6wbeivwaLUnzN9v393Own8dPnXrZ0vDQ2Cuz98e
Kum4gDS5nGZOeRMiz0H4QEaHzOtuFsq8sEb89dzAty8AfO5jInDwm4/Ondx9VPZu8/OPKqQQTohw
56tpfgZ35PvuNrBOlkC5HrdjX6KPK1byAeBdbRW+jC7YBCrRrNKSQrlcIMUztdJlW44ZJtU5q9ah
BH1lcipdOE5audcUqHwbjTrxOM4vLHH+0KH1h23ZGgESZ64ChAfhnKyRk99XOlfSLFsXk/J8fx6H
B7i4b+05DNi7CUSsIu1ug9KGhYZ6JeHhY+0lCk9r2NwrnqDhzh3PlcQhwPuSN3N9aaVdubeZ6vwn
liPpEC9Hr9OTTJ+RvgUczWSTUgHmDYGdXocwwzhh/wSmvFmsdNDwPBjQ8TtySN5zfZ8ke/HuV/gA
H+Vz4N15QkJh9gTuq2uK0Au34B0FU/4fvrZKRWwpHyoav3QL02LS+/8E+ZQ822YzXCjcHMY3ofQg
yB1l5s/lJ7MWvX+iUO329P16ipRHFk6bFKQ/YkA6sj5ayT7Oy0uBl5gmU30F4+R99Ob+toc9dWAs
GuuuIfEK1Q6R1z9+j/I7Iu0/xzSa0xm64p85lpbQkEpAw6NKUnZ9ss9qPahZMMj8vBj7wSym2Xh5
SE2sFrn/Ngr0cuu/GyRNb5ZOXzStb0Ok06QFFVhnS/3pxATJhqfs+FcGFis5C4asopq8Mf0vnfmq
lVXJqPXnKNFM4aMWGBqnsbwb4j4Acwl7dp69HtWbAYxr7ubIPzdDtERZv8lpWyCUyfpo/ghz7Ywg
LiLaMDKt3Kw9gL+N41b6okGfjEdQ8LNJdgwyOtlotzBcINh+UmrXio4QdCMfanjUv1TsdZZmFjTX
r0+yzlDD82RVcvnaBvoJyHRn4nwpza819X0GZYxphBiMALSvvW06X5bRZ4fO0ki+ND4rZqZdujLk
PnUPPxtaM7RjDCQOqalxw7XE76a+5Gt2QQyzpzembxluaIIJKKY5vIQcK9MVKK9rxe/xmJ/PQ6F2
hG9ZAepbHMe9lov1pnQFvCPWokzMhhq8bhiPerJKxEh7pLCEyaWhZNTKNwhhNUC3myOskUYA0Tq1
0X5/4CBUNP48IiOfyHoBnHV+ziAC/AgHYLYrJAWKAu76cCz/dpe2YLP8WeOd1aIIRLxHgyDiu6pE
/5Da8PgqG+yeK2KD+/O9YEntKpwzX7czxde+GAT2tCyRCALMd4KhicbXUVXWQw+OHzVsYTQKMoZ/
2NoGX45wFqzfSnCK/jZBpoJoEvv74SEi6Vdm/mr6KUohsV88F13J4MEUzl7EpPlN8vQrVteAoXcz
aK6Gnq7x4HF24+FFaEquIgBWJbIXtYLMdQVZ2FvLnHR8nm2LwmOmoFJZBEzRY83PRUtDzRonR/y9
tTcZ28Xq1JIPiM4aaCbC84TSwwflBxfHbVgVLoPav+ic6WXocYRiaAu8WlkaQ3HWmkjLxu/4p4MF
WtHfeO9LsXPIvhgj0ZoJX6SFvprbz7MOFwHmlXvLxPuA7WXBBtX/SPp5mBVRz+WOT9hSFxCEwata
rNsnFSTX58lwIVvcb8A1cvSv+n//fZzaq3aiZIsQXb+r7Fk0iQl9NSAYUZnDO9l3bPsdWmvm+TJJ
MSlnFUDKXhpae64elZCoAaX55DWvUlIkuDBMAHJNs9nAZy4LWOA/BR+C8DapE81fSFuFn2Jrz5L8
Ibt+SDByVjAKWXhJuCMYXOjQh/C/QdCYe5xpj+1q5aFBkrEr88MGHeVe3y+hYEj5x+sQbKDZuRMt
26jP4pfKbNY/aWy2I7/+bVeeFEA5E9dltqk6E6jHBigjjrkjMxFrWhPhKNdWntxvbbcuMxXPu1A8
9Amzqh9KcF2aDyU21GX+Ozgoe+ei2mGitRxIt883eMsjaMhYF0NB+i1NU7infWGO75DDf8N1/tXY
EtppDJXuAR1FRwQ7v6nsmsxrYdIn3HzG/7o+cjktnO3pXyVtvG/NIvaZq0zlb+W+0QcfetBk3VAV
m+d51A/IzlIlXMvpox+CI4cFDDB6r9uO27nlhnqmJ+ChOlpLx5bbkx8yk1UTGHOfXDZGf/DcO5VG
2EK2ARFs9tWrgxWyB7BTEuzFsqQyW+M+v5G9QTPKGhminSaexwUK/InBQpvCjM7mrtCyqHKsgGIt
E2Le1+9wx2Pe4SbiM1eliXysJNgjvhbRzVr3dxolb5v+dgcRKfIBV+YPJCP0l77Au7KV4FG3vYuh
yxpL2hGHCmoOiCKcfnOYmImAA0brecZsqnxyUXmsazcJ2oMsAhsOrDe04SyucrbfNZJxn51TyWoV
GsSyrg0e9NJn/nBIXmN8JKvEFDa7ezIV5HCPe666RpP0hZvZYFPpZIOmXJBOHnYRIBMV2Cnm54GQ
5e919K+v5P1r6XcTjdpksGoPN5kNJ8lJnqAkuKqieCfuVzh9AfJKxd3w4J1j/4hhD0AcIFAHVz71
dvTgWQzKB+wUBqJp0I5CznZsHqnir7RZhWCr9Ocd/+Y1tQVQV+x0Jxk32MeFzxavR6NxMN7v4aXu
fvgM7BTLyfyGN4BsTe73tBg1OHHFtwm/eHiNT+Z1zGoBj30+K8WZtXBGlMIG1xpnOgK4Q/qJlEOa
AIyNGeyEZjW+J4szQoBvX74dxVPp4Wa9YQ4bw/K2iHMbZyHUK3X2xoObXasXL1fgr1m788XH6374
BHbvc7RXZRQsUT93QIBP5TPsOB/8LcWghdD5bwKey+ISIenLUtsC/dr9mVG423hzIWae5USEiq0i
3/UIqvGYkPIntCrBiZQjiKoeOPShwIOD8cBouf2Q6f5nbX+371VS0Kim/kOADYnkCNj7RHM1Wg+d
jMBFBg0t5rYH92PY7jmIJmUegzWZRPzmLBZ3k9/PKTY7GRm/3lDCPslbpqNoBltiAjCvelofnrBO
TsaepYcbzjEAu6xO6gpKh9i2zb6zY2+6X8aqAtzemV6HwyghIbm7Ch0mBTbazchXBgmYxNSigbxx
vlQgWsTWP99cMFdrCKzID/5DsCiXP2CauLILuButJRUT8bgBowHwVbLG+qH1JqRlTPZAcppqP0xN
yN7gu+RvA5fbfcg6lWEDn5B+qVqEwkFz+hBy2taC0R4fqYLWYabAFCCjXqmy8Py/gm6ZRbYmPTjL
inCuU6UgA40zfYlxSddemK4vCR8mxajRrvyxveyUridRQwtGn7cLRHCmuYIxWvi9p/QA89N21auB
OpeKC7UXgDVQRRi3jjy8aYqH1+jB433FVVAPMfDQlp9KwxBVoq2ZSA9chuvl6b4kaYv24qfzPqdR
W7CJ0hT7WE0kqtksez2ZhK29Mbgmg/6qWMrBUwTMlXioXJ2Eo/jK00b8eWcrm/fYYX/fRW2bD/O8
rrpr2/IbG3AsDEAlHTnWtsaW9ZfbaS5UFFN3uX2BMLoaTFAdSepmID6xMh8kC91t5u5ylwsf2EkC
9AHV96hE34O8spIfWv4Xz1EBirUGNA9lJo80ibiap5Am4lh/AB2PYVuh6c5xDNmwHPBQe/n5jnSy
5jMQwIsljjL962sd6HxGTaQb2gZLBtIb0YJEPp203QivrUPFmJDnv0S1MyogQeNvF9Aqg7hnbbi8
1eebNE0U+sZ+zOAkXIbTXW3kP9js/wfnq+5utcQrRgfPzJ86YyrcUviQh5PJ9u4Wty2QP+goOmIr
nAW3SFfQUPCXIoDBAz7tnntNJQWaGePdkaBDF+pdUDLz1JUyomLnaM1jdIKszzmfnIO/SeN2XbwR
fDJlpk2u3FMDugShYJ1NeGfn5B+Ec3CbaGmvtPG2EEj3Z9fxCB/SCSi2fLvjHZqkF14TIrhAwFjN
e1/vDJlAMvb69qoXr3NEOBo7pdeE920b4BkkcrsNibW6JNfv5l29w1G1g6pxgEPPb+B2OLUYumBH
JqH1OMIlKBcZMNj5Qvgiihlm0PyOC//dkYuHGmyikUle1fWXTkxZ3fs0gvc7E1pb8dO1BkFXMBMT
p1WFLwvEwS9UADuh8Z7obK4GRrXulH5eXlXsoCxbAHj+h+SzG1+mrrzVKTqAE3xYIPbFvqEt5Dp3
rf/c2hQ9blSESIv036iSJQq6Kwiuv1Bu6TXNQbdgZGffezGOWDu8wv/4Ew7kTo06cV9D1kqvx4mP
DBEe1yR5HX8Rb3p2Fz+U0awA4Ywzt99f1nLzKxeeFilJSb/z/2keiY7Vsd8qXN+XxSPtFEaHbk3Y
+NF5YOvEEwcUE2KbbjpekiyFak7sC0Rb+iBTkV3ymMXk8ThptYVJTS1U6/sfvqO9u5ve3v3hz4Vm
xXJOOWppe7sTVzfdYHTLJMl34E/yapc//2y1y/1MQIk7rp94NxbDh4ebt0bCnbZ8oNbuFC1fFohb
WpV7Pw4OQIMe/+AQcbPaWM+UEsXesxuj4lOCfOuqQwHHD8l44fNtCylvsoxFdfqOuX1ElK5vsziC
zWw3tjebBuHL8yXGvuaTE51RiBCUjXpA5hz5egzofgspEUr5kou86XslSABwW4dZoTnlsd2F/eQ7
E6gi9xz+o1hL2srrYLOfWOb8PIcJ9KEMsAHXSueEJPA88zvKbhLFEDwMsv+Y/r650m2LiycS2voy
EEGY21hqrnl/zVkO8TsKGlZAmru9Zo7Aw9CGA49zFUffJY4mdYfe7dyTJWqc36qjqLxW3IiR5iTg
R0XoIpSdi383XM66OFMOzMH3zFU7YLR3F6L1cSygrKCYf0PE8gAu7LfERXyJQ4JBDntghPe3bnRQ
v/6R/mlkJG2VgfaKnMiHrH0pMWSvC8gmRwz3iKyO2FAFipPQygFefC1RQN7QhAdoV9ObdtUIY/ul
XA741QbX45AhebXbuR5WxX1ZPnzVVtN8O0lDZ+BZsmcTpblu/dU0kyOpK9NefZvXcsBIUsiC9PKV
RVVUsmBdl/oetp0BhDSJGW2JWAsc3DMYiz8COP6pKiHLWdqJUdPNVhordso9xy52rA8Ppva+YC4L
R1YCQTC8gzQ7Y3GV2uycHBwCIr+xYDHtk6RAmEBvYYS71vlYp5PQqnRDcJ8V++lRy0slaICZhK5M
vLvvGaXry7CKmppN7jULxMnlve9Ix86CEWhBTbSu5Y2v6fJGFnScChbnuUkjUYw3DeSYhv91AxIv
65Q5wYAVOJXHB8OelQUcg0QNTjOelmv7EK9O461kmBrXPc8xFj+8lWCRyPMIVCyX753mzSqdBIRi
hZHEgH3ibkxOEH+ybGvDvA1q2btuuYPzwfj1NZlYFl3brWTTCAuehBcw9w4OpVkcm8OyDdvCai8W
uyRoAEV+uZDzeKly8w6YlPCpG1SKj0LLH4Pb3ThKZ4fh3RqUaMHvaai4Veun52X1yJ/o/HTGCUip
90iczctSp1BW6ehxB1oQFjdZ9C4TLcHkQiWW1HopFeUSXdyZCB7I08GVcd/pNWXfhvAwDYXQlF4c
KqEwlj0GRWd6f0/24C57WV9+JIRFM/40jjKwuQBGNzbPRAO+0ggJ1cLFnQLPuDBn2ilU3hAeDDp6
IGcJWMRRVkBBiVJc+GC/d868kAyh5xCmffufyKKZWhAS2ui00CSxXlrC2dIg0WgxxTv+dfOejJYV
xDD48F92glmjudtvTAAne/nk3ATsw52/LBt/9KVgBc8bWRLmXzKNTIUQPT76TjcvjpkzfFCyJG6I
OYCXeN8q1Ic7flIDt3HfNxrBmCjyxSDY8ivUmw5qbtT0dac+Lc4l0/T/OoLgr4zwQet34EDKYjHk
K2BP/g9Qi8AwnsLWHAtxK5rACl05NjTPgH0MUvKJLcIy+PZ1anpfdK1h40JyMCiBuvwlCR5jXDC7
fwZ+pucDHwUioesfIpLYKHkkb+qm7tkwtGpQX7DI3V0eUeZZBYMqkd7UrvGX/o9mctvMX6XTrd5v
afgHshHZR5KNZxLQqE8k7PshBqOWj4yby/AeH/sWCkCfL5jMloI5CO71Nhlwy/HaE1aF/HMZiIcz
i2S6TKDcsT3vkB3AFFJxq5c/ZrMTSr2HM4LO8u0VsfCo+sh8HG1Z7HoYKSvUXe2Ym1Eir0gSHfHQ
z25Lq5eJb//C0RR/00nQMd+9fMrip4n90iBDar+P8XET8GBtDkVyVFhsXqbPn3jyW+radRe7sLEK
/lu2KL9V0Rzi+fIfPwMouTlc/UWoiESUO3pjzwXYyS6IQS1PpIhbHkkDhAd9EimPL5h6DQDgLl3m
32Hki0Qm5TjoJ0hOmrMtU3/kE3hNq8cKvRGeLa5DLG2A1w7WddBPBw386qQqu01SP0LJf6DjSlMF
15DHO/3eDzBQUt2ZfgZ470w4zG6LtctGnY3qaHmzhEuEy//yBgyG3Ap2A//GXoLCmsrb6qhjHc/p
nkWT4R6IjfDl9B3UeNzHWDs9/fHjN3AYv59js1clW1ReSbkJ40w+4QvFymNKia9xOpXan7ftW8rt
BXmHyuT8fEAWSQssshjQWgwWoRLdI84Np513F6HGvvRjtq/HH37CBpZsS+t9mJEJ0uMIR41BHNOR
g3NmcMCCFtoDYWt6b/v5Rd1hZq6LyJd0jsBERxAvev5+KvWPfDqTjzw7yrNM4YfZ1k+z3aTc6xB8
2EBy95kROVh5qF5IoRKsRDe64H9ulS5dhGjaD17DJnzVB7yBE3FwSOet7nK4EQhfXMgCctZuJySt
0zEW6iMNxODMRua2bRjbMTKi3DEG7VkNl5m6VEneyRvPGA3wT5q27Po5pABuXnFIqB+s9/k1J3nb
gDYqrGMAJ5PXI0dOWitifWbWITOSd0o/UmxrjCfL14rfq4cgSatGSgVlKBqYctp7wYPDm09n81dP
1Qu9cNMW7To47DsRTDMpzhX50YvErckHtfGcwwqDU8cQ0c4zPWEauHZz1oRFMgM9xK2tQXPnIiX8
KCWUt4TLVNgdaeCi3Z3pWAS9p2sopLfxLtaYxq9YJenGYAjs77g0K74DQRGX+1dEMOWgUXgwumsV
sbfVEQkiw8h9gz8oazK3stkF+PQGWgeDFhcIMcdSGKtRywLluamy8jPLSS326ToI5ZxyxI4uWaG9
2+WxaCSr8IFn+oV9y3awwkxjMQXmKOopiUIx4Q7ZyHvC+IAxOjf7Wfd9ClCCuZCJ98ZK5h1i+wNj
RhgV0mgk3ubvu4lcHtwDYaaF0lB/FMf7A6mqR17fIPdwWnUMa8ezB3xZQxReDh7opkDJIIlvzALw
q8IgmAJEP0VDzyXDQjUnBu5R/I4AAnao4bvRszfsQ3SjwXkSMbFsCEit360HtZk3nNqvbWd4QAWl
mV1c5J1hitM3Qf2YDjzd7CZrunCOzSZ4pJ6CI1Hquv1yg6VJiqccs2ubSMl/QFQcx6lULEqjqV/E
/tt3wt6ryTdJrR3MBuuRcpBvS0JxVdYWWLfElrCghGSmi3KaIOrUNZbcEwhqEbq1lrFBHfl1tJKt
kDyAO+WydToNudXu2maHuzYYWKRHJ3ak4HSYSqZ2DeU0uW6dnpRZU/CGhujrMJuFulnSseytlcar
Q/GexHOCAR20ILtfkypJZEs3TxiWi6D+/54Hc5JP4lHjtFMKRcXDh9CO/XrdwGw3xcaz0GbTG1C3
e1n+xf5oYhA3dLiuDQRDtSshXv6hZo/7J+eUlGjnK00rcLlD0gt9TsUT9vWQg6xPbU8sYH/GSEvq
6gKn4RwvIqCHWoDB4YtVf0UG7MZQH/gzhGUdkRZFJP3+6OOg8xHiVJYiGtZprEI7Aq7P1MclcWmU
E34vHoEc7GgC17MxMddIufHdKrBbpzn09V65IzdqMdC7+04/nbtD2Rz2G9y1UUfPeIcNG/byMY+5
u4SaqUSSvYahDe6XSR/5oDuBjGbCCkxlPuwxeYbUHT7tZbLHOg3AsnAGV7qu7uXFOFPPsLLdAqeD
79MJeTi9u1It8vODex4aLloY3HE777UWcjzmsXVSo6f/7dcREkGRan8CD6lkJqKz3Y7Od+aZfBHJ
LkwMtvUMoBkG1fRqwMy1EOs+CxmBfXYuS9gQrgCdXSqGHK7fHHRXAn0eD4Hgk0JCeucV3uFRChJ3
im6GrAL1Z4l7vk6NCzou9Q78UlvRDEinXRcxBt1vi93uCmOa2n3f9MJbBJpMrGkIjohD0PrfioMK
8j2YJfBqSDgnPXOO3ua4ETvHWB7pVFNRkxM+JJ1gXCiMNiHW7bOxAy4a7KV6YIsYznA5of41q0ug
+oo6zTr6rgh8OaBeYTcQlGdbyce+VnRctmyEByOepdsTc+ShwJ9k+5jLmRcL0Ze6uFi/UhO6yJ6R
xdLF6QztrVyFIxWglaGZDfJ/fGBib/W7bEBlzwObmokixk99hY8jFgoHS9paNb75BQIIO5XbfEEt
Xf/UG+2CZzYoa5g3/01J7vRpTqPOS8w95Rle6kKthv9oVtCVH6sBMCqw50a69KMtHUBMUSYIJXrM
/XbhJqn/CEoml800jfEHM9Im9sb65+LVG213L+n+2kLH2U2xSGZROJNbTucYnmwFyeTPGfaO7hIj
FraQijFiJlFse8U1shYnv+fI6KghVFO578jWMvUK3bFlgkKZwJwiJowZTyRNEeBEMIFJ7edYbPiO
AE3UwIa/5rZii5qQ+zZl+OjJFAOl6Bu6WMekf4VhOEYmRq1OU6uoa4b41AlL++Pj9wCgJh0KASVO
jrp9vDZFEC1rk9Ef1fv0FRzEIRXJ3n1FL0xcuXThwtnB5KRSp0IAJ/duT5/Vy7M9Mtezloql+o6w
Wr6HKfA1kHfkQPUjCJn/AZ+AlV3z4NFvuVHqeBZhMrMO8mCMcaXyilohAjqxEMqq69nJXdq2oGpO
5KgNWZOKOz3aAz4Izfq7eby3FubUukTrGORc/oCCu/gZscW9byuAGh7Bctxm3IDLYNPn8qLMq+Kw
Zr8SDGnJi4qUnXXp/lsu1BxOuewCB0dJFdSQGOEkTadghtzE7ZJma6oLN3FYbFnsi6puoCE6QrgX
VOZCgLErSgjVXq/i7/IXLqP0jPL4X84DfSZShF2gmF0kLcjw62/SXCT6m2GlnOBYIs7+atbFZ3OS
EXs1tNbBF66db11LPBFYuxkS0Lg9lLR65i7AmfhlgdrwJF+SgwMaHT81mqbQrM+HYa+3Lpzc0Ytm
tC2XP9pmykwnqS3tr6MAnFXIY9AqZ41fEBGmk1piykNXOJNiqrDjMQ4Ud0wZVzHllgDXApGdPdPH
Ls//kzw1/yrwkiFmnNL55B8jPE7BfOkdS3lQlPbG4/lmWjpBwgn45F0uFPlojebD305RNR5vlWxY
lY5OdmqHIc5seEVLAd7TmnsvT5C/Blw5qu5BADpqpKizbh871cWvMrpUIi2VWavQdCUR844HLdRe
htdGJIbt5JPaD+fs51opR7GbwYZICGaXYwii8Eb1SZvi3PUNwM3lWU5iMu8S6j8XqbtMoafbZiQ8
mqYs03jhFCB1vNVIa9cBERR/+DvDRdFN+EQx6ZsoAhzTOFcbV+AAvG4eI0jPJoBuXeVk+bZq+3Wn
BfIV4nj1w8Lu2iXvQ9hL9E8VQ8+U3VJxpwRIpAiPukFW1bB1+wiwigkXA6kCJaSeuPgUy18N/YBi
Y3/KfAaU7zeaFkSSNYgWKLBADoPgt//8/HzL1H47oiJmYenlKg1jGGxPs024qv/FzFRpzNQ4QBvO
N+3jF5C26YgdC+5Od7m+WDWQpuQyO6c6IVaIavyKnJW+RkhSCxXVDvhQpUDVEAreiFqGizfECg6U
EYrO5eGhwTeD/8b4b4rXbXof6HGdeS7GFN0gsLhM6EjApqCKH1j+kc4umMLZlxkUeaPTdQqTnwsd
OZTRhdcJMMLXW3EcBdpM60Lo9AILgYhwIwoLgIa6WJeVdohMrZaZ8vrMeLkIYFVSKVbt+l41AXZf
xEtfj81zxUgZWYx03z6yGNe/92c88Sa84S2lcgkY
`protect end_protected
