`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m5iOpzub7ElSvNREJKdbTL5RLQ9zyAjuJTXApD0jwU+kgItID8+J20u1MI5mjezdJOk1t9nA9OTm
vswLkwO0wA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dJXhC3s/4g99wIR7EIkz97FXP5RDA9SlZVF85tPxZ5BrAo19QP56K2FCjSgmHYm9HybewviTRalI
7DOxbDMLUF8rNwN7uacq3ayRTbCHb3ZucEvHPKAC3bgcHQ9gucN0HwA9h33ZqAn24w4xs0NNAWcH
WzsKWnaMu5T+I+QY8sw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RSPgLRh5Re0AkeSsCtx+zIXn0HOfm+S4D5ftIyGBjfD7tpliGOMAT1S/hIk/m9nrPJlKnHCOdcAi
zkCLSlLowrhQmHQYuJpWleJNhaFfrVnXIg+5XUlm8aYO4Q0yeB+N+WdjhjTfzz95uxMplJs65lNv
Ly7kyC52inQ2MqmglEOlQMbC25VulPWXrWgIn/l0v8X8xRPy9a7sbi8xKEQHUw/iPghpC77mfV7+
vgu9eEqFP6vmuW9QmpVld69fhnh0TpAWFEV5J43mCRKaxPGGBYZbDvxFgKzKaBffucsZ7BpZuMdg
a8eeWiF/r6pcljr5m8kC6vILjwLkAutaR1zT2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PBJG088JbTbb61e0vAfG/du7QOpWkcFgeD6A4cbF5MJ6NyMzlrcMczTL8RP2YNvHjg1x/LR59mlY
OcP+9xYgXyOxyBmLkEZOAWxJOrcVFozO/PUywT+DPTDDZtxKqUASR0+2tweH6lpYBID8pWYgRdDk
XuNbi7MY1ieKbOsf9WM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ozSrwMVOz5NsABAIzoggsEzn9/8bmn2KA4BbFvxP2GWmtueDJtgpu3Rl9ekreMsXSTdd33iH/gaW
OUHCntuLro5R6HYwfCmpvb/hfUnNp6+aKep/+IIf8mDSlUv88n323fv7PEAF6QdiGQGzU6CM456O
TGj1mINzbXnBSqoYxUIjagH6RA5XWNqn8yk256hScDL57lqiomE5z8AASlnFO4qHOT4xySWnpYot
zHaL88wtVpwynGVGB4290WDEULvH/qna87hPXSr02tj6fMFL1bKRAcYmUHUoYaKXO2sEXSQoQq0q
yuKS+L5aPanFZKvMu/FuZe6NC3nEqlAFtuRbTw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
cnomI0i7kR0hzx/MDuGP5eVGGMvvHQiRVyjSLJRtUblfC2z1tKr38FweB+F80xGxY33XNAzL2HP4
raLDX2jKwyAY+PgzbK02HmDqONupCFDPxMwtndSjYUQRCo38bqR1iY1JDq11MtfD+IlzVWMg0CHc
k49Vdk1Pe1jeyi0DkYihlm+NJ1+e5MtfMjU83ppRHK06tAqjmjllrkD1c054KfSHqWKjOPLG7Yyo
s1dF1rWWUyTFICOk+cM7ssDOkEqvCdx/QnKds7qsyy5lHlzt1aFhUfQ+orIEEEJ5EZoB4PXi9K8F
8PYBvHrBn+FsnFJzZdAcUXXP+D7viod0CJqzWkK518LpE6gDreIBqFVTkYP/TYwqsn8UqrP7Bmdw
FbV6nMKjDkEsSmH0FJM2mQiqJqEBRVnYE0RVsj9GUG15UtILNKLd1UowMWHmKAQlNVkyoBUrk7AL
5Ydqe8rBjEsXb95YCc600c43ZLBvFWaQVfbaL6SCBjoTzU3qVc4+xyTwegiuVoQR/1Sv8Mvy+gCH
5ktP6vIBiliaQWyzCP02gZPSvE8v0JKpbfyTH/qTvlJyzM3MPX2hPWPFqTtwxO28KP3pc8HTPPV6
Uz7AhpwOSuAK4Fa3sHYiWowU0TKGUdG/IskkPHrO60tjpAz3GKNYgMkC65fo4AVJZWecLLc3TBGZ
PSm8cwH1ZqWhZ86D9IEcLBtAYEWT6AdpIF6TB6U6iIkwftInq4MI6Jhp2mJU5ylsSahcvo8D8T0y
3dCUWE93KbhWXAQKMuNmSoOuaEl5ZXJvcxkUrgJFrX0ctiPXCCansSi4oFiLsLB3uUXQQiRJoApg
H0DgSK6fG+4sZYsK+9UwQNxqe7uSZ6LA85IzYiyus/IYoUkAWKyyg/tQClsSsavEtZI31Sf7jcOc
gmLJHTmsGk3M5A4Tp4uGxbj3EESRsHj0aylHPMg/b0mYgM+4PwAHUAv8nVfKiVc2z2bEXdDyQWgH
X7Cp+bwJMlAFXq30bOBgjTRT380xNI69LTqey8vTU4YwvYZf9/Ow0AuCFHKP5lfhapm1L77H3jg2
zp3cwmz6Zmit2j2NGK3ju4e0TAH/S9OvtkD1p+udvPytdeBYfyl9/S5bdPeIfClWUxVSmuhVydj1
Mm3MWx7G+PfcnqlqvbwmQ7+e8XU4IXVzLOu+4mqMdJvA9lc45yh9ijeS3brZsWNLxEMKKMWAeswd
F8Sd7Lzq57ORW/ovwkaxjWYw1txjDIQ5cjXJ63LzPgXBGJXWQgtMMCTeVbGjNISHTvQby7icf7ih
B7j4telWG6dJwJlqaxiVRJm+Q9bGCzZ/es3KsLQKE0cUY0uiYImLbtEVFI6etji/8lEOpZ8tmL4I
a6g4DmAwP21CDYIIQZZHgQh6ZgBqerYjjj5M2w5gHERetJoCYGPvLWBDA2KEM8opm8DZNLsv+jNd
P0oXhPG1AgUjPkFn/638OoezZaiQmGX5Dj+ViVxRNp2QkNF3zGpLm3rYBq+OLjzdgDOI+hYX+5U1
yb+LaLmLw2NQ0k+c5w4XoehfPXfWHwkcImIAFf2vkRSfYyo7AWl3xL/7K+jH11gC4QsoEktEiuV3
F1ZAGYulX7P80+eqGaphbmuV21TH5Pt/aCTW62vRMVSj/2hJUiwKk99nxF9Jb/iTwdybiBweHYtk
mTrdNE0zjx4Sehmp8DHAi5/g75PvRVZThzWFEPhD5F2LJj7nh1M2697LGwTGjo4uD9pKFYmH7PEU
U7Sdwh1RnLzHPFFE/n6pW81YteufclpsL38cNDrEtjnhQQP8Y6PgywgOjf1NmZQteWk+0yD7GGzp
ldbWo4rWYwsmyLannYjt1BOORDcQ8cvhcrd54A/FjvSmpSKZeY+sCJLzvirReqMk6lgNNyUI/pzd
IgnISuL1oDx9Kq9StJl0IB4yCsmcrpUFOYjoO7AxQ1JfkJ7DliYk0ZGEVOy3HXZDLtpZMSaeDU8X
kTyI5m1lukAUGi+tniylrhSI3xJw+qlAp14Myp0jzY0BNSv32CxvsfQrA8mbWoqzBM2+qYdc0xAs
4xASB0x6jlutGWdsjvXD54Z4UWwl3BIWAKtNzq2oYkEk+WlHYciytvwao5FsnyevhBLOPooU5Hrn
1ovVy4MF/fIXsnMZmre1clyQcPh4A7VimCmket3In2cQm+bd5fc8rTQyTBvL9gqlKsX3XYLOMBc1
s3Bm9fAkGpOSIi0zsT+zHovYi8kcJdxNNUCUyEB98ZsPzLakmx1H1f92TX5wGiwT0aljFbaxNAHj
Afs7jGfYJIROIbgenIdoamXUn/H/qdISifna8uGqxxch8bmYNcZdzNzgrwlit11HipmSjuKoOG8k
RdHs6cceEmN625QXh7RCDDCIM/E0tg7rC4U1gkyuKQ+qlMhDFC5MnZkRTRZya2+qKv4eYctvTmf9
qoGL1IhCk0aA2Cv0pu7XkAxXDkDysy2LNE00IAwVAkSBtYcFAYNjKbhkK16L6PrOwNWcQE0+HhlO
6GQD9pUSi67zm30jSx7O/kI/rZzXf8vFSqDIYcAiEw9Z5jMen8uCPE0QXDCiGAi69ywDBmw2cxhf
xo8MD9rh4MLIoCfbQoDdpLZDeyjL3m9kLK9MDvFQqG4C59tWq8IlYSuBjE/JFn/9As4WCFJ41ixP
G9XfoEAdcW0mMYsHHWtHWi3lfxbEtwuV4Mfh94ihZlAUvVy2QNWxSteMzG9+gVm8bcDnmNaFV5RG
F9M76WzBXpiXGJOH9y1SiARj30Bhl+NC+oBe/UOvroLgmmQuL6pU4rnvRIeQZi+e62xirQ+S/Rt0
fKWZt3zrHZtqfkatTTCRaL78qs/48uvBvg3ctFWqCUQGIP9ecmhbiE3bv6B6xIlzjR6plWWb/o/5
6HFOqvaXfMJ1gVtrQ9KNAbPVpZgSNEQxsCrxRnfjrefnKLcwo2aEsJEm1vGRrVk3eipnI/w/9Fc0
+F4vI1rQUpU5syWiwgkhlZNMdfhCR4LVYqhVG0ZA9KA524TflMR4pc8IXEk+tWNpxhnF/xMMZFa1
sJjikSwidEPA9/JVWLt9hUlzShCP1kKCkk9LkIwZpoYe6nhuX3EEswCXJzFOj/gxCsw5mAf5uCXm
3xSnEHJ3jNKsfx4YzWZ6PKIBPgCMmhfCMPW5/OuwSNdi9QYdhxbwOb29QO25NXbvMzneRzWNab6C
8HksX3ZjHkLlgdZ6JjSUEwvlXYON/B0dztu0iOP+aj6wIi8/alXic82UXJlkZ7mR6JciepIhgE6w
BJDBgSqdKfUVCVMLhn3kNzfO37YIArojPLgxXw1pfQDF5C4KllNuF+QrFzgMAbdS5pxRmG7vEw3A
sGr2pOeQc9aJMLIpmswxSEvEk536HJsjeekT/Rt4f9bxlBBuatI3I7SitPGT12Mri2MEFgFD7BUa
QObratw7PtUQ6Zy41BhBNLYNrLcUgUaazAQwrFMA73ZneYzO/18zHb+GBtEFo3ngVyuWeYoumTf8
TnwgRifvaFHDcqmfQxlgY6IlSt5Dpv/CuX8mCoXL7cWF3IMgl7qgeuTMNfKRT/20eT3JUTCbI7wG
3ezQ2ejFgFlcIsG6vQdoDFajSnGsAW7GmTYcYBOcFIye/+6wFOvFSZXoUUasViGtmMCk10zzarq/
avob5t6VKVd7euJymYLHqmRI4uaFAtZT7O7XGkJhyyQJOdQxY3xY6YqYbnrIDp1WmzduiI7+dMiK
83zi6nZjoH8dYf/2NhovLitfo0CI64kgCyGhhRhKQB4rZgZceHb2qxIqNJKRuhmimHG29IQSVrjX
SG2SnAvb1JPVAFNnKnJIB0t3S49P+ohvNL0nnhl+/WtT1NmtY13aqOox13uXobJpqCt0y8Lwhm8O
pUoCYM4Gx6PPKVEs3S4BRolRqQKoJWqbeZSiok8uetr+oQoYx0Vq/0MDtycrn1KScquL0CZ7b+lS
YJ9tC+vU7GnaZd86YaduU10nlqhhXabLlpLqjYSUDBpSgUG8LJvHXtABcaV0+LWQOlYzg7KJeEHg
UpinLiknPC5xINSsUTFigCxL4uqB0G8qn7UGck6Aie85CtKnDsNqSG4c/4ovY67V3Kc53cN/DNye
Yxpi4XhpAgNz8EGWnP4poTz+OtFd/QcLGYcp6pMqZd8AbZ55kRDXGvSGSpU7hQRcLd7EVI4jue9s
s97dBgbWn2OMCErOseZcoRmH1I4CCIaPRNR+nV526Y93H5MYXlB9DMxYYcKk8Sbu6rQxIatjGtzF
FFk8cE/mrrz4bDauo4GGrOHdxb8T6QwBFgb2JD6CdACHjZOAiBE5AdsHd3ujj4UwakVBWvA523jF
w2KxdA7JNSdc6TiTX3ctOagm8zma7vZn0t0WGaK0eAohgpyFkzj1JoxMvaDl1HWGDYqtLQe7CLvm
V993+CigGOyO9iqZiEp1BHkKCYkQVcCALk+4qA/k+cK0RmezWXPXJr97sktpXBXlVURHuZkGNZw4
TgUifngX1NhMl5K7Eo0my+for3nfBe95hhXq+4ngYbWxPW8CVQlKckr0M+9uuZ5KUznjjSNb4oiC
fw219lYkAfnxTYiwFOu0pe8X+SW3BgKrtTgXYgUG5gIeYZ4MbYW2BZS3q5aIW8xU9Nq3R8Cb/YNt
mr3lghOpJ/4Cy8Uzm7g+WpgvCh3l8wvwJKy+3oM/NceXpTQhP5ORY+cUTJBO5kXL8SdGL39q6l1q
/WQyT2Ak0ynBOAsK4gtrQ8IlFPWbT0jX7HJ8UEjV61W3kp75kxadC7bnAF90GQcSDkTtDO+QNFGi
z+nMOBXxPoKr5Q9G2DKBjZnL8apVnmkKfdHO6LAsE2mv+PdKXYoJNGdx18sEh+0z3XaCpZSwq4m6
vpR6Cdkm7Cg29Xtau+ucBEdrcXiF5EsDPAw+4TWtrjTpUYQdWcLFFA5QN8IBBoedGwGn1XBAhWwe
SyixOmuHTM+4F5uw0NCY0TsCbady3GoqGy/S8UXZcYYm/onGe3Rmd/qs0tBACQyFWzfrH+LlU0Iz
uzosfP2vVk5ExCLl0j4ZZSCIDd+AIZzA280JtBCaXa0hWEKWwhcZ6ykFeg3Z+XCjDLAT6y9EIdjW
IjyT7idyvHYEkgHs/q/egxBbyE+4ANv/KiPJJd2MYvdr1RRiw2fCipFvl6yFj+ts8RV8eVy0f2QU
Xai2129AHJxhbJjFp4Qa6P7qO6tVeKSsyDq9gwzRiqO4RjdJP7dz45BW/WdrxDfHrP3cAczJyFvN
yEGcfwXkQRbM5YCYkun34w9kyjQP7B0uCNCWRrYVwsMyDn0zK7y5G6d8/A666uVIJQou9ZDug3de
MysQU3YvaczMR2gGxyTOnIlD1FIhCcsJ59QYbERfTh2HGX/uCNYKPM8AjBqvFdCoIhUVX8EsybTe
v2mJj2dkxuC4iw4psGWtZgIMs9sPZoTT3Kq18rCRzA3ovK/lS/PyZbJFJgbMQu2BhDDRef6+rtAm
pFoqdZo41LTxG8ZjsdcSKtLzMwH0gZnPs/27F5dPyv5vahn8Oh6E+tAgzQC1eSv9DoYh6N1yZYiQ
lND/LxD+f+oMzcl1JyIIqtJ3ap9rLrIT1J0U9ev8GXn7hP4H57RJHBVZZCrIoUO4XpL1EsSUCTfO
zmjqvYl8+ajgb+fZ94Sm9j/dQMz3KJ03sv/VxGfA9y3aIF/7zvOvetveVlnO3pTarEh1dunDKRZg
dZ8xOhw1YG1kkoEt8dcj51B2zP4fWewoxhiFjW9b5g4Ll6a0ulsO1ZGwOVNqR2Rfx0lGJBKj2CVb
iZc/bq5gAB/FkyrJHhziinSH7nPQLYVz8ma8J6zTUJPeGDGaEitngxf5UBPBL7QmU6VOcYDzxdup
6jARjfqxAHfvdUS5ayt5QV3bavhofjbQafo76utlReYwZXElUem5a/M5ucPTV1C0CZ1rKVTFDOCt
VE9KrIZSDmMoQNVpkKjYD52HZW7tPBtEMogyFc/Fodsy5XKwatW6A2/3nqBQiUjfaKXihztUg9rf
/8dXIegsj6StxTH7OVrY/Q2hoRW2KBW71WOOvZGNHyhEUJUmtEmRGpED4WEVprkFHNptyjZqq5yy
/Zu1mHTsKckTyh0oVIu+G95L5iBjJhkVXmPgliApEgTrmAm+BaK4iKsWF8oUFW84u0aP0jp1XmXk
XXcYYyCsgIU/FPxfHhO7s4RDYvtxJuyxTC8cO3P9puCAz8ejpRsB0IWJo89KgkyZoW4Uj9qPYY/Y
Dw+AySvh9hD0S7I9Tq1+1E3NBKmRzJbWxywCHrbhr9ILNSU2tU9tpUADwbgthMEN6W6YZeFGhYRt
P7yO5CJHFzkSebsF+LxTQvY/uhSczaQymw7fgewX66/XXrv3+ten5gZanucJnEfod8ZXYHGBLJA+
lCi8a3dKoOW3uqWFZJyqYhF6z2XQTLuduRd94uMoajJhRnOrHi4t309pRQP/WJdXOBRNXlUPt1D7
SFgJYu33Pw94IUM7SR6h8g43mi5eccMlOXbccTAdsNBx9VkE2vH5+cKi9Q3iX9qzvqKwE6zzx+WA
aiPs2PhqzXHY3Ci47JcajFu1uM1y80MhlQdPvXiOoYbTacfIKmFUR9ojimyrTIIMjEOwE/RbIQ3H
R7ast11X1RtKftOU8I+9fvi54qwjD/g8IM7PVXK9LwtV7tzbdXUKM3QWtISZByn5wqX1VCE2ME4J
fhQX10TIB0KCga081fIxvplJge2OyZwqBsXygmwSgHOHcXc2yEbrd+3F+e5Duo0CFPVqUnVa5Zdd
rJmhc37Sl1AgaShP6fERhpSfzOerNL08Tf9AQVx548BPmw4Sr0nzztncrgUx6eQSDlkzAU5OLMXo
NWtgq5dotQCG0a5a8ivvZweL8DWBxygidcr+TQXOMSolR3TVYGkBCMoRdJOfxBMVa0GeHfLauN03
wTwy8C9RL9ozLTGduciQaZbOTi/3Wyds7pYMYG8DZMvJCjWRwjzi9hp0JONxnLgblt1ZE5Cf597h
jwU5OMDgwKk/GMJj33Ps1xhpO+7/z/P/CJK9NQu73DhQFRmkDvp+MW4Y5k4YhVX0IwbWDSTsPF0F
Cl7QdmhO7onjZxGLyCkYRQXB5kWCj+lfArcSbgAJ7iBiJAF0nBNf/wHsQD4dLSQdtygI8HHXHcNi
aOkQA1qGvO4PYZ4pxuzm+a3hUMdB8iXFtMtvJXSO1isfUZVWaSI1+MHMuiFqxptVR9VSQ3IU1HmH
01SZt27Dh3ZMEnJ+y5sCfteHND6j6W7LSpuvzliXreYj1EiVwZnx1hmEfWq8sZAYHWcijHMHKK38
u1RqD0P/PELQlB7PLs6nzD/6VMSGK9/FQSR6uekBKHGul5etoFbOvhLu0zAwFa7LQzOZOJM1wBCp
dnnCa5AlQi0IwZZSTJjLwxv2y7CDMlitEzUAXTwHFX16rfpB0lleVz1HhAeIHrYTHi01BXvPmxMB
tHPBGt4oNG90CQQFpEGbyjPdOmr7kEO0IoVw7z6AF/b3WtmwgzgOwFAt+HSrqYaBBQ6GjFAN342T
e7cPKzwxCKGkW2hF84+LJ0PmiiloTyZa8zRK3CKP0HgaHCqe/vEcuwZtpBMBMu+OkrnE9hKvLqli
ugQYY270qEamG7e9KKey4s4v5EjhOpxGvzEH7lTjTWTzNf7NySTqMS3RHPedzcGmSSBBgV6Bt0rz
mi2teqlVZWmCbfX0+wUC/tppy2RG1r1pMM+qBlBhOWeeJ2u2/PTOfzyP22cM1y8C4pP4ucq+WLrb
0VAi0f2y6h+ycpUW0gj9pAdcBb0DhoifkSuYDEKup6iba8UqRC0eEKzLD38UfXhRNCcIRPuCwfN6
HsLTNTKQG6pe2BALTEGLEhffyU+D8EuB1r+xSzPi4KUyb9wOqD9fXFNxak/lwDVHocuJZDn/N/6E
BZyUgde3PXFRiQ+1TqHIADdDenyT6luAZ/PEeNY13KnkC67Q4IYEA3hap2ftS3qxUDnNA936DAK6
ZfthxWyHkttsNCFa1RSoJNvdMGZNTYhPKdu+pd3N0mLgxGFjI4CttDBJOgBUA5cG6zmogoVpXe94
t/r/S+F3mFOn57TPQuiURlkp9WL2Ieo18eiH47GvXSlYZ3VEEKg/Id3/tVMkiK+vZ3h/kVtPNzQv
e/dEzOURKr1uAmlpDgMAQlSmUonrEW/2560Z/9ytTxlNHH0S/m0Xyf4ZHtioQLZN6ge8QrVGi+ul
bBajixWlHLye279DWpPbJT5e0PbXOibRjr+jv36nO9p90uuUedPHneqANVbmyW6C2EHq1AOOib0g
Mk+sBl1K3AKVPTCuN1AM5bEkf+OP0o3VzVe20nKb4GI0+Cx5cXXuhVax9wGUrTfdyJmxnNBKFjIc
3nww7LZW+umOOJhF1j7UbQbthVQL7dXuqHHFGS0ETpdEXGUomXVsoDDcX+KgX1v4ftQzpqx7isQO
LICdZxIb9zrV9Lx5SlMRGAQI3ArTtasKYBoERuPVzVQgMBt+fj+HWwMnBbHw1WNBTBeUNbf8FUh8
IF8J4Zy6HFRq1YVUAbC4Deg1pxLvpKD59msDzB7T5PO30rV5Kcftm6Nmdu/8cKgzutz5w4NwL6qo
MKAXWvY7s1/FkCyt+WJcnI3QApmL7FFZ6zLl6tIWT8fmeOzNzLvCHkNmlDjyGSogjrHb7r8HbPE3
R3mASfQPaw3eiVzQC2a7600MZOq0YsUcetBLBjwqanLJidJBPM5mcjGOCi9ITG4k6Fb4TxqZ45/F
bHjPPXQE03FXLSc+7GUso+E/5oK/cNoMlX9hUaMIupo/Uhy+DgB1Ss8i1lEfLHVuWb3jsuecN7Oh
SD3+PBlHHU4sVjtFIdGkh54Ya5GERxW4VCYCuB1fLw64sNl/kgVBw2IpJBVxZmh8zZ/zreJRGMCH
J+zjGYPQaHHp485WTSlXMTLYJ076HU5Ctuqz7wIchwNvnLb+lXAfo9UklqqtUIvfpVJtrcNIYP6+
u6NdnitXOn2dnah6MPyY4IWEFNzASgFyBrxoR4pRoy4N2rveQQjW+IGzqZslorQ8LZ3exP6imP6E
efQnMTNdRGNYqeQYCGD+z/hDZoM85peTKyiEkhh8ngp7kOHndV6zNs6DePSTP671/9VDmmEVuHYD
x5KmfOraYAFnran2vQN1oLUW1IAps/PVi9y6NK5GB4Cot/coEPH4l7q+CwyIoyh4kBxGGqRcAE/y
x5h7EiGFr1dOtYrTj1CckfEEJDKGj3WPRr3cgl2BCtPOCM+uivgdwAhKFnklbibItS8HNTiaosn7
HbqyPFEHUQLaqIfpNZ14aKaQjRdGb2MLP+G/2Rc7wNCEJgMF/i6b+3VbkHow7bLR2dkrtBrZi2Xk
LfqkzaQGcuOeaunCjkFRN+K4moIhrlXnQhPDEpsugPTbd7zh1u3b15cxKAqps7s9T6oJ27PAypbJ
iMqiIKagEFvTnzLZk/76aKLNuFLZyeOwxMupDYNfC7zNQTJ2v850Xh1VLVyrtrLSwnoyfGhcuoJP
CmHEXgNiKkrbNkaLOxVqMBbK1VibpFje/bPDkZ9iFqE1eJR17r/jwcH4d3UlGKtnsdfjWqRM/6sE
S/sQ5SxyggO0wUV0hdNZcda0RuIE+klnW56nKkfbSkSLVaJzG1JUJt3Eq/HjqZrN3933/BOD9cKq
8uYd9tQuvdRkVscOjvo5h9VZGmWHIfX8PeC7CDXZxieb2MLkQV30/fNGiPFEoPDBusfrMnwjtaNb
HxGVbZudLOyN1ar2wHSXrTtWoBs83091SYxhkDZ8ikff7K7MH2UlppQA8zjm9VH0OucwLNeNiTpJ
9Sr+TCWqbbd5w/7SW2rZAhQu/lQHI2eoy7CRPKSdSrgQ9teykRztDBk/zkWdkPh9VhnCCTsN5fkT
0sQVa8Ym4aM9ab7yuwpW/degaxlllDchR7Z6n7m3+lixHnRz3+Ttnoh71zeI4sdWbIiR8KIVXRuP
7+Wwlnr2MOXhItX9HOE+Zki2aSfHLgB0Y2JjVIKRM5eokVAXbC/8Z8RTk3GMsiDfOLf5WFlroA6E
cynXrxgNBUZ49BL+ws6yWVsPrj23uwG5NdHRWcd2Ny+XqYfDmy8HGMxcRB7l1RfG8HiXqFNKyWs7
BHN0TbLP6N+aiXgl1TULBauLrqiPJ38X8+FtVLjGoHvq7E9+nhPxiWglzVANCehLpTwF7OOLJGlM
RKBjPQFjNlnjSaN3/6zHO740x2S1A5NtWMXUUfsMC+VrEeynIB9qzPQI9jI8507M2ah7x9E3GZln
3eDl/NaOLIqgSirS6Rz5dfPOUBj91P8MGqfbx12hsn6CR4b16Ja5OgWIUWZF2Znodb0kL7KsvPkr
tMT69CsSXh83EmQzhjLGqPrvhjNKQN72/51byzNvUrlb9LI9ux9GgR/CcTgzFJhfUqYfYcG1HDn+
vReU6lM59WJ+9qEV8WS8DGzxwja8jTaYO9YxwtxHz7l1VZKWoo5gpoAHgKgT/+os0I5zGSNpuPZU
8tpdySTazhCww6eJ7pyT/USo/RDKGt8Ju1ZgFbU6FM5XQbZDNw2KNZktHcSPcgqXe5wo0YmdBQ1W
yfNIc0oOBn9de4mnE51/lFHVLnnUXe8dApeCWmFn1skqFzBuIXvd14NPU75jNcn2bqiFuMvYE9Ln
YMl7JLaI/kZ0U7uQ3p+AI5kYD0RHV6s8KJmgLDjzsFKn/9E3FW7swK1YqT4lXbedw/WG+STmczoo
wxlF/GnKz63cPbfbbLnDDyJx2r9XnoIi/iqhCbml9y43bilyuKBSWsCdUYLR7/VBop9EXuMFqgoM
VO+Qp+aK1tK4V4v4bT9w9V8frnDwzA4By0doBKmj64CDSNp4Z6mrOIwpTXugDs9k251VN9ITTj1Q
WJY6JZCA2K1aPL80kD+Ln25Cge5ur5afqIwMUZIj0yITa7/Pii6m9xPIYu6XLyFarzHBYeAgrch1
ot1MolYxfb4AlCHxycHwhdlT+p5bXzXIZi/+02XkgAKmLNEpvPG2gj7lbmsFdGugegs/+sPq6vf5
5lCxMwocVGnmagPzt13UXwGJMQ5rvX3AsnNGKk91Nclfk68fkwtz9Fm/4h5fo09ngaH07IJwlfV6
MLum03Rm642atz5gy3ljIGHYhhEeY08QolfLOJqHQ5u8huwbGRNFobY7ej5MLxmQ3r7NGxFyJBD/
PH8/xJpxDVSgOf3ThF0Jy5ww7c1NmD9exozeP9sEreAZ3l7EmVpC5OXo+VvGMkSVLTaaRSUtrn9J
lC+0v5TVikybUfKHNUJg0fMo1RejqxrzJtwIfaHjMvABQtCDpaE7/8syHmRksHbtYEXRGtmsloR8
B3gRc3PIEiOacepYqpCQ/lWF4MvWnHlbLFLrspBFYbs0u+eh1IDZRzwiUOtlaSErP/LmQfNZtz+D
m4JEEYozIGs4pgCH3B11PJcCB3QGraBr4Q0bX6rmtpYt9y1DkUWTpHuFsz5oi4bKGmKT+fjzHZ9L
gfS14YMwAB+FLjIbCwwRyk6GXCane8GaIQQemR+bkoW8seFWpO9kN8ByIVFEdBM4Wz7b6JbQMeFF
xpNwxY55wwH0aYQ28h2ZyncgaS0/1cgNLrYhBWeIlpP71enmeU8zcH7pEdLFRg59jQbQDJesQUMy
8vUNNSjdSCJV2HhnhvY7psessJLjIQowcVr2CL69/TLQsHFN17/qosZOM0ljoUQO4rOfzDx4AZw4
W6IuRaQUskfU/sOHJE/DiSYZmyKATihq+bsFo+fI8ulMBUwdXyUw6HwWdt9BolsM5b4Y90KwTKTM
YK+3hPY7QD2O1uDhgGIwYV+/18wnRnrockOiZ5L/9ETkKeV8fFTT5bu/5JzyQdLdYxStK4ubWEAC
JkSuEiX09zZ02w8PSRmN4GNlP01Xu1cEstANwiVxHOdGdtnVOw8pid1q+Y3wa2YG54Qrs0cjYFbu
kXhRT+toh0f+K0oXHu2CQJOxJ90dDvtZagROeOqVPNJhdgT4m+4MfQB1i/i8orieOpYohajL0Ghj
pq+RrC8DLVzpa5RwDcFyUUE8ZRFOTJ69LJ4sjZyB7qxqU1xf4Dd0ocNxXdQkk3PoaCG5msjWV2Mc
SDq1pbEdjyMxxV0dmfIMmRkuXePiHOqUP0wVbTiEvol/OTuiov1WzxsW+xLaATDLTrCFUsumkGu/
zqIKtSjtEvECweOoUqr5xCGRfmaPoXPYg9IFPrJTyjQOkP3JtvEspv3ztLgikivkoWJ5Ea3C2kzs
0qtbfau0+mdmvLP9qoUyBuz6OGOIMW9mn6+bgQ8MhG4goFBDPE/D6HjzOkxAw7cdlzPlDIVzRFNt
rsmUXlE/e8KFcUK3D5SGfJLhkVxzBqPfrPATv2jiS7hXqeiDOFEMa3pmnY3s3HO1yQvK7Fipdeff
jH6sgXSqqMH0M1kJxMKVN6RC7utm6zLJhk16g53Uw0cSmcYqjKfZ6VL6uZZy3KABxXl5+NfpG+Dd
aVvm7HKbbv6ppCB3x9igiPUmxhPNwGrNLQ82rMMqdRw8yzm6OE2GWwrcT3GCfh2Yw9T48des1qkU
OoAzJui86mW4nTJzM4plf+tBu/I5rBG+7NBK1aP2/5IhrvGbKynIG9ynXXAysXdo8+HVCGGeENch
1rpPUEdThMwJ7wj48Gyo2e4IW+nr3JVfQuvy5s17Pw8i20JuC5A5uuROIe5XUmeXg+HdQuArLier
/5Mz4Upx/EyAf9A5er+/OG9patRg8zAjAK3bdGxAJDi1XwD4vYicKWe8tAOR6cLbNmdSEwpKYy3R
hUPbcZ1dleWV7Qv3NUpZEA+ivupEkM84d5qGlZ4BAnMFBZUvd67J+HcDsVtBwIJkGvkOLTDN6Lzb
JnTPl2CdsOG6BNuiTSnOIA+tA9ZFCiaHdd2F0989b81oVwPRBbCGrf9fBWR/bTbmVwlzuqnrDarw
rnqbAXXd78t4ReN/PssciZ5SSlB5hTomPwlKxrVb06odu0K0MM1hHTVqnJUb37y0FKEMKRoCTCaR
gGa2gOOlnnkPctv8JjL83EQ5XG+9JdjSsQBDrio982ye88PILYSeztGlN1V/4R/DWIvZ/sls1ahk
ixD26S+SlnveCrKmjaJ6dVBJ3nPR88smaATq3oO7h8EANGERtbQLb+7/HJbeagHinLFffynDLTEm
HHnKPDXaOM2ajekxSVG4fAFIENun/SDHxQffpMxnfOoVdrASlpSxcM93Tqg3r2HbAsZM/VukjKtB
bsEIDURXwQjxlIekHey34aZAsTl7JtR1gPLgX9UyTIg7H5+VgbzsZWeh0e2Dv47hWPl/5IyO8goV
kVYKXlr9zf4nt1qgIoFXg0j6G5P0vlWHpQQqLf03ov1adW9wdjB5w6x2Yu0ieMg1bSE99e7fxXkT
qEPRTDssmD0nIYI1LRLxDsX/GAY502V4Rg9nwX/88Hsbg/0wPv9tlThQu0gmeiFcQbcpB0V2GdiF
fCvoQ80MPXwfdtDQ9jDY3jYpp4yd2u7Oi+v7Qt4dwaMO7zvGSz25fpFPPFmsaL/bdFiWW7NIIPSY
55Wg7I4OwkRRs+CL1GlqyA33bS/7GdRDwosI7Yk78owbYsyad375j13rSuRk/9ZxlGopCBrJxkHL
P/2l4gIavb8OrdlMI0R0YjFCPIPZUpotKcUDH4lNw+lkPt7ZxZhEqStMXN/rREnvh5sAuoeUcA/z
ecclJBAKuO9bPEoo6tr1QG/V4hT+ZPeT3YermlZeK/lz45kX3Mw0RfbYwWvBkgUYdRsspu9h7fRg
G/iVOCKrD9moPLZYTeK16/exIYfNFrbHnJkLuQ3ynINC21UpreDoVGmaGNUSY0OFCMV70NGO8WE6
RJBejC/y6VIN4pZh0j9p9FiS+QFjCS44eI4TMtuDTBD3jxSjsiVS30Lmygh90ExTPZWSt5oIm6vr
G1AqW7NJohHDqTZ+anC2An5+mC4KeRxx65330LkyhE6Pim4Ezn1abMSBlSTiMf/LrWaOYQX8QKHj
JReuV+eZXT7Imov/kIWzu61+2xnwlMnHLVSzy8vqbfd5vVBlNLR0XKlDxlNpenJjhmAtZxIYDOQW
FaM9gkD7eiCfaRXclHKZUUYedxU1lq+Pvz3j46MpP6YeXnHjyY/c6qVzmBI4+CeOskljzZjen44q
xAl8Xz6Yl0sSEdmZwV95foHXpIo6xlIGdn7/6W7tUvOsSfwksVl6SpcvR6bcqR8ry97rLmpo4+EC
TDA7754EQGEJyefh3w+RL0hjpuZ5VjZw0SG7THx/bv1Em4vtwxiMWjU197ULxY5p3QDSDHyldYPS
OnW/ma7OeOPqRpFPusXrmxOaVxRvTfG+/9oX0C9pR7ZOiEDx6eCkg8G1YN7AgrmKbiE2ypW92ZHq
9jlYIybgjjEQ/41k/uVsqsYmAgMvBMXUg8B69pnR1in1ULP+5GZnREQrbVwY/t5Dq7RYSwJo5GZY
pY8nrkGRfJl27Ak46W/GeFk1iAodB0WHkYoIwrSZSwWlHDY3gGkDOSW2GZS13wncx9iBYhfK54Mx
/zIB7gZIGGzN/y7mVgVgLMMneLTa72K82KTdTK6cMW2xCtm1ps5DnXHA0Ca+7YST20HBxMMxvKZu
kvtViUHKbubBjViDYmL8AJTFmIShvBEpxLPf6gd+qxMaYlLOxCqH0eTAiY/53kQ4TcvRRYx14NJH
BazgZ6DR8IgBdbNSR/Om69RlqfeL8bb58rbLQD93zI/VX5DSlYwdL7TjhAj2gvJoHbGOGEWwf+dJ
gPCNspT7IagfcOuIIuwwbBbNGZRPQcSWgGTBrOIXa14OFWz6avC0j4ws41CWyWwO75ayjWtt7bIB
YqDJL6JdVSnB5VjSoAATSwJfCn1sSWzx6wgcCSQvsVDnRM4NFNU3xFfxUyNAOuj7p1LDnNSa+ac1
JyIyMUt79+29SAyzytlEwrwRaaTWZnbrcVS9h2O7feCSbzrvmaTemPAz3fySGgAbxmZdMvIVP1Ni
+EzbksxU74g362kH5fdBrwEvdUEocjtV8su1TJx74m8FZeeGuck8eJxDLoKVB70qf+iVKMX4Aabu
AiIs8VcSihAJCSZscpeMFT/6qWImEku7Til4xpCYzZsYoP1kQi0E0qoN4opl5AsQCDI8k0dFb+IO
8FY4Rlr83mZRkuQyTETZOTGgBpS5ja7v9qgBeSaAKr9fglaOdDaZ66TtWB5M22JpAMF59xVwBhyV
r7TIZB96bl1C+1ooFOXaUHxGXK6G9SR2PJsQX3JKz4YbeyxEaiA0/4HojwXb3YveQiGYFrRxK/BU
hbVLKACO7FODNPMh6H0J+lnX38rafLuPSgObEnmstX2yyRzQzmN4/V0ZPkwiPQ3h7zhsC0WV6mz1
42AL0hdL3a1NL8pAvRMjkyduYzLxnw3unNLBToTycAnXOq29E39/WXzg69bN8pnri1yPYjYHAyfy
qsDTkLZVkIJmdvAGqMBJqhUfoZ/7lOhkbUg7hSNINTgFLs/ZWv0SuCI6WqZffRi0fYErIGF5odk9
7v2tEaOgQHxL2uM8IdKgAxSvAhgxqUVdtpPI1ImKq6x3x8eMxzYnAudQCp2aVXLC3di4FvW3bH3t
Iw0Gdo/U3X1eH8reANfVQkkd5RWYLs9mX4ELsv9Vh8zY+X+kZmUC5yc3RFMJSJ68XZbWBcADW8u4
nTzg4Wko2mDBFBy3aG09XNAltw+Dy0u7vofUPSd2mweb9Vj5G5+YvGZgjNGOPnp9gGdKmWb5kD8g
Fxq+dXRG+goFWmRHWTZRNXtAzC2zI+ztsj1Ruc0vsxtu8S2Y6nq7PA4+O+WDcgQVnQYDhcJvqUDd
51Y5R5/fMAOklzlQq4jG6sjokAG9eh775ft6AVHUdGmt2VvWk8HZ2mGgivWjT5+7OrXcb0PiJzmJ
UPGRd9rgJSW/x/IVkviCqUtDwhOWxh6Pva5BEVFMvA8+LTEEsHhrhCIED5WZwkXn/HcWz1RrpoAb
r0CAlhFeGd+5e3bcjyApPluk3cPdqxWXyUS8dUpo9YpEYSYb5HPP7sbQj9r6HYK5zxrItFY5osm2
Px2wXFeEW2bpSjbU6cUhGV1rnQnmU1acQXDmvDIAibjc+bUxo7T6VWhHh9Vs7KymRVub4q0Z4wwR
+R77SD7sYb9JdZR0BYdr1Mp1yfE2szS2AIMbj98wS5zu4I6Dq1bkBfxeFfX07KpwyPULzuq13icJ
jg+h8S7mMe3N/NVts+ZDsowszT1QzffYO1IXkNv6rI+lmBR9PLoyd5VuC00m670pcnJUxIER8k3w
OqfBoJCEFHwjLMTF3TFNmDt6skdyzT0nQysYHlwEu6vWr7Bp2Ody9+e9RO6PRVbzaQdGkcO6VAMO
dHc6bfOLI59vFmHCVBrliHHbBNshyA7DLo60fClr+ATu+ruRLLhAxfE60jWqrKCVnMNQJhzSkXWB
ZOA9LGKgCp1qM45pWFMnu2gtQqYjOdhBREdu3g6PHBUdw43o5b9hTf/qLIC0/WacLUl8cX/chvIu
LihN25Xj420khTLV67bvSiAKOrwi69IhDWBdhH9NfZbSBffuK7FPnnXTDhIfQVFzQg7BtDmrGMfj
0enR1IK7Lv2hA4NjvCv242nWeUPz2Aj6Wh3Y7Vjq1qSp1PiHRxIpCEpk36e98Bkam6PaRmdbrkaG
z/N1fBjMsMinpw/+yDPt/IjZ7+BtSUB+ejw/FVAZS1PcLXN+joa1D4FUkRegR/SRsZj3MMkMbRma
MZJTiw4WWh0Rk+Q0HG3vYL81N5f2e5wyIRVKmpZQaFDK5vbOYEop4qGkM+QVPxhXbnFMJye0Gnhx
w8mMr5pVnjBpiNrE3xw68YZqWlE3s2zPF6WBzWpkiqb/EBvOAeel4xA9DEKThSACWjFBehYELSDa
OeVLEgjQU0yyYbBMWyMhvbj/4E2UqK5IFOHHtJ58tBXp0bQ/DiKiQfUvmpz73hNbRVmHHqwzfRHh
7qxO1goQhS5S764Uk8WkBp3wQyt6C5Bfr0j4hesviZ8znoZzrT/Vu6XGaLFIwnRxU9xM4I7d4dfK
Tc/gqafwHjPVLa3mKogeVVzwrpV1YiI2OQrzq+JMNczg2ld29dkQipglCJorOhmQueHauTSwCxGP
sbLcuYrAKaYlHM7dJnT453ySNaI99FedZ4GvmzNKHRz21mc0/Vs8LKRJ2PmiPOKtb1Z8K2x/anwW
avbNV6GoJTZBqijUXnWFOJojA30D+C3QKYBpi37KjcxfTtuD7liTqndHUEF50/AG33BKGqWRsHT/
ZftKgXJXERdPyrz4tm3UCgP7HcFKtwpIG8noTLN60NF+FMDet7XtiE+Apf925Z/VgcY5nrNEVjuj
CvrfnEixB+FVrPzu+5S2qtZqQKTKeVYV7OB/YBfxGiM1smLbCHQhPvVmORAADW/sQLxIRmQZZmJd
Gw+h9RMGsHrDoFUk4xTVyRGQtpPwMzMgurht2S1iYkEX2B8n7xR7bMbXOtIAwIJPtmQG7b8skyKD
yYTZZVGKMXMKo2IcK64Su4w2/rQ2ms2dOHoz3YIH8HH810kDMfIsHcHBclgRAVAiAncwaSxh7zFo
l1+mSGf1BE+w69JtrN3ZrasaVq06Bjf28/f48nlTbWQoVQwL3C15jvdXALFF9doYZZnholqF56py
asv4tckk/prMmuSvpYuQQSa4ClQrUcauzO4/7WQgTtF+6b1PViQn2iwtLrGLRYpx/ZYKktulyLkW
st/BXbc7autJU8i6F/W4
`protect end_protected
