`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
I06Ke/HcfREfnkxxTkdiDpHDXkOiLmqh9dWloLxgvry/Cwdcrb+9YOPFy7RKjuJ7aenemnEPcJKA
t8EfDvBDlA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jyZ1bfbGRjkLmvhGXJCwpAScYeDzs53TFtOtzdB/IXBsURz5lOHiyuPeLzHZxLoeZGkYqia9Rtl4
rPZ/FntNMmT1IJeeNeUvmi3G7I8KNONVW5b04hiMFNjvEnSqFoR76F3oDYihf/WxTtwqrk1vChpI
4SD0bSeRPo8OrM7lwgY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VQDKpGQqGvNkC4qq87ReEdIwKLQo/LhNO+Ky41dL8ga9efpmqknrGhXEuwdHPoDTL82RsKAIrGDt
3T3ddD+ATYI+feqfS9mSGUJwSBAfHxtJanpEi5v8cnmaErm7trEmS/JdBVPiGhEWMmJJAQP4lJtA
2vK29IraDOVgimHczC9JfPkQ+h3OBAtaOjZU5DMB1b9BqfpJRdKqY4ERAaiFJj/Fj+OcFmvMjb+y
rHOUuOWs7T8BYpV1DFxp9e/yDrQAKDqARyLwS1v9JWS0qvJZHQWb4NBHnF3vHR39X0Gae2wQm0BU
AHyBLH0nWQvZP7Lv5Z3Vfx8Gh2e17BO0Jc3vgA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bNPZp7ZOi/5TOfRzUDe9Vrq+L9Y5/aPZ0nSqJszH2NaHZlUxrEuKGTWLxyU9pwm43PH3RUqpteUk
3oTHwKEtU2OLyFwmFRBJ/+dn/7Nxl2zxHs39BTgET9XcjIlossjI9qstrGq4Rp7D9zZN7s8TICxG
hsF9aezId2CWyyNKM8g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CEjT69Asl6fQLDA09LW9QA/0CKHuxjGwx1E+6nqTKNgV1AWNE5TUDB7lZrDyJADlWIBfm4MhdkBX
5GtHY6EWaP0pEzX7bas7n+Mb1aHa54FonXYrWKz5GI7IL/kvvuIMc4i7ggaczR1Rp8EsOzSyam0V
MDjx7uaG1NsWIsc8Rjs4ha6FVsEotLsKYCCiWLka493cy+mlOc42UztDAEYdcEAY+eTzgJR9fJvh
vUBMmetLuA3d21XYw665pSTwmB5CLLit/ZUo7ggDe/SqQeuo9+vqCCDHECn+Qa+YcTWjaqbUjrkS
u0FDz2j9+pZkmOcRQt9Fe7goj5x5XAWwmyz3IQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
gxo6Gts97rrNGAD8PtPYGKb1Q/Ylo4WwIujnVBrar8MnxBJGv4X9h0yCfVrbPnJeuZDW2QYht7TJ
MGYnTgLFhu44BjzA1yreirY+pMtkNBbblVVbk3T6kZwV3hX+rSfqut/q0rtB5hU7+W6cI1ho+5bJ
RGvHg72fBXp1YriZ78jHb4v8xQCcvaRibDjQMRq/hypXL1HQ0CeKbQG32VVQEH10R5UTVhAarSdL
IbvZU77CX2VLZqXOJCPYnJfQ0E4T2gp5GCUCuT4opQpMMeXvPg8yS0FnC4JeT09jHrV1MZ9bakxM
9IGVRkCLImzlLXEWD4tOxiIEq+7NXRVtltYtcuo9Bh+Ie8f6AXmSYbgDd5x+UeEcuspLBKsVVQUj
PTegAc11ms4smabEyImGVzGqxK1pjj/fcOpqhSTeDILWB57YINnFSN5OijKsbOrnxemuw7V4+nFJ
Gx7e31Rz1Y6PhlH2wH5oWA+e5LqXpg2ExXeRCJuu/z8mGnGiKmf3W+VFeG4Gp9jcGRg1SAqoLD4K
8j2O0IRleXCXD1XbDMZYDlcBRGmuXG7aTUi7sKvWVvziRr2Ggu2P+FcU42iBMTnaKwwUNwMMsv4k
hmgerrKFUg3aIEE9lSiSMXgK10NTZkaoncbfPOfc8AHLYybPjjm9FjyEVrws7+7F8x7R+VDmgNJh
lFBOERf6Bv+j3OECTBLKFMQIShBH2ajMpPoEwMwZwGTG+aGoAlQmCz9lCkZAzbtEMwC5KhsnO2zJ
Yw9hRVrxF6UPW4a6QhmTe5le6R9eRkiaQI4MbB2stPmB3xLxhZ+vpyrI3HzTTgHsPJzWeUvgnhZ7
kjSV9x4Am8lp0Z/BYvA2Ly22F5I6qVRePKbUroTKrikh2AE+3YcSu+7KOsa/5/B83a2c8GC0LM1I
iw8Q1fYQKYgEPJ4P5ekgwxzUzOkpsbAIoE3Xhwse2vfrVjev67POGYlwyqOuNQHAKHIdQW1kPitf
n2OGNELouVjg+m6xJJE0HwNiBRyJ/lrJoSuWCWjzyHl3Pu3lEIvgBntHIOYG2goJeyN3OSrCu0cW
8BJoJPdRGVeUb5PkIKo/loTVpIjEJ5vyLqLUZFXCC5jFcxli48GBamP7gSmVe+yua24KE+sh6VOl
v4uQHn6pAv8EdkOgwau7GFvf/Via23PRrxYfOXmCA3lEZLhyb+juxGOrp7tpW3Anfzsp6I2sHypN
QPl4yhBJ3e9RzsORmKn/7JB8ZMp1bpeFrqT7UtTkhkbqD8S2kvNkbGYUKsJ3Fjwrw8Ul5DDs5e7t
d8LpEdXsTcvNu3t7+PN/oxkexXLZb0QH/XHCsbw+XnOp886Klw6XTIiTXb+VJwRhXWJbCIZOK4uT
5ewgkKBsCSByq6n2B4G6IF+aSQVCP+t4ADU8JjP0woyFnw+ZBUdU9hY9emShdkPdcUWMsItvGt9I
Ukgk61rQg03yy2miCctPTcaHmgo+1KU+08JKgtzS0zauG9/rn7d/rL4Kv0NxMu9me53g4tcqTS07
WK6fHpg1OvCTMVIbc39koktYaqFZQRiydhAxj3zCV076KvieILTVuwnysMymhcVW2voj1V6S1760
ZIVnYoSM6R6sE9tYt+ksZZlKmAl0PU09OO8VaazHgngs6GdeNZJuMAgRou6SBMQ3Q5FaLvp6ZDUv
/On0aXQkX3Cv3UDgQSwPbQHn0eJbh8eFwnUW5Sr4nUyQpNAovFG7QSrBrnI+AqRza1YJ4w+jeWvN
4V4R12q1QYIiefvMLu8N048Fp7XhCjDKJSQHAbQJtYpOMv6Bt66n7dy+vVbEgkvwnn2ag6Volq2r
fMUbicvdsJonZHMgvd9ZKMu1zjlf9oUd5pqZp4SmITzhsDx4MyUHv4hBsjRf5JS3v+0jV1AP6XrC
/7X0fCDTB0i0QjI3Ijxj6rNyQ0SoPhD7AIgD8Ba2Jqhbtc77mva1pLG4Yz/Yfbm8V+7Lq1TKYjX3
PV1YxNi7H7hM2Mc9SPO1fdCe21992FTad/95rFx5WVCO31tAp7GfsI6zf7H/peqnZ8YaCt/sdMJv
38dEGFGHbIcO6iHHwCvS8VZsQwDQZSTpTxmPTmj9G69CgG2RR/iUnfBiYfNIX9t8fvQ+6/8Y2Rj4
fPnghmyZnzjzEriPKTJ8ucYhBjvCAxwns+2LkT3bCwNV52aTZUCM3aEwHToprde3VWeDIidvwk7h
vC0G7A25uUw04J8mZAVnOBeew6hKA94sxY+2CNLBavK4ks5fveVTJ1vqHAcuus061y3r2rqqgIt9
JB3aBCS5gkamL9oNfKAZZ/Nj6DJjDWNqLzRpy9VFFaSR4rVVjBdiSWve7xgscdX/1X5chq15w3RM
o2wiklDxUZqZcxiTb+G+/maTt5DpfdzRAM0YpLuxXKvcFnieTFa+UWK2iBlfJlULZuEFvA+kUo4W
F+Eol63mDPsrVVtQqERAXvKdQJLHDrMdnMY0a+XGv/hyULbVK78GyJWMmggOffejWdlKSCyB4/a+
w+1uSy+v2TKshwsxwlstRLwUKrONLQd/Nhkh7WZzuHo+8HyeV+3lzumVNIbN29nguw8JQcm92UyJ
gUEYxkCmEcvQQMLN/5Y/tpEwFZxypWOXed7Ss0ZUd3wsh1I5xcjjq8FKuA9/BaLWqxJ7AqAT57Z2
E1ZzTtG7PfXpSOs6DpLn+Ei+ciLB5Ter4/yKCmUZYIt3RmM00q6iNI+OqxVDnMk67Ub6qAQCbYJu
qPvlHixhGiFheodq1p9UJRlr0dD+pjGZdMzsAFLyvUNpJ5mmqDkgYwUwAARDStKKysqIygAxw1fm
fdJabQhOQ7i4HAcbbu1FH1XS04uX/IXYw7kAOq5WSJ3jkL7l5DzeHtD0hQ41zwgrC7PNOflYLdgE
YbwCEO0ZZr+PrILWPZB6ty7qHzZgAlkc2ATsKByO535NDS22bJEZ2edHh3q0IOJw6pVNg5L61yrE
VORny1eesQrkEmktoKw8/WhXSXH4gXm0B8rApr0/oWkdgPIGxULa7egRgpkC6Qcbax3QvPserztY
TwuCOha0gksBJgjjVbwlCW+5lxk0VFH9fWQKby3XhUgY3LAvkMZlxRrKYvb8ciiLwDzXjRDdPiEQ
HT4rM8q92f0sdz9RP7wFSUnFRkDkA6fh7VDdNsv5CSO9gP1eLYpC0MBALpbttbhRcyt4246cVDEW
TzfyKgC956OFCkyXZVjvMptcaAeb7wjO29tkcoUWfiWLmyk6+vGx3jyd/gWHC+9ylAulTX4hkbA7
Tlo96h8qXr6QhWA6wYGnzYLew3s9I/aDvNOUV2/KtnSHj8sOKiDOtOa4eh3cEpOW/c2uLnnDlmfh
hoaofQ2t7Jn8NmWbZG7Grc0SEz6JLFc5KBusX6hVgWo5K9khIT8E14s6F8ERDgVbiL2CeR7O0yCp
nEhkgcW6UpBfPd9MoKgNRuwlvGgYvaMOIc5Vm6CF0Ge1ZxLFk3qrtEw6BhUT/q91XstXgmxTBunm
uu5SaryPkPtI1227NnaSHq2+EKgt/RDNJHpV5TOow4AcvoRxOYqEyfZGmwWEebeBgTfwpIvXf9oz
BgjWTHIsNFWU1Gumt47jpmrL+ZsjjpgnwJ7CuPeiMNiUNLCtO3u7XwYKTdJMSnG6/fdqbHAe/vLh
vhY6VEUA8rf45wnPuRLUZ+SdxyuceC+koRrDkwP8fsQGdhz0cFjD94f0wvQsTI+ONvZOUnzTCHM+
W9QJMjEk6IJR+K3pDDhllVStbXFUZRe0TC8XakjdRTms2opheHUhmez/PtHrlN76ZTd7W/SW0C4R
VF/tCEGLvo1eIMTwtPFA8M/65goLajDbkWvMFwCe7pw87pkNSPaADNmXXx9sD4vvXaCwCnYCXI4E
OdtCEKcp8V1CGlRXJwBFd6tqjs1QYNxNTWsGZPH7EqyLI4Wc58tfjsmPA/7LTp1+hVIWs6tLG0gT
z48ffe9zrBgJi20PjryR9nMMumTE6wdz/V7KenbUp1UGqblyyHH74IuXZNzrxDsSrUgroV+FtRnh
Qb9V//6NIrcLGe47BLz/d6+ZGRuAEHxT5DxxfhxhxtEAX0mEcXxovC9HvH8vB6qczzMf+gtIdZhq
DYXFnvC/dvpVzWKMQgSHI8DwlW2AIth3Op0zPzI/dUL5DoUzTy5ExwjM0qeDNEPnUb9QCVqEzCIs
zU1y6hgH6aPUGUp5LP3dGMZPjga+wH9u5hbM11LJ8Wsqkd4vxakCDo9tGwbX7Tb6DSQ7l/Vyo16g
g7F42lJcxpGbS/bVOMMoDfc6mMDnoQzD+zXdGPL3QB/ItsvSfB/zLIuFFa85NBFnDCOi4hbZNJNC
dbjY1P1A0Esgisi/Ac/hU3CjWR8UddvYHfn53r3JIq9etWO81vZJMitczFlwihSsm9exJoDvOFGf
/phrKNkaSZzeeSpCJJkVnuvfT6ItpRbCFw+SuqMpCujYkhBTG3x7r/CzOIq5YCZtp1WghKRM+CxH
273zRk1qzGw8K7jdBbSdsTBUfFC4TpxtiPl+VmuAtr3WFVH82AR0d1d4sXe8ff1F9aQLv73fF/0O
cIoj1WaFPi/pt+6oILusE5+2mwmrcBf4Judn2qrcJvNYX/zeJvdQFfRsNPULzK0aHGvMFFLlBc7p
5C+SC6GmynQKd+OM6pdRPnhlaf0AKJnOZrB8LxyWeTfQ8WcSd+qKMyo1FT6a/noVuByv1QI8nL6c
qIBdMbuSCMKN7VfKiQlHih5R2RdRH44Hknr6KCcu/4h+P3qNrZt0LAF2lj6mtQCEpeJrQBP7X7es
b/pf1to0VMvUGWRqvPnJu90YQrX1oOU3lirvGpzPDR94KKYA27lBk3B62UvfO02QSrCeQwquaFuD
x0IHNuLGbG9WODSD4wUVab5a9CVMALEAmE72GkEITgz5wCd69pF3AOLCrSUbW4KL/Qus5il1D2Ai
rlIYfLeVA4AYIbJUV49Q600utfQN8taEtojLYAt0zVo3mgmpX4dQHAWT3pn3AGkHsjjTC+LfFMt4
WAznfI5WEg37WxT+XSqWDGRSAzl4ftZ0e7PktMfayQPbou1KIsMRhI3TSoaOFg/+GXhkNg0+SL9t
JNbvtgS7BDQiVeUKTSiBBDMuRUSmZ6fPJt8HBZW81YIFkfOqnmNqxymecl4uixnI9EHUTdGz+89L
GKc5N9doqyhrHw4fXncnVig5seeKKDXGUq+dmCuZeK2wGC1X7DgPW02NGRNPnA8hlDt81H5mWbqt
O3+LKYlsBzC1FCu9DvlfGUvd75oYD4wXxYcB8fmO6ODRDWPJYVgDaAacSTaFscFAhFYvaqBf1ikP
R65nVHDrWtPWv2g8CIHauw7cKrxZcDBA2Fq5IExk2fHI8nQb4mcYhbfRr9z1CXj668ubF+p6SAfl
rh58H3KjHm8hdAOXyY28MnKBXuSTZtk0WBk6KJiZXSNDN35/IeqPQerq/NFdUUUNYtbzWyTwH8he
uCBnrsZ+QLcR8eb/PEagY5Yve4VkCCM8BIa8ZfC+D9SYUNIW9qCj/5PukbC1+aIQVa1qLSC40eYh
w3JeMV4L+Wl+RMPRJD2V/Q9r//BZDggV1L3/vCIwdXLyybriyU8JL9NJgBAkT8aoMS78PV7knMCC
ugC36dcNzZ1xn18mA73JyCEySuAk2I+Qh4L7fhFe4CI4c1wu3hOxPOfr5T/Tw6EMYF+AU+VQYQ2d
55R90mcVycHQ8PyiQvmeo+E7ZRUsoaEMcJkPiOz/c8HHAsYxjcClJ4Q8sfxKQH9CW091wpU+Ycc9
vih1xk8Uoy/cpc8ZNJ8nRZzzs8VQEMcoy9stHCUWzMmXRjjCVuxzMw6F1KPdduZHvjQ6yYgE7Rhg
Hvmp+697i/jYgiUElVOC0kpCyavY8BFQSTPRyWwsT8Eoz+Wt2nJXMcPHi/XIUacYkTbBHR2K7b/R
ZUJvlqaw7qmyVFoU1auJKy0vUXcbgWc6RvInhRJZdBz0PVZqFEuvKMUOiPnqxxA7mJKiQc1wSsKm
Uruac0X9+dQIUJ7toMsWYIdYrnWyNbCqtgrW5LwK9xv363ZqfHFet9tCcgYve9IaIO+A6KHZSEWz
Z57QLQ72RBNpe0nr1cJu18Ors/Lv8xubpJhU55cal2GPQoqHQe8lLhYYr6YCJZpDn6RJRfV9aq5K
J/walQ7k43iG5krl6+XfBbILJZViyf56L1/pQLgG8GAwHE+TWRWH/0DsKnnLYWJZKZO/3PFYqVxE
cTzqhNG3FrBqVyfn3duXpdsNB2oYoQu8W0cU2hz6jUzK7VUGWN5RTFUQ44oI7aMuiJEjofUtcfUr
lyCvzchMx76GuLDjDOvtbf6Z7dc+meeXFAkBuKOKQDnFe9dN/NPrZDzTN1B5j2Eazlo3xZiNH3QP
CD96MDmMYaDORLjBBXbGZ49mD2+IpxGPpeDb9llriSJSRvpEdGwvo8QpVMJKBn4cR8sHQfLiPSsG
VElXf2zeSwjF2070cH+OenHrbUVnR3+pNMZENz2LoDDrgQZIlxd/2ibrc4LzBzHg+NBXjPOfr5NW
/8L8Lcb6qeoAVABwJfKp1LQqtzATdiGAxz75lb5wLvt7JqKhDkD68ZHd1A6HWK5bWtW/luOvY1/L
nwN5gfh9HcQr3Ov028GU5q+5dT8s4+edmLXFu5Ak1c0lYsdBiIpuxDOgcWUDXlg3AIEXppdJ4PKV
Ij+s+6ORnZCeRfGzEdsu1rCwVhtTX+b+XlmJmF4sPn9ZpAydAMHEYP4frLj72KzHB7gim9uZQSf5
TyjVKyJ5uO6BBP1dPLr1B32fF/+INXs1tvnirbt4omu97aaDR7odro5k/vm0Q3xxxnQwkCbd3dbN
81dhocJ1pOkF8YM8s3RAdN3E/YqKclHK1jrHYoeT1tsxxy0cznhPF6G6q36W6t7jOBwQMtPDpcT9
QIfmZ5w4W/rApE57lJasjr06BdYx36uEj42fH53hR5bVDxYE7r5vF/ojCvIMl08bEmzMFYG5c6qi
Zg5ZcZ2NHF/JA2s1dDk9YibN4VDYa5QbA8CJ6RGwCEaP7hdidTMPH4U6belm1RNFWBwTz6BDbIke
NOa6Y5l14d1l9OcTJ51aiISiFUKaE4XhEtWrt/RGXtbHJZyfAXYl7/GHYkqaRgMJ/k9qsYexaueO
a0Jmd+DHpQCzF9uZzSIZBof+2uHS1NaOQP4errf69WOZ1217LjqUDCSbyjRf42naWL6uMXJmw3af
2P2ZBeh2d3b3Y/xpyWT4sURG1bm04k2Pvj/VONszX/LCTtYyy0lrbTighSCa3sZNi3cgF82UvCx2
sfRk3JeqFKtkzcUaUTbrpvPqiOrrqhO8PbPwb0NbBG6UigvraVHu6r8PKLs0sIrCinTRVP4j543u
6FcUUNgvwcM0Y1+r5wycDuYueY/axDCgfJs1Y1XkXj4r6MouAZF6YXAjVA3DOKGa9QkNX+Ky0NyS
cwLxbjrAg9OBqVJPWbhAAbBmCi32RcCZwr9FwQ5DB2IKsnQLSrTzqZOyCY81LgG5I1v0sx/w80yg
f/IUmNSO+cgUuV+4VhSum0sU7TCkem9ev6Zdiy1eesjnGVNEtH0ZsXBwgRGuQ1xrw79fOxeqpL6Y
91GCWBZLuFP+CFGXEEgxmZ9QlvR1vtVWeyaMbGDo75nROIvi0ulc6B9854Tu3Gfvu+4YoWZBJa9J
HubSZti1OmtF934P5EoY4dgfe5sIxDqSLu10kA7sBclGkMbKG+8hTGneRU0bed50aD9trvj6y02c
qEiuasNviNPtbJF1ZoS4nIIGN2viLXkprp1rbJ1kvC3Q99f92zBSNIcmtF+0jh20TsLHM8MnJh0O
NIh7ci9t3jHhMWsdPl+J5ZyBoArDeLYKJtvZwGcDaJsBvH1w7NaPEJ9SJ2mb4kaMwb0WQgEM0MMk
/JO3F26+Xl3Ox9iTo4181ADSzZKoqktbAtJBBND5u2wRHS3VFowjBvtnxEZG4c6d5Rti2XhwYHYJ
DdH8RoX6fg8scimybiTiKib56fDh6NcBMAZhLBLJRo7ZRcYjIDoNTzs9Lxl+DPYXsdZbEfNpyxxu
epicaRlq+va48lV+SbQ/2ZEY9sNZBMWSraS24kStnCxsROD2ksV6T57j1UVZMsKGdPIH9YaIcgT0
9wYH1XD4i0PblCVAZxi4YgNWG7xr1bJRGqcGFJhW+I22pxRDcolj5E5hQ43jWLD0SABWfnsJIBkK
wrWOwHT31b10t1Ds8FR7EpahdnZgcRFyqI6gKEFz12q0j8VaxgjYawmKeJObNc9p9ZBEzsdBeZkg
T8Rx0pPY6HrdEYPjgQfbHXknvj3K6q9SD56hIEc7tnB0opDg7SqRHTS8VpGZctlmnO1c3shjmltg
IqZ+SxSCpgw6NonwnyE0iw3/gsKPhKVdQ7CHiHqLfYvOBVrjIc8x/k1bhJKU3mpyyVW/it5nGXwi
hhoUDD3WQWqCa1HCMQlnvMhUZFqQVVLo/pzbpEOviwubs7BQmd4iW7HLtm8D0wBq2oyI/iSH0uWI
HlNCdcu/PMaMTnXXnsdjvzKDoItqq7ZDfZIV5KUKuR5fI5vNLceqVEBcUfkV0P5IyFe9vzgVYUor
PvecJCLle8pv3+xcLm7n/vk8MHnaTBBb5qiwrI9PyepW6F7iUW14/WMqrjP/Uqxrd7GvMidYbKvq
gAaExjlYLbqoueSalUL/pjj/CFA0E6tHnOFxYEfIqMtN3/TwsVEtUusFZfd30VuO6DVj6Mt2AWLR
FOtO+PC+eXNV0AlWcCif7QgF3ErZ/OEJ3yHuo2NKsVpbSHiHMCX3r4vtZHc01dCh/hgfkDIAcknD
RD//i8gxXvBh8wRMzyzOyEwK1+ZW3Da56KjsjXfNoyOC8DzgKH536SUAWeF3wzR5lV/7o57O4U48
kOz9vnbhZWdQmsOGoUnWpCVb6LtadsbbLo/kTky1ZVBLN/ptZI3gM1H2h5JWT1v7UB5YQZfHHl1C
RrwQY3Vl/FT6sDDPlgw3GsGwrs1uoNaMZ6Nss6HlHHYksAJh1q9qs+yWKjYTLV64QAaM2aij7vMf
UNQsMuSqx1wMnz6yLvX0hMSSMD6laS9nLvzDL5kNUa42xcnkLKjGRL9vPS35AniFH1p3RDO0kw9g
+GeY+NS23UHs8ELYruLADJTyqRfaDllrD984t+rJZ+qUc/K5TQKUxbUgpw3YRL9KOpMP4KPBV3xl
R3GYmJJVGTSxQ2eYsmwR4iFPQj2FCY0g2RwvgETcuUCVpRWpDg5PBd3Ohq5Jk5SfWYfKyot08KDN
8YxwYnk/KNMEEetueIRO/R+M6jTFoNSQKFFJwdRFSmucNOS7/JpIDFNJ0zq4hdg4ZTjNM8GNA4Ep
mEZ6SnVMevEEHxKihxLVN2L1C4ACp6Lu5G5gANq0s2XX1RfhNb2KRPAHFfnXKzKRLi5TjKtbHjDh
Gt6BWz5Zxbt3cnLD07Q6C4cCWmT6xrpiiX+d7UiMYf7tmq/YTX8j7FRBnPtaC4u0RE2iTjx70dmq
lLpEg57B/OyWH5Yor8OONLib8cjPBGBXukeOBDI7wbhhkXiXnmFuxnMQQHqKAv/xiMCbIum0+R4L
YoDxl5GyuMkCXODrluN73f8ywTtGlcFahCw0tSAhY3AtwqeUzjbX0DKH6trZx2TrGchCZroJe+3b
30GT5pkYsnx8o1kIROmSptg/m9j0LoIY6wsrnlB5VCYJrMGX+YxEeljToNDoJn0NjV426gnm5HVL
0Rnv0tQflB9yRqW5O5uJPHpQdRQiduIF1eg9CC6sREIx9VSIDkXbkwg3z3Zdp2bqy/9UCkDHc8xz
k/KucqXuIwhw5IbGPMJ+G/+qKS4rNaH25Uo7LrqB0/an9ggKUVOzgQpfBOsUDc7K2lwhAxzkxbuh
vxnhOhmyVqPDbBj1FXBKHxYLc3C6y5ZyFWeQlDOPfvc5QK46nMcQUXnkL1FdRZFj5VkEsrdLMuR6
7OWu6ac7z18oURzQbAqg1Q6pWovpsCfeHGAYguPuBntAYT7PU0IHmRNhALCM6DdNRlKuV+SWARRa
7N3eztQ7aiXlgcwS9pkaiJb7NYx3H2Nyhduxvd+Ck3q3EpEvOAJs5BishI0jwSjYwdlRZFkbQ5/Q
FqW7Ao7I43X77h6CsiZ55idt/y2TOBscU+DPtwxB46P4hAXtI67/Cc+CCdCd1Me75zAndNXKmdPc
fwwCQbswlH/kQoSajDJpKOeOTFeodRhlE6w4Ocj8UWW5+sFfofg+JW/jgYWYI9F+B/D63MIKgaf8
QGezfpDBpDSzSI+C64Y5xOGcEtIubnKODNu9QXFiubkLtyETYWv0mmZYz6Ky7ZCJZ3ITUf7OhBNT
ZkoCRwIHfqjiF+Zclq3x6svMLjw/RqtESX0mIGN3QT4Cy6YML+/X2vcf8Lr0X+WH+hRgn5TBABCp
nLpyJ/0dDDMcwVrcRVhM1Qy5ae0ShrWTZOVamZDYOnH9IErRKzLnqBu3oJ3oVWLWWpJ71HG4veZY
pa4mFaYeQBn38W+KHzkCLE4vQNSFgQ92mrFvO4Qem2XoTMydKe8xvZYSGFGcsxSjUQvc8WFqOKNO
I6E9FsQCgEG28nHEYipDmsE0yb9J8xSbNDouimlwHIv9Cr553tNV6A7H0lDz/Y7mYFQoREWMDefY
peUHhUrS94xjaruFQs3aC80fLZyWlhF0a+HN0VqA5ByS67pIOsRqFkV4exPrkL2ajUKLl+PAtnYD
ka1QY8fCUfNxAzJ3J0VqZHZkwTu6qXoVVoC2kd/RrIcicFhM49wxB3B0levoIAaVeO5YQQPdbL2V
KoNdsytfksq77miP2xM1ssEne6AAjrPzND9d0ZAV9U1zzGX79wwc1nAI9AQOx6iyiRTzWlZED5tu
bZSfChO3CRhpJ+T9FTZnMfe4OQbIhxoK2dAMAYA85ZEU5WlM9qC1/H+dQH5Hs0LqRicNovqXlB5e
W6kQwMtRn12Eug52QXkds8XwcDWqSeY3wp5fTKcaxDD+4PcB/y5HrGQPXxTvYTY85qS4G4mMu5Za
bYytgiAA9nOwGvTEJ4RiGhnB0g1aW8NQQEbmy0jwb5fiZ25Xarg7vMlki3FByhAU1G1qh0Lpali8
poIef61vQZFsydDFyfln9mcc2E3P5Ekr8f2Aa9bHRATk4y/kZ6xrcUknmGcDp4gP7M7i4JK/sqzk
oABYSNeqiZW4I58jYXcDfzajM4/FOCY0TUKxwEMIfTWmnxbaliotBYYvS6+JwR4Wcgm2IHHUTIqN
LLfw8EXb+g17zFixsTkg0g+zsifP2ZXWM+dTF7mnQ+biXPiS25BVyQ8bWBd4zfgvnSYfaWWr7fst
ZnaBvXHeK6PTbpwUCnRc/tejlKBR+Wn8JBVEDxM09UQal19iRtvDkAoNyhsSYaAkfbEjLSg6Cw8J
30VmKXYnEaveMm+9ct1PqReTKJ8Gngt2DSrC6cBPjONqwiBbbZ5u28LbdI9V/pkWYXl5f7oLYYed
McGkCKr9h9LNC1LIYG+vb7o15z36WzvUyX/bYSRTWTE/isoypFHVvTmuhjmEfEvZgjsOGV+4hAeH
zjZ+A1GAEtQ2o7CfVVypFLvmli8MU+iRPdOcW7NxvQAwewH51n8FuqNo0TYx6NbBFRL4ZTgh3KWM
CCLDICMAzUkYG74ppqLaduFom5gt7790MUsN0Q3BHTTX7I+jKd/EPcyTEeUCA6NX3DPBn5iaNatA
2fxESuQdjIhi4zcjXNR/KV4+ImrGX0k53oDH2lMMSrG4R4HJCBVPRwqtYLkulnibGDTlioqdnEI4
6pRxLhdJu+imaz+kuhsJzpxotsNz4qwj2fqXUN0Qebzk7P+rdAsskaaEBYLkJh2j4lilEF7/A3NV
lh+vHmx9HHvAYg5pwx0w1aS5fPSj8cZ//g46ZVNfF+RAY8jTsFGALCdaiTvKgPkqZCL3eIyAbF+T
wZjhoHTGJANIXbRFXnG2wwH/dgs+AdNIkV3DkOOYuuczSmgW6V9rcftbwvTJQVMOYz6m3n7kIoIa
a41pcQkOq1H7RXyTGmIm4TZ1uZwkfzvhyPMwJfDbXWqzLuYNRD4doSqN/aMomTqhDQTZpU1jQbHl
YPfEG306DvPRRu2sp8Ul4EWNL2OI9GcSO+ecLz5a3qztoMm99+y2b71UjknySrDkbW3Fut6ds/2v
xodcrF/8hs40cK8gRL00zyGketRsIKnk5Xm8E8wuriLMumNsxmz7XMlrc+eZ/rc3ZOJsTUk1mRHY
UCiCOS1M9gvTgNc14LnWnMKAMU63Xrg1XVwEq3SGzEaJRkI3btl0P2Bo91YQnelBDTvyg5vvb/DY
YvDdP8AnC2XbuGeuaKhR1F1KPfU0u1J6dhJvuW+RHlsORyXBDW/uuIpH25wcUg1qrX2lurBalB5Z
+ZoTB/3KxfU9djLb463To6s36JYcr3Hn9EddbmgA5ylngK1LPfgDKPiokwa0IjEkObpMEE7vmGSA
f9+NAF4agc4/LC4k3omsJSoDRoq3M3a9aJ12CNNSyP3gKs6Ot9WIputM86c2AWXA0GtNjGJbKmSw
8ZV6t6m/x5hqS58kxyxzeyO2acYaALZnR4cnx6gZVBgeKmiGVSM86vd6kclJOHLV/LwQPfqi4+Gm
criPUhlzeUBnUg6BTJD1WS/E5+yYvGiec0SJOcZPwsrIZv9Y39m3ZOgiXYwiw8wjuz4B1VdqflVt
amAk/xcP9txXoAqicPPRlXknocQBD5q5UlVelrGBZuIr5Ybx8pwdS8I3g04LgxxLoFGpnvozCCRH
+wz2m6fJlzEvxdUocPpxpIPbCKJ/o1ZtGXmgZTXwDCFTRbGEJFkW/Tw5bYf89KfIUbyuQkfCIYpn
VO+T91JrP/xNBl1fuPyGUf69OHV/+SOT6/ykDUn3rt/PeE5R5EznMIkQBRO0tujd4+bv6MjiBB+o
E+dItY+ZUoabLVdbt4l46r6/lQOSoxKUT7dlwGWJD/6dctCzFwulxFX1VHtAr9hbGRPDwELUq5a/
oLrfF18OvV2bfkjXymtSUFo5POmwmxGsFtefc2xNTCIvrJb8RoVhmqZIZG1ylKYRMbMa8hkc7tWS
pT89oLI/5CA57DSbR2PlEJc/HVymMwBGe9v1GgwjXbaqYN6UN564+s16hkTXbh61O6g5x8MZU2xj
chR/WCQO6hrpMdpsQpPBL0bpo+xXjxFu0H6EVZbZwn9nXY45UDDitF6GLL2fjYcM2T4yNGDXJOFx
yY2Y41yMyql0+zaiffqh4DrD8gq5+QyZDWGOO/432MlbUTpbDy+nyMgGmBpiOsiUIPTU0hGomPEC
U+kqhpjP5vCGMjc80pkzc3k3gkcEj15h0ZjcSHz4Zwu2IIie130gKwUfSgapzOFHqSFSICcR/3L4
EfMp/5VkaqilE1S2lcU6lifHjXKYkRfXUb1S43Mv56PLpMcDrkDNgbYxsFl3htbw2Bq3yF3BjB7c
XNQcBIQWeu7CCDvqRtlFt7mOcyiWHoe9H2j34tno4A+3+WSAgdD7Y2yzHeEnLJxstyC1CUt9Ct2C
t/h7NqxCNquXeEIVtaNS/9DtpQL3LS8ahxP8PQyyBUyAVUdlDPzuFWExldIHbPwfJ5svvfc3NArL
SfNtVwNyILSoPtt0Fg53AIx2uH4GSFaUddhKFX08EbF2LkQRm5JFHQ54X/iDg8Uc06HFJkYPArHW
HIw6jjTND7c3gK1sxCXxO7Oqt91H9Ugr/TeLChM1B0GPnuPbD75YN1P+P/bv/dFcQ4X15g29Iho8
bl3wVLe0I4phm4RyBHAl2Cy09HcDk7sBoM4MYkvpW9ZFjx9ogg8wXoQ/tn8soj1dIfN2bys9vzm1
7qp7GBuiHCyKsApi0zmZyY91GhVCmzHi7ZbBaDc6gvi1z9OcchEzbecox7cbf4Mi3yDI7MG6HDtg
7w43RtvlQuQYJogXoAJUME0q4IgHVft+chVmnACWdZXrTRx6QYDvZBQA2fYX3g0cdPHpMzzu4yVz
8WbEeqAQ9Q4HGAtf+9dYJvc/QAgIcsw4hxmCZXMkXW7IvS9AS534ji2pqk0uY6JfBwsVHcu0bS1C
W499On/88+xx2r0QFGbcWqIYmkmfn23v0u4RPheedV3AQqVSEh3ehlTPGPtNlLA3mOsFd+gafikY
J5F98Z7B1lAsm1KCxzvXYabyqpqjMtXg1mr4E+1ir5HrZDi/rZtOOna/blVUYPIjd83lm+o4+KeL
b/DEkOxuyxO4vgpWbjpNGm+aYE+uuSHlSFJYVHxUtdCt3Dak2ubBBRvcoc/VmX1NxhIaibLHh8LS
jyzZTtELdPWfudKZueD/j08I7HBetSO4i44d611+LsMLaabeIleShoBzCCtfoXqbcJf7sx9uD14S
Qe0Yx8HmbkEPZd7cTGtLXAqCUmczrD8zET5qV98Bc9YWfmUcMKZ8jf2+nd/q2T9IYE9B6HGXH+SH
a9jgwEu8khT/vh0EzSf7RYnlSsxj+Kup8VUZvIFKEj5XRVrSHyk2hIhQm8L79PDtDz7rBLTiVnsv
J68vuxrS253cTqZSWSdpuLzCmMHO09Nquq6E+r55yssoK7Y6JBenx+mudil5PPEv8LTbNN3ZN+OM
3qva8dSuBsRnwW0hun1A2Mjs938hmsB2OT9ad8gfhA7E5R/XX99w0VOZbU6wfP3yIejtSs8M8Er8
QsCwPyr3X88q2Zq9sMyNMGZan1z7eXfDCKvLUl9v5lTCyZW8DVcazEXlT9BMbOQJmOJoN2HQQZn7
ORpSvdRgzU+uPOyhlyk4z4if3O3J4zUggYvCDv4s/lbG77zAxjugxuyCu3b71s3XcngjuO9n8PR7
K8zyD4hIgTPaxLh3HDjbw4kzTYssC5AB2VkXEmJ3Mb8sF43FLnx3q8GnY8Hxnwpj3vtbFf2ZjkSp
IERu6ffdcvVBUH7nbgnH97YglK5GjST4rfjOkouwXe0pZDADP3bZWuOQ8U+6jail77/xcehhg6JX
vAMdrTAVP7RYpJO30Vlzjp8T5sV5XtPQp3AJYiw6qDyfoXjBS5ZWe2qhQ3rUK3eljgWCHwF8zZz7
pMEK8mpi4ZlbRafnRW7dj9omTKFxpgWyqVertNjHstbL3SIsDDiyhbo5YhjzhiIgPuTeSgTllwAg
JLKUKx0xo+sJfDR40+XDp2nhvaBazrJ/75ZHametv8siWjgmT1MennW7S7PMD6ZRriDDKPopE2Cw
NMiECgdP2lnxzP40UHfF+AYMbKibHr+PhsH+heMPrjGzjWQop5RxE7YVpglqXEhi2JXUdffjmPgZ
QyZjK+xd3r5f3SJ8KHc4JidreYQAOxKIZMU+7PNkp05X9fE+ev8ChIovYiDw5UBibFhIMhmw1m04
UCXjMKFaUKBSYY2zESiykdaXU5KJ2gX153wbTmFuTVnwKK/7aqFN1Lhdef1VhwrmOamz+zGpBYdO
19KIO1sbyhiTBh0WudKRkfCG+Erv+eZ5TBosoOu6y00Q2xJHCQJ2d7uUrJ7v6cwV4HR0ciZdpSLP
NgXSY+w2LUBPJzZmfBR5jNfKVSjjwBwcLCyc7j2n7WSw0a8XQeVEfXYF1zU5S/S++BK1Gt5G69V7
OnvUnRE8ktsa+jZ59rVFSqD/tED+y4a245THboGJFofNomp4BRyZl/676bq68uPgQTiavKl57g9/
uZm4UqFKF6n2K221HV/n6ZmTR9/FoJTW6WEX4/QYLE5nO+EZTJwFrtT65Yv7CXkKeRJnlYwQn1ya
geg6NKNy5xxRFQPCq2Rga1dWl57UozWquHZzw6FydevD5Z+i+uoCWXPWybD2pYn1/2+EdRbp9j+S
Wy/McETY2QNB5vSm1cmaEgtrjivqDLACoJGi8wVbt8e2AhVBke5Eydqc/D8VbFe/dGJxUEjbiaOP
9IuggiUL2EcdJvOd7u9jyVIeeLtk94wUTdYtd70bdZc06Mfq/4Ta7KZATgYLIKwGlSYZf/OdRvm+
EZtVP/XRbzedYxa/2HGBUzWSOh6IjcWOPt+j8JVlsXgjk0Hm3PV6zoWIymMv9hlOo/l47MietDKq
3OLb8jSAiqCpbfWNugfwMmGf/0S8S7lAumpynU2OfddsxjALfxDyxgHrCWx5pfUWW7hJo3jKpIUJ
qZgtpn7JLOYcFmGuI63t0HjD3Us8kn8z2szXUKh6fFSqyLAYn/q+a5GbrGhvFT0qYWT6dDRSyvOm
LKCBeG2HvyyHPB2II28OSjcLz2Ne1nsEsjX2xNjMdX4BKxGj/y3yMhk3NEg+tjHUA0ZFUuCBEme3
F6qgZ3DUX0EVBeCM7hTKTTCIUeY1Xld8P5/mIY3pS3pnfXNSzJ7/Lv7qMzHyhi4kuaYE+xoGoAuT
lZrqQ7ludsh4NvXgKvzesa2zaYY4HbTlx8KKER0Xv728UwjAFPxA3mIe2HccyfWNn+t07+wgogXJ
Yu2cZbjFnYZkhj6IRCe7ceNASPuo+kIf/Mjw4/YuVQuqcVgg/Dqy2e2zX9VyZT5nd5wSDBQf8kd3
0s2U5XPNgHzdTPri9i7pBvYvfwBVazZ306XkAvhBBFprbCct8l36wKQ5V1bPipAo9Cj9mePO8pRU
lyzs/5cO6ZC01N/cKFkmcTmsaAkpKURl6ySK+Np6tU7n2V9Q5Ob/b1Ux8tongePsyTGWm/FsgfRi
AdQOCr27eD93uAG2JQpzHL4xEaZMQyTn/fQEfyTo0/JPfd/gsZX0hjqmsQkd+QDaoi7Fb9qUlEnD
eksL35ii4rhxAu5N7bx5R6sUYIoyz+nd+eYsAS1sZrYogtBu3idn4Chifz69vEQqFyClxL/8zh9m
yoZUboT5lBKsvQTG/wEVVRYxPMDjVq3xu1RsSCY7oGEmxvK5Q9mr5BMfPQDnskhGAvPeefaUI+oO
hbzfMZd/77uszXW632L3ONKz36dOnFChKFuqGBglDZlWU3PW/E/u9Ya6kGmtcYTsw+LVZfN54Xyj
4cVk0Etpo9xGmIRK3NQ4NOLSiP/9UudENx7DC9hRBWBjOfaj5iPsTm7hOCv2Yiyw8BRrwlwlssXe
hvW7GrR9jLB4HR9ZIfb8JBlLSck4Zzw2z86YhiQHVTlOaC65aXWazvu+rKeaURVXbsHZQgz16LI1
18oCNHo2m/+J+cHtIPLTys4aCvqH6gzwxalcM7Uwg0P0oceX5vFYNFXos8sph/DgRb5AwLcXv7Es
Mtaqj/RWRPKwr6O4YbwIi3qlU4nTzINA8kZJE8PeGYO77OJE1SNYAvD3rzuZBQlJliQT0OzSqBzM
etQFRSlFZloVmjGc0KuySLvaxWDywWE5IDZqa9VyZsVJfPBUAqY8s428aAFtDEslCy6ZBmGY2v7y
zKcIzbQoihVoqmyHRoQfUrXO3IwL5o7jX6f8drlVQERdx5heGraqfiracz+lnk41HzRpjGGmm+VH
cB9xLK95hh9nN0LrOA58yjj8fHb0juqu8f41/Jr9vSMMA+kNH08n3TRFfsz0d3VL3a1r7QpSs7gb
fCktQmVJDlVvrUd5wnjrwGS1q8LANl37PQ3HmLXNm7fxzTjubKB7bjhk4gZzkhBsSNKrtgQUmG99
2apGoE61WV9834AeiFU4RMI=
`protect end_protected
