`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kurRNsF/116/axtOvoikRx/B50modjP/EHmNfOYGMpX+1T47YinGbf3YUT1nQFyymGmFynazP6qg
CZKl6AqmEQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WC4npYuXDJf/7SghrKfefbXRWo2QbJraNzzR1mDcY4EmV3b00/FHWB5tJVoLfpIQVgdYHsGkneiK
iuolgBV2SCOnO4ViPg0tJBdogfYOBUSAQ3fuRuIcZB8ie/IQn4+PrXgtd3PVZSFJ9OjZ02bKnWK8
6KR6OZ4kolCEhNzqw+c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ckNs4qLJXHxsAWqs2aUVePAFGh4NIGEIUNu1IWWZPPva5K3fmHahWF+9AOkjQeYsX2G5Wts8vHVj
9fyH9byLMWz+7ep3K9NBBybAJtUuWdiiQT0Eu4Rer9zRswlM1RF6b7zejliX9HqpUdKTtnTEEFkQ
dT8RxpcD1iDZIY1eInKQ3Z4vrj9cdvZZllWQ3aySbQqc4F813rLmgdN6SO2LETSz8lFBqKOqB56O
6DIn+DhP3iJI3ToksXrgfbhOoIRmzk8Voh2ApVePG9HTXoIFWB/A7JbLJQtv9uqUTs+h5FoWXD/r
5dLxU2Kd22z1tAbRg57vC+nNkavx1h1Zla4JUg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mvsZJu4YmUyrhRXG3fTIENvQtQjtW5Gb1qettc9e5Srqr5yrsPEHT61UDlecAKihMgQUi5kbDvt6
3XSKHhfxFQQ/8/tIp9QZHGK0MQ0B10K7p3RRVFcPS0iddElFFFskFDrppASQv+OFfyjG+1rtwSYF
sj4f1rY51rh9dktsS3U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVwROVVgGYHl9rDneuUOMCckhBq3hZSO7On1WKzLGK7iYt+AGTRtSJFu83nVIL+wgkc+cjJz/ZBN
tp0QHhwstS1UfPcP/22b5qL+o4s3ypDGuJ4DvR+HcP4w5M7I5v8lqBp6V0Vx1ueuV3eT4aM7NCuD
/wtNDGZBs1O0dw1Ak92BqYs/IMgygaKmpWvv+io6etTmh6JihpscojfYOcPBmDYm38HgMfqCO8Fo
ENG8a6NBYPmjUNmmYpHh34ZbvuAVqZvTBszFiWOinF8dJbYaR6jzGLPWL2k4iW6fGwgs8IgioVbY
hU4FHyqXvarcxIRx2n2qSbzMbr+iBbxEPJJ3mA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
+0aNGQMeMJXIrgz0P3us7qk/wiFv7jfj25dninB8MI7dGYjeYmvAZRUvzp3MV10CO8FSN8LxQxfz
cilwrbnUwbi93zwme7kDRXFkDnmNIDuvfv1RSjbr2wLzJEt9VKqt/wJ2xG2/8cZr8h39Bf9DeV/z
MyubPfQ4gyLYOReYTjBZupZCrmU9BArP19xbwrR6/gaTjBlwOThR1dbiql2oa+5FMa3NVyY3VDke
fTXn9XaO+TS4Gx5qziVNUJdfLWmmHCHR+ISvCNOPGC6+pt6HJRWE2ZzSFoFv5gj4oFMXJon5Xj4i
Lp+b3L+rkctL3veTtuEePeXAeWdjPt+D3vQ6lVQ+IRvvx1V5S1qnx7uMj8dvHyT/DtV0qqhi8rP7
vWMVhH77tx6HCeITU11bRyHsftVBLFlxh8JUaftflYNvoOzKTfQbiiUREAsEZuiD8fvRwUqyIW4W
KQOocL5rJPyets968sieHHwacTwfko0E0vPlaPa2s84A9pap/tYJ/3H0lh2CSzCg1bdjXU6KGpIt
+/Bfqw+aFTjVKMuBV+buCFzJS/viT3a8aZ/uCdryucPIalSdDWaAY0InnI323R87weTj18gIrkzO
yKu3uNnHaQV7pJEK/qNvYix/+VzHX8riJyyEjuq3pXxCbcVJll65ia9Wx2pb/FOIbP57sAfrBMAz
17CZjVeTHgAvwDWLYqY+eP74mIwt+tKBZsirVYkCZIBn2HvqZ4l/3AbTeUddxpVRC3+JgetW3FcD
qZKAVAdpvKbUcIPwOYHUO8t5Wx1YQKuQSGVRt6l1NVuOp5434v19HL+gR9haab5G2kLleHqLfNjS
fJLC2A6+SiKUWaQcqSKquWkMwR/x0NBSz7b/t2r6HwOE5W1B+sWDot0OeQQWvhHLdMLvm4MN9K9t
F9zEfvl8cdH0oPo7q7eY/26Q+7ngSEHS0GxJBHsj+kdcBzIA/RVrb7OVcdisdThZC/9XsSr0Yqtm
rMag29dqzHfggKOLBEbx9ntOS/3AbIPy6pKo/EQzB3UQDX0OyWnp/LCwQXlPTP1lNJxlC9yNILFC
VqjLSOhm2Dt/21xLLgQCIGT261JRSSKYutvsVSPs9Q/umZI6sRiV5bR8+C151wCSwN49Cj8CVYtn
ynUWOaEcQYuRl4hAPezqFjDYEWexvA13x+mvLUZXdPFzsoTA7TqUorRmaqAnLd1Le3Nqdx3TlGu+
uD/pGHtkZhHFCwM7yaAnFQG5ia5JrDSFq2F2H3LkDeNgkum/yAyg35hbQkmGdMXOWtyXHf5bxmny
Svxvl09IgvZS1MmGfrXJpy+wROJx6ct4xiPSbncmC0AF263SlX32ZVBVaOFa0iUq8OfOvYOvcEBs
eIvLKM4RYxh7AigJ7YsmZm8PDqrdSeKLCxMyBMNwJ5+cT1HoMcPWeURpWEhr2Z+RWjrRDTohVvrV
K0x1q0iD1gCd0cdqOGR9zMfrqOtfCKsAIhgc+UG+QUyAj+aaFKOjFybVRc/M1TctTVpsR5CDClKN
tv7ozXsVvKkb2a10RAxvYRuoPJ2eli02uFJglxXZtGpc+yINuynoZl+/AA/MNqmrHTMkGCHr/SXK
RUF6qLyAlr6o3FpnpyaKEALVY7sysLLLc8vOfu1oTZ2Cg87LFXIiE1zNMLOgieooKrFKPr3w/Tcd
9ORtyK6RQ5vQdY10u/xvuY+LtC2vAqO2AYhYc75u0+cf3SZNfGU91KvW9XznibtA/qvmFsajRERG
8+pEd3XrcAEl8+9eiBGUhd3JlJRtbqkVShG1cWIwjCrea+j9Q24Z7lWl1JzRh166HRm3tB2nL0Ws
9pQ2o0LNrT5l6scu6/E6aSrdKysbWhO2hFVWzWiUlKLTH9UtMUkjyMESL/hgIKRuiU/9n76t0/BI
RS0Thx+fs/MpH+dZz0N9CYpBCs3ZVoCKaY5VbVjwKqqSt3Vfu/8ucpLSCknHu1Tj+xRK4GR7A3ZC
0T++YBjJzk9fWZy/no10k7Ez26HGPAmgkiDdXVEWAW/yDhtEOZ04REO1Mw54uNgL+FH/FPqqYxN2
GaUITbutuJizWaqkLCn3gxCAG6f3tam0ujLLV/p7zfInDjYsKpFXyVKEbtZ4Jcwi2+xJlaIvBD1b
QixFhxpt7spDo2Ku8mylhhMl4RUzoRllifjPC7Ua0XIdWfNHqMtewOWWPS+byMpwjMSfcxqUAu1L
z+hPj7xp9NyuEjF7c25xzh3a5rxsQtme+f8mSNPXUS91u1l7O0K+I2EPH6ulBX0bJsg96/qu9nTI
wT1SZJpaWAY8qgJeeb3IK9imz/tpm3mXjs0ZCSFk0Srq7k3i+kEhlyAVcypOa+kZq1lWxfRbgVCs
9xr4160x/7pZxiyaZxuWl70UqxQTxj1YvAcgyZthDMWYeDmBqLcj6/4iOJ8bbgqqzmxzcRPN4Fxg
jAM71PpoPEMJ6ht3WKgzxAVHzlCOTVka8C5HHhDY0CkZUynk3ahTSDna4DW3O/zllt8UCogDbPs0
Ic7nysHgYufKU77dbY11m93sBeytcPghri5kB7ejWT5FGLtvcz+NwGvGiM66c1gE+7bZEZv8xsG3
ItO5nk+EMygE7+c2I84Wvx26s69fBdDmK9Tz2UzeoG9ZVUNxCxWhI0L5AfPocTjqCOWOJnyy54uV
8EjNkvGxhvdZdTUizMsuQwa0LwU1aoM7VWlCdqs5Ma1/RSrKsgXUfTMF1gZFlzhLVl58vI+UIiOy
O1aYgfuKH4WJNIzFWaAUSwW4CxLuUUu/9ltBMh6kt//rbmb2dIiE9vIAe7bh/9tvhMstohGoun8l
3GvX01JcYwsZLOl/bJ+rtYNjU0LTcSogvlYTKm25VDoguk9P0/btBwRSvulCEIPrS+TRlRn+AzaL
MvHSyyfuWWKarNQiKbNFj4+18QG2EQUDX9shus/Q6bcqUlnBH6UNChCcoA5KwOlmdKFiETQwywt/
brAi2wMhSJ/iJwDHu6AzdrhCpvmrFU308k5qj9xdYybWk3no9DrKz30pjl9Epo9yHI7cCftnDXbG
MNRfCtrmjGRwyc3F/tRCwsfs1VJJK/H4SAd5wAGcWBNOd+rAAp1E/MyBXwPaAoaOfRhZrStTGWeK
x2Z39zTMXklZhw+BGUtQqXCu9XeTr5Ti5g+9QQ2V6NxiDaBz6AXdl7LE0+vy0TiPHX8xdBT4oSu2
9buxJ10Mb+ynUYZTnI3/nZ+8k7eskP76Qj7U4NbEk5XnRwQ4zXK2IKyrzXSMIPUN80lZa042/E6E
t6ddpfCWvVlcyx8PQbjp+2kbnGNDr/AO9kUqXpgG0MhjTQerGHbAoB/qJ6mpb99U/LwBv9GIxUxR
Rn5yQPJMY+SkUNkuqdubyJRhkqFa7pfys/YtRH+SOMdaw+xWTo8I2bsIvybY2MjKjHag0s9zw5bT
KyVd5sxgpEK741dl/a41aqCUZ8xN1ccgypzLWys19IbMzlQ+t8+QT6ocpuTH+TH6VXGD0dIF4y+V
CfwM1Vpxy3w8abol0k0fyu4EfglZRfITSo5WugYGLt9vrBt1vWzL7d5mvIR14ClLeP8Tt5/izuqM
iUja/ewzpYODDdRJt1Y/wwt4WkRrus+GPq7D2BFNs2lNkMQ1bRIJmY4y/ct1tEGgyM9NkN9NTokh
pnmeRdfXWA/Zqg+oAhyxGziktyf/1Zt+USu0a6CMfHawP9WPRPp3oS81+j1AntzxsXoVQyza2JqD
NMqpcF1zONjBVasb2yOr0eAF6fyYtYofBn92nAJLLDBm1CV6QygJQK3Ze0Xlp32uhPBc/OeJSFYY
y97UJ/20lNYK0pvVtBKcLySCoUnEvi6NfsSIIV4uI+xIJv09kjtJPn5HAMJ6T4zsLSHBLDxTbHRQ
5XoFVQoGJiKKwiR7uLneayXGj7pf0x2nGFrLbnaBeR+54bbNOMZrSIQA36GRkqze1CCOc8P3tjuU
8UnfymcgWbI6NcdCPI8CefjXZtssdKQT8oLDEatDMf8Snk0Fd4U3PAalP4XLQK22/lVqTQFfjbg/
c33KPu3WSGfN7kzNJPZJgWYzKvbqe20a67PhA4G6q7GkJby6JcI7T6dEpyLCqH/M2Ve+aE3308mc
2bW1td6jxb/h2c0MCEsDeMxldZJObC4cl2Xk7l8ddMsrPuc3fNsBjDO7p29El8Dt4XHIwA2U806B
PQh0F+QDSwMR1W4tU5llceWgLlALqFBcHkZ1oVRSR5E6XP9HRo8/fVSSjo7FGwMQdVM/N2OGGxRu
JvWOMlaJgOBCYqBLWBNjwClfFxWYysWBeMcUREdDc0sPGBh852xg/fuqVaYopnxmvg6Nc6Hh2Xf9
qPj0mM6beaDSiArha0XY+kEsicW8Pv9nUOFjMrGkVi8r5N3UZijAFq/AlI0ewh0mRjapzxahYdZ8
sw+yKaAuR+jePLsUUKZM99q1wuHmgLcfghJAQw4tzvX9HdxjNuGsbQQycmZgAt4dPKyIPmh2vG/u
KRIBfMXAUYP0WGPyAVMkHoQ8fxTXJo9d1wYGDVwXebsFrXhnGr7jI2zuN82T6y7ZBoJx7zmlU/MZ
FxwNJv0QXZGKZWcBh2DJHF9gWwCNc7HBRASR8LIuIG/49pg8PFCWA6ORoLnv6QYyZibcZWI/6FL2
/AFm60aT0R5GrWBjFSuXB8x/HD2iyROjkbGGzpZPMtxaX7Y2X9z8oOnFXgozndsOk854yHvvIjRH
WSJO1KRHFVz431pY/p2J7NukE/jiDZqr7iNKJcJR5q906t8BGP5g+iub3mT3QiGknjF3zYBIxSej
ELKwa7UuR+zuyq4bD35olxB1S8CdvjFp36GWHYNE7sL/qMcR+/FhYTERWClRKefVNC0utK9LeGSl
X12PT0WKxq2Kn85ZCPUfTf6fZw3TaidtymYProA2We8/v5KAJVOZPcZyTjH819N63Q4mRFkgwpIf
t2sVWFFe/p7j7W2Yi6gG3nqZS3+OFqB9b0W2oaMyK68JbY6jVoERJJwsA4SVfsKoxTXUTiOu3bFH
r5xo/pJLo7bXomSiFQUhGTpMSPygLV7rnonxoSK6zf+RaBOQKTA/qrGW7KgiN/Hhau4L5QnhQsDk
y//QIsoNqH5K04c9LF5eAlrvNDtDnUInv+NifEjmAbnvIVhMUivmZ7G1XDtq1v8YDV+856iX2Tl5
QPC/XyXmxGFkSUrbMJi9HBV5DlPSEIc31mwS/1KlzO0PXIfQ3iV2djQaGbote9sQy1MzUd7IMAh/
sgNyPLQURW/ps98czCKN4oG1tb9/2RnW//Z56YS3eL6S543rMOAf8Rkpn7FJev0yM9rYbR0kOKSj
0cVUg8XV0Hd6sD4NEzXJkJAiga+1L08csHcI6gBnc50zq9+fApF+qtnO2Oukp9Af9ZEh/L2c6CAz
WAe/Pm8wcr/jhdfvkf2ACWYFbgERniZ3JzA5NrVmS5UHjAeb3dN91+tdEE37B0xe6WpXo4WcDqSu
rigPKb0cS7LF/GEvc4R+1P7N1QN3BO/C6eVWm5HkghftbvBGcSTdLUgeJic0DloODDjrBMQFFwWa
0coCr24WhuwcT1pMQaPgboCZGM2xuw7bTaC+sHx+DW06Mc611Giij7t5HxTAVxv1HCU5ZzN7ycIP
wCs1KbfgGmSEC5EpDLSiyUXAW0G4Vhmr+UEiXw5166jdfFPG7uAAmMHNQDtGDGRDuhU8f8E+sbuI
UtWKnWc1czGBnboDYYpI/tAQtnA3GD3p/zsza0RcjWvDnPdwjJUopeRoKHml62CwqlBg+71Holan
Ld+oQYkx/QfN82NOYnI9o5D0TiOqWSYV+I5fQkBxY7GsZC+nyiFQ5MjvpnOqJ4THx/Xbj9MctRuK
nJeIWAZD88Hqa0DeVnH3yasKKoHxYcMvJaOJNuUaVG0OcoDgNoX02PuKKfe3swC9Sml/wXVNzPjH
MycdlvjdMSd8A7Bme6pea3rq4sQmaFFxp5doWAhr+ud8i4JJurkqpbZar3EYSiaGEf6ac4oDiTlT
nCj7yC3X879PhJs8eBCbjyCn9YV2QAuBjJkp61ybEgCS91JTfuMUnA/nSfoXAGNRmxd52YebtJEN
Kzlm+YRISmmIa3wVSFsMsvmuVp11lzeDosip7pSgajRftr6rEhkXA81VeHaU6iymYrQE0q0oTOgL
55j4jfbGzGJOCw1VAitSbtZ8eOoo7FZE2iHBJzSml8UQRxNHJ3KokhkX1EoJf5i93ahuXZ/KQsgU
m4PI51WinKnoWopoEg60dU/9vRMHJr8ZATMLSaOL3Gz1mtVP9wAUJtgNBYdA4Y5rmZfKa5/HglWR
bruNgQ4UFNp4ZfFWvXlXRVJXVKGodTqoPBjSVEpaMklqPXft1OAVKY2joVhlGn1CZh3ldaBUCrRZ
ZYlmiaVQeBtFvI0haoTY7X4t1y4sDBcKvhvy/PVKBVo8fSdnUEp3JrR+64QQSSMlJyyOIPl+nmUQ
FzrhIoe8NI10xOFi2/X2T18ZfCuZ7a3TeFbiYlordIqn+HJD0VDp4B42F/A84pIH2maYvCr7TIl0
4ASQLVh8VWZGgJPgwvBhrJ/E7O3PACEwLHbQU5H9ZtHNB0xGSms7MDsNqXTRuHzxM00npgsKtid/
TahEQwLcaNNxHgayVumLUMj/HpZIq6lZy7DOW8bKaLD1CyecJX3YV0/JwgTTPuv5TiUXSYdxTDdn
r1s962RxEZLojuozyp8wze7lNm5COXkUFu3CUUSk11BZhgWAAyOADosCYPvbxE14UCkm/3c77oi3
t8/VCnq7qhpkncb1KnoofXp0AKIg8Im4FoCFqEh2fnVA4JzIeUtwMWT6ZYGN253hQsFBiGlXFGqZ
2qPAHmzlRPYwJmLrESHUe4WJqGiwjOLTyN3a5tHHKHFK/8W4LhMzImOKz/3nOYft9Kh9MNAdZ3Zw
r7Fw62PMozH/tegslML9QfiVPebWcCmjxw3r9kvphwmK4inXi4WGVvjm/EPo0XCrhTr0opFbtqLJ
JSed1OwfwuK3Pdx8F0pjXK6V/opLGQWdOEEAkSFo0fV+O/sBRWCxgRrdNkvppzlxrGo7cxcfYyz6
kzt9RkwON0lXXdRhnkR3mFtyBvtCUrv9AHhoyk3sBNh4DHayG8G5plw0SAvVYq3ooDVrAkSBrYNG
p0San1HBaFS5LJS3WLa7rMiDkS5isPhC6AZKUygEcF/crM1/SQMiv72uhHcBGx4Kp38N1OF9kY1s
j5ZkGlq6aNsf3UdjjHLrtklaCxaVMoKvQ78VYGhymYRQYS9arQZSaB1GAHCWHfOpK7+myNHT/Mp6
wDnRqhFdW7xVZTADpyPZ3Hew/TkxJDx5wjaY7upN4ghwQ9IdqK+z+8foEr705k1vhyDg0K37+KiU
2/XcTELv3lxZkfHjOE520JXHxzrVaPExT07ba69U0AAs6PEO85SKpoE6FTgMlPsZYa1Dbp5L6H5v
nLnD4l2UQQvbDrD2LF7J5PCOfaRCLLR8I0fblwXg+SbJ5baOOVrEFr1pLC/AoGQDoADx1u/ByCvY
X6FxwNy54IIHcuwiyGBq5Q2gELIT0ACKaUqbQLJ5VpLjtSKtZLaPwlH8Hb9x/cN5PTBls4u8INgv
wMsg0rcrth/a48ff04CjfX1hy/QDrbRWu8F/8H6pMCZvw5dU/e9Y4Trrku+eySC0PBZ20FvqY2aW
js8XEewj5BB2wFI7d8LvWanx5szRwD4fRAcLFSIXcNoJnPHyhaTvq7zVoVBfLsR9joBjfhc+BYZ2
T3guD/U8uzFwq5cw0rkTKuEYf33nFTHLiL3FgN4oxQ6iogD6x1V05Z1k+A60XF7EjcDARKlVKvTR
aRRSSUToxX1z3pWUTcYShKuOjn+CGmG0vr0Wi3LnfP6TuL/EhXjyJjKzN2Kx8PGKwSqGVJjSRgWg
4nqVP92yKpBF0bPedV1STVT+BN5JB8qLIM6dF8E7g+h9ov2OtIg/f5OOUpSBjO4uZk1kaUgAlhKd
jfZE8tHptsPlHsu/13AU3B6W6vXvcQsMUgHNJLf0ctMgMgRFYBvq66WEQhXMtMOpDrT4JWs1aXFN
61uK4URDELFAc/Fve3nEIGQb2biVgbCOE+Ym81JMlpRC8j5H2ghttkmarnPE9XYE0TkQgw9hgQlW
krwL0SAkkD7C/2pM4SNY8jLnQmGIHHLYn21CdR1wZnrB+aLprEX/weccMrNr4Kd3WGFO34sCVNRV
GWaUjxUDVFNU8VnqIvcL2UZCCMNfKgfij9SQlUeuUFeb5P0yGhxeu/0SetMyKusqiOteJOwNch7V
OPVI4UC2+qqVyPu3oAD1gEfosR4NlqfSjpIgRmL4aCeoYxXJ8GfqqSk1zANtOWG0pgFCe1sFekzX
tDvO83287QoCJR0G+vPilOe3U1PFtXSyY0lMnE4Ob9I6QwxWprwYd8iItgGCr3AsVcPtE5/C4PJ5
cpBSV8DoygVpuEmAaO8VwJc+wstK6ji+OC1Bu/CzExFtKwGvG8yRPtTfz68MkRXneWYJrWExIP59
0FbWGcA6Jn28pLnd2eWj+pJk+oOZ2PWrU1hJ/XbbyK7DUBYXmGbIMkqYcd4ZLzX/5ZHmlm1Sfonr
c2QL+0B4QZ+zdJ1k7oCw8wUlx5lmbaP2a5h+Gi9CFYe6a2SGyeFuUdRFFBEVDE6Otb2HpjaWupht
S5iIcWWL6Df/sM8SHSmPR+IiLRD02efdybuMfmJdanNNK3W19ueJtYDBVnd86iQWlK3uRh+5dZgo
17xzYpTMOU4qRopbka6LV1QTOT58TT2jt1Nx016ldTn4KEUm9XCJuNi4m1gyTGinJ8uZOXOGSe3M
ohk6qvlEu+VZ4CEkfNAFfvU6Fkmn17ltNOFS8BsREMQQE5daLS8D7vkOdqr0v7wqVwvjTf/iU/cZ
boq84EWsCcEY2Mng6ocFHAAPbtHLv0TBZFHoYq0QlrB/7ncTxKOaicrrFOTpGuIBkM73cgUQBanD
J8zKg+UUrLuQSwQ7gUuNM1EtHpDAjMAjr/9tsBY3gaX2oZ+W9+DTHFNRrBAVajX9/MTaXh6aN1RX
bLhf18+0nGyA+88XpRNN3iasO5FSJ9D1gcc0na4hBXfDEumXW+Kl3pz14sdvWK3RQDL/2Rkj3dq6
TfbRUVAh8dU3w3SCSpOL7VAyw+ge65k6fxIdX5O7gWKphkRgItjOEDBC/Cona/ru+62aouw6HL8c
XJmSl3RQtJFWVYjWg6qPvmK0AYLi4URK53oF9tkeUT44HvYDslTDkrPHo8K89wJPJxQOi/Ir0Avm
HbkpXSqEWsc9giyEQ4oMlxAgluoybcAicGZmZeo1bLtSfRyzTmobUWmSruYIBVI6c0OM5zdAb0zJ
zPfAawVGHiCC8XIkyCiYPfoe9SniDxsxPcmiXYA9Y46dO5UqcURDfjd/w4VFNBDJ+13ukq8u4RzK
d9CR4Fp66Tp3AhP0BDARrUfJTf27lOYBvwngjUH0jTY/nubiIghcdOD0eAtNa1KBvRV6Jn3okkgb
xTvSOcr2VTAb3uHkasWs9CscqumMOOPr8yUqehQ2Axkj15V3m2BwcTao5GK9B8xbyHeop7rLmtkf
3KS9pnEZHESMLsQ1IOCJtiLAFgB2IRAYm5BztA8hFvjg46ec3AlFnGW4sxqvvUBuMUoOHptUdle6
3Oj1H8uwRDcOoc4kh/+cfSrVADLhgFF63jnyUmSerkrxlxkReugNK3Hrs9cTUzEoEzmYdf/NuMJH
5O6dbJRL3v8DUP0GzQRUo+EgBSCsCzu73X13lBbW7zoIpTiP69J6kyGEY5XD/1BMPEz3k5lVY3me
P4AnkSGgEaQ7HMfo765lkna/dGDsdQE2vvRPzu082lggH1DpIuZI6wVxGo9IugYyRClxWihh5O0G
iVCYs5Dd27IlTXlvQwBnErjc0+EetgIqam4pKrAb78lqvfpoMdICPFY0cmnNmyniXN1B+QOF8OrX
hh7lZaUYr702h+mMaEiT3cN6mIRNLr+uYiu0jeNnfXBUYWpSIORPBTSt8zMUaymQf+MMYgdJDNZH
qAldq2t39S2mu5wPA8S4w8S2C4rXlW1czg7INYDGpdcd/7NOf1GPe6YZKT7AXYBHmzNyg+jkOPqr
iEKCSp844zjj0CJVkzycz838hRmUQ5aykbgQtCh2NGTg6VzLAxEKGoNZttblgyNofk3rAnDEkLAu
v+MdvUH0i1Uu8yGWxaleW6Qd94UKMTPci2thUVbWVhwXEXWzTjdqUMK2eq9cEf/agrPLJIMdm5ti
1wE1IkwX6Z7RB/PoomSJnK29219U2U8rAMJrLInJWDvZ67X697CPlIv6ydIH4/QFqWBb3aQO8xpy
V2rZRKzk37x2V+V6cj0WrTxy6rRHkVWpFSH0dviPYvTC7OqRcg1wV0NSCckmF5c3Gtv1V22T46Vl
mNITPVBd9W7sEv16u9spMJIr6ZTQ9h3eZcEUSu80/dVlAq0dPOhnr8g0deoDDxUIEVhUZIDt0nKl
Jo1u9nWeWr/EPZ85VhyXPXZKbBPfIfNW/brAnLAtte05ligZptOsfUMMv/+c17JzLiRgr8tB6aNe
fysrIacloBjVPzL2Pf2w6skz+TTUyCNyiUyginAzT4HUqjPCDJP2OEKJhkTYXMBGFlFagTOXd0ib
+xzlmEdx0r9X7YRu98diyL6wKU7N2YGLu+ioxUtv86VbUlILWip9pNE9PDohvChv8qoqHvdWxV0W
UgqbnTnV2CfzQDbl3zqGw10Vmv1/GxTMLJtXJGNGshR5TS6rGsGuxjcinll08XDXF4+m2UOEq87/
KEu9ZsjZ7Aehl0JeWcdhiS8wIdGmBzZc4dUDaf+WV8CvdvaSMoHxzWHXfGY0VJYOMYdtctMlJ2wd
PL7O/8AkWB3wLctZn98wIwBcHfLsycL5wjxAadAxZd/DT442EMGZ3sSxC572t4xGJFkOasWuw6o9
bDm6oco4lhG+gCus/n8IW0hnwq4/7JNr6T3Ys/KhhGlGIPWmKaIJ0evphQWclOkk0tBgnamlOfO2
cSEemCei7HFONBrqqHx4/2zWorIH9m1FRUrbDQTNQ4NLaGgFTZjtv2TMs1aaFnnCaCWuyixZDyED
2Zt7IJ/bLxYAlKcS1/kS6+xrGt8CAHykKUdzfZQ82PyQykcdw8ft5DLtMJC+WSsUAKt5K/1Ziz5t
ZdwN3QMXWCC3XoB7/6ZSPiw7o8sjXwlME3RqtwNaGjCAOH7EdRiMGF4uCANBs6uAbQI0fF11pKj4
DQ7pdK2ptJc9q/yz7C/09iljKhqvOlnbQZL2PKatQ871ZvAmRp0jL5Ijk+ll6l1tUfmhSt4Qza1G
KF/+C1TSOV1M+WK+5Jkt5LRhHESKwWnfoxmLiZgOoEHwuwPlzoeyvT6H9nhhP6hefgn82uTVBcTo
T7eG+0ljGRTJz3H67HCQ/5s3zFupUdp2E9/30ctAnykXucdGrVTsOMPdYB2o7KiKWHTT8hUNoG+V
M3q4kxzvlGe0H9XzDrrvhgXUrKAjFaX0NjlbsOKGbK5l3cvrF7DTqkuUSkyrNOLhLetc/xY+6f+J
9LsWGjVrbqsSFFxnWNVy7vVjoXaNVo0yjdM3PTd7X21cjCTt3J+eRIGpHeFbBM9WZglGgraP+dBj
fRje3EeiulGsfQ7vBYoBLiash7RrOFOQnlo9ezimMelVsUuFQKnpolDOkLg00W2LrGaLOi+WKxbK
307BKkQivAnFcxplUs07hii0OY8cjt+YiIMGuX9pz2mYh6m+qJAdofFHE/yapIFkRgFd/4oW74Ax
dRbIE+8IdxokgnbmDP781v1fT1VuRPR9gQmszhLurqgau+xC2T67Ni3fVWiRB2AmsUL225p60VTh
wS+w2b9P15lRxyf2DpaFg/7edeWA1i9Vky0RycRuXe8OzLDv9jo2MwkrVu1INTb38ASPa99Q/Q06
joIwiZHBul29v3iidihWr19vF9hGCO8CuKiVmd/ussKTmFwBdz7iBlp39QI5DdNE14rNtEazREeD
48+vOrCP4V6JbsMI84OyAUXkVXTkqckCnF22VSa8fYOclfja3WBuN2syquE8Bw30Bf7nazieSr22
aNHY9IrOM9q4itGak2f8boF+42PbVCH3h9lbbEX7TRc2WWgxYCTxrwNiwmXt8Xw3vrUJdJcMYks+
pCsqRamzNPwCHPIYipvefkt6/X/nBIHTv81u9kEljcE6n0UWSbHMcBuyawSsczvQjhmnR5nxNgRv
tLa9CLxqmOYv/zIziAN4jUuAyhUETPor85FLFmaS5bBB5ZFN3eVSBAWSeIyJpJKv7JzzpgNKdm4J
+EEaazyk3CRet01KSThbubs28JkoEDgA8yEReEM3rtxOxby3BF+7rnof7oWVEbstBRIR2G1T1/UH
RPjQmhqxh5AFM1+74C+ggYb0f/qgRxSnv6mxhcefDDbF2wJkm8LMB5IEoEmEvqBHTnljUonKqbqc
1Aev4UdWP7Z4C3sLJvjcZ7JcQrFeiheM+zIkB1jMd6qmDCJb0I7/hUsaRGzCgrXFlpxR5EQ6wc8V
KWOJnk6HoP3X6QpHGPrDe5LnKoDoYYgKwk4F6ZGV5IttnmfJ6Yb/ti+Z3SgjyFsZkrhez//ekCt9
9JpxZ9vG4J42kaRdkQRTmsgFBjOxJXm4WIDaZIQQF8E34VRQ+Y5o+sRMqP4rXDcKWQUz20IIcceo
1ueLJPbzC80LJlB4u4QR7nlVwpxAZpFtJwmVvEc/UDZrD3IYAtXTnOQgNdDP2UVXwEUeI0g627Ea
IDy/XTIHHEKMIdpCEnnfGYw14J3csgyAZmXqazhfmCLp8CSFDRzndohy4m32rCfl6E+itAdVugic
SVv99JpziUu3df7UGuhjC0ZBQOWQ2SRfB90eMkkYnGpOPgQ6R+V9WYpGxycYaXA+C1ocS0BJlp35
hqqyS/pSDSUZ9O+Rnn0Op/pqW2QSd0RA2hWg6vVM/zRNr9ookkCXXyAI/ZYN9nR0EHb+ADmhABFP
vGNAihz4pHpzIQ6JP9kZNo0c4uxZJF/iaQPCjTQWJLiUtx4F4+lcJICNKThyr0qxjhgTYQCaMPnG
33kjAEw9cSUFNARTTpVNnCooIxrfGOKtFrNhpu8FKsUMkMLsgzw3Hg62RJ8BBjqaKN3SJc9usbf1
yM3PkCjAmcTk9sNV10JgQaCKbRWH2Ta5Bg+0dtHt7xFcaztgjxo8LnOXVZ15gUULxL385AbgMLaz
SPMGwuAFCLHN46y6WOH30+bVfSPJRVkHKeYWfG2jOCepwM0bctYQt5PuBgL3RJdbT07ARafHPgmm
WbDbVAkaiRpg9yauDN/wmkwxt0eEJeRkA6Fub464ttZXnVI/XQ70HiGlpn2nAnSdSYULLKbZjgHc
Ji1E1wfM+xSjXHh5likbk07MMeNkWLIbvC6FO3cFThQUsJlRZ3dz0XRmm1vYOO+yr5F+zB973MqU
i57Kl/grqZwivEvUW7b2wnzb8kWCBgC0D55ve3qWxBfvjMMOaE8bFDjxpNgVLvC5oxPKhfnIz0k4
oMLUFLTNv8rPSjIaYnxsVQPFxDNILTV3p5VEyO9qrmyX0BinozuZjp/5XJxmZW4ZyQOPuxBPnbFk
wUBUPoFe7LaVd2p7ktKEtbHAR7MbHRWR506C89kXDSjq+tMEKec2ANCbz48ZxybqRbED9mNjJSaj
C5ZFXYOyVeE182kkFimVJ6Q/rDzOiVP/qm10cHV3mmOvenzBEqZGPg/9XXMg8xJelQkWSygHgOP0
D0ffrnruj/XsdSRKTKuSuHtkaQOM1jW3gYz2vbfZoPxCW4h+XAojBGc4t+Pr+M49F2AokVaU9cZT
wxfJbpXhBe9sigo+P50rTsBlev9sU1o1x1/qEnrKh8kriispLRoNhf9swmx5KJRje0mg08qmOv8W
kjgCvfkcyXY9rDb3syWmjYFW9PjKz0uM3x3y7LXwpOWFyPCxqh4bcrD8kfz3O8rLwHPwIY07QNmr
RjPlPYMjuD0LE5Yv0VFT6UgqVxxhnZ83V8Z1Zoj4CakY11UeZEN5xRvaCVzX8g5Q1gvEzUOLWk00
9lZJs/jUJjzo6rfG68nD+eEPPI6uGFApf5ZkkSgikZ3x5MRjlEOc13udMIJHVHifnr116qjqBoyA
QCoIrdQ6gU1oX6oOPkTiigFDfZLu4jc2yYkPzz6SWYs3Vu/KhusE4tJKytyhRBcuNXw2KccIHlxF
zTlJYM5CSBQhpdtRvj/JhB3/3f8mVcyyVrgE4jAYGIM5XQaZY2faHQUmfBQjpkSc59xzInenxccv
ABzU8DkSAoqJ9wmgwxC+XITlorzREiPtxNdOs+Da/RBtsnZ6IJVkornHiJFDllkXjMurYOdUYKdA
+wKbzbE9BmkiJDqGGKMIczfPIGnE6/uQa434Xo5W2NBo/KI5JBfU/RQc6BEZ8l0XNNtl85R681a1
RImz70dH3y9lckU3CmuYCUldFsSVCjpwkYkRLa78ksZYC84CSONAVko4RAxrFSR6aZDxsLsetQmw
GCFWw+L3dhlSSMUWtE5nZYCKqvm+f0ZDNJdHJKQeAcHM+SxRJjtjYnUy509uqd+L/TAIcKdkj79N
UdfiJIE4zmHDCMnR3lzg6ZO8cN6ZrVVcU0j4UEk1wz+VJRJ1wPfYq8RPJV8bVTNLugISYoIw/vMV
qX34Lj/sQmaHcqzzY7DzlqGulx9OdSrEu/noWVfuw5jVEs5iXb85H+PBVhHFT8M1/NvY56Ztct3l
SeX4RTjIW6okziE2/zSDjduBgtfzi4npG9QakigQUgitXrb47WYLxN4RhfL8png0zZ3ZOGNlfWwk
HuCyLXH7pBIJ2F6QAIP7GcVv7FO8j9z4Z7TRCzzsdk37B4y+cSKnoy2GuDK9SKl8fLOYwjOJx85D
WNe6owBLn81M1XTW5qgptQ8Dy7C6x09pOB64n8Qo7IiBBpITWq8AtuXqfgR8/HmPuj4+OqI6NdXr
JeSUvA8533ZN2U1jWXD96v/8c/LhBhG5wCEFBvvDACJltdvhvlOcXggOpTmb1XTf97ec9PA/s/Kw
mwD2OmQAR1RMjesaDLEt73Mp6KePWZjPGik207PqOme+BQIdKrgwIvED1zaVrCSKRXgAtVTXtN43
q92ngFSk62IGWxqE0x7XIl1pzWel6iAf18eWq+ITFVpFude/DbuWYbkZ+OX0KhehowGcIu9PMZ9c
+X59S3jR7AzJaVb2QZDVZoD5FNCOPctmxiazf9cZyHmVod1ndMJag1cLRr7nkTBNoSlzD+dpmqJh
is1YVL1qExTUfdDIYcr5u1qva/NxV+xsSmLBCeksGs2GqtBPKm58NLGEeOFBIe2cHJUs9zEM7jcr
FzS2japNK4pLd1FMriOsXh9AZ4UkRjHQ3YQKV7hQ8l/tFmR1xfwvZUMhxIjsxF0/Otj1TeXkUheo
r3FYBMNerytO0uIs+jRV5jt3LmQa/1Rb/NbpInX84puO33gNOcz3MqXUi0ze1KVyHcSlBvZvTkEp
F/wjRFKF+MRKdsUe2UaAVPjvTZJDfgkAS9ZE6f6DGNQUd3Jl2espL+YfTbIqeS1RXlsm7y+zpQBn
aCenQXvE0JL2ZfQT/dIK1G7Mg+iqwLUCe/SPthRWU5LkvbLPxirdu1VdH2bD+kCdxOq4v/fFa9en
4h8ETP9WwvT9NBEryA2oocvLghRzERV6d6FCa2ZoKZjudlKhv6yFr/R3OjHcVmDI/k7SOTk78JXY
aVmDiHZAjN9hsYLBIlf4DWVpOhkwnqzgdkQMBWtauH/ZXF5CN10g8m1EB6PTpDnrxfP3LUItFlnc
aOFDRjLRMKcN3eq55CN3WeO6BqaofegcaorKf1fhQrfMQi5I06zRwFhz1yEI2oRLw4CV7aaPMaXO
Z6M3ct8Y7bum+AVfcqMt9Q9t/w84u6ElxjagGDTwRNJ6Wm9B7OcJ6h/IKqe1rv0Te+gsxkok9vDb
Ip90ZOy6z3jQlJT7eaWJLQotPnFS2DeyWnLYKgBR07Sd98hX4pbXdFG1iHPqbcitFGjK0LGydE0A
F6NtYkBKugD03yYFnpqbf/4fEE0NW9FVvKEg25aMCzH0JceXW2FsGYp4/UHF9f9jcbKgyVNrwsWE
+4IA6jqlPkf3DqkjWlMQwo8mqjtQr8pauFYOCNMVdW3xNgbIJOfgBG22ETH93cw1VHd71TBVzXfx
3/bGWHMTf+RCF53yrDiWJzj/NAPpV6Ox/XlutNuLWb4HAHAlutopIbwWCUhAFv6Fycq9PVDdx1Zu
35b4OOxKczkFeBD28S1r9FLDX09hN8o4nBxdlHo3TNkhZ5XfS4nxjpCEeTZ8hPdPRz48qH0e654M
1bM5gSRME7omBlJy8OzC66aBwRa4TOY11LW4zzXnfnqdELg/NQr9Lx9Ykd7ThwWgGVRXGiKd80X5
+doakfze8XKxCvveWIZTDrR1N0hq3wZ34QDOUcqUjK3akuTn8VLLv+0TFJUx+8Zk8GiODXpnM4Np
OqqdA1YmZ9hNDJUkA21rbaahXkCyTiJUnO5xH2Gu4hizV7aGkk3Fh7hf1Hu8LwBAZV2u6XByMlXm
WqpQHUIEhlAOppcXiS/q6LYvQghJBjCJwLpt3qqIK/c8aDSGuuHnVyKG4Z1paf9RKVvGA2o3LQp0
bpPj1BYhU13mHSxwjDFXCts4TUwlAIJ+TKGa6+bJ+16aeZUqQSZ7px8MWYxHtu0U3SHb6tTVyy86
D7X/OkYssmOock+uo7GBIw7E+kGQvWPBhePvoANDdXNfusQQQh4sQL+Ne31wb1JpWKvKvSXYA0oj
D5rjJ2eRgwlkWxGotgoTAZ1HzhXA47I89l/BPk1qqBtq1Eu7xtP20pD1E62xGASi63ZqVt5En0da
ZlqNgUBVB+UjYHa5swbXYoLt7KiWaqZQc4+fnFcWbsmD62JldQmYN2FBI/+m0/KJeKDEk/PUt9Cp
MBxHLcqoGgTQhRaoulrUv2O+Lak5tdlqXbp9rPueEs7kk6e3tqJNSKNUyE9bIatbCHmYIXUtvUl/
0YkXBdyHNQ0UeY78DQh24y5el/X6wQW4meRJKw7UJE/xTTOJn6oNWtbWun4/IoORp+WSsqlXr4Bh
JfUf8XxelPTcJ5HF6Pb4NtXxcZmo3FuxKxbmilcio46KHIMrhJ/ZQbOgXydvT1zYGshmzbY+vsBO
GVu9JrIh3wwWFfWYE8h89UB20G+rlzQTJrhRq5RARWkclAMcDtDtY1VQkOpzXdGMfh+ZYY2yp4Rv
byfj/8g5yfHCqOqu7qwBlwbEluRE5hW14QtBeIdcMZOwMyhrSuT7Vh/UBEQImgxSRizWPJmQp7IR
qagUR+92PtlyCf8JAyfV+Sp4mPW2JQ0N+T/OGGfShJfWwfJqGRirWUNpVTKsSz0jvQLMOKy3VKwj
9DF0Z+7eZkFFn6P9gdNd9ABK9F4QaLful/sBCStWZnN6EKmlRhzoUgkce7uvkbEahj9HcwHer0E5
lh1Xuaa++kAZaRbax4L185qGrD2KItXAD4JF4YuCSG8Y6giEiFSunhu6V7ARNsJJTekGlu7F47yU
MsW3CFoZfeOgItBZxNZVTp+8uBrwNc8WgaTzDmEZpR+WY0bgxHfGtaPE5+zb0s7RYvmsHnj7mp6G
WEAPGcpGUi8x9NNT1nCdxRfx8uEp1BEnRAH0hLtHpL1+DwDfgYZlgEHE6FTjD+R6M3wjy2tTfuKR
daRk9y+frSX0VBFpO4uPTVRV7c3eYMbAWsnyMqXENbt2HPAxLleocT6W6wXxJcTN3XxQOTw1Ugds
iBNfgYJ/3o6Jcp7Yfkniux0YWfmyPmNj39/AIFRUHvmtiZo2I/lZQXehf7pPaVGmi77mBL5dnxdT
3oEd0HQe/uVYyFXggh93KgneNaV86EZkvLU1qC6g7zaqHVVjlx4bk+B6BH+x1cEGVMQ5vjcpML9g
b/r0c94/lqi4YiM55uenI6noWWXirz68Gsr5SQ+u9gaY3zu1zNLl4fif7z22QRQ/IRHJE/kUpueV
tModS+JJFJxPv1TI/eUuz5byD3/RQBtG/I2uDtEbW79CJPTMVz1h2KUBFQdyHvZbeuToWykx6oYn
Fo7XEb3h3Q0DVK5lujC++SlEHrOmFwZ5J2io6fE+fa4Z3nT8YmhC0AUm+NBfbkyS6h+1C7XEPHxG
Vbk9L8DQrAzFLR4kaZJIFRAYdJ6N/7/lyUGWa7Iu3n/hBshkbI3mwHLDBrDS+9ZaFZCHcMzX3FEA
Res7S7OJT7VG32P7TCg5HUMX+zUaa0yO72FThwm0Nqm0TOK0jUESVGvCo7ejwmXKWDa8G3JrCvh5
ty14hTgRMcYwqP/WvrvkoMDIE8HJ7vuDOi2MAv/exNkOW5/Bb3gi6DG4BZ3QV3fhWsPg8eVBIaFY
iCs4R0t2IFoYqjsKkf1bnB2CxUy6XzonlQZh36jxHiSGtFvfckbojN4xcJzXsdOdNtqOQi2prP4V
kNubrImAvSQCEIFSnzzS71WlG5jNpLA3u5mFU82ZksiYllzowddHXyhqv5daSLdOGBjRVN0BCQ0+
ItLipWLkH+6VeGxcH98kP322KNwl18+TV3IOA7zYtg/2KULRjJsQRmyAJa6g/zQuLGmXFElFPvrD
tVHWnGOAUbkjCnZETwuJB2ldeGRphq9xGjmDhYFsPjgvKUL0cKXiZYMl0KijgkyUUH3rs1+JCHUl
cOI0wXA6phy0KHg8HcqcjXKtta5vJWPAL50OWdS+3a+Net1agddUR65nosB+HfPzbCxj9bm1CVui
0yTT69zcRTrH7bnZzFCNL+YFlkIhUu37g6VflKmoJQNReHB2N1qKR29xxW5qBjmOoNDVIVnlDlBh
B4L/ITp9217i4ALzhe4OBgwiUDgkFvVskdDMNuUBmKVtTkxtXJtP7F3Y5iVCJ29kvqp0oUNWK97I
9YaP8vTL6IwdfrJ0E44Y3MCnR//Si+EepbxMQ3c5OHggsvPvJ2NE67tW8MaZylxEBAetxmwaBDR7
crt2JlAuQcPUfV9yNCgZeN2Mw8QwSyXPAcOjZFB02xbU0c/SN6t/8+ilTLclPBuQ+348ctJlyo5y
ufxYw1YZNUNOZM6N8vMJicVLFeHz0zIuXRXTA//6+z6yOomctMdUrnVCdrJwgVuphmWCef17/uJz
FwIYKKNQ2BhaPr5mp6UfeoBm1V6lr3Hh0TzvauQsVa2/3gruDr0bajYcA0GA/nzqTEk3H+XMWOsc
rgFryNi1H7iF/bDvsmgib2k3XiR27sQhi/smvaSW8xD45kTOWc5SGd54h/aoGy23+k930Kdwnx0c
ZllsgT6psXM7EEXjkO3eF7yEAkGaiNiZzuTfRC9TU5ghIjgRu6TiwiVpb6GP+LieMVc/ssD/Mr2e
crEjpmexUjvDasPKQvKxF6TP0TJGjn1ln5uNif+njJOv+x2JHZqyckYM3Btv3Sje/pIy06AFJW9w
U4hF5nKRzIYvQK7qLsfTnsdKA7VnE7RqUxY51fhrUuqYg67UIB9rDFpV3tAAe0dOey2OTwEpSBlC
R4nZs3Di18Rq/7ZxBPvTKQoH2lvTFbhp1FPrXhTeOAmhDmmLhFilBcFWQvaPfYREBqN0eR/CzR+0
WkCnbg0wcchPZAbfGeB4Dtdot1+m7Tqll8iJ6maXFqv3/iZyul2VIL/AOMKgx1u6MXsWiDg62vk7
5lxqyllUGJgwlRMYKBJkt4NbBSbSxhitctoMhKmIg436ogEd4rq02dJDLGFrpy4h/gAxVBTSzA+P
Sst5UfCwC0QPB5IvmrhUn8KxqtnaU8BVBVIHMWXRoM2sDRR3MfBz4p0D73/QX72yL0f+UQfeToNl
XHWalE+r/b77EIDEpCN4aRSptfMI8DlsdVIhX+vd7jv31mvM+p1jQ1U0FwGmIBYz9SwDu6fT+/u9
rjPblTX3PCc4cjYnf++GMKCtOedP+D8vV6RvNeo2pxz9nFNYHRgpm2t2xoRCH8lhrEhWa6NYjdP5
iGKH9pOwaA6f7gsVm3MaZuBR1PwbYE24zzyn/AMZoA/VFuD6kJ/DHcJah6u/375N8WiyO4qQj0ly
MglTX/txmYhLUbuDx5O+0v9DocA3P2tBNMtgx8eNyWYAuVvzXhQhsulvqMuhW3so0I06lJM+QvJI
qyqoeVWKt8A3jyetnZcHfHdyVXLVofgn8eHM1SzuyISItWHA0iTFYYToGgPbbdNuQIuApgdbHX2r
KS/aohfIbZcGgC/g3xTXwjel96AQqRg675owxl4nIJi0bYwyDCB0myZ8mciBEYbsQRVJXa4VZOgd
EZUvxKXSwEPcv3RLL9sjk0M9GwKx5ddKhKpP07NNYznXblUELi99WFEBj30eCwO72FlWZVZybLV6
tmluNKLJpOAOu5vTlaJSzZ7sFgFzu3tdGEUkXHVyhVhodZTN37IGPqyMp7aYvTD5dBknFJC10f6g
/yhFWPg8JRyzjx0jXSKQl6Q+puP7+u1wZfzfiYbib32NF23wmXXTs9TIoQs61zALBTPaukyNQf9F
0K6IVGyQ1WZ9M4Fg4YSERMNGriCxKOUtQKXi7jyaQzCPFszMTIcklmsYlpGG9h30q0UVuvjd8JSo
PP9grDzfxcU8pSkvUZ62eEh3ScE/jekFasoq0ZV6/89IJOUbEDtVdg23lEKYb/y5EfUWga8Sd/Vf
XP9vLULu4cOp2LOPvUFdzulbk7WDQM6kM5QO+JlopbEeqUqYLYGd25Ofsnp6abcEj9i8aDXb6ocq
Q078Uw21yPvhgJVGHbx5sxhPrrEpfY0ehL6jnflnbCx8o3+dHYdrKqRyf1rPVA0CDcf/7m7w56le
GbvaK5K+HLF19VPMqxdub3rxZuuKtIKobYaShkU6AGArCP06fLf1ImK0Fm9Ql88UDrQpEHlRQ4XJ
W+NpdQiMU3lMOQIUx4vSbT5olF5fgaufzuBe1394Ix1XVMGNiPVb0tL3LV/wFHH3fU4s41I/7esi
gm9KgwfjMhjPH/jBVpKTO5wj21kbgQgizOoMAqsF30L3QM1IN9Xqbee7dbkuHpA2f7eWoe2ZOni/
+k8sEo46RBtoqqf5z1xowqOKahU3e+dfCQdo73bPhvHFv7tYYrNc3Wd0LNDtVsdiz5haEx0F/yLm
YfDHIVYtNgXXFUNlX02qtmsSnyasJK6GRbfw6ybs8nhlIx2+ddLvDeWurkDfO1MCDmwqKbYzzk9X
1v6pCe1X3ccmLJ0s56M5u6+XXvQtWZcebiz9QT1yXVSRa6upjdcz8PtNEznaGi9wo0lDcb7lN16k
phIt7GkuZnPX681IGc7IEL0R1wVNoC2I/aC9IPLmSLq2+kqpEXu89ZifobieFuJFRuz1df4C8UWw
Wjk7nKd5Oi7tDo7qnZS6f1pUaBJnKSTtUQLn7IHofkv2Yu5WtJt4XFFLUtI6CPa98e/J2l4GYGBm
dCCRPzzMg2iPyOA/nU8YWZL9IAWmx2Rq3jNMDnry/CnB9pAk/+NuqH+avZOAQo7+bRld+qT1rcbh
IyLtOFAGx5O/w1GyRmBfS8vuCxo0zdQUCzsbHVUr0KwIwc+Nr75qF+SXFHO5OxazC6cQu6eigA4o
E2pQLZYPfBCY2yIwFnt2t5wzXPZ/XBIyp/Y73weZ2Ha9alwUTI7NQRmM7lCOVVQwD7v8KYlazndt
0FZ+DtcKUFwIOQqxmpE6/WnJfGzuUjp3ci4iuPqkpMRFbD9h+QhG2SObTnFH+h1Ivewr2lD5xrMc
f3sOVY4zhhQxHuKVc5/fE/EYYSub8wk4FqC6zvVmC+HBGxkaqV8suoHn9zl2TcfVuLujeMVW9FYz
iT0/alFZuUP5wM/K2df6ISoXHQnMTxDNUQb88dGPM2UsNB0eGH057HBbSeJr2HyJvaNrbjg8G1L5
aUVhH/o/MWuMSL/qPYc8bIC5Hh2V7qoi82HfOJWhcajGloElKyb0x3MUCPIZhmlcEbjSeSucgnGy
O8pl/N/i+2TK5CsnnyzmrGXHAKdRdffBVFHcWoJMfIUsjNqsmPY8sJ1LGe5JiXTKIUOMyvHXi/hb
49xRfx0qDsn7xr3xnkPIm0+J2OW8rgwFWYifWxhln2nY/DCqF4yp1KlSg86fw9HoaRpK8oqibu8m
X85PC1Ss0k9/uyTYhSyPkuXvYHgZUau4+Zvc7FZ8sweFgT4wKontNq1YPE1hkIgQFwc9EKTScVuO
kiFFEno5KJFaCb2UorXeOLwA7Mll4ELeyovJKblzfv6b7WPweWVDJT/dTYANLH34bVvBAUO6VXzs
frZjt4tqbM1gpGQBihiTfH9CwJB+9DfhBytDlfwzi4kbjNjmc6FwIjiZ3rcukQy9NZk2KlbttMEs
lLu3lfIaGDNBZI99KO0rc8A7G3t6DNJZ5ts+VQ8quJi44BkkphXMmnmxElf89JzTlk6BwV/3me97
6Urb+7xZys7yBXrrt466pexqoC06C8RT+wTwK3yo7Leb15EHymehBNaLs0eeVnQoSOwoVSXxpBF0
xJYi9huNPFl8boMsyxKlu0ddRw6lmQbhPU4Fx6FxBYX8xG3fL/dlx/myxmV/cIHATz+z4ITAwiTA
n9PKrFhEpw3CIfmcIO1D+YcEDy4IOEtghTY5KXktxLsBSZLUukvWCcSdqbs6BTZrbbxUTk7+CRoO
wUMZu7/snZBdBnIMZbVvFhN5jeiopAqr90INlFn2A6J7QiWLZGVXqHtVQt908e+S8u5VIPhG0+/G
PtUEw3SVWZUWU+LUTk1a79n95TWIpabOm6I+gxnQ1lITQMFXRBSfL4C7IyqG0LAnUmZ4pu+fMjlA
h6WhdbDe6PPv1RXFkzSTDY90dHzc90rTFzUvbyr+iNkQpY+6MS277uDwBBgnllZuC2zioMuMbXCD
2SPCdB+awLRFC7qn/yLxCJmwjt6c6NYXv2eJv7zMSLgDDuY25j9PCr+jAZPIVX7ub+DA7/ZN5sH2
+GFPvWZk61szAmOVlBLjVMLJ/4g+eXwAf0BisROeNmAQSKLaudy5h5zRo6inbGPvnxujtjLymZ2c
9hvVFbkOrF3v+NjR2mW56qotoenDWTR/Wp3//ZPQnj8FUBHh3DFPiz6zcsgT8FirmiQ5r2L55LYv
vhwfjjMNXZjiLZymmCv93yHOV2Y/lTHB/OM+yWFCOshyKk9we9L8UuGz1+gv35Ta7d7zZKYo9P06
Dfx7zNCG3oqcXGcezgy2L7tEpHAMRiTc+88/onCVIIXpLxX7KotTmRzXM01XKKMxwLsXjbW1qA1L
9XfObY1/krC+zZz4w5U9qXvFRphKKZ8Qv3c4xHqFTj4oaM79lajkdpQA5ON+comBGjepfCeAUlIz
E39P019NCttwsqhldGUNHJ2aGtkEReGcrLLvlhF9vdIRTmDOhPi39+AtXgaUZuznvcuiPYij7/ZQ
Ualz5b+XrZvkUgjtkkfhpetKJUp6uu+8UZRmvCRssYprWgWJS53kutOrm1VjWiHzuLga6lZdzC41
OSMTPNmi9eRB4IjOTCumPecsW7QJ7NOVLqX20P8cmq5zo1+EHTfRYqqYRPhGrKFTifiBcgexOJxp
U1+EE65FEX9vILTSbEV/YX179dRx8LyVEg3g7qrl6qaZtTGtSO6xArDxpCjgw/S5/m8QRa5jEqGH
VBSph8e3rrrDXLvskggRMfAC9WydWt0z5J9m9tw8lqyaTYy80nHcJakahQ6njI/hu18t9qcdHw86
MbC+UQCRKif6vCTbbUBWy8jsCrUovjsR5x617pCpON/d05LsE8QeZ+0A65pblGPle1CRg6J539Cq
56C/MPYKub0+hpnILqZOffBj/y78QMfX/exEScDGVTUmUhsK/e484w1Xfmgac7DUi+huqe9TwQJi
i9PMgd/RUI00DsO+V6i1x4ujDOhR2d1aIogiQ04oTZ1g7IDSmE/8bGJwYMfdRdHdRseGN0KjOThn
gaAvqovugKvxgoI54TIqHGmpPejBnW6O7whadbFYRM4/DRGf/y2hAhYDQTfCGi6o8pshr3K5jvSK
CTeb2v0twc1n3+Z1I/YS0/NAgxHes4BGTBiPPjl9MG5x74RFS0ZfXJQV2MJaXaxD6iBD+PUTlOZa
5MAhIKi1nD41gZiqM4RWH9s14U30Oqwob2H6z0EhyGUlzZr5UQLtYBfQLMHxy3tuND7h7fMi+nYZ
WZEq7vaywKsx8IHg1iieTzKEYjKTZWVFSnqTdcNiVOynyFcrEtbSIGRYlhQaKOjM6fPWTCXafgLC
X22oYiXio03LeRzc6Rn+hpK0P0QNl+m+9+8NSUGectzCeiagEPuElnQv+9FKGj+CwIpXBHUuZuBY
0Z2INZaw5pd6p1hHWmB9NnZ8nOSpdpQ6XPylllXQ5MCevVlI4VtGzo4QlJ0uSDMlSbpOdDNRhIkA
Mbsf9tB6Jw2OaQP300IGkRznB0ZFNhxagNiysIjP6t5I/YyO9VOJgmGfBmdMMGtBnqxXYnmzSTJ1
KY+fZhXzXDhOgDRuJpnNTP2Z64ntetyW1VbqV5UZv+wLzqm9rBJHDqJzamUy7p9FpwbUvwz06Xqv
86s22FeI1gcUsKYpHvkzhkDAjwff1a6J/TIhucDcRlU+Ms0gvbPaEDjSFjZaXWegRFhATqQSYNjS
AWeqCpsY6QnErwyLGPETuJDGdfHucTBH0fmk2XLpQUJ6u771Nc6CAdhYNn7VHbR8pUGAsFQMcPsj
9RZHOVrCYWlTqj1SqGuEUVilt4J2NjI/wWyurM0g9Q8HzLlpbCLzu9vBgnKC7mJPFYk5I3c1eICa
8NyI2SAsy/QBj5RhepnZpGOWMFEfFRwX1jH3gmSnRAQqBgguAte6JCAXSc0lsIBeUv4HwizqCp3D
1/gKALTmRs0S72Fy06AKiaXD+C9pGaO8RWW4RdAyspq7OI4502fvDUKYrP5eH8nOi0lYWjHhsSBJ
BtwhOeA+RHztTicKjxbVFTmsXIABrfj9jwH4RAAoRe99vUaHipPEwtqIRQa0wMY6Z1xa06fF5elw
U4xC4UUaz/irl2XdNtcSKQs+ZYFxTAdHs11YiESlfogSO+ionoWh9/LnJcMluSdNsMWsQJvJJYd+
J7rtCWXMLjssdwZ5AiyX9ApwJNlEOKU2sfbsmSJvI8usS4GRPG7fX1EZgDQTpZopjZXfBMwvYVxV
kbVAl2qRGxMUbQFqTKx6vNBYEQK6TjsKYinXj/VQcUvxjMNHGHTZSWXg1JtVpYrrwmVW1dMDunBF
LkLMYdAwmXZtQONxb5ITE+y7d9J0+8tetr5NrQVpJ1sUVnRLBtBw9SVLae33J2E8T9aZ6NCeRT6u
18/EO614R7Zsh80eFpfd3hR/K6KKCrEoVRM5atRNAcvBsfGA6dpRboVTJEGkoQjKAbhwxCPd76pA
MPqZ5jvPpIugDCctrZ+rrlPD40TBA6pDPWNvJ5HWkajFDdGM1O+vrSpXHR5+56/IGKgA6gFnDHNB
sRLPyppCoTlyxfSRyVQuPboEDMfIVCgEY0nayymCu1ZjXl57w/KYCw0gMiA9g2jPqWL5bKyLop6K
KMPx/Y4ugMi7PRBexnO6sMW17ehGtuJv3p5g1xbUvdCJsunYeuMZRdIYrqX08ac6BdpUnngCvQPV
mP7p+c2w2NaiYWkYia0ZQ1tmeMpKmRj8RmwDuORotxWSaamXk9OQmGQacB74eAE5h5AIwdenBYBa
FkyO6c+Blw0k+fCaPY9vaOvJMJEIWRAeOMLBL8uFDyjTSqBzx3kVkFIWQjZPL0MeOPmoObAPOjEl
5RYUnt5gw5xBEG799Kc2qTz3NbZSYSmijqh3kwZ8ODgNjtzHkWEerLcFrj1KrpwJQcmXo7jHD46x
TaD9yFXD0Hn9wD1IeJr+aVwVOTBZHBaBFFRMDoc3g0dt7zsrbFPFFOUu5be6wpqZ7VhshXmdgarc
txOBaw6cLmNkCBGd9ySu49ETeVHuY0nlIK6HJ8vDOrwQ1QdHci+FRYwp8L5hJpYz2XmZ2nRH+o+G
Ou950uGUmJJrkV5/hJUx/a1KvopVJ2b/nroy5cYXH4cGx+nX4ckgzHGPfmO1pwb9FOYBxXD/Y12N
ibqdOeDbABWoNkitzsjZkCTDAT8WJK4jPtoCqgq8kogUqzf96et1KOICT41LVLE0wOjFvfuSpKYr
M7MvSbgsbWHQgpKlM19czThAfJiLLaYwQAMlgAQZeh9H+RfMV1n8PgO/pdgAsvCT0V1fwt8xl0mf
EWuc3p8vIVebSUO7oKnosZ99YnYy/FTSNjlkw9YxZszXVEDy4YUJKYMiUM2ND9JPAZNmEbM0QOQU
sq06eISDRzkyMSN52j2+rFaSzOvS7Qk6oR0ZLZDBPDd6FwEBswzHc62v8GsZwQskFXr3LpSxmFOD
GVmbBXDZ7keEh31Hec+8ni5jYbVOQkIB3Q8wv9nL2JQr/HqGKBIAHrfcIEDkBD2uWrpmcGNR1Qb4
G74x06U5jzUITqRH1E6cbXxk2xfZekCgB7sXrPfQqTPt9ukOJ5pIbsliqQtS5pUpwmqGbgdxsToK
DW/okYeNMejhGTv0byhQso6ud3dTAoFrSxFGhLhR3ZGHMKGsuC/acZCwx4Y6/o9LBg0+QBwT17pW
5zr6EBVk83mX1pMIsqCUvfamQar3bLiCavb0RuYsvckFx8RQiznYCXBttqT4DnzkXxM9cLhHGJ7S
6R0V4Jfk77dAIsAIbHYyDjlvzJbcB3ZNMpPsJea6H88dV/lyU9D3fJ9D/BAqcMWD5FslM90tMwlQ
k/+ZSoH2RvQMpXujPhULZqX7hbRaMGj2sE1P04+2sTgAEEeuDaewE/dS6oUCQ2J67iA03ilihpK2
4gKZUiFH4RBQ7GpImGW2vLiSJJDmrHYwvulD0OMrL8OKTGXn2gxcYLt3C5LjWA2AT+gJw1rmTrKR
KvjKpo9fLx+iV9dk2/40nPylm/ebW/SwXULUVJGp2Cms6quWp7LkOnBzYDHLTEeu++K/DHIzlEUK
zfZLje37W5IibPlbIXqQ0dYVD+ykeTXUhRvsOBkRLj66p4Wd8cxLhIy/mBa5dGpBDDxPV220KK3D
GUwftIT0U6GZWFXGIbBATlRRW/ZS/KEEVOFjy61VN3w2KOvSiYHpurzsbVSIKHwxISJFua0W5un3
MOxlZ9PT5ELuvgBH5G3RibhGWyotXqhRoNepSkhjchrjH/V5TLivwF5g6622mba10JoUQjugY8aO
x2S+VWdtKC2cSqJGSBXXF9SkmOrJMhNK32maBM5PcwIrS90QXPrtrLrE2VKkNriO7V3ATxcYDA7n
kqMQbJXADP85ZjirCPlGDQ47raRNXmzp8Uu3biIF+JKTokY6Au8KyTOVRqGKhCbKeHuuecB1gbjb
TxIYbtEf+RZCfeXNq0QqDkO+8m+XiaeGeo4QMA/+eVfiqEnC8LZADzfA0Spa7tQU/s8fSihjE/nA
plK11TPeB+DV0zF6w11wE7YlA+ZmcVKRLgJIr2CD4Zvh4W4RuDF/FSwNI/IgQX7WCENVaitqsm4x
grrtTVifeNk2Y/uZAbiJlJhSZerdfPa9WaCrDAS4zQoKpVmTXpjg9QA/F+GbUMEeltuT9g1pgtqE
Wa/X1pWtiDf/urIyPao0pMtOwVDOmZgsk17T7e//vxe3G6OxszGUjkDxpbtZ0G6psyi3rS/LaIpS
N6l71jEb4fhtH3CJvJGBPqaiOg5HJ4/mX+Bwf6Q4kIz4Ev1snx2uyvCWhbp6jyIF4rvysvqae94f
3bKYRfyuX+z+U8dZv0eB7I9fJeg0inaGNx7JEd1epPpj0gxo56UUwgvufWg0ky/l7j+Vn6tHpRiq
YsKhCWJD5GJROLGEvIzg81X8oKIqSDoMZ/qnEaNhOrN3CnpSZonqo18XZrfiV6yUvSJr2Yq5pYhI
IlnRQ4AqRtLPmKT/FMDWXFScJTUpqf0xaXUWVGUiWoQB+UF1xww/QKyvphlj1sDnrZlvErIw+9dE
KQXVjnOxTzKJ9z2+4v6hfpKQGugfFQ95WmQDdfD8N8EV07Gzhg+VaWYmEkX1Nu0/LOBBnXu9RIGt
z4YefQXyXi+3A7Imozv7poBCHFtd7t7cS5Q1I1Fv5A+IRngzf6nNGURIEgRN26Cy0aXJa2H3433A
gBIeP1Yn/sfoUzGQYoGpPRa1Au67wfuMBovXpREeiXRvpBtLWSeCIwY+rSfDZzMVtadaFDkj5NGF
J0hkDlAe7XR0B6vQ6JNN7dhmZnuaZp7g/CqyZKY3wRXsLcp/aaH4L0PFnUysx4aqg0Dm9QAD42jV
eLcpb1T8kjEoBUht7TZjrFMXyYxAENrPhj1lbuAToQxOPsfFiyButVvbNcZNWNDwiol9JmKlp8JM
r9cuStLD4pPUBiP0N80lWt1EWxaopVVA57s2kQDx5Tn6huFqYzCTHIqSNJvakQ2LhZCvX5xfny+X
pnvNa5W9bb8KD1/wjEA1NLW/t6UVRjKe0cq8KhUFodb+IQfmuAaULdvd6g4oAZStSQHJGc7bFEkl
BZNZdgG07TRPjgpl9cd68z+0jyOU6nuaZp+A2axCulYvqN2ucKyK+v2lBPT/8fGepogPWHgDMY+W
0Ce8CdRtw7y+6NQpQQkhp1Owe5T3meu4BYCUjPClmlR977RZoKYu6FL8faOmCW8uEuDtw09LDknE
ed6p1P1o0CHRp4XYELlmDfu8PPZThTmjbjhTLF/yO0giONFceNdfnuQrQoADkrTnToEfZWvs7Q3p
AUTRE25mD8dg6VYK0GXeIfzJxF4CrGa8L9ou7VkS5LbZDc6fwX0uJlfkmRgDl3gwM96tko1iHY3M
2SVmw4DpJnbRdYgtUKbmeIIZLY4FrDzEiHpwcZ2LwRv0xQ1OMHY4O2KnYonrZO21OYYtWgRJzZTf
Dkcon4YCAI+3+ds4LqKAjpQnA6BGiWGj+IBsFV0aMWPUphzkKxkS2jd5+k7BXCGGAC5665aXpnGZ
BEodOVpik5APm1afXyMyAMKduY+PzuLqja0Qv3+40l076NgzJiAVnEE1hj6yOq4pndgV4ALKF7cQ
fNvpGlVtFUPI9Xjp5vQRi6ETii3R2rxgMnm9jSOTqctzi5esOK9kp1daj/MH/hgffhTe6Ub5oTIH
kcG8d0UxCkg8MBKsEal3XSduk2tpCUNE64wnEH5ladnAncU2lBcwyjvqr5LFXhzcAZ2hESPFZkCJ
76A75/qTDODKBrgCH81fbolz3p+kuAtcIJjnMM7wq95lqhtGYXz81J7y3km9JOyStaukwwBaIVaC
iafUJKQ2joKjrDj5gDz0L+tivSKuV6rPLewrDH13cWQcO0bkNZ4l4xHO5TEmso0gQcE5CKY2r+Rf
P/1825QCQTnYfvIRGS6qmXpKYEamQl+D8C/vO72vsnn6425FKIxYN5m1cUNEXUY421As8lCLw+Rl
16iUB/rm7X8z7t+FrvpGNV1nCIFdVUeDyMfCuDbAyCdHeyytCr0hG662HKFEXE9AUcgmg6ijxEhB
TXrJRbk0QQSiMLrUdOQBY+AiZbfh+OV39maFh2IWlbm/2jV+XW1EfMsr0K0x4CpF6ehNo7DEef5P
TEKI5h8C9mAC/YRKSOkn0oTNNnzOyhB7J0pKnncsLIF5/0JG3/U8TDvAbteUvGwlp9Dqh2ruzZIQ
n2g2bbZaw56IP5PcW/WINtcSFrn6qF9I4lxFeWroz6MR3Dzo43/HrOuM1V4ntqiSfHgR7NrbBZU0
10P9xN6UXbuIZwDbXC2G+NmzolPuWk+RjXgtCQB7CmPyTyA/USTxJJpeRrAYCddNhNWumCwCLicU
RULoTB9quBWB29b+DP5TxWT2oEjN9Kq+Uho3bkHYFhFhv6qzcwRVmm8SiM0v015TTlFCSpkPxUi8
ekt2KG6qQ2jV3tjOijvnqdYzMOBvuOH5D2benccd6IANnfwaddp2er3LZxrp2z/ZHLPGnmf0LWOx
+qp5APhqzJ8OpRtXdCGfD7O5aQYJs5+fGV143Ef/5yYPEIOoyOnEiDO7cq0ZyF1n3L3EspTaLfKJ
C8t6o6Ri00L7d8uSoZMor9ZKpCs+J+Gv76cHmea/5Y+SFbyC28mkVsJHxMvSMbrxBMmzaOn7HjsP
Bxya8nVOHznnIOnCH7fmbOyTv4K0eJIJ8pS4vin8FZNPo5JUDTkJdTJl+xEYquoWHmmys1IigwTd
K0bf1vAVfH6k4e07exEF25wZiwxkDgOBeSTHUK19ygGXfJnSMYAJkQ6Moqyp870YgNR9sawP3a+g
/NzFc1C6kM5hgvgTU/rSnSXK/LSpfHVNKUoseB8k9S5cqhrJMOIVOuc2Z0jGoHmzuZ6k3LL0B0As
Ej28eb2EXh4MCXE3Pc4luiIjf8EN0GfNRfTqd45dFBN6BYAqSb1i6YwlyrXx69vZYFRM9PtXBkSN
+rLBHmg3w3B2gyceFBiTPJc2QI0XEP9Ui2GktR8GqQPSMn/K6IRfvLUjUHcAa4KwqNgwHaPek8fm
haFk2+m3MVFGRPVf3Pd+CrhGHDpQUEhNP9kFEU3yl4sni+92f/mUKK/s7SXrkzkFVTxX03kGHM0g
0uyCwUEn2wref8ClfGGawwbvycPyF3GMnq1PPbiCyylg///g4ngddtgkIpNZdEzwxon/0HYIPkaK
I8oDFSFN3stietjJubJMCBCOY3Ka+HSquTcsb9HtUrOQZzll05Jrf/U4tpg1yZqWyJ1tqOxnpWsp
4DvoMIr5hul9Eymz9WDjp24nrBqEBqUxgyn47YXNEPCsABGWDsxoDeUmoOF0DFXW7z6jBtENx6Jx
cxKqBy5Vzqb/YjUO0j+t00MT2kdIMWv66Z3pXnofbEWhikRAjSXkZkzkoNIEPWWIIMxfrLRMneJB
b4z+lAqLCSwbrwbXKBCUSlSZjPcm3tyzsUR2W5CRB0POvy2cc4Mr9V1mX+jnn+dwHH3sCXwftwT4
RHLqw/hkwl3Lz0MzJ4Yn7hVZ8ztAz8lGvgc8vQZTMhEaS7eAHd9ZwhPu8svyMgIUPWBhbsdlk0sW
ej/ZZpncoNlAc1MeOfxEaXVbvwOHdzkYPSS34wI9CZTPWAed2RJi67WMnZu+a8naA9W8BWN3/RRc
clL/fxpaTUVuT9Bl0t9bXJU9bpv60esABSyEcdteBmNZ4lU6ubhN0AopNHaEBCUsEMAgSslLkViU
YxfHTx25j0SHUMhhVi12alk31oSqxMmBavN3b0tXK8ZkZOWUTz4fvU7+e0ko4l+0O0CD1ehgRPK0
Ywx8At9kyRTmzZT91NDLd/Nabx63nmDqEZPu4Hr31cWA7wFgNQtdZL6e6kYofNoqFbvDaJIn3BLP
IgxSr7am9JyCDYvfIHUGSi6Qj60qmtNDHa2TswGXxZ15XzUsu/1siaEHwDfoo/hj9TpfiMI7mjt0
A7YPYzyjuNY+0DbjYN9YFlF1FtUNhl9XLmZ95vd9qz62YjvNq+yhFmR90lyTXb29G7ciCAnUtJhe
N+aTS7Fl26aFgimSeDVcLHW9ulubBch898RfywLtl/vu5or/jYol7L7Js4bAgA8YxHdthda9jyH5
WLd9kJ6ZelDpPl8brVobSov7FlUJiqjN2zGWzPQwQ1UzIt1NNFBwMklE4d6xWUH43eCxw1I5ULbE
MXL0Kh2zm8RTawEJOb1BqP7vf0WfZEuy82pWFj99tBlX8dWtEmiXE3Mqu4dBTRKa57QyRzzwuqsw
71R5FYDRFPwMfaKhaFtr8uoBqneb0XhzRmVQv4ZKM0rK6oyGZ8RZi4C25Kmc3hlF1IGkq4ur0m0c
Nknlajd1EyiMSJ8LFlRJx6QSkpzzXFMmmC2G/MWnGHSkKRluNXYkKOkit78G4xQUx4zIlZPWbRCy
fFGjs7YC+cliHtMjGJfS0NKEggw4pFCsKc7cvGhWCOooHAuNv6Fqq3pXcQ7OnfxOYOcBcniycPBo
UiLZfrGAViaS8WB8h+0VxTy/vbu9rx+q6kiUnlxYJiu54vG3Uy83reyV3PZ5Nx5wcCaRYC7KAkCL
hm5t88ltG3BJ2swZY64Xx0A0ozFCKs47AQG0O2Mn5sRCpJA+zpSes3dNEnzZbF/JTqxh3sTwwr7b
HguumvUO0nvgTh4V32wBMfOT+8LtN541V4ljsYtwyJI7jg6Fj4e2jFwBSULIgxuxJAXo+SvDzgD8
ws7dzE2DLhNcUAgnsEf9biGQL/HkqGE9smh9n4OT5gayPWhTxo5uTo4QW4YqpKCAIf8srNabhdN/
Stpv1pPUCEIo9uJsMFMyUHqKkzBtgyXnbPCwA2cxvmHLI8hzE6lu00wYccA1S0QjCZYMQeXzAOMw
hzDOVrRSdxwqFlOeQRMmkz9gqOhgeLFAkrE0XRdNYrUGhAezppIueXrOW99JWR2sgNy6X6pywscI
g/30JAO4ceF76LIz9Z+FBYnaFXXW+7+b2XsMCDfuhF7XIkAm7E91sKOCVpah5D2KocspYvyNjQbZ
VYCN7W5upRnpNdNIZz/MmEJEJnkkZolzyUpPAl4oB2+oZyk1SgM7p9Hm7w2mYVgxelAqLdjStXP2
NEmFwZWQ60DS+mUb8Udlnowu9/U5EAjG83FjddwmBxvn332O7h1ayvhc14Gw+YeTBq0btJjFpg8o
qNUQFGJaT/fxNRV870APVvQgQLyzpDWFKFZsGWY+WeE/AaVsHz6qIp0cDGxpBcK0MYd2tupIjwmw
HiwPUhETMXV+3HrI6BeaxbBSSKZhF1Wawzu4jLnjo2ioyqB+7L88KnzDTzRueH0C2sU+n5PyPj7a
M20EZiDRzufGz9qwKsB0XbYkac3ts19ZbEckmbcbagtPU05hyneol8mUg89nWIQ9PivIGuwSQsjS
mQHpyCyJIZuMWeZWm+cKCPz/JMMITv9KrI26jH3dPWJqzT+X8HV0xTk2owCKKjqUve3PnRlbwZUb
wFYowvRuTxGj1UfT4hYuh8AL/QUDBtGAVriJzP2kVgP84pT2LRrxxvNI7rq03afyBduzI2IuqtCX
JQr/cp5nOwELQjXO6Xn7+CHx9UdN170oJ6iIcbFLp4Qhzj9N7ysz+ncw7uol6HOo2hTCnfUCGLcn
/5yBUHX1Y/HTJlCB/RwBcWUAJGSNaDzKclXwowj9FRSoGt1uc9nW71G9odMMiPcJHs8pNqnO0k/F
ZwUGAaFRHAP8JiALJTIGZYwK19vMzHO0jrRttJ0PCGk8KsrCMzxt59/3L66HNmPHiycBLH4a0w88
pcbRbjOazu/wzjos3TliweUFonSDiP3QlP8/ADn9i5M+cl89EFyIu3CnRxRyrJL2o0AEwgu9qG94
GPbGFpjJgVPqDhy1VY2IDRaTOi6FWJHauxNTSBMy4nl+jBI6aTM+guFcvvWkmNH8cWJvwg0FgWM1
Vsebczl+qUQotCRk1r+NI0WtZe9hbndCSoAP7Pxd2OvKQC5ycHijvJ2POaEkTkvPInnFLDhwKZeS
iNdXJ46b7c7wnftQZoDC3UwLCysrYysV0gsOF7X/wEOKV69HdiunQHnWU4iul3tauhtJlAL+BDvw
3sqIdDeUTKv3JY6Uuovda/ULekHRhuHbw0EIcA+eVC67IQyCQamX07eeMGHai6KQxcWyx+99pmK0
Q0TSRwotz6HHQinzY3aY0uCh/8plJTrFVftSdMmREvLs41T4cOh+aXFryAxpoywRUCVFNXUc6HgR
xQJnYzbC83jusHnQFLfYsMLkyLbQlu1m7/SvbFCTue3RmMyY4lHZnSQlG5GBnAU6DTH9KHL467h1
fNqt2CNXi3XHgxvsAbKzwJqQflT3QarKxdXuzBZV9l1s81v9F2yw+UH6fgtK35dnQcfZulihV8kZ
SGbjUc41tGer8e27zy2J/oT22NeeIsKdQOCTUUP0rkBkR5X09B22pkwl4Bfaraybb4G4/1cE/0Ww
7hlcsBddUdrylvHs5xFl/Om3dOmIxW9BQyt0YxPtRcrwryKH3/JaONlT9/G8dRq4M8hCfuCV1Jlm
syLIrXYJ2L8tydCrZVmnYy05ePmqLVbG1DfuQBldecTtV95b1E6tpBDNKQsNFhdFUfOP5d3ow+ou
B0fM85z0j3Cj3kW3mXnTOrAefhs2krytOp1pJ6/bzYJbQB3PjxaMCLE861OiCMDSr7y1aIS2v94N
I51NeSjFtjFUizpqNVpfAxRoaf4qZHY3OILZk/MAHcQPQaqYLfn1zB2aaFp912OnuXSnx6j3iX21
EA9vuSSMc0HHAim3tq/gcndUvEgUfY0KIKndU0dgyVeTfk3yJkwe13ccFQ4A2+uw6ORUsrIe9jim
VV0ptFRYH8JxlUbveGiKyMpjsR2aV0npLk0Fy7bQcgWjfUrW7b10atHztxse0+lFsKNAY11qCesf
XTN3BJ+WF2DywF2kHGvwtrQPW8ELp6seT8X6QzYthaDXYHuPyudWHFGplWeu3MjDgXN4bfGE5qEs
qVVpLtHcg1zx+mwVqbAe62vsqXNmiC4OWt9GemRWY570FykbxkoTuYcYCjILjHFg4LHV4lQ3HWSu
P53FXEdjn4wZLOpprjtkoUE8ir8MEZEOfaFEAVZNse5atuutAYGXuSybl7cj5NepwkwMsWy4cdi6
l1bM9A8NryE/1aHZdnzwc8eygZUYVvhhSN0oV3hk69PwVrR9lVUjznha0TkzruGkKhbZ09ZvU9Nt
hiW4o2MUGXJXol0t24/JnlzvjcSBTe4hbHrfv6wkWxUEhY5AQRyxPPvREVzayg6+/9R5r8mp2Wth
oeT2TYGpUoYyN+F6+SurrQ2+VaoibF+4EWkoabpoDdPMqIap8RU8lWL8SIQYclPN3ldJSYdUPcxN
MMo67BceV8P/qas9HKwugS0Hp5UlcbM+eNxxr6iJhkYL1LAfcwbm3HNzo5Ca9rZhjCTPghQzYYGW
UaRxnow0l5Ra9MfWKhvT5OOxmGY5C3BsLIGMicuPFm90MdnhBqi7EIzDwfK+h22ru1Z1hQY/RHft
GDgAWPbnHqR0SqZTFVCbAm0x0aJJVmdYICIe+z6pLeVaqA0AKgGns4S+gyQSUjtgH2Y/UVEzOA5D
lmh9h8I/BmohkR3oshwkAsgDSKrd9UZtWuTPA9UsEAJC8PaRsNt/dJYx6IJ7K/a0D9O07doZ/x/r
ipwRcIFInunHXFGll5CVXHHlcvpxmcl1X0XvMKEceF4+tT5Lsngf3KnRY9s7kFRzsfvizrwHFXDR
Tdc12CVF/v1XSH09elJIp705nHcJD4lChvOhFp6H/E4EJ3p0JWP9fYKbiWx7PcrFtJkhSpaEXbFt
vianpexpmhVVVU52CGob0aoDxQiCyfV2RY6uvxrUy74ddhjG1dAhPl05KoH9uoyHJHKoQDIYlE41
pRMgsa1/iCke/j689rrAJ3E4Xtn/mMH+DCW1FjRGYkTHnbD+yYrcF6cemhvcRk8fkNZAQ5hJaSjy
li/+FgAh7IBY+/JfPDOltclQBeaUq01MVAjWUMMHh5e7s4gAs/22qvt414hEOwLmLpqt/lBBvRjZ
ZthrdrvjWtGF53t5ZCpMigFVsgIfeRbXCtygEuBnoG6aA2ryu1Twb0v+8PsHMZlQzycrulRSdp8i
bSgK3y+shZiaegWtJENn5OMLee4n4N8j6BUyMcCAcrfytlYC+VsWLexAbtuLNVe+wQtbG71m3XZr
jF8FpUbn8Y5bD936lAo5OaZ+Qme0B5Omo9JbupfHSMc79/luOUOlskHaWiF9DJvFiJZqe5J0494b
aVSwxHAW8u9Yy5y+SOvrIJtamMm3B435DzLy4WHYgG3yOJxnhJ9cQ6P0UHCgkFkW4+Mueu0GkEmc
Fmrna7W5B+VahqNraj51zQkQ64RWXfyZ3ZPzcPGjlR3xZer2GMkQLmivkCDPg/uyb7AvU79WqzDi
KAtOKoCfDBUYkVLNJRo6wshaIPs5+UFNHhQYLgQeHDjK11W+XEfCBc1Y8ETwWvbfqXkPaTNKjTP3
wb3z+Iz2jIhTPhtyHwAWFqOdZQsl/SIxMD/Sl0QX9jix7oHP3UNYuXumFEc9gzDFVt/rHMxtgcEQ
WabUW8lF0RecePK45WIzUj+TlxprK3dL6dXOxkZlWRn5s/ycBuQ6OaTixQYl8T+m9wv4q0//bRim
IntF6ZAIcRW/3hAZK4j13FAOiYQAWLLfOFeaDWr5ArmyGD0quXSBiTWGmhvg0yT2BDLGTd0iEPAd
9iFz3zDkf4/fdP6Eda3I8ty2Aa0eCnOjyAItrUMl1UkZgZSBmMxu+cyej5CC4tkk+nP5SRij5oxY
ne2bU5uxdH6G/V73v4usaOS2VgnJN6fDxJMqRE73QoGd92z+yn0dxISAoHDxyAwkqWc0df3wqMiJ
R9GWMmQu82n6RLIRr4k3UeiNRuAizm3Hw1LxGpnppxn+uK6QMxetP1bzdR1T8bPJIy/CXdMnJB7A
MX121C/iHic8IVYSZjULIVsktxEOxjcV//nm7IpnwlBdhfvRzU22uzWhgGXHG8GhQ5+fH7+qtCZB
qbDpFUXRDVgGSuIud8hzUCm0m9t0A7ABwSnHSlfpO2348p+A9PWOw41Ny8IA9sZKxmzWkc4ffnyN
WcFcFnKE5dCXscZdtLqmAueAm3IIiOl92Ug0ux3EqTgwIvMpIqB7eQnXie7yzQYKB5EzaUrBbRTd
YBdpynzIC2Puu8FZFgq4oLPbPWLVosyu/HM64Gjs29oJm0ow6p/iVuREzSLD1tMNjmu/tBP9Eozi
9q17Hnkd2Z/Kf0ESlc7g1Zj9jkoF+OvOzP/rBuqA6gqO18pRVJoAooMLNui6YvogqwkhEWmEOG64
4lltbb5G+05QIyw5q9WpNSuBpyCWM8TJSX9foH8urBS3+BbmfcLg+3kOmiRXxBWnd3nZY/oaMrb9
NvPGDUD8XzA5DEQZ8097+IOvI428UKjHCuIbQP/0qpH6LN1YouiqK6UkY+phcH6XEenyHFRfbJJG
nSsW7xTzVZJwHSekr+7FAx+gnRUYt1j2u36ye4brFIjFD1GOtwvL3Lhlc+FUO20yvWNZPh29N5KH
qlsPVSTvdZblt6G95diH0L6zIG2pyyKTBq2V0BN9975zgB6gTikJiSXYqsy+g1/RRlsF2SKb4wN9
YPZtUJyxu9NNCJLnWpwU9lNWyNd6o2fiQyu0oxOHnj6ywgACsPP9xSUe8+39cbsx785I01m/Kb0F
tUlnOiMYOWdVwXUD0QORfMb2ntHCgb+vcnM1w34+vGoBCYMs4tvyLRNhhoKJEvIBU9S/yC+DDOET
iHq32qC/+HF/IJUstMXEHHU27Tku+ZO4IhytU7/zvE4u+Pv/YXcW/T67TvYa5m8djm5WKcUJfUnF
gMPrvcUFPpk3NCDn45BYr0DzIM3S2cirMp6M08Fp17R5DqwdXrqQs5HzhIyEUZkGnKHFUzz+P0lk
vTdIQ+C8rUS4Xcep9Ny07fv+vGgeNVgNWb3MTM94NrlJO3kK8XmGhzIPxCRVErYGYu8VX0pduDvo
x64dt2PU6M6+6C45+VsvzFftYYJTDDIEyagmjt3DkvqAhkbql4yq49d8UlGRgj7FHMDTQAn/Tnt/
T9GMHNY0fKfGWK28OJD5huBgFx/IDgzuVNEcP4oeV0DEq2eHaGsPMhb2v5mcPb92hYZ5EFgVP3NZ
BEYGLALun0X8QofKGxumphnBHdodr67M9O/M5wPuBAHBZkbevnv6vo/6Cw4PEbTk+ItXv75AGaOx
7eNwsT6ChRv5aJnUVZltMXCgbWyViVuvfLoNy8kRtzo+lNusE9wM+KsV92isZ4fIAzTaC0+KwD8k
/xdrD2JNYKCbCxJTewBcxNALr66a5hCNuFSwDny5RvwczIMOUw3/z7o6uVAhtWSuFOJYRcuSx7U8
hDgXPqDrjZkSwP0uMKjre6kykgvNS/YIh2/diaVHoCkz5nXA/mbF4kJ3jQjNiQbn4dJxIx6lbWhB
4f1srybpv6Ki61BgNcJCpO1gLoiwCEDoscQsUVPPhJ1oVBwBzUy0NojgNtnvYTOjppLuZqV5JGCO
uWz4LD0iX23StpYqqayBF+4+bbFW/rldLXkYZMJUH+a/olTkiI2iL2Qz/iL85wxdpYe3M2Ef00Wa
YitAg/VP3PAdB6bZ1j1mP+Br3MJL2b83JasTpAm/7vlunKEV7aldTe2vuWh7iEH7RH9DKpHd4kQ8
zYfRc6/zqrax6To799zUqyEpye0g5cbthLEuGOUeioOiyc6EnQRX3rInLWfrS7NCvSDjuFUpzxvx
Gd61H5H9TMIWtfveoWFvwAfdAkngEeuUNYJ1R+UMgOYSbhOdDrBAqhhYy/Nx6kdImY51MO08+w3O
YhNhbRnH4PqGtDSWwLgPYTs5KTXdCRdSEXeaRdVO8ofj2aYQMFgTrLltu1mWRTkgpgPgXenK4XR6
oH/P0TdcTDkrUrKqOWvL0Nnm6PboJ/ba5vnBVnN78qxlqjI0bMqRbsKdC1upOy3QjtXvsj51ZQ/3
VK1qn4n3FMfWLHxiHxKses1CSLWIFuV8Xbht/UIGzb1CYU0QuuD69Q3IWx6uH2rJH84uab7YtUsr
liJMPEwQlN6FHQQvT1/f05Y0SZy4yMIE050nxjRa69RaF/B/pf3jSxt1xPw11wlSssGo6gzkMQoD
HK2+qqTgDxTAtvpbYYjc04Eaw9sV0ITSB86ssbefHINR72ipxbvS2A/ZnUR5xaagZrxXpkAIxIEC
mRjLFtKDIZqLO5nrosC9dlU6SNJVauNc6RLDZc5wr3g1Uc8czI8duC7DSNKgbZafzGOgPyvJEquN
+QrkMFccc3ApRbQ2YeLSukLTyhvq+T5E9SwYhDraHneMY8MzpOUllVOEGim6ZzcqFwQVldTVIH7C
XrJodzjc8sb6InEpM98P/KMJW7wiLHradLzAsbBzecPzU0lvby/ObwJpb7Px7CbJamqI+TTfnzjU
YFk0aRzU2QP6tgOM7qQleElA7ATG5ukci7wcF2dhykj5vvllgB9EJCoT7IuNLuDzAf9JaBSuSD0x
t9jAEHTo7oB1X/B7oJVPOoq8IeFPaXgwWwcCAJ66DUUykQiZNoAdQ5htnVzy12Iin9RBhhY0+XnA
E4HVt2c5/3ikD7SoEQoCux4GT/s2Y8pC5o7aDPnuS558VffboVQiLTXWmE1I4+6NMH8et85ItE/E
9iGUtEnbIzYzTC7OFaoW1ewKPTA8M1O6oQUPH9JaPnrdExMxwBpKeQ7ViAGz5bU37AqJjU2JzBev
1mpHST6w8XNFqci+NC2a1hS7q54f5dkwFxciD2ndqu/qvhCFAVuQJOEqmVPbRi+OKIfK7FC7acDw
dX1HVU8RafAgwnYeF8zrLX2uUa5ZAV9/Hf9kH0UcSeA6/gGJZWdaS19Jr4rkHcd0RPHdHSelfE76
kvqHzyxc93uFuJBKMfEY5gz/4LKfiTHBuYeXh7Ey4xMWSM+CMGjgK+tImOIajY5cpDtl2ELl2V65
/HWlR7dowjKny3DX7fKgCWKNHiI6a25KhR+KycX+gJUTzLMcNWoYs+ncSe8kQ26aMaiexWxkkaxc
1bVTrdv6UjYCkm32qKyLDghrGGrDT/3Q4hHzt9CrQ3B4LSE1iwK8hfD0eubj3d1UDB1nt5y5KojI
ydN+X0QNJqn+/wgl81b4HmNugl9W9UaM/amvl0kQ2WZND21vS4Q6iBHh7SJ/4liEEZlWMSZQugBx
v65txjqnEm8ntensBBDGAJKljXJO6+2oL01EoQ/dvhgXKyUHL0O1NWcHgLsdmHnMbeers1E+p3n+
jkW7o8twlzCJDxQT22ozkUWdeNeCFFVgdlwd69Fnl3VuFyD9fdZzfoRb4tBIr8a7Bed1TOftrmqI
bUMmnyinCK7Y3fs/no2D4uxqmZIjzim56i4Ny/P2WywUnBFbzdJszs+OnOvcYukHanSsUMzl+bP+
Q3LBjosaVX33mqMSQxQ+0XlpdOy/A5ZG10WJqpKLnNVMdabhzN0CPgtRZakz+/JCYWIa25xe9to8
sW+AwMY2h7SUdmV2WxTz0ui7yRz/4UoFBuV+UCvKZaZ+esPjXgbOCBUDlY81OdxVh07ZbRhS3O8s
LnA8DIAW/3jomnaupjxWZMh5reT65NSmT4U4n0vkIFwz+e0hkZdwqtVE9fypeLCKXSp1Mcee1+tD
15Q3D1olmmE29P803j67s5YotMes52geWNvtWR2f/9X22Q00BTNFM+kbjx+JB324R5398g1k3Cfb
Ge7FhECgrohVATfuNBHf6YR7GOl2DlLfM0PXquMjPd9Ahw8q3E6t9Wag4Atzoi8yaKXi5TBV4LZg
3W59zuRvxpOeXN33KS98+f+E+aRG3LqsreYiRHQnVe28pmsUAox+DFoIF2i+OnemEJp3KLvcOh4N
M25zD1zBOfzUARBJBqqytHgzdmTMf0JQWbFv99nql4Q1B0RIdBt1Mhzt6fL8/vpPYpSWuFF7nhrz
uAZM/jrS5aDimvW8+f4pZoQz71Wiw5M8HpVZxGTDttiQMIwHH0v5jDMp88BzUXbKr9NSj6nedJ7X
29/fBYPy5Grg8TXLYIym0gzroRRO6JT1emA+HFWsLS+NwueLXosSmXxhjXCXYtVi1oLGJ2RHkXlX
gbY36oq9Sa08sR78dVFlc0qp+W/5RUIoT3FSdaJ33ms4BQ0isk3bIQVwpmPwHHFhMQ7rbmJuiFh/
iEr0YfWSyC8Z5DQVkMr4sEbLHXBUzYxY5M/dYlSvLSgYQRHWAccSi/LefkrhhBKgiZQ740WSZlnt
v4GDLhCEAAiYgY0qcBdHPn46ZV6k0hprn48vkdOj/Innfrm6yu92ey9QHetcYxeoTGLi8WHWMqw7
lnBDQpevcLjLe8mrBCty18IIj6xvMp564yyv2HwgmeWlqD6sGuxL8RKaRfTC2im+MxvcjZmkq5/t
KX5sqxIMGu8x4b5o2oT94PWY1Fzep7Fpa0iouiM7ElPiWBntd8zVKXCL8mogAnFCxgue9giddIaV
hsEJTpXyOBSiGB7bbRBOf1d3zkuSK/xVcvMOaKy+/OoI9XzUuKGVCVSztEZ5SSKJSHCmkFSCNURj
vUpVdWZyyGLjcdiaxrrk8RP+/V3gXBL/C6xqlGcqoIeeeUCCpCmFaLun3crAba7mf5F2R0bWF3aY
iViIk/XR8O9erb/tilF2OJbbqPuL4r5U4tHb/ycs9Csioy32F3W7Nq55cFdf0I8uSLjW6AXem8Xj
P95DlW0Qfff3zKr7/WL8zWNAvvdTp0TtZU5lE3S5hrAfdeRYSrIuZKKFuo5RSxso+og4/tSVfHBR
DmWOGAEymp97QAJRvorOpZfj65IaKTXdpClTXyA+Al8MLMnU5ukWZnftfr5ktJXFOY8DhlFVsmtY
qGBN7nFlRPLxUIMkvraBDYvHrUO7BprZjrrHN/ZkgGuDOoVvfSpBtYSxIdrFKWGFvpDgKehj8tvc
Aqs9oKC/yDhpLieUdBxPvVw4nsGWsvYHtcc5yWK2BsaCW6gqj2KiLfmUC/ic1xSQBuhNnqZRYHlQ
BZv/kXIVvcwbgVh8d9E14LsbZ5MHw43gEVG0nSrVUI+ieXI9DlgHPDqu67ZpYfGaXweWPLHYhQCQ
Nu9sJpgj5HNe1tETdOxS37ExXQN8CvjFqf1Xff+BI7jY3UtBIJpOOa3AAvN7z5ITihSF91/3LOK+
ss1vNwV5ZM6n25GDcBUKmqdB2hCOef+qoQ4yf5S8oHfXUAVi+xLREFyDLmn770ineH79/X0Rzc3Q
QDnhgXz6P2Qy23TqJcAb1n3WgI+bHC/DUfQHEYfnmr8pss108slsSlUydymJn7/yOThpyU+amed3
ApqDDWqodD3YbsPvBwyoHCdDJkAVfY0iCN3ZMk1RE2SRVQ+OqfBWVfWVfHgPGRQPUgK7tQBu7N7R
HGfVG/ktYCTfijIku2ZL2M0FwNpIii6C4X7gA19UXofGyRmVmbLeAJEqZQvOXJpyUzZrAaMeNOtQ
B+trdExuQP/4V9KEHdUzPJD2frH2FMw4VhDjkpap7D0xWi3wvGQflOQkFuUKpQepiuo6uy+DMEoy
dBnc2aYW7RmgzqGGLd06UuLRv6Nbievu6QjTkldzT3EgqcL90PVRRxATvB3unabonEZgK562Mrah
SFIEO8x1GW//+Arp5+0roq3EkQOWLdflyBv8run/bn0Z6tnUWeerC1gV8ETtjHEfV1aM2FPRK8IO
WzkKyeiH6gfe59UqUDEDN4NnYfrHm1b5V4TS3oTgOcXSudsiZRIfW2o947mlGLnaT45TTD1XEzMS
vIAxpFc1poXINCHqig8Dd9JYABCcKG/7Wed11+IaWlwHuhQ5gGH7o9R+sFOOrnEXsRUSezQqqrJ6
NX64DWQZH4GGyTX+Ho3gjLtASyTzYpd+RDP7T3rY7h51WV/LQEpsyPEHNtgqi0pl3xwg6QSbHIwD
LiDIfiNsXkD5s9OX8XjVVHwAs9VU5gk64U4+LOzYTTeNzNF5OK1JveEe/Pu3tP3fe0d8IFjNl9Zz
7kyp+UJwHLiArjhuhakYTbRGO0uYng44wZ+4RKNXTIImbmTofrjTCf1+o11dYVdUIEXa8mlYEAM8
uf42N4nTk4DoCNrKtY7MeTMikRgKh5zx9aOZsUve3u5YcAz2CoLBogZKEP/fw9rpg2UQ8u4KTtMb
TIMnBcnpCRo5DFPkczfZK9J1jDK6a34qpFS+fjxzdxEcZWtknmoDGdNJnayJOOjzCgzA3nBE+e1k
mju0KHOTY00fGuDnNJQdUpSIV4s1tc6V1soPwVA8dOwfAiEiFY50IIlocPrXWaw/V00ry1dwNpXg
zTKzFs76QnxUWaLnyDoXaP3/bdRBBXpYpD3avnumaNSev+TPJ8zwoZVZuYELgfYCQCT287esHcJO
T7B3cZBE98QcJC6zHrJHOIVa0LYHFBwVtnB+d6a0KLEBfaMI1nbjNTCCGyhO/WmDK06zC2neoWcR
1BHW/z5cDAphPYFVlEVNx/6ZqN3sqkq9iT+KictuWppTvx++DpZfIa5QTizVpiyZ4pjo6Wzm5UNS
S94AxDHdGjvfQVB3GEZCWBLrMAXzV4SxmqbW3ZhJ7hVFLfx3qu5IvREPd04XLXVG3Ce48f/psLYB
Lr/aeuMHz5K7QczK5NdKzGarWOwSgVka0O10qYFvV+M+t1e5Afp5wRfg+XhIPP0NSS2MuLVrFvSL
Yj9iZ+pPjgLV87/FDtSk49bkzWDM7M1KNtekJY3UboA5ekYskwlEUb5g8Vw8K5O99P3AHUtTuwhl
NV3m5V732s4qj1Mi1ZRldBxi/uI4UhTEq4Axxxc5D8yU8NNTm2cxc+oB1U05oQ7xKrjhVfLHiUpT
pYtL4HZlcAnvuZsLMOjDv5uCs2NRTUzklqMmmj6YU+BSyJyNecv367Iv4xc7Ee4kEGAdx05j4mf3
zOhaCnxhkwv1BhvexwV7DwZrwdZufSrjrRCJtoWevF7QU5YKostPAmEazSubD8lbFGX5SabS1cab
2UWDdWpfxWh9mYLDFRbXEP49GWfAHNo9gQZ6OinGQbsrWjj5lylGmtiIgZNP8rPU0a4TO8GhLs+C
MXi0hz8zw7Plx7aGiAcXSTtyJf8cBywmtNyFHCN9UTrX8VH1uAcyt+kSf31pMcnMxBXjYD5uIF8p
xMkhyHfUxrrXhO/EWUU/bgB66U3KRjdBXKCot/Bi347Fy1BBBeSj8uJRFVi27Co5srqz97y8L9SP
rvs7HG/ao1xyFIWGItVD5A7vd8Tok5fURzqHMoLq18+LKRBHOtuO2dEyQ4pubCUF177iJeQHGETy
zuEvoVMh8Am7Y4hk6NOvxNpsNpJfC5CcNoxWAxsf8/5fNNHVXBMkRDllROTQ36aIVaavtphALEJl
HTToVPf1nYeNsMyXcxAOzxgulXnA9+FS8t5pn9/0oXMJAsanKI1ARVHLUS27BD9We5Tqy8RTmdkX
yNTf4KLSwAp5yic9QK8C8OD94fFY88SFjJBVjLygg8iSXgBq4cbHvrw6DweIvWuh+WRBkxQYxbQx
eVWE+BpwQn7o7SlXwNjE11Ph6yNqeVlwfpQhi63xoZ+Br2oEdP7MCbwkQ7sQPuZ/mRlbQDaWoI6m
IgVK07ShFnC8iASgWfigsCe/oUg2MT1yogoDcxrUQyNCEKne4/upMcdW78LwSMjCwQocsGTFXasl
AAd04sdS2sQjjPfj56anIRYiU3JhVBZKRItd3CzAj90YrAFU6d8f7yOv86ichsHpQfqi8n/bzvwK
VjmzOVK2KXmXBP9ozXM9KE//4NYaWK2F4KKs6J7f0OG7zLziK6/7rKByTvXlOryKLFGOYcxXBCMu
zv6dtf7STfK9OljQIN5gwpRAjAFoQniLBjSDDfLoqhzfZ+5W2mUJl4pgZqnBn9QAZ2TnyVlh9ZAO
B87N+vCyxhFQYJiCBh1oCghg1qA0Nri9uy91WacO6nMnWV2cKMrnR/mjFijwSn1eDqVvwc0HGvsi
7p3OHg5+8ekbMuVh53d1/y3j7jPplnW8ienYGsNliAI4gcp04dIIC8wIdxM7lLCBvQbQWJrwJ0bw
wxGQ8CkNLI7HzNhfvmv48tsEuB87zM81igdHCjbekTG+7NQGjDHdKJw/c07Snmzq9DYyNVQ50LNg
/K1ylcGUkBaA8UPeodA31IIutcMbX/GkUEzYYqcCQ2u8a+blaBKtEkxifG7Mmj1sxUaQz2wqIDlO
1HIcclCgUIr2IUo8RSgNt3aIP062hDfuhbvpNpcom2+maLHNY9xEYilaBCcO8z/7b0JVPDar+ewd
37B/0joWlFkpo3/7k7yUcY9A8rZql2b3+ctkBbi04vvdNgKtGVpd0ZaKKIxxJ0HZ0Brn+s2MhdX0
FBNskOzC51hMrfJyMMlCuayfFcT8iVH9SVo0Ltfqk9qzP/BGogY9t/6kze6ZRzAtvDN9kHmRkbEc
Aaadvp4ENkynKU0Fk6NR4/Bg56iqmNwCiBNd8CDpJzD9T5zW+GmEcGU9KDR6Vkv7dE5jS2MHlWt0
IPoWur4EvIDDCKXkb5ryKVpW4lVrpraaak9vzuU8edFxwiJy1CeYKefVPFaLPgOWYdq7IwcJGmCY
XuQk/yz2IS+pkX+MhLcdvTmHCDYRpB7Kaf0iPV9KeFN4q3F23bZk9zlRBUaw3LF7wfvMNUKJKpau
NQT9YUZ2Eejk1jNN1zOBC4pUP4tcieng4oYdSo92Ad965apdxPLcaKYQB0HHkjqS0tRTSXt+6RIW
aqDxH2W7mIVU6sxf7bQxhrQl1DoYhj+cBa7ct8kh7YeMAEfGjtXlSJ17u+2L+DtKoO45MHaSVd6+
UKxJd8yYAjQjTrA0sSYEcXAWmzBrJrGrF+fhctffTuv9y0/FlbO2WxuSKo36s6sfzst8BBLdsSnG
BKxc/SEz2Ldtz33vWp1StjswEfACiEO3iS6/y+GTYMuSR8kP5OC52sLpmiXUBSZMiCsDM7D4gu/Z
1PYYonAhKOhax6BhPMALpNts9qLTkM1GUscRrwwBSJoz2A+G3fFbC4dlpZdgl3YdkkANsOLW6eQr
9vpY4CN+vTv56nCuuKf0iV1Ix5kykIULJyIZUrAuyp7PUlly7uV74MH6bZ4rbTNes2fzQhkwXqLQ
T2sGC0YcXFyM1jOGLDRalge69sq1sxSX0tL/D9vs4HChPWLegbqLuHG6jetwBU1pDC7jpcTnrpRc
gx5OCL872Rb1wZM/VqSavm/E74Gfb3T6QqJQRgzwJ1Tv3IkyE/OJXwTPAJh6BqiSdpYwQ8WYnXRp
7ptM7Q0fw2jCZtqvHii0uYAprC46FyY0zFNTC6DtOFe4uGTseMOw9BkCF7fY+WkndDAJKYK3IOdI
48iMKux4QdQcCHBee29JOz2vuSRpkkya0cSMo5P4KkaQvFlKevnh4Dslu+Io/bwE4qWQmkLsdntw
5dEKNdQC7HsatcTMGfBQtd32a0u7Itr/sWrZ5Dxlx3Lw0E5uI7JxfKD3Hq1eaO1VGNvJOpA3Jojc
jR/pfQ6j5IM8aiRx8rkvc6VPr9jTnuzP36ROsSoLg9ismOZgjXQrww90lZdvyh+k2UZ4wTyIg4wa
eOEOPz7dVjXkycx9V+CZwiakiBGvzJAo5G2OUf+KXx4LENMW/0j89pszHVLJc5LnxsVK1IRGyHQm
Yc9IbbgpBawud8HokeVic66ge0M+chBgp2xwXYGETNrn7TBikJA9LlNyJy/+7WXVR20tB2cpkNM3
b87/7vVKuIHLOzp+vnfvFVnnwu0AVENDIp5W7qJOP2b3D5Bi4B066+e0xAyhetdhs1Rp2hO8e3Ky
2DxU7Hd7Mq01ufoQeej3M/9BcQKxo/Bs89eIASTlv+Tm7YnqcCET+eYimDe+179VmIayE390jJ9K
20MNze+mSGLCtUFBbxYO5CDXYUAhKcsBFZn6DzgXTGEQYTIPz7xscZGXaFMBRX0PYMGnktoHALis
YqsQxtlVW3Hu/MImsfkldvldBf8ivntqoNWNIYSPvvnJdh/EgetYe7RjIKlXdcHnqo/Rhf4dDH5G
X7lOS630pBwwyZeHxPkhndFvegPNWZre2d0J6o6bZq5FsCiYXYijKOcBBsHioKQQ3cdQb6wN/JSn
1GCRdUEJJ9TnjYDZcVWYyljwL1WBVOvqcGoBZTLZfVm844W/0zsK+WWve3/GeOzChAA3W7F4Vncj
/0DUZ7iGc2n1njS+Z2e7yrdQAis+VgYrRKeZS21BKsddwtbVcU4eh3ElA13MYe1klebS1+S0XXTY
HfdK9EWj/CVsXylzm3YVOl9G9Y5tmayxgIHx5nehC43G4RcvJWUiBNB436kosLKpXQUKrKCrjxYm
tW9XUu/nn64Us+xEwS+Me1KG9US3e7aOcvlzGzWUJVjP7xv0AaYX4Uj32ShCIq3/fc6cBEjKxLn4
k0a8v2z9xkzBdXVu1E6HBkVdEDiHobLgK+5oS0S+wCKSEn7QukIPZhcpMqab8gJP6BhevKycIAIL
+ctioizqG6jS3pSiD7fwKpTOxLnvX1czcrJm6BuIue4OrPC0aNlS3Q9bA/msq+iE6xrsKQF2L6BJ
LP9s0x7Getk7IaMrKAx5393O9YvyoDp9x7k8kn2BU7mprGpLo1uwPjPmT/PLreRK7jRbUdSnioVN
KJfE7QD8EwiaOjsOObLZAMFXwmWly9DTMdWYzDoleKZpTERCtnOwzTmo2pUMREASI3SIS+rdGLSm
Oi6dgMGpnkY9FYHkAN4mwZ+s3odx+UrPglxaJA+XgPWkwKLlENV8vX5cHghDK+XG4zo0zZ83Y6J7
9Cfx9mku8qQhwSzrY18C+Nj6nS1VZEERz7C4lL1F4lA75Kh6Ny8RumhEqJ6vZ8mSsD0Zl239W1hJ
mVfK2xNYQESa4Q6AkXv55W6WXOU/7+A67wJmLpJkAiT7xpMQUaPvOeb/aiRfn9TEtcmxZkPpbzuB
ukagWeyn3oJoYcSAExvlC2y3dBOO0q8KdVJlPIFl4nsrEWtmE5xFMH+7qoCRlHz+K/SGOdjlxg3k
rr2//D7ecP9LA8KXaober9o/IFO2mWhgNoGLkTyYFCN6iny8uYoItWt7xprHASEI4RQ3ne6ZatCj
03TNCT6CSTGIpRWjIyPIARJKcy3P9CHDBJ0WnLsGPsWqpkXwqKR1R0OilOd9qe1zIqUEJMNY5A3Q
J1oe0gfDIcxLBSIiF+MolGmhWm9LL2enlMtZo598w8q2e64fb1xueV/pxmsBhNNZa/EsDq9iC7WN
qV6pElW5fdUkdZBmjiVnTbaBz0/WyhbYE1lyoW5dAUf6CpBPasoP8LCQkKvQ9HafHQ5ZNLko7+32
wgSnSR08aq4Gf0ccQGICl4xHJWxugG5htVG326jHTJEFdTGQQIrNPhmwBbqx8lMEA0hrKgk/Iawf
JmsgDczpo7kbgmzxjengi8yUixXw0BRhZN1MIO3NlwZVCXLpHbA3ZsZdutE15JO3+qayafsXTAZ7
7/eshE4wvb4tXO8TSLFGLHsBj1litw4fdqhR1fL6a6F8qPix2rsaUyRwhqD6O7Rx/EaQ77ewgJTQ
5TBv8BCKWxnLkJthUuJizpDp1XHeVv0J5e5hrYRDj/jqE+2TRlq8on9irGdn8sN6HL2xL+N73oFb
rbIMBSQeAzJnMskFDLpZj72LEymcEAsXjJDGrdDhiiGsAN1zx8sw4b6alP3ACLtIVnAfSSoyohnW
eq+zGv4NSDVPYw+CSHB/QUtJ/cbo7cN9GSpbRZRy+rFbAIV3e00JE8sPgVjq8ibZoE3HoOLTCYRS
YJajcfabr5HUhkjNyEWL4MsO1XLBy4CYfWZdHC5zwhkrkRvGXKTQqqXygZPJaXUgAXW7CHtGVRWQ
SFTIedxUcyoxgt8fenQxyZXPKePWk0FTuV267CId3X7kv443u42W6kaN4ulvLES/rctIT+yt+VOH
mZH42dPIq0W4Rb3m/1aSTilCvPT0HPcUHluW1yv7V6jX75y8xm5mP7xGMRjc0aH2GaPHDXJfv0Tu
UeoBdTAUjjrgA2WdM4Rz7YOQciVS/Ron/ZSwOmS/4kgaVzdv42WETC0RAFbYvVL/s1Dv/DgzMBmt
eLFy/bP0fal4uUWprGMJGOzp/D008Fb1BNswAGGmk5djwnkdt/udbeGaCJTrd9lkaTgkM6JBxzxX
b7kyMdg/sDEBZ5TqlMov7NFyLL9V6CswviKdyH3MIOXLOkSXAEg4nouNekM9l2LmpQ2e9JcuqgMC
s+7ea5uMXNiQVFUhui2UKwktaF0Y1oxx/2V42vKFk3jzcLtNFjguURc9YkajIJ+sT6NbxLi8aya/
6oRby++XdRu1wPsEWjAXQKubvYGESIGsQw00Lf/OylMGqOEm00fdPBoN8jHQeUfy4j2JYKfeDVC0
yCefrn5WQsWLtzrMAe6totA+j1wWBeRRusxnc2uJd87RDpAd1UyfMUQbPRotYTak2DZSdbI4Jipg
lOPpI8dZU/vJ7U4nPPZP1XVZXmxYfEfmRuDJdyLO0Q9nSIFmOQQ7Nk9Ii0BECpN7ycHJr/Gdwi31
+/TjAKt6eNLTPQDmz3JrDU1TseZFM0XvuVSP/9MxrdkKTR3NwXaWLv/JdvRe6dsvPY+NPVIz6MOE
vG21mLIXkwAZ2A8a/id7/jOXjDudMbkTmzLaR0dIfvTiw2TrbkR7H1cmtEz/cSow6LzYwqJ5kwuL
ZDSmoiOTjoxsqo00kX/zNsFDDi0dKBvf4xGzAtzMHMw2oce7dPVRSgYHQ+pQ/N+F4SMLBIuX12sC
77jNWYwaGCFGlA5jr5VSQZ9doyaOwMoZhyOhGD+9d3eR3fxy8szqyuqbBJdTXUraJLv5kvSJKrMD
j8Dh3VwuZFS18og0W6uKWzhYeUfPfWAYLtHBunxB0VzCk6Qqi6WqQFRe9FPtfvAiXMUNXHFC9zTo
VW8A5GKMkkUb+wSQNUxmwuofNjQoS61mafL73hHDwloqjj+bq6SK2bghO+T9J94UxF5beZOY8F+Q
1bX6vGHmmOAvUXSzsjnck/nz0R40u1f2/mPfRqhG8bfj1AEHTmuRk8Kh0rN+iltGstfxrbiLzomp
sCQro7BTdRD+E2g/BgSoxpADZ3ly29UHYF6L21kAliI0zqrkZo8ZheVK7oepUmVtAtzrOi2xrkyA
ck8UnCaKfgejv9NxrbamgdiSnqrW0S4poVb7mQuJ4pZ4uTg3Lyv8jmXU1zpD+WMOolUO2tIHcG/d
oBZUffQ/2zUaDcdnpKtnzjI7qUJJHknhs2LLMvg6AvIoGXFkLrJTv0D/G10uiaBfJvmkLo+07gsd
gKJcl/cMQ9E2Irbc39ScgDugsyB3tmsW1evvY4bbmtGYSRhiXarWdDT3JjhF2G1d6a/eC93g2Ilt
r8Ao2NNHkmwfAAgKWQfc4DUvIoxbj3x5894kaTLWnLuVDiZDJ7a9SEoCj8d4YKMQWvS8TVpOvj8C
qaTE/GBpqoGQfHt1Nia59co/IhuCV3CXQpDmZ931miB0RzT5/N0S2AIL1bLgue4KdYHwG/R+deZ9
qTsK+pEtm7syW6dVDAyeMMHSdI9W9jWoMPte37g9kK9Xp608B90oWNjxIsd4AyLC36R3Knkhy6ti
NmZcY3ZMnqpsThYNRgl8ELwFrWoaruyJniwNrngZUDanRebPvbjr2ejrOg4J1jA5o0PoYZiR6qTN
gvSBh5oH1413epLrP5poOTem8RQ+KkRtMC6U5i4RlaXFuLcSS8gc8mLpBjl9YVdiHK2K//8xGVeT
nyRIOf4y/cTNRRrieQ0lJcAeP3dN2sjaWHsZLxtrgv7RZ2q1ugtVET6RvkEUpRXHnFsVrcUEuu/3
Z2xNycu/MQsW2HSBduy9+2wtxH6Hcv1o4xL85NxPgYQcnlw0FBqjZPaJ8vd+VQ4A3RHcTeXVsYdq
o7QaUAnFh/4SlF1pStszS8NjqXBubEUoG4OVsR3dpDXg1Twj/de0TGsxd/OrMJdoOaREhnNiR2jJ
6whTOkKveH9t2hmMeGyIoBqXC8W+ZQW8huLzqHL5cVCzfMxATo8kMZnn/NAL7/cUyfHN833vrP5M
wmVQj7ktdUkjnCylROe9+cz5FX7zoVyXFGpKK2keUXoVMzuXoA1LuUwpgKvhdK/HDUikELRLAUCN
543ULSBRCPljOq5YKJSJmw9EL86y7Z28w4OJAKHsMiyKqEGsF1EaQycPFUGX9dwf5lLhUJJAqTAj
t7WFjosIX5XDCt8VOSn7C6xc+Sy7INpenPSO3MdnNqTEX5CFpbHlwXpJez2XZOizKDyaltfQh2Cj
2T0Oyk2c2zMKv6LYdfHmcDAq0QuHplG4Ns7GKyv8SdVj+JCDDUEKyskK43Z/N231WG4K8kg9Yhix
Q90//Eb5zMzR4OdOmMhXZpwNMZ2dBl4ZUrOeec71uPegHQH2sRoQQJNUQ4e6wiVHZZ9Tl3xUPFH3
fsfALQ6fi/vwigCEBMGvTbwEo9px+ey5qqOwBZUVHv576uNUYxCmQlvS4/2YQYBmPQFhLHH4mEdd
mv27WVgyPr1T9icagwKsMmNtjANpwlt7ztkhsMgRM1I5GRwgAjt0enkZ0yTnpvSqnOjgEvjdCIuA
yrxg/AlsQpFlcXDoOLsS44pz7Dq9N+qgoNQQZlG/qHFIGq/xIxseAWwJKT+sUPkhyV2z/oMxvGBw
xdxrfdsxu7jkiuVK5eYxGfYlE90ffKXf29X97qZ0aETVzvsaVi0JFv58ayd88k9+FueN6t4wV+4a
PcncGwUvjKHU6bs4eNTgHAwLKVFheT7mEiNXEw/skqZIGOAlz0IXk71CWHGg3xgOxt6qn3RDqYsl
AuD0cnpyZYfenMFE+4bdcp85/a8VAslqvk6pKQEBIgw3KKEhLdKCqNIft37KyOzmgfv8srsBsnC3
u5fugQ3iX/FHDQaFe1qIUxeZeUh6VBb5y4L5GdaeJotWu4pTn4lcMNk/GMkZ/lZX0S5vdnvgDQud
dKvrV6ztEO44BUcWJJtPzLDI0IEj0emdvUlNk3TIq/DoEZ0H3TIyIPlKBftGwCo1LVP1KsXJp9Qe
W1Kn8LbXn3uili1t0fAnCAs0A8G5Ze7oX5L8QvhOPsD0MPWsywebKfKROeldNiG4Uxyp+hz5lGzT
Md8atqpI98Skp35Hogrd1xoWxczGafaQ5/lQOixm08n0s3Ab7sSIcLTucQynwgUAnqk8LBAELCqm
rMDrWDYLtbrmMw5IbQCpC+XnoPz2YSeUyte3K44voHf9/K9WCTwVX3gLiIhd5NjA3ubLD2tbYT8b
vp2RBW8yCFViSYZabEkyJO3TJ3MtyG6nQRcVKiqn2UQN81M9X/OjmFp+NeV4EclCu6fTOLSeEnZf
bzBERvOxIq14x4JgRnSMszaD8hnmYrHsbAVYFfxgpdjs5lBB9qYpoj6n0UYSLihhZLBC02BbOhdo
DJ0c1lSjzpF+iagu5AVnuSathrRp/xk7+b5rH5/3uqJ75LOUHaQdVn6owpFOo5iWHSKARCL7XskI
TmI44DoG/k2k9rr5WBEPdXZDYsgqrvxixXcMbTUpgx83Svlza+l5HC/GDBnznVLHj5MVfnFPi4Li
XoZQaimutcsQdarmD8UFM4hvi4K3/KS1ut6Cp0RAAV+s/cC9B9pFgz3lhQmaRNnq9xkZnCWSiDeD
9p6Iw8AK0k3+6Ebqbi8EATNrF3jyEHuRyqyClZvFCyQeN54/Tih6Htr1igIjPk52JeRUzfr3B2Z+
TM1WNmQnRm4+RGThgo9anSHI9utTCX/tQ1/ZdF8WvKJIHnMtDkqPHuRMDphUFRTAmFhyJV432u1c
zvSlfg31g4lx7z57BWct2SHyPCCX5z8d+V+lbipK+ZYNWgd9qryRNzvw6uodDAtE/OxnVVLSQ6fD
YlUacBI9aTvgxG+1aAL4wnuTV/fFRZnT2I/0B0Vj8rmL5SJTyLbgesVxzClfInWzJGfDujeR08cC
LJp6cc1T8C1LGbumK3dZ5+BeMnaGBfk0PN8l3rRe95kavme55z5JA9B5ZMuyiuD9pXuSc8evUVTs
5n22bQy617CeZPrK8acTnU6boeAxVAB4xQkK3PeMa2u8vUhcaSQNacfVOF59+vJUfHGPaoFLCiO0
iiY34vg3s3JYtQ7846eKlsr4hjReN2rhVskZ6TeVoOPMMw3culVTbs9gR1ZhETmDf0jDkGTEDzgW
cGwWsm8kUpX/E1SZbawLud9+bCKqua120Y8KPOPfHQ0GGxShEsDe/wsWnJUhBiEac/y80DYjf/uN
6XEfGxiVGFqeKmY4dDLR9isTzu5v93iB/RRcw6C7T9lokFIid3GzH7l3g3wwCeVoEgaZusbSoFKU
uUxx9ji7KminlElkhGDJQw+naqCOzLrhzpmGFdygDAWYbbkBuLScUiMEMXmURbZzOYN6YKU2YMey
V32WlutXaKme8ItOQFKUsq3Kuw29DdG3CC/Nbij5GjbR0NhEGo0tBde2AkX5O2I6dapS+dxk4dZd
eyKIHJW8x3Yf9tStsKcBroFZmQE2+IPNLC7BA3kN5xDWtq3KUxQZZ0rPzhsKxBDC5H/VDlBGIy7g
fcRZFluOvsI7OqrcgNdAZZpa2KzIjsIeQkiC6iTpFZP52xZPGeMHCNLdR/HVvb4RMQVA9G4TPpxe
nHXSM/cBo47l0u8ICOxPdt59+sRnmMS8ssJgncZqGfCCrqF1m0NpMel4Fx75VCU+B1iKat9DhgrY
KZWintno+sTmseSOTqkC1ujC3EELAnwooLzRBMKGVajwPtgNjTtWman4GWjoB7KXB9Ir2xpylrBJ
eSyDGRZdDOJey1JvFnIWitDq9ltDnbAVMzI7cQBx2YS98JeP9Vm3X/xoKgWFIjfjCQLNiutJEy0k
ZS8weoEYdyXUnr7rEi/QVLEVkt1wTGCZ/1TuxWAt7lI9DdClr6zS1MrphziF6cMExi7Iet79wtEE
PfGBZgd0KRp3KOZbam3Aqeg5ms6FD4RwTIMtyQytUmu0WdLXsEszSKwDqpjRxh4uHkA+BX66/4CE
xddMsOLvoogaWXdPNK4X9XNHhZhzbKEdY9W5X4ePDHs8B+ihWO6o+qr5zVQIsPCwKfVmBtiu8Xyx
CxPH5ALVYH9iuDcCWJvdqgD3T4GPyp/9AMmUHT9fn8ZwHCuUe0vbRwVUXA99+YHTuadcLhEHGKUs
Irc9qr7T9jhAyB+7H/q8XICQgUPb6NnouNj3tlK6Hqwgp772qjGrzZqfeRZ6oV4rHLUKUa2idgos
Z8EaYrn+dnvfnYcdhnB46MMc9f6JPjmKk/cXIZrFYkZI6TUGiGk3XFTNC56wM3niX5L1Y2ZlbWiV
G/hYiSEGf/VHE9ejw+DeAOVqDV7oYx4A95v+OMZG/3oHhT6qUDr0Uj+ifOCzJq4s6pHunlWvNGX2
oN5OapE/OdpXUAOFroeJ/Sf64urhxXo2hfDC9EPYQI/fOGYjAfA4PA5Ae7sfM4KkPKbv0XgnuEVf
wC1EKySaWg5pCs4mSTAOf8qr1gLMFGT15upWPudicsGVTQcMVlEzn1rjWT8J7ptTniD1JiUH5cPA
N0yz7QfuUNSW2jnMRMbPU2EXK9AsPJKv7+KWi6EHCi4mLWpzTpTUH1/2hm2MO3CzDB+xOhbu2Mg2
vUpISWBHQ2yo/8Dc8okJRxUUraQKcnbWhV0kkfYFpk9JWr8QskJfE3u3i+/Xb36TOM0Jlzjtd3I9
wTPqo/htCFkkqGuXgsw/8+lxYo+8gGo9vHXmjbuUn8Uc6ccDldeNayn6ugvXia4M8QBctdkE/7Zb
G8DEmRkJ+Movq2HNqq0TkHtsnAXCby8PVqvk4buobfAFfriZU13AZxgFZd3CvFmzwBgV3L1AhYTQ
MEdgNFbZemUIHizdGkczwJ0/cjvc3WTHDuFQYW0w+NnL88wvyR4Vq9pGcIcvPWcoFXVtSWm1pKdk
BNyDGF3Z4w4EujhkUHOt7kGPQvvMlHspaj9WlmhNawEP1tbtKeW3Ufv4iP8NdUnLP0CXafZWGVOr
fT7yGE56zjh/UtL5RcMWo6bJw5cvt0+eJggTQYuU+crpvYB1W2i/BK17gmAn6GhHY9ijp9KxZyfM
Q5U8Z8JqV3OgEyNS2XRBCQlRrffAtcr/U6G6YFVQLylr/HqW2IemYepBIrQarLeu1RqZ5v5YUA5i
Wg3RxheFzNGJNgBvHdALnxie7BirhRSjmY1wx+Ci7a2lIkYjjPqi23Oj+/qelozBqYJCpaQD9qhV
nk8BO20Z6o2JRUNsULN+n4Bid3oQCxf7mtW3v59t4/n+XQy2XqIQ4xCriDpLgV6VZCzRSXfLJ+9u
Xc3tdStfE5bYC2zkebxejUtpUKvntmBcL++INoIYgS6cyALXmNSQQUgQYHLtMpGpQGaYhz2x9pWH
B1rLcKCF5SErnhtbMqTMyGVRXNf8xboVipshqreqd9MThO83HyJEX+R9ir63cJSoBbQlhlBpSPyC
euzlj6TbQvE3kbMht2ryBjFlCOm1Zfx/ZPDlyDr5G1R0n+FIf97MYPHHVudbSPj0xaIUGErjon0W
UaG90XCEcYhhjAsFFsqTfAhobl85roB/oLGz7jzAXDpPDfwcHgSQwtPIHWu13/Hhq+BXjcC/7H3m
VEAny3UfdtbnKPqa118cdPxcnNDPKU0BSmwd1XeIFZSWmYZEWGDe5o/ZaSDMK8B/0J5ep31UONZh
KMKWtgf0ku6PDqljF7LeIuPjP7pkz71hL8RuDJBjgqKFmD4nbWs1vpjAocPgkxBp73xAQn5gAVJr
CbWCl4etSEV7cCD8IggEmLleqKwPywzUAmwGmXYkx224aTpRyXIYPFEtYuI0RscdrLCyHIibtR/Z
yZ52RZqsCFpVWp3qV+Pl02Q0UxBJb63qbtvneB9owlZawHGAq2X9tRihaACsG8scDCLGdQR3wstK
dgUxLqCJA/ygbUzhXTcjX3WuXez5fMGXjU6mueflBy4pFUS13XyggyIZ7UBLqipGBMD1UXd5sjL4
u/0CEUe9Juw43A/0DcWPSleyHo8VHFTSo714VFEEhM/MPZVvvels/L2egR3/oiDSJR0++Le+rD7R
JAK4z1ClZZ0Y0vaqszQVgccF04qu7ZaZJnz/sEyK8sIeMipkh1mSwRcmgesFvEUYDQyccW0RzV2o
wGFdh0yk/9s5BuRubsh8LAZ15uKFaQh6SPmZBnBv6Fkvqoa6gYMPj1t4PY+PyR9RXm2ogQvYEfJ9
GV3FfozzJf9nAQiX8oAgRAj2sV8yVn++j5RHDG+W09eNl0MYsAVHMCcPq+1IROSEqD0WFBk7KbqR
ggKH3R11ChuIiYfqFN0uNkzSDO94dcQVwmfmyyZ+6MPeJ2D6jf5vMsDrRP8z/VoQHksxLEVDCRJ9
r2Dml9aDMhc6KCCN01BHFa1NJA558LwMdwsO5vT7fKRaenMF3ksooaMoklJtdWePnikLz7IrZico
rGXKfadi1FbVyZJiSRhtu7/V+8CWw/Vzm4IxTQ28sGFjlMwrsw3fB37RytLqD6Lqb7LWnCSSoZ2t
JQxKDrHTdnZrBv+D5PoktZ8BmiDl8WRBayFwf6J2LhikVCv8YGLV7LJQyi1pcgOT9BVAwmtxGPxG
V2np6Tz2ROsDvrYtahifHRQy+CsOm7dK7MPQFBe2U+mLdq/GhCXE635Su1u/KGMCojwwOd4YiBVr
Zkd6KOoLt8eBJTc2NFrvW/vu+aXLFO/CKC3UqxSIZwiKSbzVLomiHpYG0nt333VqRGPJvmPuDylW
1+yJAdJuxU05rO6H0kOGcQIhxxjCuGAPjhJPZmXfBaOHXetRpvxJhD1doohZU+RSn6nrwXIuMCu6
+IZ8JBqr0FbVS81sq0zTUKrhFSRdlQov2iOegOU/3G1+qsRi4ZyhUdpWOy4U3vqeq4oGviHehRAG
t1Z8h0IdfPcC5W4AS05tSrjYekkxrr5IO0UrwV1MXfKoMv9pjEwS9jMdTHx3KVNTi3XE06UW/FLU
vweP8+/hu+tQiHsKEtQu/IBmp/J0cbbkLH+c4MNMO4YaoHMUmbkWKcFDkQnFKWRQmXrE1yA6pkN5
ATl+cdg7CbQbLAGv6jf2cmDhTUtK6Ggk4CnyBUINAKNaHzNtQDMA9gUQZ5HLcx3UMsokwHdR7K6f
15JyraLZrYQvLj2WcvwUjwQuhOKzsBA4J2+r+ZZTB4DIMw2D1GGmLiE678xWegIMnyI9VCDJhlWJ
NO1rj2lTg3FMQWT2atnqWszqthgiJK4tVAmU02hhNzBejDZ6aZ1yAC2YVKR9T8Dg2AS7xnNRVfUx
wMzJERu8zRspl/vzdR1I6GmxoHQgwipOAJ8YpX5GW/A5A28kh7VPw0m9uy8gtu1nEd1Ymg5IOHsB
Iooq/O8h/SgbR5QyFC5A8dR8TnnOo56QgZITQlDKwHp/Dr+EaMCCK+1iy4kNLzP/vWMrF/UoY20n
mw4w6ycS3ttnNrGkoprOB+UW0zAfvzMVaxonF5wk0oX69leutY8ITaz2WCtvWVxmUe7HkTtRaK6Z
dyUi/+/yWgpeVOprNeVtkKMpX/5RHWLW6447NuzgMlQSBA74v7lZ846AUul3coU9r1bWMqR8EBHW
YskoBS3LICWrRW0AGVB0tbeDPvSHBggAiHna1sGGEqY3Ihp7aBhMXG65m65XhsOIHA1qBGDAUIMv
hrIenbkEeoWkNgyGPt6TcVDGNoOIl+TJYvgHIHTbkkmtTFmz5rCeUL7w9wpNchTtKP8psacIj/Uo
zth2PbyG3O3FvL1SLcgarxux2/i+FVV6vV0DfzzRhCRH6CWyilFncEonK6QnJINdTagw4WRq9zsW
iI00LsyO07B7d0NZAPzSV4a1d8h7IYNSc6l4Uc5G1lMS6Zw3inC3X36yxY3IHTLTn1llm03Pje+/
W08OQwtMwQQud1TcZzGa0579EunzM9kt5sDlYkZogA4a5NSvrhY8ISCWmP5dj11+oynwRkHCXMNW
3L5+uP0VHGpxgXksi8TpZuhw7PC/+WY3C8aT4qomFghzR8yzi0scBtvyIQZnSnIfHUtG7I1viuVA
SsZoo7U3soej9HunVMsWPg63aAHvbG2xQHrPiYKvKWdVtvOYmrV8olXHzye8QhtD7umn3Ve+0pVD
kIhnGzGsbXKy/tInepsEj2RbOw+25iyUxF0vcBB+RQJjXqlWn2frG+tjikhBYZnjcMAYCwuTdm37
u1I1b5qjs9AVxNEVBexV+fPb/rEztoGxupepn8gdp0M/nzWFklSmnQ6lh0OOET47KVS+xyeQ0cuV
HLveWdfY9Uetf2LvAJvPi2OmA2ttXF15BI/ew7DYVG1UCg16EJLqzk72nIK3Rk42sTRq6AUGaRwn
FlEWfzmqoWN//owr0k88CqwiDGjoIQH9WZfyYw9nWBSfqOAOAdfp2V6usUPhryhhyHUfRHVt+uEv
C77G9BhYVdvbXAwkdPD0fo0hNXew/EbuWWgREpo5m3kmmjSPTpyIg6jYxS/9SdeAMGSFQ3VWjktj
48F/651gqFQT2tK8TAXFTmRDN3jAGdrs+0RJiMws+40zcFVsS/Rtq6qg1370v3DK//A3dMmfDj8X
JnsIUVJEVWXqbIJcUay+O7qrtuofq0DBLpEnmVQeDIWWMFJ8xVrSEkWSWNYSr6bGTqDVeaeVC8MN
dDsUgyKh+/SZqAAN7SrCl1TQ8bn4SJEUG8o/UVqbSSh30KevFE2aTz9IwFEFjyzX91MPw0L/56VE
I+70AzQcgnx9QBWUtoQcuIeNgMKgqxr3+Rb6RQUddp4hegF9pHNNoYtanz4dlp38OLCTS7XxzB96
rN7EGmMs8ZywoXnOaOnZHA1XZ6x2RQAIhcfjjeOHfmaJ9RdAscwt5mE=
`protect end_protected
