`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mXNSQK/SUn5WKu9di7tCsBSbM99q2TTxVpP5AEGWSbTwazyo6ryKJe/G5BLBgJIedVo1ZYewauFr
td8zI3B0cA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cco+9BW6/XXIPO+Oj+K+XVA0VQ7DmqELy6EWZFcrQLE6fEPUOY0qPkuw3Yrz5/rsWX1ocp9BSK4E
ghI+RuPiLB6+70w64jza73szQ+9gce1kYZVU3bPYDQQTVi19ZPuMMb3rnYJOlkP8tkFekqZzLnkd
PKRjDpHeJeFLxfpAkPo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UetISM2Kj+dw9fPIY5/TQEnnpkHTEi+uMEXpAUbTzVTW7uPntumtxjhtT+ZeahOEpu6dhv6X4Zs/
gYxZBgdnqkhJ6bimynlyp6/QbElKwcCKPBTucFG7N6e61RXEJLZkDzXSr2TAch3zIYi35eTLoCVs
PGOV6Mu3nKqvUxyILPxa2DSerZQAjl+ttl8r6fCAVe+QWjvvFOOfhr5RvE0ORQrGJk4SRvh2hCP4
oNqpMajnSPn0Xf5x5WHPME2y1miL2a2hMyGY8ftLJbbyun7r+hxCnzXj8zL5lyHn8+iSUCdLsi3q
2N//o1cYWqYEoDrck4ivX2MmZFH56LKdUfFHfA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
upvKKrT8hRiwHK62C1Wk6nNnsDQTLaEnOAWHueoenBhoveVXgZejlDIIIwoZrpH1wJL0oztpG0/2
QCIT5iF4kZUBAMtxxN+rqT1O4kMCoOCpGNrtjg3S7waMZL+bdQnBoz/cU6+3pI0Tl6iNHBmapUgN
F0wZ7hvMbQHoQpFHp7E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ERkiiA9BwyoNQXx+u/EMKBReJTLMCwGbthvKKEBK2YKZev3kkMLBngaP/Vm0PwXs7X7JC7TD4W4E
kp1/BbetU2fBf8OJ9N90OkfKYA4A0jbI+2zo5VAdQC1UuGZscNO0YFoz+kg8+DPoB7LgDa/SQRj5
w/PZRr/P1U1lILkpgL+j6JEdtpRiQxmiryUnZ7sAtHttPk4aHv5bgR9NTwT2RBhELYNy2strYjpz
BWzTfphZVDs4ErwQtnLvjfvpJKSbruIMJaHkbq7HDieM0egxMc42A6zEKBMBonvCep6BujJM8zTE
utTL7KxYKEy+2SzcXba2pWK0oH+GTNkedg2TSg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37424)
`protect data_block
9BzOXYXM0gbcoJOX83z7Nj9FHLTb7lOu8gouFNMmMY3ybE6HZR+LqWt6wfgZJcch/5oiAj0lICSF
JsB4YCcr88fB/uXmVIw20asKtgZNhfEbF9NBZLg0QxPsA0j7PLH+1YQ6SGKF0zE6hrdGMUfiBpcK
1yiwlTavmM4oDldPFTCZPD+9EvnA1xMvmYJqnjNWsmbG43DLhlYpiZwovPHy+uKy2LyxufJsJh7+
ecW3RSEfitvZW8CI+mgXqCeb3062GxFzBzFub72UIs7A0BrvyX0cG4Dfmj3cXXR48ucXLMNz0BwM
cI0DpPCL9ZvJzkxofLgii+EOfF66CgY6ufy5v360yhqCmuD06Gd39HcFoj6dcVOdsKn1vaxs1Z/s
k/c0EHbEb1h0ZIuHKdg90iQVO6N90Q+6TUlFHICeWM/l1Vxin/6TosyYYI+Yr/H8K6mAb3nCa8Xl
V6cuDwAtzZ1J8FYLOWjR+rjPX1+bnNyxPcRytthXnkVggrXRBgZXKGkq6uWyI3Z8+/Zt7wucs10G
izeFwXH4LG2Xy6WQzM9OqecAZY5u3qZtm9jT3PG7kH+PDORx/sbsQZkexAp+zTvTayANZlfLJZIo
Y15AellbhcrAE+TFJmYBwIWbq1fMtxLmiwaVbf+iATJgSlCR9HkXjKuvvnULZuD2WnNELKv2Xf3v
2kIpvMV81dB945W78BTU/tG2ZcgAMdk38nAuelsAN72QRhDY3J24mkbisVQVSwcKTECrACbKvyi3
Gn2wwY1SrByZeP2A+gWUVZPJ+tzyHY8vBEbRhtHVgTrmmkC0Ism8L4TtSjCy/AfMkrGMQzm7AlV5
m4EFZftQI1o5ysc5UsS4XrO/QJhog8ba/5BFXEzfV9Jm5qZYNgjBKfscNHUytZs5NgbMmEMK0YLc
AzwX1sjRT5obGrY+Hd6S7pZt4mD4kP7nk7KdCVykZhhGEnQhqMQcVdRM+5T3lx/ZjdBo8cyz5dJG
AAxB1ClnVyqzEYnkG9D/wC7Dt/fB0seGZL8NHcl/B2fDtMJmsbD2Kmz5tVXfvSBAxMI4NhWdWCoc
18gyTUuzU5kD1k/YrrG31Sapl3G3TIsTnElCgaz2AMC4vvd+vZFBUwFMjd4aEH3SzHP+WNzxZsbM
7c0ms2kH5EVJRezmnu54W6uFsv7C9eC+aGOSk/16J/xnsFkVWTuTH7XkWNKmdC8r4otztT3oKH4I
2mjQI5n85wKfixOs0xz3GiERRriOEkftOSj4CxlnRqNKanvOl6wYjut02lklKYFzw5z3qcSmKNKJ
9QtzJeQnG0k8e4LZYFMYcXG43FzGdRbHOxzKUQ9fZ0TRNZHrZTITE1zgdwc+OOFXDSbTJSuB+KNd
bDcDrlu3Q31vFhGqke8nzq3WGrWovC0Z+f/7Cm8F5YVhjaRDl1NT87va1LBLZxfY6QpIu9kfJWrw
1emzHTongqaPorSxLaM9TjjQ+If48F7QhuAB3h8fSZTzucr7K6QUq2iYTrdNakAzoSMcjyRyrWjF
BQZqvcuhecIC2FIiXFvP15Tsv9TkffNOs72LPty5J/Jxh9fwHUYLtVH7IIIB9q0homJIaDufikIp
A9TdupvKSP8c6D0GtCLP1gEBI0HzpFyW4jrBLrsHlmiLVf/a2ma/HVdef6BSbjyDoxwYMQoSznFT
Jfi0p489Eg1YYCW/YYeVixud5vOXHvA6iiemjg/eU1Ss/o1CQvOnL/AaoGf/Oug0aScF29IiJZUQ
47prw4/i/tCEEqjrNBCEUhrn9k56MPrSWLNH+faxBAOo8Q0bkURDh2uafof5vbMNfJ1GxA8HjRVq
GDBG0C7FlPzfR650GLUyOce3W20BGy1yTCVl9ScxGbSX5NumvfxQq4nbC1/6epUld8OSIcVSfVXb
Q5MvUbYl1y9Hm5YRegqhY/BmWm5f4c4rimkAzr9CojY6j2i6KZmQlh/5uYJJ4eM78J0FCg2FRAsm
mP3ALnUg1hLRBLxGK7Td+ZT64nCcOYMxvD1W+NiVZU/78mmdD1ho5uyJsBztNcJBgYg1Nnh99qyh
qH2U+sBpVTl5CuCbUcHXKVp1be82SsSMbvDVCewhb6L18eh536ySQeiSdmYoG609H4MVtChcc9et
XvZ2O+T1o9stML3/PcRGm0q+HTxwUfBrthkByajuj6DUDk0ucDVOfvPzcWOOMeDUDXLuRMQKlnJM
tni0bObVai5tzDWf5EJ5InM6oFFvasAO0BnwHNHUrDGkhHyJNtVVYlLt2sDvARMaOfWrjWBG8I+F
d4m7pAVs7ZD/QN0vS6dblzMu/7q/p/OmYsJyxkUwZytizZb79vazrL9yRMD6wKZ+4N80r+6MbxPb
nA5KS0BcWNJt94EapjkhrLkgUaHobqRWsN5eRtluUU3nmzstMagMknGZ0JSpAD+za4H+wA4Ju6yM
x+7CVJWExIe/PXGkCr//BzmRd8u4kpNlmmu8AUiMk3PhVmIKW9MioPEGCAVaMYwUguOEG+VBXXtW
wEGpmSuybG/5QoogKdhooqx67AdxraOIsM/TbDI2rXoFBYNY7I/8rc86R9p1Mz7w6q98576cgbe4
5PF1CYYeYiLL4VoDBhF4ePFaGI3AODWRR2v2/Ra28CShiEV5MZMSSUu/G99P0YZzUXkc6c08JjkU
GrmM+MgXpVCeS3qxKxQ3TGGS8noJUfMYD7H3SDMS05SrRoVu5KduzbdDRw5fSGx4USJUhTcAulGt
riSgn1xXDa4RBrwNbco1xBYMGPnhv/I6yAO8Ux1TqaadHYD2uMqVUjsOrpDskm5juPf/VMrPhkW0
Ji8tMOoVu8+z298+pKEJTBPmoJg46jZc/wLaQQVH0H9WRZcyfCKh1yli+ILC19JstXv6YZ4Q5wkn
TJo9BWyZ4mrzQxenWh+e7YcOrzimG5c9hSDQLS1wmM4HL8NFik7ElsxXztbxNCAAfQN7kzrdIZpt
/TzO7usnXqfTOBWFA5G+E7gZjRNdrFQmR3LPDOZfJi5XdyY0wuorrWGhoH9IE/xieY1YA9HO5TYv
sFsJ95ObQL66jXazCDytoSQBkEIsvwCo1xZlGwi8Ouw53grDmJoSHgHHwoqQqfbrQ4tOUrkjh5gl
qs7gQ+86IO5qGPKheDBKTFcDs0X02y1X1Ii19NLFKoJnKOAhTjDT67zbuYn9hKIQYPa5QWca8quX
zjuGi9k/cLUiIojueDjTlGI2M4bM7nlrNQCHBEDqONpy/BShLW+xWzhDt6DXeiKK/D0mbODOWL5I
3cNtBRxgxTCxAcWlKqhAex9dPfwdv+uQbiUp3+BBK/lzxUkkqsuHH1lV/AysuWLC9TrjN59Rw7E1
zauPnMtTREbnT/7UzEddhIVbR9S9MqzcYD6XO2IBLUd8q7tIg0g6Ec2uOayX5HO16o2WdEI4SzTG
BNVvalDGcIKloRiYu8ELNDp3Wpskmb0S/ler40JgZGVcde47pVKXWxv1scsyoIEuFedAIIsXbw5m
rWAXWFOEPss/kZwVpGAguhTpowBHaOFHOHdYv4+xqOgBrKJMdRzzg4l8w8ljOWcHPW5TJu9PcJ4J
VdfHtC+Pn3v5apunXZwMUy0+uVwjiRFxHQyGgw/8ETmIU0+hx5Ldt1guf7BPIcMHBlzqR+63P5M/
BqZmJ6McPCDJeOaPTA2IJ1+iylFXCB0sOR7NrgMDoe27cPlrEf79CIuPGmLctPC6gu0mWvBDVK7H
woyiKO7YfczvOUtu4RsfS2WMRo95ZGJBVnXVhwvk9irXtxG5IuNSeSRaMcEMoFravBKUNCrov9F4
GaOwasZg1n6IXUmsopJRRvCkpA8FxNgpyiRvn3Ivd3jF9TmtMny5II8/3NKeWUVgZIIeCxJrKqCK
B9DVkk00OBjlYYHAhHaKQ3O5fTMsL+G8yn9b0YgtaQRJsCHsVmMMUyvIb3t/N7E2lkDrPU4DWlj+
OmwtndEkoMDxuzLNOOLj87DkNnmSBmyBzNmIjhTeegJG4A+tnUb2vkxA1nBK9W/Y0Qm9Za5ux0gj
2zUO/Im3sGhjCId+wdWlnCvwUo/W5/nupJH8wmDNjipsRfiv+1p2eLPt12sJ9S1gkDBoVKORUG6O
jWoWeSuKhzWSpgGHNtOOxrdltCd/4vEt9e+xLzvyN/674hqiq9B5kep7We/WoXs8Md07buUrdesT
44mS0/ulZhefMIlAjO7wq9IzFNF4uFPwBTc+E0jXLk++5OavPbasJ+iBq4ffnxlOxg+tRn3vDinw
gIuuNKGBUL2Pmwcv1HOgQtJAKouAtuw/YtIzD4sN+2u6bxTg7rzm+MtjGxn0GXv6A4acCosbl7uX
GBhLFskmtB+6U/DCeF0l8/uvGYpBLaRnFU/erOCEd9s6YFlQYcozgRQD9r5hFSzOwHuWFpGq9Zi6
Tna1gIKhVHeZBAXNsAXUgflXY+MvJernLimz+g6PPZnU3gz+CQJHL9lqcYaG8tH4J76P4uOYlFHc
McrS1E98kacEJoscoBkQS/Rtx38zl/VDVWHptUDotOpxMU8cEBm83mKyXpmtXGKMIcXf+qEbSjsE
KcqpjRzP78Y+B0Fyxff5Ujo9m2wgI5TlkpCUQF4anZRGP8sQQNxt4SI98OONqJXYQrNm/vQ3voun
vKnCd3am3QtL5jkUu6GbX94aukaVVvbfQTj+o/+xaBIrB4vu2hOI+vkEE5QfNHut8DRbSaBe+lhw
oM3FczJpbXeoTUh34bFjVbipxPXwOPeD6kN6+FJ8/2dyQHghs3IF61tZZ68DPYvr74NgeCBW8+MY
VVC0sKjwFjNmG61p4S1ut9a6j5Ud/xxIo2kGc3rxEjj/F0qrF7b6h7MRLPA7vMlQp4l0v8YQNJXz
1dbJ6cQYEPjQCy82wYH2s1houYzNYdCDKgFftFTa1/ywU/443+SF2VHPhbRskbLaNCGoBMwf5+8y
+ban4jq4rxIBAQer3yYgxH/E8sd71zw56aI1BHjZvXkDzZmD6253CplHazJuImM0wL/KJng5Ezq2
GHkReRpueT8kdKRPJRYhERRNIIjnY/kN0DA8KbC+BFFUDSyR+CxZNPwlUJiOPSOE8OlGRU/wPw7k
U8wDaTZPTkbAsFm4Hap8oVWe6DjieFEnLhF6X7PyivMEmEPYdBgqIzxs3mMVFPpiyvtKaapdB6nT
JuvOudUWNjfag1g0QOTNISOzgDVuB0abI9HUEfJLbNHiA99rd+j2iqxUibsiAY0Jv5t8pZOTUE4m
rt/g1Hs7uXKCnTl+p+zzIaZn+xpePHjRB9SYMM2Y6meLyKYn117JiSBsf9hfug5HVkJ7kfKthWs2
DUnV8j28juliDz34DZDPHfgpPsVHredBLfifzTckvvKE+Da5Nwh0Whs50iz3DOmQXM4AjYgVbxc2
pNkmtQXsWRPdVIc0JaAxp0fR4gy+wq6dTf8k2LjJzgTQiei3v3nLemM7PiBDoyhT2krdcgqa0mXG
pS9EC1LRgvGuGAyPanhjrCzEhRviKq9W/XkJ3uLQTZffYtjF/ofeM/f/ZGGScdzslxSUQQv6UD0g
ey7bwjxYpoPisgsAcQf6kW9UdsFYblkBgzLc732hOVwoVIatfwX/OHmij2J2TLhod763uLYdnmPN
Z2b5y7G5YtEEaktBZ3D27qiMRG57bctwvU0SXiEVG+AocMKb3YvhSy66SoDhLu4sunvCiEPo5xjD
VUiz20lEYOEuXJV+G+blhA9RbgY3FVGXjacqOpfJq8/tWvPFkAfFo7BXVa0jIgIY0Aiwn+Xc5sP2
Fdz+C3c5ivBgIDQEy6Hx7HOBw2cAQ8M7wV3CMuNWc+EMzQxAIKKeY+32tmOY2j+yeGzB1S+DvH1D
xtlG3w6o8Qg4I+4Huw/tTEdxmrFQYz9ZV8iyaAUhPsYWG073nuX2gij6f+WkhxwlBw1T44jC7O9S
oLbF0ROAgsLEJRKIG5BWKv2V4ZcxNIKOzbSUq6cm1EoMi+7kQTKig4UwKSsdPEfftCwxNzthJ5By
jXl6d56/2//bUqvQ1PXYWfA9azeBYIqfJI6ULTKiHjIaOYyl+ofAQSbSKC+IiKz1CYztaFJj3jBW
q/Hjk1xH5JTdLm/39fEBrkoXcK0mq0cgHzhu5Fu6mZXjwOQ2k+P2rWYtkiC/8kOKGJ87+heyO9G5
XHbDTUQuzpYUWrALQlHrsS6csvDhgU9T77ltVwqgUK+ho0djkz+7gSM7u6IRvYV9s7Kaz1rV5PE2
g1638Qjw2aTH4wZTHp5sJljxRuK4ssUcy7TXiYej/6wGcpj6m7XwoKDEYqD8JrhNVUYfWnt24ntm
yKlg26znwoPLUdjFP6Vpor/TJA+7f5KjYNGipdPExvF4EvQVs7qxGgLHiO4kOYdcmRfphc6ogvbf
wMFTXzSdSWvyjB/soSC5Awo9CJPKEWTZB1zVFQ8EAti7+NCApOfUJvTi2JQN7oUQ6Sg2eSawxx0v
enojGRa3GJryHLAU7WQitGGcyF8VVEK90VXYHMwVCUrJfOeNJ1FFT1lBRl7KLturIm7876PMM38o
iN7r7OhAqIWtF4T8bMy+NJdp067uAbrgvsEhI6VbO/WZOPfzGP7wpIqdZyC3LjxoYCmoNqR2JPZF
8Eol+xetQ591sfNCjKDPiCH0FG+hFwzrIcX9pPlL9hiF6Ri1xaMZh0zebsw2Ly2XuZmU2008cvMJ
GcbWaIVymX0poDLfA/dkr9MbkH1WzYAKsYRZKbf1Z1J5KSOcRVJRqsPLrPiUqedUdPzWJmHoXA32
vMFb4XHabIqZ26E4z5EKMr2PGztJAz8+hoDRQPdjD0JaHlFlOZSlQdONfMvKwwGmPc0tQ5+o/TA7
l/4Xmwv9tf32il0glitjjY1dezirxpojCVhPj8gjD7a+HYBu8VlKkg/Uas83RjJ8nO/0utJPtepq
JC6btnD9SR3s9obo7X7E9pNRLprLTl4ITaQnRwXLfSsWYhARRnxX71w03S+M0IecVJgbI7FvcT1R
hkn3w+oIQIOd/ASglRx2TnHp13wLDHi74/a2yGnTsqAggUPFlgApW4ed0tmXTht7mifdB2QIYAIU
ZY+eVPpZQ3vLiQDtWzaX+qTWU2g6vnqoNUx0cDkcuPc9aJOP/HyrZ6pZNJrTMwG5w6zYB6GxwJnw
EnnsWBHEMV9yUxV74bcNvJvGDspWoKyuubzSzbkKjm913AHb1SftEa5gy3JQX5Zma6H1g16dO/ts
GlZKqVVbjY8GaDdU7grktwF2c3cWBOygaDSQoqPZmrsjoBcTbnPvJz5OYdbVrxNQ7lmZU18Jy2gw
XWC/5IY7IrWIvi5ieuJvoCOMqdWri2+tiVQ78S140i2jq/WJUaxnYDd73U/9eELwIby887mOl4t9
hWVAcn1eFSzYcZYy8Ug2GkHtqNTxrIHc0D54wxm7gF8vGWbzm0P3G7L0LJqLuDDH3GDWrFXwb60U
o21IXEY3vJJEGoZVIJSUu923RO+4XtQ27uH3DhXbTRhWLjJPGl/HpLTtP41bhG2lxpU00ASosrya
E22Ns6F5S2uyXalOTldP3dtWMCToZ0Nr+kccJJyTDyBT1IR6lZaVErJ3y9N3NsAepQEF7nTW70x7
TPZKAixD6z8WgZf+6uqHODG+uOw3hMtr0V34CohHvHHOZSphCLM7ov0scAd4ps4jSR9/khCQ4RyF
9wzZ4bs3PYFNXPpEThf/p+QwpI/8tTPxRJ6R6JiaEFCQfy/Etw1eJ7TMZF1k70P3A0m2JG0INiOL
yeI3jCx44IZCbIRjfnWYM9PLg9gCwiIzaiFCMJJUCyVv3Miqj+ZBx5SmrAl6/HZP5bB8Wc1wk6Af
U//neSwqJfVoysFT6DUFKrUum/48x9L+24PlBXdCy03A1j8fZ/Z+be69Ivvpdh/P6YWNL50W7T0k
7Yh5+Pm9rWZTEpkRhxq8DwCxBjMTI6tTMgJmz/CEw+xJ0vg5x6ATW5+ElvPiH6UxmJa30Ud2vIzY
sxlkurY9B+tPzpiRuH4rq/v4stzx+jkLScgh1D56EN/t7gsnRDdCvAGTYiMVd0yIYZkHgRXJRKTN
RGNv2YiwnOrkHtjSef5Yef0KIzQIllMBmr7M2RxI706tu2tUutF/In4p2CcM4TTj5Mvky+BwVE8p
/pacXvW7GwBfIHFm6i8VaOpCLHdn5s6D0dEc7e9rkGzoS8l8MNjbjVq1OOtR4QNbJmccLU50RFlm
B+8aAlz09c12cUHImOLWjyTtVOjHHkOuAdpSTUj7+Mq0nRdb1UnMQy61qm4f8PD/zjjsNd2ZZoPN
SF7jDDPi9d6gPPoBP/OSuy7abelKarRwioZDZE0v2DjR6nUmc8v66MpFTl/R+8MZnq+XTntgNNTu
vES7AFvm5wJzAoZzviBT7GPe7iYvWxwirIWJ3tFAVfiHtaUR8kJhbb4go8qoZpDOTtURsIGoMN42
2/u7ywBeJO/3K/JZX6RO/0/R+lB4xQhB6TVMGUgNSpmPUNXJ0d35fUdZpR1mwMNT5l6BVaSukFqA
KIei9Tjp+ggLM2m+UkZWBIe1pJN3j0p6r2p/s2PhoWO9FcoSZMTEnWAJMWXoyWeuOczLB8lmtWgM
5xnbXjF+4lxS6Tl4X7G1aauetRj6DnYgkiutOTU1T/4TWtRZnmRCqXnylR1FJetBRRVC4w5AUuXn
K6hQrq0T0BdOaI5iSNvLpEdfUcBLwTlBp3kjIYy7IVYA4UQXFHp9Otdobfit3slFYl9vVbCvcvWf
g12A8Wv5UPxFbTVuJuChzc5lmbriKqfloNdTMx0zR8+YCqjxgKtE54XA/CN+uo8NMMZqIAR8KkkP
mFmHIqR/e6c1smmlWkQalgsvAyimX0I7qiMKd+jSy0jTmrR4OZQzN8BQTd3lgkHxTbEh5XyCoyFE
a5IU24BhEB94bediTpsTI6zWYfclCJ28ihi8AQ/r9gB6d4bmDNduaTV6QfqZvLE0PYnbcZ6qOiNW
YqPBpAVxuaDoOianUvAka+vtJa9sfEVJNjPM1K8n/L4krgEL2JSyaECGWvo4/gITCDpaE+mGYtD+
7awFWUw6P1cVjVL2A2AfkACkqsW5cXJb9tw/Q3RKAh1KNyVbLkJReSK8izEJOP2hTZwB/hERbPqR
5pA8kkmimtoxiZnNpWyM77qg0oSMe7r2jvQGuhumheTMLFpmtUOE7fDQrInQE/PWq5bOd/nuDn9X
cREsE00VUIl6hvVoreVxcLLzV9l754bLkQ+91gp9B/SSFZzU7Ecc4FBq7BljMRoascsapiTNbUdF
mr/yyaA4HzIvS+liAmzx4YXza35v32RWhJVqqq7Iqa4Gr8jkiCNpJRgSEMn+OhNBf5mMaot55tS+
29Pvwv6lTXEIwi6i4Z1TFZpyIAeHIOEkKP3uAZwSIgLKvzRECD2kL1K7dcY75kRpGU0DJYT0nsTu
mUGfmzWcAUOT3WkycYyJaIJQvxnkZHKp7XYflGFgKa1xtF2QCs02TYRqmkFnl3JKuli3I4t4qzKy
kHRfyx7VBLcodcD2iq52QHemnkC6QBTD5l7La888ZCMRlTSMjWlLCedDVeQkXKXXz/PFTDJlN5Qp
meCOeY7lASehze7HXHXuRk//3Crm+fiHKjcYW8a4X/psGL3qjjEeOWXZKurmbGIo2tywa4B4kNlT
r1RPnWBkB8fyOI18ri4kAyLB2GaAW6u/HaQkmV+kTHwAv9LO769YBjdp7A4+A1NMrhUzZ45+9O0H
UiyQS2dzfqOmrUdZnFVGv3O5MaRNj03Mwkx+JEAEFx8NvmAtnk+7iZ5XkTzGyqfgXGuO1b0ZQteQ
tAJzYBnpSMdj8a4lIGgpvkNabuqmq6rgVQJweXCJT2LKl+Wk3OoG1n1Jne14z/PZBVFzbjVcUziO
fXv//qaXj9ua37lM+Xje689Jamj5PmJtSDLXa/AkhQj9Bgo3YsO5BOA+MTQJElL71kvtg/6zVXoy
a6V4PwGtmmdipiIx2rQiuDYKvlpq7nrJHSF4GYbZsxasOhMG+HA1rIEwHTUuo9Lz51k2O8s32H5A
d71YrfJc5bUZsUD91E9Cy63E6yNAnl7LlxfjMrpjFRVh6CQG122ut4jEBBwHkAuVG3mK66Ycj4cB
BFI/9rzJq2epreE8y7UHBkEloMRsYY2ms/sm6j10lcz9fS/Eq2MN+x+NO49v1Dg1/URXWm7m+cnD
cSpO35x2Hl8ew9MvlnAdVo2SuWUSkGA9/lXSW5K9Z7I9bWfD2EPyTRUEMOwygm3Dyc/Qb1dc1BCg
qw8fLLrPdkCkfOCyz1SNLgIzjfsjYHnsMrWF0/+UrGZ3pDMNo2WuBLjx6AOWorzw+FJNDhA+yv7a
c0trSP6yFtNU0DHNmBbZbwJnE5vKrInYxDT5YsxAnNPR6sc67rlY8U4Bb6Q6qkdWTSKLUZpcjzyY
9MoZ7CdLQFGdN84KrRbFwsraHucNRrwGQfTGS2VpjtFBT+QbRr3UDEGUtoigWcdgAXPQxhiTO4ah
mBdtyL8tKXeW4jzBaqgNjITi9XEXqvjAz/vlgPMCqapI6GBjpOZt3N82LkA1DZsR7GE1Sb9sD2sR
8x/m246ZooMOJfVWEn8/Y80kDLWeH9q7Q9EI1Lc1HuFastqv9H1qs4KUC8c6w9f2fTurQRKigUKT
H0SSUSZQzdEpnPuKYZr7rCiC+GF3vl2hGASXCOK89ibE+rohAr1OCVMbgp59gyNQ1IETmMTtMlsM
v4dgEonyA+TX46du6hS5NhQ+e+iGC4zff3lylY97w02gaxPILQnjBOx0kBAo5dc2ZrXH4Xl5foH7
FpNvNDjQd0nG9wedwOJPmhcxS2M6OzO/yjujSPT86j0bAc7YRY9JCdriOdDBAYx9xFPBc7MATUt6
ffh0hAvMfO93TV7s9leDVmqOTt/gf38ab+WhuiPNaNfFDNUVtq51sGCiWMKuu5q4RNhUDaNub3p/
dhwYmIs9b9bDH3Ac5kMI3Pd6qXXSIJefLePTUkhMT/MCqE97kc8n6+k4/Ud//qjzZk3TGohhk5kk
xwfv9OHTmWr0kqF4gRMHxs8ej4IJv//247XlZe0KJcNCbw2KHgDHmzJKwcU3mRzIXmP7OPn8z57y
b39oOudbvB37QcMfuZfLvY+wjUFu0Ff3qWRbycCE9W0mbK3LObnWJT72aeHbgDF/rdmosTcDI+yD
V+7tY8585HcjbHWBo//s+8W96gCf+zvFGH4Bdj9/vYXXFNGiwDdGjdtoiCG3Se4gM6umL6ecfigg
+8Xq5YehRe5TCxK6lsaILAB0FXLTWUtCmmPhut5qLLDhBVyezLteo9mzXfPTSeVMxMhR0rbdU3ba
vM4XTMLue+xab2PrFoqSxwDe1LGmtV0UZcBqEKeFRtabxRh+YqSLBs/twIHXVdsEBqZeH3fr54cI
8ybSBoefjV29Mlydo/6r1cskRYCgQCz0s+lu65cMsQbYnUzrgDf5CZ5iGoMp/8tpy+4R3kV5KMsk
98KFeL7RxW7IqDCNvguNcH0+xI5J6SDb2uvifQsx2OBga+qh+2NBdhG68Z1Ks1EZ8kBiR0y4t7uj
2FcXUgG++uYiAHkN840vqYc9SUBVA2DtdcKQ4CNHqetxd9DQxy0W0mm/TzuPDpMGMogjsvmI5FH1
+endCXA09lmo4dOCQx51TOjrVA5GLAj8mP/5wQbRBlTim5Kh/yD6lEviVa+MRQYPzFxgRshvAjQ4
/hXMDyvMebH8Cmhblx2aYcMtzxFCKWI58z1llxk1ApDktJeZUMGxZ7gjVkWfv+Zilm3+B2p0ae/V
fptYBmkzAI+4C868RSY7glZqroBIcAX79SVPU0RJsPQ541HnCyTtVoQdnCm4yPpVFl39gtC5T4vE
ZBwiaqm/+O4ALIo8k73Dt3PLO2zW3GXa+TdCYzxSmOs8KrM3M3YSydJP5uTPlvdbexknybxLXMRr
pMyWM4f2vVEiZLWr6lDUVlM9zfQsmtkVNtU0/cp5pXKpaLe74PLvo5ZHG8N8hk7zYkXKOn0ThylL
kV4/J5PnJCUsbP5zCfkNQg5iXZyt/AHvNY+CFH6CRGhLR4r2UidN3QiNXtamkDhGH6EY2GN1jm9f
kRkUlxD9G6wpzd2NiSWQnJ4o3CB0fzHJqxbMASHGXhG4BAJZYuMXtjnxCCb+yWkS5DN2r6e2s7Y/
7AWjkrGU+74x2h9XUaR5dEhCKps6P9QQa6VcfYLAA8bfAhXJ2yfBGqPKim+5e3OZPqCxhMhbUB0y
VySShw+bfB//6s3xSqcQF1RcDQYHusRcIHgwTdSs7lv0BvwhY/L6WrT7/kM6QbsY+UEP8OwhPxKI
Nsj5JhFj6d3Dr6qMJfvH6110uXIHjiowBTT6MKnku35Ox6ZBRHtwO+8HnBeZpMuimQ0ZZPDf2QeJ
B/GKzBiOpE7oee6TpaNAEDo0GRtGustXmOXlGuz8SzGDzpFH/ZIb3C6+gyu1PAflJPaq1qxrlTan
lIcQgPU1ojEuKG7JUUzWZe3U2h5AtFBONrzM5krpGPSisqucA9HVABekvzjrJIZjM3GyHRl10MNm
sJybkm1jdSZbiKACAmYONKoXEjL5aJyO4JUCNVRXsrwxobwaL/nTPEQLP87LxokBWyex+XCEat2O
Sziv/fhz7PXV4MiMb18eiKmwJIgo53J9L74APrPUkDHmmM997BWjF03/L9lcBQ17DGYulR31awXZ
X/sqrpEPxzctT9cRLF0IHNSehz6IMUK/CqGiitj7mqxHrXtPc3VaSBzZnpBZD5GG63v1memWhXn1
DsvgoxNmf86TTjl4GZ7HfSB+FDh6D9h8quocKCX1XVa+1/2qlRGjIsaqwe2gcsdOwIEiMned9zU+
ipLb/MhI0vGSUBeFtk+rObxUjrc9pYWLhv7zjJr8HZZmq+eK2vefvqhYDTqAPpvN6h8ASZm8Qyp2
iLKdy86WNNdMJsUGrz6xIc2TCuSVcm60MwoQYFDqe64tEnoehKNbOpC6cmmgspWvpzRai0ST9wdt
WZSiGFkHbyABaeXYeusnINkN1JNiJCyOIhD9mohOb2L4D8JdGrlPVmeH1cvxKIdrUb5m+aBMcV5z
RaiLBQxEuSb53i6sy0Z/fuiQWiciMWAIJuQllA1WZ8mdL2nJmYRcjatoybOvZoqSFv0axRxcKGLM
w1IiCAMDuI7fPAWXkzSfY2en8zbl1obC8eNkwUWSwxjlhOqLJG5c7beil1gufgGh9Bu//h5Jgnoa
XCwtqyO0701LpbCyXTNtJIOXsDeuWoucbW+MjoRgx5KJJd0jzpGQ7CZQ/fYVaxuLoyByg2Y2gz6i
ZBtzUd8HkW9cZUrWc4fV+9jQR9T3Vqysf3SN+3fPdluUotdC5PGh9Wi1kR0rlv82bn+s5oYHyJhJ
qvdT3THhFcIOXtf6mz6UAJ5Qg7GlPPliTcuIyU3ZhUa6Reb2KtT850/6Asv0emkuLIXFQdmYrtkz
MQTqnycq5fiGf59cdd0YbBgxlnRA8mW6XY+VwxCgmt3r4Do52ujn1odFQsZ4xV1F1tFjokgZYWhr
rkdM4qzA2KHwrCgS/LSZub0z9aAU392pHZKasycvc6CIsKzbrThBmqMtUweAHbdojbty7Sf5EX0j
PMMO9zFrQm2x92h72asulTzmaXVfvP8LmhJxVHm7JvoL1llWvhcnJuksgXasAUS7aFJWWxPvQxsn
rcT0KTTvi8JX/3Y03+x98FVjZAswEYoJvNxoQd4vlMZGAvoRMlRi5Y0aEDN7m5Iu2cSn/NmzgzZ3
W0WiBkupAjejobqGWBBKtUIojJV0EG29PLNNiG2emZENUR0w99xJadN5JypFjfPJnKwcx+4e0Ivc
w8gR4sLsZKQCWsZeoM5FH+klgJ9Mlicugn899yc/1iNBPDSWBWeVfOCk8ORoxMqQK4ZJ5VU/NJTv
e3KmEyJsaFQXLAlbZpvqnAI8qFdnCo40v7gsQZyngsGD/U0SPcfkibQ1+LrPyDnUgf5JOs8X5cl7
ot5oeucnJdIdjvBtnP7VcryEVyA94KXTqGFp+Sn12Xzng/NMT5z9xT98XBYXwQgroK0npsLNjMDT
3X3wkY8kln1W4T5M+59n9T7Nz0iygauyYMHnUwa+PpdMsANeblZBnjgwuIJN9PxKEQ1opdrl/T8L
GDBjVJx9k+TAOq3BwOimdPhtJ29jztEN/J9X0DcNz1eYpaTjQwJyw/61UQ3n9DNHXzblCmZTKg92
jDkXxb72hKgE2XKEDIxVMoLZcnUAHA0MWCjXO1LW1fmHcFXsDaPQKZloHj8shGVWt5lYHZ1IEYqz
uOpNCAhrkAX9azE3b3KwiCGxezZR1Hsqdo8Bz9FUUCGz3VeTI0zURMIEtWQ4lhgvcX3+ucDikyUD
TbY+1e63ILFrlbCG98D1T74D8s+g+z4xaAsLE9ooUbZvMOtcyBnMdZ2mQmAP7MNXSi8/dES1aPbt
YcOPOz02diQZh0QPYraEjFookpKbNoH1NfM7BVohD8qfrAiwgx/EEtuu2nUWWge6a2eCS5D3jfWN
9GxCkxdmKf4FOVa/vp55tnhvVMy2YCS/XAYsfpRKvvlvrINktBLU29IVdHTY6ovVP2o0iPuWb8IT
p4BeOSyen3XoaKIBSDNppkxW2TKrHX9nJKYi/GQx3s1PLenIsEdtGl1M4gQ6JFNe1FMxEcpXc9Yu
GfDT/KscsRtuGAagLMUNpGXYBBhkPBj3f0v/s0lNXJkpfFZ8WobyUApbBKlMMiTcIDb/Faq8wYPg
SA4DKbX5tl6N3caR6Nm7cathnNykXQme2u/g7rKPFOpEVwJf+g9MMcGQSR4BUM5cOP/B+Pnyb8QP
wAqYYbj47fCdbmloCY7TD6eYFTwq7uzw/UVq+Cbne+Mlym9SqfADQCfvBXTWym+ZxmnewgS3NZHS
Dywpa4tvXr7fVrzrIFd3D04w6k63c4sU1zOj79KKasrZagwgYEuMVBDHP7yPP2G6UH8dcr+8yvMt
AQLGnRGGsgZQHj1B0d6tVaro2zafQifMPNXJIqcdkRHxp/CeKZx3D2+s4rJ9Jf7UNuH1bNMB+2Gy
2x/z0mNiNT37+X8oVfiwdegpDAOZu1jEgSDgvZ/9MBDBDiuCax/VOZ+Znsj+W7T2NnIxTi0QRdhV
rpq7qn/cvDxi8fPw5cyNKfJ0elBQkD4lY6XFmb4mLHLdqdynkSvZn+2i1jiuKlR4nApY5xuLVXF8
yo1LuDtllCk8e4h5HNbb1iAOMHM+JEMWZT7DAnE979EDE2H/5gpVCwNLBVz4ICbO3fohRenqkg9v
jLB6ZPTw56AyAZPQCLw+/kEHAGj8nfX4rkPrp/T/jCq+cfaN5cc4lbn+hcGf7JYULMOOZEcg7peS
qbEHQc3h4Kjx85EaX+eBHqsj5VZ//jNRvVNRfRfMtbb5JdBdjATI7ehrW7TG8nEvKdW4EKiW+2Ue
GEh/o06UDNvBq0H6cbP8q3bZo4CCxV+c/uTTQAMPHpRsyOORto2eihlbIHxj9ORjwFG8GcS/SbjB
ejj1aDEKSOqgJY079Kir4/ROQIEBTIRHle3PMsjQdVnru8aySyuDOzR3AYI4a4IHkFDKk+y6OJRI
LUlu4EuijK3RxtjX9WDNTY6lHF2oJyxUGNB5RKPecY4Q8zCak78OO7PTzIpNxzHonUTNX7weSP1i
7jLvhuRlsAG6UytDOL1mtmjz04M/DzxVdJb25xXnnDRO0Y8AyA7koF0tfkEVhp5AWhYhLCjx6FOY
LZENDjlyplMV7buAahqYM+0YXZvUxLkU2fX3fHuphZV7DLlWRSirOwpPXPyZOLaqw7xjl5LroAH+
eqg5XCpFS+4wABuEqAZUXSRzJTCDEkMo9fpxc55vMGm1pClgFqeYUDTQJSO6BEqFiLoMgqROsvo6
5QfMY0iIg5GeSUA311eV7zft9pEkVtN8OdF+JENBc6MxgyV8K7W/UxGtGrtGmb4EMAP4hGKJKItN
AWuRblcoPRNlravtL61bH/bXRGFnXfdCj9xRgsu8H6EjeOGsT7y0gwXcA54HPRMu+3Of4yFZSmBu
fHXtKS0QodTcdo0FSLn/G7IW3M5uGnVeDs/NMvLiKFRHr++7xn1NYjyKsbN7t2o9SDb+u0HxhJNy
2HpmttUsCOYRdZpWHt+Qk5onG55Gh0+wH9bgepJ3vm1QwFYqlx59Gr3rV6nieGAzH9BwIXi/US6N
apwNMr6A5sJRkqO9pM3KZc84jzAVVuqPKc/vQlAus92kHJzQix+O72u0250upFq9rJaSXSEc7syj
82rDUmpG2mSwP/Ax07nDBAygXi7/tI/yYautyxwB5n87KP5RRYTcvi5stqdQPTh2ir1Bq7NXYA3P
ylnmK2tAX5kRmZIgVJxurtlIRez6RodJWZM/wvwrGLRpVaiLiVoo5XQoCIjzvPdeVIzFRDiEg8TF
jVqfroiKOh8GsE+sSWQFnvx6sHDB0i+NmT3M0Z7F1xrL2Ip+D0/8td0NxnRiLhnUymcSc3emoUMc
Al/ayngMJgWJCiZtc6vsewk6AL69JCWr3p1N3xRiXyjTlRckWzpxiGXBIAAK+MO/6SD7f5EnPob1
CI9Usr2hTcVIvxmOXoWWqv+Hpg5NTIYrOp8braYeD4xtxMCUC6lttftZ7WLql/0BkDR8i1vMNcoI
x4Lk8XRhb2efcqSVYa3zlMoTD9+aE3cNbvqKCr9GfP59UbMQapLr8NyEyc0a+JhzexGHFdQfCXwX
T6wNv3byFIy6rmvPKpcar8TxGW/k59YtOJtTv/raXFZ+SRv89EnIVB0D5lEmCZT4aken4o7fFi6Z
XdSebmyqDinB9WhFroVBqlRaWimPfgOzeU55OrbpRTXi6hmhqv4DvV60W8bsHjy4DFdmr0WiRzcg
e3AXwMWMigIUmaG2u/XMUo80s2VCgcoxwkOHeN7i7NYEJU4DZsaeuJkPGrZin1Q68g5Ktot1jbuh
TTvPRCbbznq8Y2YosVZWCdG6l9hnjHEYrp1Q7ZeiDt7jJ4y5KXqBv8VW+9lUPD+t3rDqlbSq88Yd
2Voj1Fvy7u27PSbFVL9H8iiYztib1yF0S1r4ZYtij8Ju2dPFTJ0lUOuvccm8qh0TJ8fuLzA1jxsX
VJTsmG4MlT2Tq3Gbi4XR2t8VNMMmh8uLVJVqog+V0BbEkk5/KttFxSr3h0JvbmROrAfSmDG9gsNP
RGSlA1pEQWT3fUAggc2KiJKRr9OL1w0NZMgbmPUR3369j/V7KwzVO/YSGdIZ4XqDt55KHlGnEl3Z
01qxHb6u8bYXpjptkjSFT8Ueb4G3S/zS8oYT934F1haeJpPZNq/A9vxWM5dxjtlQpRAkK6QG4V2o
hrwMa9hwe8BPcR0xTJ0uqmjqqeMN5xJXYNbWsCm51fswtJCVjMI2y4fO7fXyL50hPwTvuxCFFbns
aYcK0hxDyYOWiakWEgk4FfXNcXbQDk3dECJAeJRAkAFuu0fTWsiaUdtQIDnhQ1gsrEZegPfW+bMI
nzqOoIQBVAN1rt7kLTZXeLM4CZHdzJe35WnhwcieHnOWspYhQrRdOnsyei0NaRMWmRLYmDKX/TEZ
t2kUSYgTBAKobWnKFJowpsEY7JMB6GJVAD4rktEXEVSXKk+EGp58IUGWvuM7kErlCM2HqistwDfP
7YrQk3cLb8xyEUHytfgBOBe/gxbLSgZg3meK6/Uvxf1rk690FW6fDozKxKK7oJG+ILu5tzpFnZwC
PzilwpvHJSQx8RaCXPgAgqojiNE9mZbazmZIbokzJWISH6bncv7ZwOV5AEXUldit58QDHhr4dtOm
97NiGuZ8g/+vp0UYjCjFso9wKu2kTN+7jQtobGKHs6J+F5uZ/nsI+2OFvOL/5SlOoDeTyeEyX1p2
ovlg3nYW9A2a3L4k26CLbogGlYM+6qi3Zy0esjVT55dfPI0zk5hKVWHouy6+78cGI5yBBYTuvdud
buWpWlvYxtPOC1byYvM5fZ1Rf5XqUEcLZDtK9EF0VOfCMkUAGwBdtH7yv4d8iw4hCH5PMdXtk4tx
qkElDlet9/9m+dJSvfwuD+kxb0sXP/I51SDNtH1RJb/VOft3PaQpXZoP2/uWOJxxjpvxL+5GgM2o
y7M5HxyvwjzZZAFUA7GQiA9suT6a907Wzn6V25rS8J5dauGOTruEYlK4U9iOm6V9+HQCFz41R+x0
LB73Ztw7xBhM33fTBr4Z/3Sxvvx9rSUaR+CkW7/3Rny82U1Bl1btS8/XtJUn8+Pg8+ZqWD7zouuA
uMnIpHfNiL1BHqoSAbbMWdl49ScajFg4PVh0mND4Sb9vdspOZZAoB9xazWf1m9ur2aHZCYEDVMz6
36absiJCHXtHnHHIBHmauV1+YetZwI7dyMdVAXgX3LYZd+ytTodusmBsEZDwYEGGtvxtKU9+wawp
dB6hr9WMMQ9bpp6eWsTNNGHwJxorW1rYbeILSXpj4OW++iu1jsnbM7UIKzJxEI+s6IoktK7YUAsf
i6cxk2o/wEVSdWdv14XDoV+iQ2x1fXPaeZFqJ1Plpe1XeX0+VvjvYomCtWSKoIag/Qwm1LR9oWk5
2lTdrGnhPAO2OKxooNBXsLxRZ/G+Yuf1KpkpE5jpTW8ooYRwnW8louc+ZReswaa/HhvqVwc5hi2C
zZLrC9scmyX0CwVctB5fWz8URX3663/FZkmRmtDz+C9nSpdAfL21mEmjWllEScWqbq4vS/MnpAmF
gt2O/UKR8mJYYN6mVIdQSig9jt4t7zzPqJj4WXytOqAmuH/Gaacf6R+az1S/tBZet2vt9uE3cQZc
WZJozBJXEo8bYgD4LOlMlesvUnhlZ5dyb5T36Cu7UhGUNxM3r3flLpZssIYBxwc22puTjBNnJaca
ytA+NzsXeS5svaV53HBZWqRBpwvefkOAhIsrsZT0wp5p3/9OK0pY27XY4XJffIqtAhmkHzo4+K38
o9ZyELzVFXqr+htfeLyZ0RgbC6dWWEafRhzL5M5ej8Biccw6aGKc90IYKqxfKIYYNG54M2wFggRu
epwG7xRzxGkSFPXoPvB/EuCD8MgO/Hujs152lnKNC1fz4ukGPUjq855G2l4YWajmAL0B0Z/vNJ2c
177Chv6OVKkZ0iH1NkLs+A8+IDJemp3NyzkoUzVXFyOnAvS2xYNb3m/Da5CMS4lnaCm6BNiGL5PE
2zXO8UklRueMri4cNRkwB66D1WQ43DYs6mb4BrsdoncusRtpJAigMxc7pmtXa0B1RoxYwmZ1/gQB
vPYbrdjTXFEpygoblClzm1pVrFEJ0kkj9etoA051XcEgK8G3AbWesSZJtiWA1/Byh907XNG/Ndyn
+zAVP/CD3TgsjHta0bxbCdDr6HTQqBGXVbL348/exf8uZGnytS/JtqlPk7pKw8JHPJL4aF09/7dQ
FivYKGL3piiV3QOlNGjnsw3eNegDxaNWOgr2j0BmL9iP7KwQGCR7+44nCettT7eMnRki/JzmFA0O
ijmlRD5Ef7FS79UR4dqhFb7HPUygsC8V3VxtRgd6OKYRKYrlUPIYycrG5ZgZDyZuP0stfSZMLTfy
hB7eUjr3pdIoAkeaZldLRjlCBwWFtkTbqCXdzzSPqLvOqAopE1jjmB1cd2jnELVmN1zWZ1Jq1J6q
Q3wNh+j8JWGVpEHKyS1K3dyCrvSvP6taVkc71bYdqMom1h8Hoc8UDbjmUeSm/3Pzoaxv+kn6byGa
BM9J8Mlm+ATf9C70ncaA5SeyMzZBcuCnVqvNR4feiCvsBxWDbQa/7kBzvz1vdopNMrvWyzoNWYI9
Dwprgq6HqhgXQTUhwqCEJvlIxdAEG7yjj0mAojO/OliTSEpCJKU5lfyBY5x6ibmTbnzywD8x/9Lk
y0PIuzTQ5BrISzllO76Ce8pz99XGOjjhO9Z7UvflJBJpIA0VZLLDztvW+vJq5T3AR6yxgPnGCnhL
qKnMakWp8c+2/IH/C0+iGdYg/4xmUe8Qv0eJAj8NKm3SnQfVF3lDigUuvRj4hTFKV1hmhH8OSdz6
u4nEF8of1llV6PFkJr6A7XClx5v5oiK+SsvZWvxe9mGCWPGfRw/VB7ie/f0gIJ2yQ9KrQBBc00Tk
otmqKAxX+Q6JdFFOvnC/7p4MnchnZ6YGHmaNasi2vFGKtkzVFc46C+Oqpix4ClieXR+f4U570eOQ
OD/0ZJaiL9rg9iDH66qTtffWI3GvbpxqnGdSqwxDSsqL6LBmAao9STmebVzOwb+Az31MPOaVN0PT
fF/zFKtFMTVgmuq119SPGRL6/CSJRNGCiX4xx8L2ezMz/tNcmK815oW4j3gQPg7a3uraJmu+xLO6
Fo9hzAutuK9AM1cjVQVKb9YjFbBjSRHAnvb82K3as1BBVOvS+dVeBb/qgI4fu45T7nbBaGEJYKm9
vEEJCmEUAEMU4+Kcu1RUd3Sh8pG2q4UTyBzFejZyRkxOKHU3wF+0PwJIN7BwsiGs5WdnjcLUi1ZA
EgZkrst7mBPcQ7OC8IlCiZ59140qqnG7EcvkIWRidzjOfetO1dy9BF0pUwv5IotrqLNHcKCQwaRD
2DYHxd5fpgQkwJKf2svaEjFZ5Y1VY+vyOJCzfmJMiT1xO3zCDp61dS6rPU82Iwhu8vjw6j34ZWp4
UNG7ajiAKxKdNkwXFoV7DK4N/i6iYm39d61wqmJIug818lsBNIcUubKjaG9B4T474f6YF4XoDMD/
3p+Gq/G5Ok8r7XN6MPyb43BCe+2fXkzSneqSMYr8u8qIKm29AZM4IOGNaxp3Glk6xvqsOIV00U3k
kpPdjRwV2yH/Tqg5GF7sVI5+R72XCYi2hIalDYn9att2HgtxSwCbqQmRubqQHi8bHzbAknR29O8O
NdvXxcnAXr0IinubfA40UALHXgwHfi5HMbdgS9BHTzrktvjbWYSp/cinEksUSuLi0QYWghdfOBmf
jL/p+JJDlCvZsy722n2SLkO4S9ak+sMK2DN9Xa1oRttOHIY+4OsOWGcBaffsKQZt50ktw5Ndkp3Z
S9vcwBCiDoerP2AvOLyELgyulg73pqaGDzlp+1M2cnmQOx9+iASvELvIB0CyqSYQh+mQhkIuAXJR
faCdNs6iG7t5pJbrvmWJhzyh/svU3Hp1n0LBNptZCRjSYO/adtLglnMe+nqaEggcGQxUva7St05K
rua0UmGnVAjkPlBziyK7/Nr6EAXOOfQtNVQPU+PWI+qdCKzbbPiKVzQGnrGWwQP8H812GfQiLPmg
G0TMWsa14B8QNuwYPhRnVdicSCHHBK1gfR4jMB4IH12n/iGClpHTBdHLbpv+jgP1/ijex3mKFdDS
4+Htv5hi+pUoHtbhk5oPNGSHaqFtydp6vGoMYAHOwyRLUW3bx155B3EQ7jpsQ2A07D0p50PBb5Lg
3yPxhmfNL+jyIQaWSSw8xzih4m/i83XP/ZqgGmyvxYrvreaq4TR+S7ju9xQbbXDGUlOkVqzMlg1C
TqgOc1qHFquYk/9LpZvuX9jYqRhoG7Xh/wC5Pop1NjsxlRruqYhm8O/pl8bEd/ifkRcSgTaTsZq9
lj/iQQr9wxkIRF3d4zcjErCihmF7jfBcquYnMxDeNLPSHF9sSCRdjQT18bM3fm76GDsv+38L5O9F
nTr+I9Vi8Y0SvKFQgADBqS3SQZ9ARlNKfUiOLd5MyHxmhsbYHHt4PD4sziFrJ8aYWf2Rq+yyMwCh
4FBzMFirf1NaB0Ee//u22FLODPjQ3c55NfZ6gefuiMTe9GQRcIwU9W5YZCIiTwJPewBsi322P+Pb
KUG5WeWyoWADpKTZw/qDLltOE+TNdwdNQR3D2M8obix991ai1YhhgxOfvi73zZHJphEeST6qhv0W
/ZSd52LJIh7lM6t8X6Dorr6u+V8yL3wrPM2pLVLVnYUP1/LYl5yzR6jVMbmn36qL4AzImHuTSzU9
pNoa2FfYWEI+7+dNvtYPnfw72bNNF3zcYVpnHPfiQ9HBf4bOL53ksaqPSNq8SnlKlpuqzxLBj3xu
gFjSK2QJ7CN+ly7lNEIp+wKKWDgGpkpdSG3EEvK7tXoiNDdjRN3yzE4WlBucHkcz1y40wpKa47wQ
hhVT8bYxfq+mgaw1yNm++HLQ4uxS9nWWq2j2Y2dqwXyWh8v7LKBW0Aac379eKn1QudvOGUqcPZ+d
ZkbT3wroZmvhJy6GxDN7iVmgWGbQaGlniMgMNmy3rE8x7rt008Je81UcO4ykYm/LkMKCAjXAKazB
DUKCezG8aLIxc4spSwuxYytrIVmpJyx/BY11ARdOnBlMBlePbkH9CkSdog0t6T3ldqNtEAiXesQG
UmR89Zo3w3gCOqlprcmpZyiBXU03D0yPUJsUsy2xBKEMgz5Rih0tc1l/DZ3dO3+LKEyL4TnbS7+L
+58/3KbZl4RuEEDCqfoGTYORM8oCkGG5et/AlELlLM3xtYDksA6f/97WrPYC6lKBNSdbqEEfuZ5N
XoPymvWMusMjaLOVnvnEDcNXRr12Kv1PWFWfCUnBVnFGv9ks58czvIAdNREoUlG2+RpXVE5nXAFN
7N0uiCBMb2LgNpyHV96LZILfrv2MNl4ALF3I4TOewPmgyE7qd1nIXQBfqz8yqN0GlyEtib3dcm2O
Blf9xMXbYwo8bs1lXz8l2ycKQsuyl7cyEU/OBcjXj4uGmuEQswCJvFQpMbdBt/OXq8PmazvK1qJx
LJe2yPuuVQ2fQWhPPL9LozRjsXgmFgJQxCR1NHBnjVsl/evqZDStNWXeNi7PbqPYOdwa+wVyyGm3
sBzBWFrdV0LirtPidLGRZ9LhfcaTMOScFIj+3ps3H8SL2s1D8aa7GdRGrUsyLzYYBvS4UweBnw/R
TocHTHEyIXbS9zRdyqfWnLr4iWyePoHc4U+MLd+dwDmjxoGE5Bq6ZogLdh0h06yAN4qp0SDC9pnR
SsDvZxR2vNIAXbkFyflrPp7Bok9qpUKcjadAY1EbjpMPCXjP0bWnL8eBgBL+Uya2SXVu1cJWrkLp
mAA6OWJ8X/QZAUd2upFSEgMbxKvwMBoZ3wSleG8t/qFR5gcvoO+zplzOCQyUoRc8Yr+GVVnIsvzD
hMTb+PRZUQoAcpsT4OkGykRpD9d9eMmxvaIFKtGNKfORhWzI5L7uY/y8Gr54VgxHfzJKETiuXDO9
FOEwu9xivxd0gF3lCjyfq/JvRxSU2X8IFkD/ck8RAlVSS7fIL1NdhYEaShVnkG2dFyRGzj/IAA23
SQnfXu7PhvBmobkJ8gZKFyifMxgbEAyjw/8W48hghEgJzziO/vkRrtxIoGdGgVNDP4LflU9og2dg
NEgWujxlbmRjy53AxfV1M39xpVqFPoucUcR3OeU5CjdmieioJszHxUEOVlTjKJperfVQgLGLQI7i
ihyjtvulueBz0TEzXh0+xGKIObUhdpKZ7BYnvqj54ANTxg8Zrvj3KqcMliqacqESJtBwMlFpNvw3
PWnEd4mCbNKRvCTEVziGlM+LZKa1xJe4hoJC3J5dDzU7b9uWmY5y88cfguY26RXIyHD56A3/lR4b
iHFNppP9eN5pxMRQNd6qSEmv2hz4UUfoBUU+uEQpp6+KjqIgV6DUnVSIZJxzx+y5ka4FAry3vYYq
/AyOJkb91+UwNIXrbjqBphX3nzwEuQmFZ8wJH80AEtRgSWA+UN03uwjr0yCgE6mbydxSD9Lnv7Jy
lgSl138k29JFHvt5+f3MTHVPJ8t1bsme+/e3CM8Gk3SNbvjAL3Xn143JXT23o4sN/tBqeUOmuVVJ
inqWrak1aeP0vdfQ0UWMWLv3+F+GZi0m0M7bbfBXsb+7b91Gm4Sf45GzqvT9G7/HKjk6LrVHHRB8
i0M59j7jgbT+6rFc5WATjDWEbAgx6JAH11/wJABBZK5A76HysIp+Q+pNF6S5lXDozWrq1NpSgeMH
JHTp8ig/+6QSL21/4Ito/xWZRkzTDXhhVmd55A8sisYCtVBC7HNjTwaPL+eij4GKiUfNqAPs5A+O
oZHEnud4aGdD9DWIGwau9a8a7SP/DEFbATe6BVxhyM9fzEm+RAWA0NodW/F3wgTHV4x2krUpZ3bC
7d5XRRtWz1Q4kDtpO0clNolrrRWXqOFLG/q/vlHBgjWrcgfp4D+xpr1NOf63G8mvPnplgAgcww3q
GnqLSIhsexyp1R1LL2c89cyZ/jvWyCqh8cMyoatebfFJ1cyxAB8ZfWXEwxWR5aShUNiix0a2Tfi2
X8+T+TnPwR0skP8RDspSHYOYrhOOwRbfJqTkOq/I2xDO7eNjiTXnkpO9G/nHVaTQH42uHZ3VrFPD
LFAVfj4dU/srpejHFoJ0WISR2KCGYQtyZ6RpcUDzmyDVRc7j10DVMEXrene+5jjTfW/ewEogY4/I
pXoFdpGThv4Xs2QwpdV3IlainBd9o8oFBxo93FUaQSoZmKVgr5mXMPKHoedhftKvM+baE67Tf7yN
JRuSLqfIBIScLQNq62tuYPyUtiKCP0BOpRW/7TugEN75/BFPXWPLCAhCpCqB/N4KGgVdujtwZoNz
MSkeJxh5CkwmsN1HSM02sneO/p2crKNk6m466oD6izIMjhAM58bTPVluW4xS22Qz3KOmmJlYwl3l
v+WhFkCHYTOZ+sHl4DOUWYiyP53FXR168yYemKhPh2sYQfu5HX3a3OnTe7EfXkYL4/dkfU8/XwHC
NEY319DV3+s4j0NEuyVlD0LyOKV01rOVYEyn8rDg4kPTRRzkRvTepF4XziRxYqTIpVTNKpR/GoS2
mSPYGVtB59TQnubPS/XDnhfCmqMRDmwovGu5CXhV1KWBB3QtawENixdfCocOEMFl4+h4YqCAN0S6
mCh7RKBDxoIad5/pKHcMjVGV0h8lMULVT7SprthiTZLOHpV5kDVP1ULNSt/5xIgihe7Hqc8tH3gV
tJtgWU54DABRitPoz1rpTWUz6HV2mipkOgWR/lBUnK8HVU8bMgvA8rOOVqioWZ9PeLHTq+Ep8s2m
YOAq0848CnkPIVoDxi5fk8zbIYQZVxdwdZyAEoOyZUfgXtUHjPuoEeqU2+E5KF8vG9+uKyXoq6Ou
sIKTvVXow0SZ76ZaZQj0kYm1hIVwstw3VgT8rh5I6AwDL/zcYFO+dudad0fVWiToDykGddfBXdlh
AvQgN31qVYD0D3x9ALF5FIxzC2JGwvyeOhHtfo8rOKHlCfdb3Wv5Nv3XrdL7CX7CFNfizzHbG59q
MegrPLe+7kMOPjb3n7E2LGVirDX8YT8W09b0VcbolbuJZjphrVfTfc1iD1QLZIzkBrzkKn6zMujw
6KK+kHcqtfMIPeWXgn4ZIiPFqtKJfUXQDzpoMPbC2yxi4lCMp5MI2qeXf/tGbdRtNwn3AF9tD50s
D+wuASg9khCvd79xpugQgZuoAybK2YKV/PoffXjh3iGp13T88h27mjdbCnOvYqX+2n8VPZ7Ltgj8
EnBuzvQvggiZbjdQCFsDyALt0eargi3GnxM8/cwkZ8olE8Son4dfhV1dw6185d2I4HtVRNJGXkpE
IGubB+YvwtMHLVGYW7aX2DrXhuvUJIFHb9d/RiIono6DBveOEIQvPaqWVnr2yc8AfhbcHXV6XjAm
Fv1duXNvJTrdax75CL6ABiAuKTRkpE2EEvzdxebhzbZE7eYiwFrkHOjtephUJreAIlW0ptEkrziZ
GDckrDYa6PEGY7ul4eXAEsfDGUVDY6SmFm59EQK54vtsfWy/U9i5pTsEtWDl8RU/Frzo1bc30OBb
dEzz9ERjxQ94bhCW34+cT6YSWBWcmjDSatxo6xAa4/XCa9nbeDQ3k5yRRpsWNP3aXtqOya1UoVod
GVgZ8NBD8l6NDfGUbLdCfCGJHkDQfhTi4OeJnnkayUlzn49wUJIks9fj0j+eUwB3dgu9FYGezhBb
PS4A7TVc9OCsFyZNKdv19UJ2OnthcuqrQII0/Ickags7uJ3TPrLdVkJJMOF1HyO1aXp0zQCalD2u
yLemhLytFY8Y8fn2qBGqJDZeJ18LNH88PPgm3bC25PhSAfaS98dIuPsowOdqGmh7flKMIQqyaX9y
TVVxHxZag2ryUxlw6rrkuXhqmBTvnWCbS3sje15Jnp8niSP5vytVdjtikvmKWeSpiQoU2fa8q2oA
vX/dRjLArg+iL8haIXc8bvjqd0Pw0OJJLHP5phdvfl2nFjeMxK9kDWUNq6XAfU+hS7VPBLbJYmCd
KptXVx6JFNT2cTx6PaWEFjr5kiNnsG40AzRZgR0bxKnkdnGrOj96csYcxAVt32aZcrKGMMzXeHk/
UPx/vWb+bjnS/4oB7FYmzkYRplKk82bmhS6GI4JQ9gwRmPqhP2yM+ZpFKMex1bwFZynhxQRZ9lTw
m8Gp6TVgpRjEZ+2IfavhVlBcnPoqkL3EKQX0y/LFmOJ9mDRbR/wRWDTF7u4oJO9lcTT8iecGjifr
R2Ur6kwxKF81U2/FZmqAR1QyvV++Nu3flSglGsymGMS3DTPf1QPJm2HStmOwbokWpLUv4e3YMR6G
KKpapv/o8EQcacHYbQHt/hIPorgnPvrmAe89T0rYyFsMWQPSKwFhnnQtMLVL2yA0gRQtSvQnBCtr
DTD3u5iF9SvwjDkoS98G+L5YkAoj/ziMGwu11/t0Zj4FkwTJKzOckm3LtxpvxlMtF33HvufF93Wb
+XbOHgnzbeHFy5b+KfWOoq16rSBQ4mVUEXnVuaD3UyJQ1lt8I3wOe4k9AecRD/XVjepOPLSy0AsJ
UtXLzF1Mdj2J0r5JZnf8SnVOvITpBNRBl2sPCjg35iZju7wOhtwS5ILRQz7soLSa3nNKmydVersW
9XGkfpGG8PyjnZ8aId7U8SC34PqWTjhnXgOwM8Q5x87/ZTlaVDN9Ze75v+o2fMMk04winuftJkH1
4t7IsMlN2gDihZj0ecbF0Rmg9TFU8+6h4BpRrhmwVhFAaj32eAEgnsaqw+UuqqkfFdNwL3uDOgtH
ktplX9CgLnH1y3AfV/k2JAN7S78N3GLYrjpdhRGemmhJSeT+ktVSU5ZyxQSVG6+1QDgiGujDD89f
Yo+36SIPMqpkRKHNUVuQkzCXITBPJpaRIleXMVMMK99Z784YLibP5S4zS2pVpA+bPjmZMf4Vf5e5
rzPIZVTR0scTe0DyUADWPMSBm9y5ak17iY3MUnxrct9Yu9GpmA1XIlgS/Z9bk6arykisVXPu1syy
pyOzgx7ghdTfDrHSqqjnfVkMBI+sUWx6XCaue6jOHsCgSYmb0uus18y7Nsg6ho9128h8YR51zD4a
iPbteiO4PnqXJVveBBfspYpI+5T2/914rEgf4Mf7QniO63MF+nS/cAS+6rZCJhdIYmWjuNg6ZH+w
PtEHk2SdJ+ql45YqXKalIktNXpa8mintXDlnBCSuyQEyOa9HF2OPeL9Y3H3NFfnLxjOzUUIr8hrR
ldWkV2GpU+o70HQtTQ9zkEznp44QyzYD4+z4U7AWkM+Iiesd/2i8NWIrMh+PcQyoakTFcBAwZlVv
dYIvtgpgKfmUjQZzLjSHeFEgRJUWLX28ydMT+1LNY1ie9jI3tTEy/ZLuH0bZDwh+ewIwx6zuV3Yl
ZgoeHLIDSbgKfm/JLDbOTS7CGfoUEcrOvGWysNXLq90uUZJmMi+ITLzyL2ChzMQtW7mytqDtqA+g
5aFPnpwLUN33syFf7uqqFFihPgpN8HdoG+CuuIl2hUESqbIXkIfAYW+fA/8/ZRewtv2r7Y0Oecco
IWa74PyIVNxam/rLp54WvOn2YH/DKq3XNMS64W9hLYFt7gGZ0PT3hYVnA3Wp2xo+a92RPmZ0N0Q3
nmkkwpJArXstD8kzK/R1BjCDZsJ9t5MUYpVeGaSpUsRdTEmyDwuDsizD6ymqRHgQSA55G2RhotoH
MYAhSxxUA5tYy56coJFH/hq8kDYjA7+P/ItR7mPOPKBh+1/z6xw955kU8UJPUYjW++niePSqPQlN
ur/4Yr19VMLhWmCftr5bGIRwg3+JBZjmM+z+TkrQmdBC3opJjU0O4dxEAFQMhB2owruCFKNEC5Ep
FTdiDDekJI/JH370OB9b45kkF/FO7NZMXkprlKCilveo4L8Z5SVHk2s+ot3q6fYOZYrLF4QFXCXH
F048pFoBJdFo8smwc2ecxfXsH6lQGD5fRV1LFsg35tTseN49TrApnmKStA7oJmQatl46jieO62T3
nJub3s89wCeBOYx6KeS3NwbTQgsH5c/Qoo2jPpTng1hai80zmw0lYsmlzCku9pZZhnmjNABn88Vj
p1PMWLeSugdharvROuXr4wygbaE3P1MiSc+LhQ4kne7/A3Pa7v/On89/dTfBXTmrlaGh+7naSr99
qi3Qj8Te1EoJsv0KyIPOkVfQkSZiL3a1xj+zQOzT7Q3xZlvSdHQiUvfn46NCfPo3PUObkiznGwYB
KRtzFgmCWMsQMtwZ0AoISJTSJw+r1L6umBmAIEleSJDTEVT79+kATg+RbU6T42zl5OzzV1OCmc2p
PuB0Jb+WhI82wMaJAVAx7noaWRwin4zB8/qmXFGUfq3oS94b3ZLor/I6FqsmbdU+4tgBABVUfoi8
w4iAKVc6ZnjqGMS5BKV2GHIPmyDGCAxGlKcEbrAxhD4ySh8Ipr6amFD6G8g7PmSUwVs1jhJGn+Kt
H+avB8rkkhfhNTmQ9faP3dYfwBFIuO7IRohNGLhPW0uKybBahi2Gz3P3R03nG3LiVPlaDdH2/CP2
BT2LZRgR9zQsm+zhPMv07kryUz4IV66I8awodc+AJd9rdYnUjRRTq0BIvK1+tPTCl2sXGP2BSMAc
IjaRYD2knyOeAzXW2OJJ+88RJ5oLeILl/VpvntfSWmUmjE+cA1LQFLTMT74T4KkoKoJNicNCP8r3
HoTY1EdLGzoEC/xGTh1iCTN4jBE95ReJU8jc/YZLMaardO0j0coRfXphx7v4jB83wh1c9214PFip
pS/5t6gpRXy4Pmdp7R2cM/U+sAG50pA4gv4Hsw69sF7TCVAIk/CSU9OhjawJjR0IUSASloZxpX9U
jhVUdm3Xp7O78UpJ98+ffCe1zCRmTxdii4S9tXFiD5IakC7CMALm8F4XqjzAirGahrTe5/AJpzJr
26zC6p9CaMNKnXznYo5/M5KbraszB3vQuA6ZnZX1Erc2vymT9Rdo2X+8Ps8hqM6AnUWq9CAC5QdU
1x5jEIR380u6Jk560dESMK1Q7X+ifbmUJUfbuXguA98aQNx6otoWFpL3w8Iszb6srgUYs1CyZZMG
3oh7/AjWoTQJh7nGJNI394EzlbquI+/Rmh2B4QexMEknIlUuY7b6A4+EY2tWvzg97Bc+4S6YzJLx
urXBRheOkQ937VYuQjEsvMhZihkGNUPQXUAGpp+e9SLYbAMtQ7heb4UDlR/uaZV8YLcf52gNEOMV
tpmIwwHrzefT/7WLbceB+nRd/O/dYh1a3CRoc+YzhCuKH0pLitIQpWtcjNuS6nQAXwWQAG5h9qTv
PMKIokWuHjQszM7gVG0y1AU25Na9eYFzKS1mnwQA6cZDHIIx42J/a1hxdtOJW6cDtMPPC38c6q0m
P1ojri93UHjSEfePZ2MF/ohM53+ulfeq0SGqEqbtddfE8z9BJaUvnkis8JDfP+op5HqZPPgv6Liv
0k9IdA+2EBFnlRF21ScV3q8Vi+xp8GhNFKQPDbWq5MOG9MSRAHTkw1yGRCSdq/X77wGWv3fZhRf7
d++KzXRWlK5GCCIgg/igiUgNKQF5B46F1D9BTDbKUOITLzlKZxYo4tJd20fKwCcxJ4XGDApP4Xhu
xpJtJH5PBV6FMfkMqJIsx352+zJKEqXBpHibbay3O931edQ49/yWpo11+rSIdiq1ThUheVzPA421
nos9D0gaRSL9XILTnjq4DaOHT4YGuzZ3rgldw2nlhQQ6G+iAC+D3xQtWZ62RyjwwtKix8lUPwyrP
cac3FcEDR8RhCiPvDOT843pa7coDyVj9Jf0xnF/M1zDuoAx/urVwyrFLQIQjmFwvtydwbrtbA0yU
B3I4eMr1A+GCxPZtJ7shHB5p/A64rpbM6GGCPDgZrVn4I3YyQYAsMDcHBuOdSOyWf+CMYYhpM4gM
ubwG28WqnWzUWQwOD/pYLx0pRiYRhXB4NxyoX2rT7tlefo/bSui0nxsN6o/U3hXLZu0Vd+MATjdm
O2b3rQdU0n7rghOgr/waUHQlNwrQNw2JSTUnbEACKm0V1ar16CFs/0gowskWC1XHPS9SDvqkW262
0emawDvQcPOWK1B/PaC2scSGMuvcFbJ6bz9fptTcUgkIliGlSySp+41UTRfi/v87CEobLFTe30zX
jjD2m1Uxq5X+lGuhK/y4Ub5epUfCSvORVhTqDj8Fdeqv7W5fnucja3X3/3N55nGHG5duxie8v6he
GT9ir8MDLEqF0+WKXTXjUVnmkLPrVCoBKhxnXiDM7MSqrR20UYqh9wfwsJOu2yJHhbnBk6om8zJ9
d4aYVXc91YycHSq6aOlMk/2NhebJ+kGXejm000OAlQpzmeDVtX2lSdwC+mczu86y/nrO1l2fkcpB
G2CmwOYyPLv1I+0dBEzu++BOquoZgoue0We27UlOcNGaNlyNq/a4jBS8LbA9zlQYa2Fjdi6hlUL4
XlVtRxUhfOFuk0Ry0uPhn66pFsCyo+tRD0QSEfj7gVfpGKs64ew/+Fj5YHAb/WygxAa4jgL3lO6W
UkCV9WLoCqB/XQXWoaHC8X/UyfD4E7ufEgWdeF7/Ns3uF4HnGtBrC/hgJUU5XcrxCt71x3iFw/Nz
QkElAx1aU/zo1xpIs7j2cNaO+dTrjb9X50rLQ05UxCIk6CExsXeWYh0Dnmrns29Xt9MjvLi21pn2
YrlKjloJ28aLzl7nT9ovDqhsILFyRyTbyMj+iL+9g7bBh6PD5eEjxvBlw0eyNVj8PFTH/fDGAo6P
64JCe+HnJBpthiUvQEWyy3+GtrCj1X2SIOy5ZmnEhgNoMIfAOocNzLlGV1S5eoFDgI2OWq9rmFTj
Ci7Z3jGL1Opwr+pqr//sOkML56zZoo8ExxFRL4LyoMgblLhJ4iqiA3E97G7hM8ZPHsNmsttdGcxt
u+7YhuDoi4HQ885unUclv8e8Z+jKS7vSk/ImPI7s8H7sLiGDIFwRwa/amqC/ghHHeVCTwBA6DrT2
vMUDMKw3cDGvZD7WdI76ZTo3+o3RiEirTkyoww5+pn2bdNhGg+sx9yQmeafbqdG4Fd4gQQUAaDwP
2cK8u5GW5sFUT5/ZllMacJRaCLxTakTPEM+wddDIykvZSeiBxKypZ0pMme8EJk4l/vL1UMfEeH2v
63o3L3bfyjgQIvJbC4CWafn87L40KEetx59Lsy9+AJN2a/yy8fW7KP7t682mnlibx26/Fq4W+p9q
43n9W9aTzXGC0UT5FRG6KS4w6a3RYPoiKKq452wu/MCg8vymF9pR0XStVTKEVGnCyRb6LYG4LshK
2Vj7wG1hQdbtH6aO0WeHFdpvELUT0+7l1F+PJZr85/1pwkxQsdM2/reDA+TCFOF8+lnIDSW/X/c9
DXxSHDmptvprcaO6MvAG9iGXo//WV0xVz359e+dI3YjQwBZRMgl1OHPTdA0rPQvAxGpsBdMIh36+
3QweXl7maLSUKZ6McEmYS7c0+Z3ingRqJTR+8VVjMfOCpSfVj/E+QAvKk7Derla/Zgdv5/xo7q10
ZLdNxOsGS4HUm3Dlj/dN9WDeCq9CjuZrf3jGb8HhBFX6+F8dE+otGIzp2R0EYV6TVQmqFwKqqhnX
wacroR5sxkwguEuoyhM1w/jB3QrS0aKqhKy1SQpr/VSsTfitHlEUDAuvr5gXZGWxiBsEL98+U+Cl
IPVFCDeiM6+lNze1fYv6z9W9MUClzunsYnDDHZhJTmvHa09tsB7FMOftP0B2qTxHIhNn+skVC5IY
kwOSoBweMHm+BGjdZKB8JYA2GJOpnBIgtP9Dvks0ye+Uw3Nh+b3X+LhdosEmvl7GY5Y7CYqCQNKN
nlQH9Mn4pXLAoF1gnL1OKv6Bfm1sP8n2Rs+ZhV7S7vbd0kUJJ4uoUO2jUxnW0z/WCv0Pzgf1guwG
SYaXGT8NgWfHWdLw/ZrQn1XS5zZEwR7pBKi5Q+aL/yUH5DjRfV8FKLc8Gvd5os12fGpo6RKGSD8z
xHQThQxxnKRxHhX1LqDpTKcN8eL2+FRFx0Cr5nZV7xzB7N5wXTloZ6YF8Wvtz8hbqFkDmw7uC5vr
+lsvzER7RaOnDDbZ30auU6Vp9DTYLJUjg1ihhDkekXxyLy68Who3xzOujVV7IrvaEC5Q64DA8SN6
gKP93a5x50iHSYxsRRA2IY16Uo0dHjftkg3NW/BgmGJg7l17xI8C6Uu/Nvk2wQ5WHNHGuuFKecJF
8SUjvUdQ0mp+TE9ZddoKISYnIPQCsN4PiungVtKina5bJU1YjS+uack5kQCF0NM9qpMtr16EVirk
dQMBZzjEKg8daYmHpGOdcyHUhypDx9vlwa6QAZusXpi4v9dFVYoUfErsaUVWi62fC2Yq2In4IPh/
PyhflSn+LjYyTJ//OCKWrYurrnL47AAk29eiPOxBuRhf57PNQeUMSAGhnXZL4g17ILEoZD9Vid2g
bKFBm7JWmgikof+w+W32DSmDYWd0eyNwksH0v2142xzOOEM5ONHTNS2RMMYcVhHW/5aGMFpitnI2
UNPV73MQukyDJ4EU8fuCagKJ1KWsq3SQ6k3382d3vcOvpuyAj8W0/7AmQURbOsOu5aXh+1J2ckDf
Su7jucEX4h8KGtAMT3DxplnCJHUGclU/M2PcSZLuxRIDs1eWRYNG61DZLLGJ0Ls+++9j5GyCZPXX
MnTWO01Hr0BIYZo926cXveQjv5CP2sDpPXbvlmlSQ8D5sxj8D4AbnM2rXGgNLprym4EMRr8ypQnL
HWfHQoudvU+BH73u21o3/4twrbc4o2gC1M4q8y9/hrCWmHzuj1pZ6NZPuIctaQ+nkxNE0zIwkNYE
Op2xu4ki4XDmFXuDVOLkHMq1GDyhYJq0PqGqWpqXDSid/4uKKi/C3+FOdme0M0DjhNRD8avckYhs
6yOubfxgD2QC8RA4A3qjW5ggooJ0N1x6uxTVUhZby3W7JvLEyV/Ij5eoQZfR0j9WQitfAn4+SDkd
h3rMslww0Hv6ZxIAmPq7q3pZU0KcjuyCUWrdW6pUavRRXezChZHMkM7J+SRhyt2Kf/4jLmlGJZCS
Zc/op9apZLIo21EC3rhfWhu2LrLbnuzAEUA7QTOB/12uSaViEDgV7Dzkqk2TxQKPjInnLd2X/Zsw
YLqAAcIkqq0keaEb5UIb8qVThER5/p4x45NHyxOcEDNfHLJEztCvBqZ9dA7o2VRIuZbHZlVYy839
4DsOu/2AgNUTwTmkIJ8mqhHsj6lyXe1TKEqoTqU6NSjiCyDSoBwMtOLu1+3U3yQoSW4abEl9nbET
gpa3LHjqyl2XUApTUIFva9Nir4oHwjihLzu9A7r2lb25A1ucQb+h3xapvXdpuZpAaWRdG7DV+AB4
EM0TDITgu0Z1YNp78xUgh7K7kOJqVVWmACf6sLrNpekWNddc9/IGcRTXhL/M6bPbawFH5ylfq9AA
pe/XLhzlSoXGARsn3xje4c8cCifasv8iE9+YgXL/SNhzgwXhRG6zu1gKEKkOxCVDDuyVaopI6Ol0
Yib2Qu9mV+QXaSOoUAIMpqE8fXSTMnHZl0M9rKOAOs8z0EcyIjs7fKvEd/CD3owIxlnEc8lKqP7T
mtgP7SVZizWc2cUElPW6F6YqyA+IwBjOkaXsy24ABI9RdWMVWYVRENwYiY/jIW3lGBRks5JIi0O8
jyPG2XQ6OFxvTVLnrYt7kTk4W7M0MG+IxdoYIIPSYASkLmBhBbw5fs9jWVsx9QEad+tLfhuMTojj
DaRn8jaGpYVQewdzeZoN071Wl+gflRsxT66ez+ojGoV4LGW0BPgIXiL1NpO+IfWnO7oZ6L5vltM3
PIysxZiCXlru+xM/8Xh/0KGSoVXoX7a6epWcBwzCilWdqEKrqWSiAAZAHZalG+zPQkli10MHFGqF
ICEE8lPbszqksWwt0FK75mUsWnj3H7Aks1H6G2/Jqz0YpI18GGzA2e+jL1p1ojlC75TVUMiYsyDD
3vmL1Ws//rI+OiEbacFTgOepB8eH5EIfBCQ5b32jF7su22U8AQeg1jR8wpJAaNjVCCX8/VWlRffc
QrOWcn6Ao/MsKlAUqbvFiIwprmE0eQ77z+euGkQv+g8FwZTqAxTytvsdAfNZ/QjE9gLsdRZoKj6i
EXL60+70Fvff8rxcXyr+1wPKD0lF+Mu1VphrePqlGhx+guua4lDYDBwRCPEp/rI8+8nhPsibHs6A
URHv3d89aAghDbpiCA01Pv4TXPp3PJyd3hfABa8oTMWcd5yCwvgBT4S63F4okMfD5lZRBzSrowIn
MIykYzr0eaIQs76KbAAxTZ+szOo2Xi+yOxBtW199+QCO5ovFf8ZHfvz6V6cr4c4maWXB38q0IXBa
FMNONQ6+W9g4uzURD4zLt88IpkgD72f+dY58DR62G1eSJgx2Bnf40dxqoPDR9Zwdbyg3vv6/kIU8
enPzNRkfxlGCVyHqpSzWUbD+zPo9ktCrYsWBT2lA8XKwLBNzlK64H2ij6eR9vYi2pJdKvIdunq+D
f42uhVPScDbiKte/LCIEEnawC5BzgGgiyeEXFugBej9E6IVURZMOPcgZ1drovYs3IvrwNtABeQu+
aYJqL+A+Shc/VLPOMZaQb2N+wpa7yJgWKiPnMlho2p0Bs8mHmm1jX2kMf9xJUVNLQogU6j0lAukh
0O3HPdcH4pWHpt1S+IoS9Lv02YfhlEFzENqDjmnHWlZvLISJiTHFkd4NgJb1pOpHHQRt5FLU9qfT
zdmB2nNsYrz32L8hsl8dvl667cvDyRvfQQyFowPpLvmPTDlOV4Sd4AcGZ0IzHuRUej24RkvWPwjP
aw1DrSK4klryjssZWT4s3S5YCxUNTk4T/mGhTVvJTvgGYyjXS/SvqIZ09M/ZTl9BJc7zT/iUvfRZ
WB0ZMjgGpi7Lg+0j+28ix33YT7iG8l6eeHOAZWXQL6JhdsQGbMMq8pwxUVf09PKu+vLUL2SxcoUh
XAmrhx+FQBxUCrcfbeTOH00auhU5RDZPqyriBFwfy2dVSCcg/yEUFKCJ0M7r2u7vuhzByBQhmdnr
SA7b9c4K0+z95yb7lMwwU52SNEUps1KoJtygmgOzArkChbo5rOVFu5BMHxxGw0zfvDpXLq/nW/BS
YGpWuBFQJN0UtLtq9YE3HUBqPThhopATI0IINdJCY6CYqP8ShtqiCXRZFLj3GSLeJMiRnQmZYu5z
Vys2+sVf7YpCQUI7g/YfOG0n//Gi/0NtswJvG9jbZNxCmGa60l+t0vjqHGZMj0jpp27I42iQKpyy
JbTgkv1io6U1T7djvWZ0krPIAFs6iGYoNnbdYh+oqZwi+LaAI7jzl7lcUR14pmWkwbL/fnol72Jz
m4DTVtR0OuEc0Gsa1ehgzo0Yx/OshxyCC5PV4JW0n52mcA6ne0IX8aA5nsm7rr8daX/Rl6UnZkd7
13NxQ3ZCI2pMgLMom5GRw6uJ/bXJYBDHBedcQZHOOrX6pdY7yxkCuvhYpO8nYi0ZrcNIS0i1Yw6O
OcYKUw+o9nu87UYC7yceKaJaTKufDZfcosbZvuvLYAg+A2BW7HYevaqGto6S0zaPWME3WcVU81g+
E9v4O9wMUnLSod7Q4CYD0T9ReGB3WplMd9Pd/tSjzgHo4bu61xrHVJmsNziZdstx789yPW+LcIql
JGdAWGXRjlQYEHjnwYo/6BHNnGmC4l1dkyHiFh1UjJeN4bCduSAMrd7poTsYhpTbTrWE/OLYXNgB
SCABI35RsmNccbp5TXcb2uc4HdniDYM32l5NAfQvgV0Efcca31SawQjyzrPF9FgsL1dWAMYVt1y4
CKa/ubux3DuwzinFqIigsiT/B6nsOvueC8NEBeXU0KnKQKTF2Egq1aaCnIiI4sIeAhC09CPJQUPg
lJFjnryzUVj1CgA++oOVTcZBfIRK+T981sHr3EaTjXOJHCHoRJPA9obZJDFh35Xs9d7JUuXVy/Zf
7FEFlw8Ucl3G3rA71xtZ3VouqM2H4efy/AWsGBiw89wYmd/jFjx8Q2yFjv0q8TBn+ujPVvyGc8tY
ghxkj3E6qmnGZmav5Em2K93dpTRZSSjEvJqAZwiwxQgSCsU6GpV2mm4/e6qMo4y+DBdKSfZDyInz
qoG1zAyrZ3/BF1UCfIpHk3vqH01L6MeeajyMUKNtf4edFNL2vhRaENeCpn3S/BB7OWrHysJWHwpb
p8dBqMHXPWzUKc3jZyYYiGSA9E8Otv90S7kfwoFjHLUdT00A9mgWYSzG4B6u+c+6dse1Om7VNfZy
EGmO9RbDMRYEO1o7jBxB6FMOmkJgIr9C7UieTsQbZbxHJidyTw/XO68Jc4+uNC80uyJmHZZ/0uEp
xH/gMwrMcLrhO6xAEgC+ykJlyQxGHAr5AV1CIeLBeq1m2cl5fP6hGYU/xd+KsRZ1kmL/BvK4Ix5N
zsWWVOpY95SiBuAkQk63wZIvehaFmkWNgxd3d2wehm1Fg4r41kucN4ftVkoie/pUWqICU5lvP0jn
MizoTscI+YkeebtOJmXMUrcRN1Z9g93Cj3R89MiOAbiZcLxOnePtTuomk05tGrpDgW+UaeYVXbbV
50NmXYC8pK1DTREH8zmpAa7EmrOqBP6GFxJPtwL656Cwdq19ewuDitgrYFrSYegjuB3vGA0VGQoY
xmlUrYyIJOAcgCl9phpsZjzmBjTm1O/NHrKu2pns7YV70TKeCplw4dUsofbwPx1DABN6Nzl/qTPW
YUQAbsDQn6x0P4vlIyX9t0Bnv0rWNoTfMncr+0gEom7VSaV4j98Dq/gwyVjfFwnYjGe1z0VKtiw8
2zuLkVKWqFKWc8UY4MH8N7l3wzJ5Dd2lA8TJdWJAOdUcZKCbXVsqI8Z+skF6OlPfcbT8B6DiRwGB
hWiwCdlXvOujnbGAA4dJHXtULJFnZlnwFq6SdaI+GXwNmuTVS89vfjM5yemxB46QjEce5IsIxphp
o3pxf7pn59nwCz30Dabp9HiBRiVXV8+lBa35FHYRiNLQNN2Je4jOEd9zxPjM2/SoZiLh0SGHlEvJ
/becfuFdNAFJG6bV8weqVqr0zcGaoP/95+D1fWpeercfwpGf7mmywkbLuaoEikZrTT4/4py4Jw7z
KVvTjFp1KsPH9zuKNx9WpnAoRAVsfkqR6qg7Oj7WK37hv+78ydmb8FWJtoewd7cUYacCCQavLXW9
ehhiqJRZ13lJPWF14K9p+/Bh9Uoz40/J39bYtjYAkEcpR/jA66j+WtC9U+QM5DXhhVphAGaIRMrz
KUFMJTHk2cwp4Qn/r7RfIaowtuh2B0zf1Kw0llrztF3hHy/6ZvWWOUamOWPXj8pd4QqeIZam8E7M
lG8W+h5w5z6sCPqfPaK8Hg1pNCnHWYQpv/p3iZvEPyfdu2FF7Pd5wQQAx+pinUEpm/RQStf+Zak9
XTVeR48ec3I2ELB8TXujbv0cStducC1kPSCu2QSu+zHApKpE1s9x7L5n0Eg202hKnEkU9JH5OCh3
HB5ZsshAtItZlvsC30yphkry6BCmXHG7HuQrU3ZZkCxXTZzidgyEAMg2DH6V83pozpK0sUWwIsXu
kJbRRJibU6nPTX3GFB1GFCDJxsc998jgyCy8eTA2tR83lSe60yGTxoWjlvfET4jSxxnE8vZ+nWDg
yh8hSoFuatRd02qCIw6sz90wAcgGqmd2TBy/NGp/jVIxR/EZEibAd1Pzhto4YazfpA3rEGA4Wo1h
N+Nj3j/eKDIubKU476Ec32NmbkolX37U9dzmF/yf8UIq9G06NrnAmGDOfLie6mBigDbkr1h0BfdC
e3VaBTeXhrlSbb97pirTyy/s8UvnPMccIWlS+K+N9gwcx9DIjX8qMeeYal2vkf1GkiY9caJF8FzC
BvgrG7H4Df432Yq6v9zkwYksfAGblhm8HLG9Zo4AszfZeixrGrK4ZtOvGUdktPpCM+q+x/SU2Jm2
roe1K+tJwIKAON2n+5MaoJ4w3wKi/M6p6mTXf0OWzv+e0kTkD5TuazDwkuWpQXkpArhGPidZsOQs
dpQZE/VcsGHfKlxttKVGqQi6j/z9HxmpMQEGkN09vQ2OjctdKfsuPOqbD67BusMyQl8vRjunBRcc
X6Ns96UPGBsYqGK4gM91NknRlJT8cJun1ZNDfhIaLLsqYMH+6gtK4D6xvpmQguA5IqcoRFPZD3Ar
ZdoieKpFKwxz6rSDRcfWiWfrHFJPqvbm63dtoy8+PUG80CFBrMOeMQKpJuFo5BnC2ShA3BAWaKGT
1KIVHk0EwmbQvd2I1gaouaWXWujZh96UUhri1X2cCh74ID2tbvt/OQaqE0xPzGSg6zAxOrGuwYXm
5UK2KndU38Eh1XU/dJBIgbxJTGigC0AMpoQaKSt+pF/bVS1qXdPyY4SktFHGOKuQxvycyOXwz+Yp
f8YhK4n7wta4DtA4rLyxoUkp1wle7hc7T1ER7aBUyUH5awmnt16dFtV5Hy9zs9KVKYQyZZDw4YqU
QVkTE4PvPNyh7UX4JIXejYwUSBBtAkPwUcm/oJLRx/JbnuC7gMhvhE9c/H/sXS3E+o+tz3yOZ0ta
FQBU50Pm0Q4B+OkWN3l7dc3GGNhT5jE/toY5Tt5ILQW/FhKDL9/pq2P7H95IQUy8gxE2vFOce4If
kwBEhM3GgEnRnj81KhIkabQDXfQydVVHLwNfAuY8+iypSuL0Qa+s9pKoIQhSonY4kzBphNQKsyB/
MNRfXb8A4ujy+WatcnckAK+P1/5ZM2Aiy/FnGhAlpUCynGB4gxeIpgFPS7YCKF5R+AagjizqnzUc
m3r/Kz9YkKLT5R1JS1DuZdn1PmLo4DcQe6lk/baxRx+NXgTQJPLOfkbCFKjvUMKcbYKPHDCtTo2h
vDNcGLHZOCfQUKAX1RnNKZfLY05PdAsnLFKhQtVFgGGGfQPWm2WCivOTFyGIjNDr95m37v/Ukr4n
3pk0UYPxa9ZW++HjZj0xKVuglUARgoXQs9JWiuQ7YxLjBazdtm7xktBkamkHuDIdi29jOX2RwJ5c
UcGBsUjpFU59hLqCf9uielOFJgOcbAu/Y3SFfKkQvUAsvOOhIb/dBux3TLbkX+wSTu0xP+3EBjon
ceHKCytqfqleitX+Ft6NsXtC2I91cweM6ojbTc6cAFts1Fq8cymfPliVFvLdmYDF+dxeoH/mLS89
zmtGRBcHvZ3OwvMvoJg+Ukvz9jqVgqs/lXBzUpPWhH1lwYtw2c2hEe1/idcMSk1XP3SqUBdJ5TyR
61YaxtX72fmQcQAI5ElZXh81XD3UugKkuG7FJvtWyWHZKKDn1H7xfLiteyAfTwqpl9/Zw8TWGLB9
0CGrKDoHxt71/2R0UN3LTbVdA3rUr6K3E/N0NMd8o/e1TkJeSgsthIjibLKFCa/n90p8ym+bmRps
XNtlBmgyHZ50rvUAx1Lwcgfnv+cIVkzqMoBaqslqlztGIylmbT07dZGGwcFP3TsVuMPZcdixqNaE
qi0gwOFJq/Ts6XvDmfjW6YmzcHKdEyf7qqdfb3R46y5D8yql7P2TzqNwakCyVugXMjyA/vbi1xDh
8tJuuuYpNi5VLZ1EwXib0E2+JIlJcZ64tZ/6JkT6kqED51jyZU4Va8P90dIVINimcgyCAvZoG240
1Vp96BWD+ivt4dDsfN1fQ6TGxh4Z8PqVZmpPrZeiePZvJ3RNSyy35GvUkvr3qs0UCzlNpp9Zbd4Q
vhBvry84iNUwVkXxspHKm6PREVomf4Apy+bH7iuLL6JJjFsDzTMEEWmv3QXsTuUSkaXYTrDv7RlD
2XppxaLoosCSdQE1KeyI4nLYkNPWnUo6JsiStBx5gu+Gk3lMXwzxRH+HGDndblMUlJOsMblM0A5s
Cuih+oEKM4XX5TxYgQOohC6XNztz36QQK2+oOdmyYPB+RRCqVZYDyUTUnhPmCgP79zXpn+w8bFPi
NFEmikK4/X8/hCPCyEGFn50prNvfWAWUqW8Hvk5SplWZN0STD7CWSzNv/N//sTCNgKHs28xGyVoW
qJ0AVHL2GYS/2GkHv7xaOxZaiLU1QnU5hHVf+JPRoTvefq7kfW/W8IyV23AlDaMJcW/uu+bvYeWq
WwMaq5SOqdlZ7EEQtxVBzBMFWUwvRynd8wY72DQ7QdAcDEFVzunRxQOXv71bnZiKiSTvgPEsB09c
SVhKCsiYJNayEl7YEqqH/p9p+SFScKEmJnFYODqu2vsK597fP7KSTc0QvaTz2PdkV/JQILcxpKAi
37pgRwID5Kuow8EgYG6oYMPPE4DKYxlsF+gXi8rPVevCqJPcCnG4EA4gqiy3yJnvM8ndapsgTgo5
zTny2YitXGFS9O/3WpbKltsMIUqW2bVJcvkMNjPkDHfolenfX7S4tIsg0MHsKo5nqNkHno35OKJk
YYzOc7/+V9DMPx9GGLFmDEjFXkDms3q+dRumDLpAyazVT7fSyNrwJGsMuoMKi8VdBdAS1Km/1G9R
HALbz9VHGX3CxP+VhgJg+qMbwVR+HmVcHLt9RENuU/qneuCapoNB7iOlQ2JiYd7w9vfNN2meYTww
7vqCezFHbQR7Dy1NF70Mb2ZYbiB22hRIdWEMdkCrpleQyhYaz4Pujva9KGE5SPXiumrLEIkUYMQ5
rl29Lv/svNKj9hnXZx7VI+HeJWF6vp8LWV1ix4QihgKyiWBB9XwelCYkUO13Wr6WBFfmnEgc0Mch
94qnYlnUkjLXxM4shgB14Qhez202a7AH2FwSSfXlf5jMspzl+hK6QyTO8EKUs1o9+ETZkJUAUmJJ
tvdKGBbSEHVrl4MYT8NEuddycgKLoBzn0Zn+9ZVkd7gletovB+k0clFHRVqyLFULILxi2/eMg1/p
F2oVzUoB8nUShvx/YizmRIwP7PRjY4p217qjcE0Z3sA4WdyvnTRYS8zKr8tKviEhq6h0T/zVzrOu
quiI93IHytmUrhXe6RZXMO+jtahEKJuSHubKMG4QKFTQPR1gx866X9k8uSHqbePj6PdqyBtXJztJ
31ng+VcIl4CvcBm9vKXwJY4NPAUeoNRIDNycwPmMNIh+Dqh15i8SaNzLSTm79EK9HpquadhIiui2
TYIUuSWQd5Ep0Dz0WSBpQ5ICmvSkWKpcOCQRfiliXZPEzDnlZSE5Gxr1i3wzAG1r/YItv/JDFdY4
aGIS5OLt7URDGPU7DGsXagLNwxRYB9Wt/d/GStue1y4cCyCfT9tG3C3QRBeGajnebuSjgND6qczs
qkL/2Ooyq9+8lNaRU9ADa/8D9Sb7tkMVWbub9TacJLwZDC+g6NczYElGFq22dwPCW3qLcY2xlxRu
NGtDTiQDiEgoynR9LzbQjslwa2BOmbx5GoePUGdTWrHMj3gOzGwV+fQYQu38fKGrvSj5vViU7Zgd
f/AG82Zwfjd+Ieg3fW7KL6SJtjbtfCKLm8VVe2JYjssy3qrR3oRCqBbBhIvOmBZyTjIt2xirlHgN
w50eoSJ+Tlihb9oRhXs0n69GdcP+EoJTmWUbxLhSo3T9TfaDiTrHMD/zTZ+bzzp143BKLAYpMoDC
TX+ILkZucfWyQrSk5EW2C9WGRQ8qr4Ufp5Vu52W+G80TSEcAvH73gvDqqUCUqEVdOL90Hfi2PahP
aKcd4B8JBZbU+ayVlRMapia0Ehsv1Y3mStjWOpow5YZsL+no4MxWK9kz5tKFtPDcaC751folqc3V
onbVnj/hdr80eRcXT8SiJ0pV37hDtUOOi378x4igS5XP+AEmYaZLa5B6JVeSVSakMQiAebPrBTZi
fzyvxBFpna4jGUxWZspK9qNqAZUNwWQyJPrZB7cqYWJsHcySims6PB+vQfqQjRg3h77PfUT4LAsF
FwZ41752DZ9WjTsgUISwiZmoD7XuLQjtuusb5KELFPbDZy0ZWSx9aKIqL8sKuyGMOM3OSbHoUvvx
ccY8FW2vTgBsbh8Ta4wdgyXa7CgOuIvIVoyJRW+3U3xkQJqLwtC1o9zsx/Syh+RzGSdjhDFIFwiy
/mKdJ2bRnn2LBvjsjXKunjkpbdvK8ItuAACUZzaapPwkwZ1Sj+2rdBq8pN/+LS/B0lf8sramAI7f
AaX0qcrV23qQx1rmJLbzX8Qnerq/dRF73mTbH7HRWV8jjpGvnq/B0Suie1pOEHq9kq5KdeYdp7JY
NJOXiT9sL8p8VjpJ5njlPLnd8BA9AKMZc3a1qVL+D7lbtVI7+sS7TONImbHQDsI2YajGALbNK9fZ
QWPrQSABTc37YMof3tqMl/gMSuaCrXoGgIdgj6s/nSnHVMCPKK0FJCGnp1ceS0GcTThwsv/9GfnR
uQAQQus4WMMBHzxDwJs+nLnylQB4za7U6O0PuaVCXSJMl8f2PX4NlPYAXigizukh980wTQt9Oib5
/5PFTPefGSLthHw463QzM6hLG7c3vxZ67o5R+KNNKSQGkSZKB6w9y5SE/FGajDIVtkvZYAWsGiw2
Hg8/SWNAWxQlFubv5PBrFWfFHtWOgLE0pVTrIDl8thVAC4JQxFKjglivaL5tj4aeN3GFFi4vQkI4
js8z4+WeISZZ9cEInOOh8FGBJylk18grCYLJIbPetZTRT2wbUlE/GvRK9/3iWpNFNMdCG3RQpbxB
TTcFMlLow7r71I/7H+HP163ht1OWEpOLBPE0V8IM8x2UwG6UaajlKptymsGKDgoG1G+VGTtKFygv
mjlAEfHYsOadS8joOXAjyOyhHecxX/rDyR7Evv38MJz/jbrW4KOZG2T1GIPsRzdourma0nIq+Xn2
H90dErE9OO6pxwHCZaSdJHAfBEqIQsDXhQWCslLEZGoxdKm9jTNz/0J4QpqghMO8eeD1vrzetTyA
jFjtKTynKnfTePOIjToTay/0lR2WYdJ9WEsCcXfskzeI1ruITFwwu64BugVcUlBmctUNJjvTS89L
uZnewAO6+P4msroW/VfoX+6r0508xQt46sOaDNsWkF3m5ph2U+2fDeLrYifQoZ1/h1VQSDE+IKmb
x+PhgpFMpNT9kbCVcE/vtc9WGNXyxmmik/9Ysy00z+3iCmcAed01P6qYBaHh+2r1F4TSw1egLq1O
Q5viiDU60tN8ZHFxfaB9wLKCn8qL/vVNri5s3/XYDydYJBKiQNWRSZwBedK2zV4yZku+4nfYTqnu
zamWIfvgUA578bflTO9CFoGu7mEV22wEYdL/S9ipzJ+wX25GYt6LE+73o25mzb7tmkavIa+EJZMk
ooN5Za3qXV78DRSrTApUDad2W+GtUc8ZumLc8TOR5EiBO8zxENUUzodWc6TaX6hwakMzm9tDJMW3
MvvCh7Vj1o/JrlDSRkVGKXJLm/meN3KIw4np61/7FbwR2CxDnUKmpr5Zzn3cNbKB8A9S5wLnMcmj
hpEluT8FzTg/i9vjH3WjxsJ4rmMAT41THv2niCUkIjTsRcagx+SWJ/Vzjp3hU77OObgzL9rzbEYD
UNHGf+A4XcY1+6GbIuzKl7z9j8+QmdXGZAjh1ZJ1q0vn+rjwQCDhZKBrvbgpsKisttgiiXlG4Hyn
AoxQ3tE6CM0E2Dol1iD7u4rBZm6/nmbiailV2KMBmDBLIPOXfg4mvTeQnfndbDTH34/7UGXMJSsI
Rn3CTh1CdMGgsW2D9175doHpgyvSpezbbo+2mUblddATS1fKGCG6/PlF/AsLA8NDDoGv5KkNjOUV
IMOaincKvFkDvByCaKnYmze+QdKiC9hkMbp7Wr8palrveDgaHCN+FvTvhRdFLV+l/iFciKCBD9QK
SjovrfywcTv6UB8W8RXp8rh1U8/WVqofYO4MKL06iCccBHLzP2QjVixQiCuiNoWKZboWhJv9I/dH
HjYUMfqwNjGGKrM/3zdJVJJbOvpJ/qaPeyXHBYZpS0CYNHmPj/a733gMtBHd8RPyrX5Nfnh7Mc6a
Q4RMF2BvBt7pTJg/cx/Lw9kDcTwLhneqoYg7SdpfEIQMnL6/ksOTKmrGIMZorR+Kjxs/xgrTdf1v
G7aNakO3LiapnU/9l0x+61BJD6gLSWevG2lfaKGOphxg6wu55/GZ9ws1QEXBamM5Ib2rUql0a96R
PAJdz5id7RMxE5bXwinexzzg+n5845IZAnu7nAdchUBlcMP+vttDyrEdtNlEzrV+5jZMYkXbvHKu
6AfCZOmDblgjNfD6BZELnwryZtQVL9b66ey1b2dnlwADEdr5/LpJfW9PVjk1NgswAhaseLNXDaoA
SU9pgn7lx1TuRGnavwyTDogGdLUP6FW90wOii5aDzTO3H2/jzUI0yf+sWH1hvaC4/NMH9ej4plxp
yevxQ/9Q0ctDvoSi/q7v+jROsg5Xo3+ojS8GpxKOp2lziDQ2C1zXbY4R4myDicPAk2t/wyGqxosZ
9BZ7MF4hbgtvlwFgqoI/B4V3MeYkC01g6MrKlNHf2X3442lHKLGlhSBMMNRZrYSm5mNjXk6rYOwQ
FZtVdAhcNwXq5FqMfDdjvSN3wtlENB8jS6/IlfD6nbGwx4c2wkgBiuombNvhpKryO75yBSNcLhRD
EtZ3IlaKorh5VackClKf2SFG1x5RgTukeAWZuaD0t1lM48sdA4fygu+mVUUkXymUEO31HYyllcZm
tV4gQM5DzdfaI268SuSi7Z9wn81UOwfqZp6pVGZH+fxdKIwXOia22E4f1MwIpPxl/X89uHWa8PsU
Nprkj+XnmZpBR+JUU5KutV/dJq1WWzW7NhF2d8Q6WqzaPOPYFw1fxJxHAwclR/jqVcV4y25INTBy
r2+80JDMhfJCeq4xgFMNrbJ2HFVlYbgsAJ2rEv/djDH3tnDa3qAbCOHvWgaHevdjwJjrzBO1xQdv
BEnn+aPGQVKXfblVXy2ITaH3nl6aHJ4ILBxB77H108wY/+BHIYge5tyUpeHgXphZoAs0Iw08GUxP
S828oO+DHuebnruvGrgsVEKORniJ6If8oC6BjPW28Div4IgkyGzvE0hM3yXBJ/Gsdq+TxfBQxNIw
m0y8Jfg8PR9jej6YWvmnyrOBBkXI4CwW3As5I2aWv/e99GIJgKg+WP8XULnR9EVZi/kxmEZJRNYX
HQ7EUQo+gku0pEENWhpkO4JYrrrUzbH8rI5AzZjfroJHUibb1/PP4kTNx7AAM2RKA4pCxel72yP3
9QiV0leFqofgat8hYTiya7EQdkW7X47dpcXygIsWysFT5FDVNguq0JI2L40YtrI2ovCFJ58dULrl
fETPdh/OyB44CGUQqFFrmCKkqdTQ5Y9tBC5YaBaFrDftOdgsOye/0Dq99imJCAoTMVHDPEPeUqau
TgPEMF/tI6y5CAybSMmcEBC1ZwppbjDXHict8eZ+sn9Jj2Jj00Yh2L11ypWlJFOZ/r3DE09k/zq1
aOp49jUQXLuC6rwwKxDeHvjB8gO/eUvlXrdzxFM13q5q2xDN9mIKi0QChfmfU4V6cylgDDVIALUv
N1OsqgZylNeFzL6+gS6KiBkaHeCZ75dMYviZESZ3Wy+ykIWzOOISQbaCABaoubjTk7a3+yuwMDh5
q1AU4oKPHOhmd53S5mg9G2mE5h/MUyKETvNmbDE6RDPRhBi7P1SLOqnHZApboIYAlIClSDNV6tXc
sJwHc+vSalON2TeIIGiDuzmRiaXfTzquAEdGZy4zap7v3EDUidz6A+DRpkY/UMGUAAUz+zlzVCkX
wOFca0hQPW5YNXrIYIJ9e530hV2gpa9QVxDIXxhDZC6uPtZF8aTdv6O4QhZ5DKoEAMcJ9+6W+Urh
xOW8C+F1UEU4uaLQU+VOZVl7jpSBQbRz+kjhGiIP7ijQTrTv5Uo2bu0FZKtToOAFC1L0CE0gUMYi
lxg9GDjUBIYrp8z8Tx8C1dHjcv+UX7f+2iFsIOpKUAqt42+PBnqiCCu+Ujz1ZRXbRh6g9xFKQ5SD
cT7z2VSFfMFPvPqHDClTHRQnPc1yG9FeDPYXSQU5I3CtG1pOvbbYGFzZbVgjzas620wevsVFxm4V
TP87g7hGAXopGTd9Q6dV8etf6BWf+51Ih4o5rm4ZNNya6TSzS5A2eLSoWNPMlO3pObTuYo8OpNom
C5NopYOdgOLl5wByz6C5b9QrUtCu6uLZphAsd2vH3GYLXFBO+Na2K62YfGshT5qv8slTjHYqOdr4
Z5Y/bMIf++X1gquJXbv7sH+WdFKZ5YwOGu7MucT8fCqmyBgSLVxc8Ky0JVGMBRD1qmXGdIUnMBHT
uapjbyA0stiPy7BGc/1HKNT5SSYLse3DXvTXYNDi8pxmCuatC+N4A41bI+qmIBGEs+PN3yGvCcHy
BT10FBMf3j8TEhvpX2WpPqfqQtZu/NfqQzKRo9y1xkRToSVRfJ4h+YfK+V5d51NL1PskU6ktztNT
ITmQIIa1TWdDBFAyO2PK2tfBfh5Tk8ugbyfmI4xV3t4wLiDEcoieL3grjcxZv8F7Cjq9JACeOMug
73F8jHurrhpy4E0PkNW7a8qtuumCa2YhYpQ3skCbtKSrjWUNlK0yjKo6MDTTC8IiJgYKXvAcMI6W
oej9lfvfu3KQVGG8PMzDYkgn4pcJlUq756DdTsywFiFt7sTFclHiA02Zk914ZufpiFn7JBwOiuHU
ZfVJJVeLfVDRqJ72WNvLC/n7jmZFJ/8KPtSHOvjSi2JbGL+1ImXcmlmySk1/1Sxk8WRklekrr6WD
YcOIBcUMhBDhh1zxWiBWWUZwK/zQDUBYu+3I2QpidM5VUzKUFgSnk/l1nGCbAMWZR7PmqR5ad2yI
wLmcOs8pYA5LJwMjw4m4WDZcn+QrdwP4NlntZB3wPUGLa41JSM7qzBy1DnL7rF1iVZX0qUu6bzSX
XtaamJNIcarCNTYSXCo72LXA5uZxs1MCyMb5/adKPAqJocmEoW+MOljZD56yP4XdNaGnN2Y3Ydq7
X8HxnpSAd1za1fyiy5eNh2R/MEN2PHSOC2g+OmWQqBBc/LmbcXVnq5tmvdW0aTAFyqkTrhasFeKp
wr07362kDYkQ1sWgsvyPPP5TVLrPob/jcMlSDimLpU/vX7pk7IU8ll8h69CDvnmyB2q/BA29jn2p
I2Qaxrlen5R7kgdYsK0lBwbqoWqK40dv+G//Ma5hSyHwyvHU2qsKv0JheTGZYKDdZWW6Iv56acMY
+uHb3OI1CL3vR6kza4Oubg9WXmmvt6r7Wjw5lArViyalZDPAz9ywf6Aaa50j+WJblsvt4it1hSbd
AtFjeoyop+ad+wRKD8pINGXJ5b1sxFlfyElK1fBwnSL56JkdfeN2p6ChITozAiwxs741DLOe+dnN
MNZwWLcd1Pr2iUzB9thEeLmHstXDa7qcP0y2JCxoM5hGgHmrcGkR6a0iAMkGzToApibi11LoLzxk
tkNk6op6azSIDNvtJ8JWkm6rq8e7hxDoj4Hm8l1nggo8exZudGC6/PgfWL7u1c4EWBVLAvYbZfaA
M2/2BU2dol43YK3BoUdBUQNSV1isNQRFBjLI/k8mOLh/nVHkQpWswej+6PzWKOhmM8m9qrhXtzV9
UvfUInz/vZgnC0I3l07Wp0vNJwarb1Y6Mlez95FtaftuCp+QMRcnVvkehDPmg5j4TDxP0zZjxVwC
W8HISP9Th55q+qq/5Do5e0FhVgRiS9NP8x1qZfZCp3oRbt2mhyhkBMm9hirqLpvNZf+S14dkQVyo
NGvXshT3YVn2ljBeMqnaiY4pFXmLI3poNcwvZbx8MhbWMkMQA2pae2GUrUZNYeicdNX22Rq3OAzc
/dxUBMhJIJlTrEbTBESKn2Kmf19WxxaTKh10BIYsYS9Yy+wPLQm/WOqQUfvIDTP6HT8JlvwVPsCJ
y0A/biAPasZCVeGG/NKuzE5RFMqJ43IvzQ+3//wX1SwrIOEK1y1QZTVHO2IfLgBzO0Mec2/rLSq8
tCEuQAccfvyDpb1bo7l+SvKiCa5l+7slTeOugZCEs3YCeu2wRK+BFpknriHnL1Scbei/4g3g7+SS
VSPDfxeS3ym0bWmVaB9JM5B5aKjCrEjSao2JUfrHKnYwwv3fSsdehwMPz08hDBnP2/8/rvFv2N7F
AYTny/m15iP9EaXggZIAeLIabesCUW14Y13biv7VMvqr610CE8L/DFcjWZKTWW1bJ/YIh6gbTc5j
Bl1t2XQLak7Pf497q2KWCdtyewcM9m/rgebnnO5iBOsEuGEPwvxwHFi4IniUfH2BRqShcvmwwYBb
PiXgzYsrQ5aJFIUxuDuB1kLwXcIJHdgo58CqK0wwJn5S+LOQ7UgrLmUmmtKERlEjNgG7jgfAsczK
xekHpf83BK7zT4NMXPC/1QjXSLlMuhIS4w8zgD2+dIo3SJ5UKqJlHUjnK1VeNSIEG8fE6X/Jx+HT
P1O3LIUZOcLx7Q6td7Hrz/zIIrOHaflN8ObgIv1jAt++Fh3SmXukt8KDO5sh+vg8doJWDHQrGb3x
dY0oG/JiuT8yRoIY72dCwYRc4xJ4amHTXDsmU+eKpojcKRUi+DC+6gyvHQS/VPkJ6s8cgKSIiy6K
3+rQeEWLMd701ez0/yirDV3IrAvB1WKUPtC+SPZqnLRMK7PtkL2YsnFgBnjlwxlq1Z3kFIan2U3E
8/bLT4CS5mqFaU5FyKCmwzIc70n1ncx285PM/xqwDOKC7N2e482kLFfjECLXc4i6vC9qg2nb0xBD
0R7rUsy/+NlLcxI0qBZqUooPexx+r7gZMi5mkYjAJhL3ApdSkDITurWldZE5S8ijJD+yQjmNlclQ
CpG4+2EeQK1/0CbSdqJ9WGynvWpwGdjemUSQwUnz67zbYi/agt+j5wIejkJ2k9ssTguY8Un3/pqx
4VY8ntvrtA3qZXL1tCqfJoKeVJrBrXue4bnagzWHvKC7Z6t+Mj2cZTEBoVh4BObJIDQfPxJgFB1b
wcAbt1KbWNF5g7XsZp50AVJuXlcdunJpvyOwsN0WDOASeePYjeLJ20/UJGekTJXnO1zjey/cRl7c
twjDjmfF/MesqQwDqiFWgNUlJknDUnm/bl4UiBvOIARi5RcDhq1bNVLs+oOiL8hvLIoEn4plkfhd
x70QuzAn153XC8GUqM9Vf07GR/W/mPfEfD6AaQ6EwSimVApZ0MkIraX0OVGV8sFsRzsQMLe6j1c4
iYdrOaWf24u9zfXfVW8TtoAod2hZnjIPMQr3LCPPPv3zulHzRGME3TknV0HG/BTvW9yuRAFN8eoS
nL+Gs1l7lyh7UJZvFgKw7yLq/dLgNnh+xvlV+eZVCkGgzQSHJ9/AL/PRyA6K4bNKvrMGOQzQwj6X
y0FyCvDiCZ0D3FiLa+wr+cYoUeERbeZKi/85SjfMuioH3HGRqu8bytaZcHEcd3oYv0r5KdiHLMal
hcJOaa7F4psQ4S7uRQVB8yKZOTVUwAHI8qIs4l2ufrBBrkXyqN5uGmCp81V2wsToGSR6g57CxTKK
l2mN5pTXrZ34g8QgDeL9zvCGvaFMi1n/yf3paGhlv9N6Ue4kvdc/zWfEgCRL+Jjfwm2eS3VIc1cE
s5T0wY7UufSGKqilAfGMm19dD+9taDOtIX4hiUN9k9oaqXdTmEaiq5970ulzLoHxx6VJ0YP7bW8T
g5LKAFbea3U1NQ02C+RtiNkdtKAN//Z40TwEFvI7m6iIjhgI8BGGdVNmA71RxcLQw0zq9NcEki3l
KiZhT/+fjfQh/2m7DaB/Br1iYttO/4tYJW/o7ze4tXXfOrTBBYGGYRojQUdv69WYHyUYUuxxFvTu
SC4HcI1UeIJ88Ze+MMBhWRvbAQJcdGnzWjaXttFgrOWbQUo+0QnllUWx07vtJL8AfKkg/haB8aal
FFKK0qDqLtcwXsVv+lXQvbPzPWfQllWegZZhCwLcPYKvDYsNRw7W2qV8NO2QBUTeOBjYLlDaR2xZ
WnldQShOsnfgg5sYauG9PTnVtpBfefb20IXj9qQTIiI=
`protect end_protected
