`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YqLs8luoVD2LOx7hLHtumeWWjLsgVYZwDzNhcuP9ppuB1zekOAbOVLgm98uBKeQo1HKdKN1Ib1d2
FfyN3T5alg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SHVUJgndtshwUv/pYQ5e5nU3PoYWTAxANZeYDXWQtEfdNrwBd3FxkD0UV37/Hq4Wqjo00SALlJ9O
bjlG3fWqCDCJXeemzliXBvXbwc5p3JEPm4Kj64TxKW1ytdbquoCvUqMRtjFC2281qE6bUPV0Yx7N
vNYO3Uriyeg1YeXRr7I=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SmIAZg4+ZL3/Q5FBXzxTp+qRw6MWAhXcZUDyiIgoJwLlzQ4jhkw8MZYroUxwmdlUWQTS4gdEjG2U
wPsf/C1w2gYUW5KmMGcsMrdIt60AmN+4/pt42er08WOnLAetspyTXiLzOUMPcEYWOctUcNkj3wJt
Dz31sxqFu6E8W5zInwFODkt98N/sBb7gr/yKmoLw8pxm4L7IXpwqbboWgn3zZhWAls8LXLjORq9E
FwrrgI1V7kH5XgCOMWDjKpi76h463pH1DIb06tIEzOMVezTKimdwjhIGqmxvF5+qFzFMnIy2HLAT
ca84by6hFJ/AfmxtjxDplAKw+XGUDfboE2GIfg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VsVagsSS80a+xvWFkXtXcXs+PiK/k5F0A55U307sLelkeGBRQjYsjXGIKCNxHLDCva16Kt1637Sp
duxxnmAIDnHPgvNDWi4rmh6C4KhlVEw3oO+GV0QA4wgNgsP2SxFSqL9OinZ5vjHkTo4QQMmMQWyW
TRmOG27NUoLnXexpmvk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I1RqihoX5DNeyTGlmTYdJDyQxTwUVKenNZKneGJgeDEfnaq9pi/V8xuyN4wP1+lb375lYNUlYpnT
eyO1JYpe5q2bKlBmQIQs5Er88JwJOp2J3wNn5oZzsIM2wXsIKwWng5xLUFxxxcTHXFlqwFT7mPbe
oQ5ZBnm+Aw/ROZMx5JTG8kjvAQeCILXiP4Kdk1GrQ7Rfg6FAHuMty00z9NpAAogmElrLeGHMbb3+
588Pbm1X5j9q8he2g4LU2Nv+gteagJAUjrxFmFUJ5e4Z0Cw/5IP1cXjBk46iOtQjqoSjyYa3w5gm
ouO6vyvoKxv69isxhAclp9J5n6YuC7S+jvamFA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25744)
`protect data_block
+IfSizmIIiHcz6llzlkv2P+SXMT+eU5tCmVG+s4w3sqA/Izm7LWO5Xp9Luqd22CuuukMfUmpQpXa
JqSiBxTxvPwWC0T8ydsswBN9wcRcHGiErJwDDyii/7dZH2xsfT0PzLJVzNpNyWxhA1eW9nwO9otG
lNC3CKL0sWcVovlUJOJCAc0BnB74c5Q/4Cl09S4A64F4WAGPxOAVigGcuHNUZk6/zJyXLf9BPMVA
+wEOk7IDWc/+L4JscLa3obmt7yI4SJ1BiIhyeqDNW0i6FLww5ygvlw49I7n8UzPGUHV/rb3+rC92
+XUi4l3DzSMC8eZkyA1hw1Ed8LZOKIWNuzQIBHlElNkjSspc4AIdXQIIRnWyK8N/hYcvvgToAASv
W0FxiyyJiR1zWVDBKWWEIqXUd3aFCFcQFlQUNK/rRMU30aNWeY4u+q7JkbfPX83XhhcIBprxbAKs
/OBLJ3wDfsnFcybWdAXg2cf1umlVTgS6Sm0NA/uq9Jh6VqVRnB5cOd6pnEGb9/pcPb6A5gZjSoDk
JOkP1VlCKddnU0RbWiAMLkqJVSuQuFWkJNO5vip4okfz1RwPm1O7+Qi25b8pApfSI47XxfG43eg8
bF9FjFDXmP5L70gS1GlztalJhWlthwd4mSxwhoi+3AmZ2GftDD8qhXSkGolX6z5tKzJRcW66A7u4
NRebdF71Le3cwMSq/h95EIwQ3UomU4UJdv9D9W8dVHEerQOUO1Bq58Sp7w1EQmc0EmE7hrHl2WCE
iLgGxFA2jVQz1g+Mai25dorkapBzhmn8mkgJi/CkOB7o5xuN9Kph8+PhPEVMmAvdXomiopR2g4Bb
bS2UWDRVBThuRED2ll3I6O+C1cfmAgPlsUN63pvwzVje2ktTc8F5TklgdrEtJKWnY1JdUJ86f3Fm
XoZooa4A2MQj7DexGMI8Ws1Zu/ay+YTzytwKmeZtD9iElwVUATz+cNsUqVNZ6ziqBMv0HkWeZJuv
/8+tPrJfd2PCHTFGLPtntV7Kb3ah/AHGdao3JaUnW0+ZAgWTh4pEA1iqm4GyVDKYfUhkINpEyG3W
h7bQJ1j9gmLwSEuwcYI4RBCcf4GBLSwxblXqJppEVtQOSrSFEbnzRQ7gRTYxvzDuxX5qoI3SPfjc
v22QT5o76hsE1EORkJExZ59SwBo6L+uTRRBucKnsChIknvgPVDyJB7l//UnVm/yd4w9Fsgks+h5t
8YpWatvt0DcIEq6Cu0iWcEGsflX9DzF91SNeHHIouWQYegBUBGKBX5iYlLcUgiaqM1ss/xOIwXyt
bVCPD6y3wG25o0mBpxnmolNwBTAi/DzzJLALQlyjD/H2DeXjFXVcsv7A/MF7edKEchVAQ5RLGAve
ikUjK9IjeVkVwXY3E+c7K88ojSEYso0XT3HFpwpO0j8iSya3FKSOKWIMU+gPPCZ/kwdqiHok+tXA
EYU2H95B05CU5JITuE3ebOKd7vkkJfGeAP6gjvtocUlkxSOLxMecTy0AjVk4kxjUIKA0B1ZfYBfe
OAGFHy3a9WwyoBK2XaWh+Q9pSbnoMVPZgZgKrYK3bBAhubKMysCGF5ZqgKkU0ohS/A2x4dh1eVac
0rvCVK0koA7o4N4aizS8ngJ4Gn9AL7aWQ4jfyNOyZxn9NCj8VZ2TlwDBO92tL/XC8rw6wOx70nOP
ci47/CYz90Br7MGlG2uZgUIbx3zKSu+HdrNgl/EgOaWGgmIdO9gqrZ2CWjo48/B2ZK2FnaB9APDG
djb1PsFVUfEEfhwze/Envr1GmbWprgUkn6fmlQNrjzZy9/BF7aoH50Vq6GQqu1tTuhYoqmHQ90sF
Yfmgea8w1aAf4j3hOpytmT3oOFyjQeDWyxbkmu0MQkGAKvNf92dDm/Kw6rimfTBEIsu5C/AQ7AcA
PiNlOEN8bibj1pdze0YzXAdoJ1GwBBcr3FsEDBe9sx2toix0a69N1LTm4hfVNjSUliZHJ66ZUi12
W8RwN9rFV9/E2mvD8mVfp7CE5mhN+AAyEWPZDq4hSER1TIXnb1XNCNo2zAriWlI6aR1Qo6tgEJy5
tH2WNKUdMw9SHcWFaJ5yMDunMXcQQcBxTa2bbAS4sDLJf3kP0EM29/CysKLHmgEfUlOA/vHjgEb7
tc0rfD0f+cVGShqzPrDtgixDDf7WX0lZPpNgq7ISdnJ07VFDQTzVwCtQj+rc3rR+CHeea29xvjxV
v/XllqbHsFaJdfKeEVbYgFzDXt1DbG1hq7uQmULuW01Q259/8AwbP/2IxLIdBqjX4lPB6QwCcFwR
mszSKFpbT7Q0wTPgjlO1oOYECB2mE57ZOCeLM5xPzNQod8+weSTWMTU51q8Q3F5vWBeOi1NATS/J
MLbgXOcuiPq8qiB6MBUZdSzqFUXEgVDsGppxDdWXAcIeOZZ4GeR40aM4mfY1hKLUA1Qw6ZoJoudV
SEDjZ0G+XA3PmH1XVNmi0znwcUokd3SQSEEQNDtXw9OD5gpJVzah2LTa6ovz3LRab9u8jHOPvXFA
oneR7SHp4YUvZORSSuX0hWgDBns+ffJnAY1yLWdVWyAnhtiewnAqSoAlctpFlLdYdhrehPDHHHhY
0cXB8kVP/O8xerVo1QgVOInmLtNnFBODy2iJpvr0L5SD/aXhY2RET1PCO+PZwCJXJq/0C98BuiME
tpqtG8bCzfxQgo1KOOYxXgWSZAC+L5fAn0itBO95OadyBghwLNziPLEGjJVF47YaoDk/raVY1s6m
ionfMa07y0Cuy4bWiTvGzJWh1Rt7HkyjQ4v5X0U5yMD6629xFqzjKJw80qun6/hekY9DiUll5TXJ
D7UnOS1HAn3F5Y9xEbTzRqefB3XYwYpJbA+bQwEDAbSIyXy/APUWlqE2ulsQLMi3ks2VlEEw8b7U
Su+EKmj0zC3yme6Y6hB9VZICdjVznP/N7chROWXWLECzaCZtBMzKfuqJUEor3NU9d4rXmoEj+ijP
SOvJFjjBhKGfSMXQgj3yVviSHiawldnWTFZPCeo3ZxE2YQwKWWJCMDNOel3pO8gpFWkn5YS3zLdK
AmPAYSaQYmpr80Gry0gVBiKgwmk7dbUDJU6HRO0K+6SsWEiG91y6Bd7ZRegdoTd8AM6x4mXRBOi3
gCfAnEN3SM+yXpo1LRCESPSpz/HEYC53Y7EwybSe2Cj1TyLs6e58EACij4kCqGRVLn+8toXXzJoq
okgcVeYR4pW28UrnjNu6WCZrVXz/1sEDufaX5ZysRxN8ehgqryXr0dKux91ibjCzgmP7ZGajjYS0
dDnakPx8jomlrWptf14fPfoD2pMtiezCeVgm31MYt716Dr0t+F5UZYPW3OfHnXZGkps7LIMHRQJO
ZvoUIQF8ca8S7/6BVhj19hfetQV0DXSH008fRBA22Rw9/ZIM86Ra4em/OAWv0oNc4kYUyjS7+0t6
WObx5rLsJKmaN51XskVxt0DghJj+M0Kzi5FB0vivC7T/GpOy2UJIylwwfnD0L3IgrD0sd7vHOHjm
5kO+/L5/kFEXViogF4QypoQn7B81sdumZSjW1Vv1FVu4XGQIaw2JLciQkUqtfINPicNH18mhUx5y
jjKPCLm3EQ+AS+az4OUryE4vYsi8R0YoJ6cSaBz+YeKL9h5S1sdZPKZJ8lEjJ3mO5PO28bjwoCbR
NoNCkkNUXGn5tghPNxKaQs0jHcYgajVGfSOcTGRe3oZQr2OjJcowbJMfI0SEDunMbhCNgSZPlFrO
qQ6+o61zxhVMWjgZuPWJOiUjK1Ju/z+FAzDRwj1/nG0BRx7Y4e084lLTRR86UaBN3n2X00XoRJbd
mBp6QCkhSdd9W1+W+4b26Oiqo/Gjwy3TrVRhLCWSZx+EGNXjro2yjd9gZQ4tAfNzTFoVW6Lszb/x
6A1G7nN2w6Urzg5cPOHgQsB4J9SJYrU30e39svjf6uGyo8cuPrQKU7gkjaClD6DZcUWniNUDblQk
Tw7K1408SxEZ8G2zdwuzx5683xPn6IoaBPc+zTcrpcFyFlLW7PUYcGyCjBgUaYKsSUYwEgHB0xTJ
UEQyNGgH/SMetiTw8itHJkheIEZ0HDYiXGk5cVHEVqreQ614IGT1Cp++CmZHDYj+6Jd+Xt1l+HiJ
Ia/pTPcbhaEcNWR8PqyL2EbEzLST9RESB9974q/RYUXCrRlsddgOCkwwWZOJGEEg7umzZialYi+Q
WBqXeDjwQwPxNfr/cRUCqu6QZyA8miU62Fpss5QWKpn15FHQdL2SDybRDCrq7/6zgQqioX7rYZpj
hp/pW81ByifNf6yCeBHRU/MQ4gNA7cQVZmekt/rPb/DDTU9iyiWkECIfJ9buBEJEejqcdNgCp6Ws
lQkMZPyCyKmo6WauK/vxfpFC2PHfiwMgf5yuUR2ydoCTglEWL3u1CyF3QmLJt2b+7VIFVFsEWOLX
VGzFsEL1d0b+cTS1ufQr7qQpRcK9cUJqwa1aA2JPS0so348S8/SgzE9UflKULwQVc7ezCHNqRGwl
Uqlh9uzqCB4dtfW9m1nGjXJd7LJhm89eTE3TOsvco8r72z41x19VZl1opRJgJWw9snE2ZYWp9VYw
n9OTvASVgEuRMKWas5Xt2QfYrpe+jz7/rX2PMUjvNBnaHav9aRMKcwPYKUwBWvjp78odAsIAN9JJ
qVYKjVyz93ww8rXMx8Ktusdx5dJijqSJNPBE1DHBYd6OalAi7tsD/So8sGJ7Bsznm04DMbHndMFX
2Lhpcv3xRP0CF1LRfQyXtYfh1iLdxwtYs+RVZcKGUWtC2WxSdNDqMV51+pCpJIvip3iuiJVZFLM7
J1jLRKv1t1iKayRcCQ+yx/qL/99SDC77sBgzI9Y5QooMj99Cz1ZAqv65/bX6n23ZqtO79n+MbyEr
8BVNMEByZHgpWlcySzaUnOcTkt5MSVv4xbVIrf5sQNxOf4YfdKkz7bnCA7YkmOWJTLju8lGfOphU
eSD4dGCzRIZqYAOTYwZ58Ebf3G0bQ4RS68AqsQj43hfL+umqz+Hhfel6Zfc4xvNybO9bDOwH9LF3
DNgf3gBXTGR1xKUG6aBC4MzB3SjcNB7hWlBL4aPioNFNLke6Te4l/UuDwtvzD5x5BtbEEbpJLw4+
w5vLcH+GDN5l9KnuPYUS+F1iSLgJAwgPJhAwVRq4ttaDkgDJng1/jB9MRx00zcfTWKRSvc/QR4Bw
uzDeBReaGgd4WCFopb4lc8GML62chJBC14QxRNGgDBIZn9E3XmcGtI0CkjpvYdKviESzqfUCeb6/
MSXFYwbUxxnEgTMxrYQnywyMa+UIjlLMaa8JewDcOMc3m3JsgItlSbDdKC0ZRhyGpswNhelsK8Dj
qRcEAvxHmVb1mw0/ajLdUvEG2FN95tihDgAfc2L76+BYwS+BrL/XgydNlSQM9OeXqV/ZOsGSAW0q
giHsb0PlUL7oijE1PV4MRDVpCymFq8A+EaaWi4lTwKeVpXYr8hB9QUYib+e4qMXHLerNVtU08X4o
SHBlXzkinjM6Ux7bNyWdAwmyOUoeEmZEMW5iOMJQXiGQNwPLh/ujcBXUNljspFBxpAtltxUvtYFc
4e2PDyLnTf2z4De3qU+h6xoiXo2uWhujh7R0AVF0tbBWvkqVXJgDxIgkna1SJjtgPdFEO06KdLwk
3ApsG7xaRhz0/n+fAGjrxbmCpAE1PCEJjrpm+eYpXJO7hrZuWuhfDiqWWR5BocRb7F56AcWRE/lu
/L3igmP2GCEks4IFX6GjAQP4gQJEfXUAol2QQ6nMuTq/JhY1C7eKLuxu0q7iU402liyaE/07zrdU
+v/Ik0gAnV8+ArdzJAlyjchw4BBVJMpfCIiPlzZOjh3JXRR93PdwB0NsLWtkmgHxLTxEDlBaQymp
Puxmul1qIgZzOskhy9PHvpPEAC9I/z852ouMgj95oxZYitEeIowpDT3rkb8VoYNV9Y3SGkj0X9Zc
3C/lDyeW9mUgRDSFDPlCSQV3/z4q6C1OKIsjgAkSQs1GjZ4dHEQXSOM/jR/5U6uOmMBDt4tudBXD
1wgnK4yUHlrfXt84IuksiYgsNAI0Rx46yFcGFI+e9D3noI4oZYgizNRtq9Fkg7mxCR0CY4DMo/57
hYeMn9aYe47d83uW07hbOS4IHB/PeXTSm4POsXL2SKfbBbuDPFIjPfafpyG4oL4WGwzLI+ZzhqX3
wX19uQK7lL4CeWOB9OVZjm2s3VU0Q9bWUvavlkyOrGcHfSmpA/uGSR6l5VHrKjCkdH3jNUbFqUJv
Kaw/Bnj6uAZanYhuiZSj8Jm6Bx1GUXYfXWziM9iRLs0SJl4096mv5AZQrOX6bFU0p9vbKP2+qebu
+V9wYQwtdP6Y3qFA38ukcp6+PNQjXLXy/nuWGj+bA8vlPOHzCrCGVG14n7s+H+E097IcEJ28Jwup
KaPcjMJG3+Z8fw27tDpioZXmZIgPvbMmeb34mSg9aXqzUYNr6oOGAg4kdh0rfrPTCNQId/7mEcW9
atwlLjs2dpPd0QEVGAnnpTqXic4VVAifGEo44SZS5kAfbDsVWTbQ+QlQPWqqZJczjKWDXOb0fc13
avYLSm1tfGIT72sqWyuojp2uY3a/J9CicDZnSMdVkE1INfAuIaJViMjRZQGrUtfNpZ8B4zLIPNTp
j5thGznqQoa+E7MuZLfwVWXLPaXtaj/4VLZFdqM5xIf+Gs1SbLYSkMvI22WAbjl7joqr5WTOcd7J
EpLu+cdp1xYmCQGia7o9MmP39dxben9QLNciPkcho/BFB1FvvkjeZwcpeTUUWqr69tS4wxaEUmpu
KQs4uBl8xX8Nhscbiqrq/M72sqaUUkl6FwdcIF9cMOFGhDvBIBNcWzF0d4IIbIJDR/Bv7tGbG8kM
SLz74oMHUevI8HYYZhgPQGfVsttynuyLwjDk6QPhr4Dz1lLKH5Hv/V7q1/htea4P3tq2JTexsnSA
9LljacPXzw4i8VrjjHV7+5C2C1hpyklMX+1pSSYIBPGdpLdASdvPtWa1eLEb3M3VyKHqSmU3ClSp
A0ZzquP1N7+qmb21xeEAbMZjYHQFO7A9hF6LQcnFD3iLu5I2x0T0Sm55Ft4xK7QSWjxGm/NaST9D
/nSFDLnXplG4Ll8xAeGow7gyJ3AOO57VzrVs6U/BIsTOYlD5CJXHBdx/o4lG46vDOST03dxwIYJ0
GZUXt43/6/NjOPCcT0MEumj2CHqmMRs5ATW+07IM8YF1qCRUh5+EQ3Kt7BQ6kAwU2GJdVlcIQEGc
3T2QqXbr2ZOg3JW7H2jTeoyqWxUjfKluYyhKNxlJw80N6HFaa/04tweS6Rkg3yK8X5zYc4RLdnRi
diIyWV7XGSFoU8ZGXhQRX9gkbamyQy9KVRPNdZYJMXJRB3zsicDPF+YRjUfcW8AB5WwhvZLBFXJu
Qw8CJXLjvOfDYk76Zggj2i2I7RkBusC4texIKKPBoveP/68jiRJdMHrohFWsXqzzErf2zoxoXyi9
eKKVdLk7VRuELyYs0m0BDMCT3j4oIE49zy8lCsywqNoBfE5kUuHrHoHaEOm7cYEFoKacSvCzj93E
aTsnuhnuSGnM2kKQRXLbmuZJALwUj9lGMxNHHM4XdaN9YKutCSQ0EOQi56mT+0fczGYDkneKGYe3
pSXqZjUbVOUNNimHTT+b/b/fR+n5vfGRGa/fFI9Oeo2G9drn21KRe3aNCN7MJSRGyXhFovEiCC6w
/O1lhsQSkJ8dmbMHAi01p9QxPkdR7XPaFgwHpN04RCwS+omNmrn9EGjggH0xRDF1l9DxWzOTWTOQ
ACv0jQlpsTUyetZ2i0XBXS9unDC9e++2qXLgiWEvCHsozj1OrTn6u47gCSNgX7NH3Mc0+Ykbbkkq
Xbf+ZHHLUvPihtJhk0lnKvSqXLbdxHKJ7x18X7/jhmTPhC+4O7Tul6VmsG/lspAcaZ7o3otVWiLM
nBLgFHRcBIocGLEGIjdIiSkPmq+H6I2/d/YZ1fA2DlQJi1aUdvQHLKMpHdOe2yPORh5iUnnyq+aA
DAl6D6EpVaqefhy6JvvbPFPc0ab39HbEjr6ZeuRoQibMkRudu+SsHRINw9xy/aKTvA9k8R+VyN6k
S+dlBAvy9sp2Z9zfaIDi/Vt7a8oliA75UwWrnxTVTc9p+5Dpi0ihwn90YOWNt9I4HPOPtJiiUO3L
R54GYjgQDGSQ12nQcnPDaisJe9wVSRgBtgRIG1/3F7OnMioOVAPjUD8pyXkAUUMdc6A9cSHjukPi
kUnvcRV4Lp4AAAmSZJ89R3fzBfcYpZx42xZmrfdw3dKeJM8slJe2/3TH4Ks34HE1DmMLLaD0yrMZ
7jW9vHGbKvcwPiSu3vumZYm3sJ8OW+U9XOVm05Y4vPh5eSKmlil3kDRM7zMwhLzUp646OzWKZypD
XZ6oSIrQuomHPJ2FJVRrXjqNF1TIk0C9Kg2hfyvqraMySPV1VoGii7qk73FwzCiL+pMzRIP3LRgh
2Dq6WlcJPZpyNPHNXv/n/EgWbusjTyi5p8h1EiuSrZDKTp2caAKGovz7mwerob8xP+m7z8ucaFDS
5lezLgKux5fzWlguKqJcAmZ2juMYxHTrB/3ebFGnfTOUrEIqXI7tOVW0zePYltjhz5BcvLnecNsm
TplhRsLEjifG9hEWnxQQeULr+sYFy7UaMdghi3XKBzBSl8FvfGj/mrpuCwfk410g6RKRpDQdeHYP
wrDtZZ2cpRLFQIQTEnU5+ngb6GIKcRjhcbHTQMHfjhewQJ4//VvU+wuoNtQiJ6vqAVsZk0iDqS+J
tDl/C3DNfoNqM3j0BcNCVQp+spgGKQeAok2XJakZiJYH1AgHrwoJfsV166NKYsjIinvo64ewOYLJ
9YPYf7dikf/RQIXwWNm7HAIib5EeNdby2732ZH6CxYeSbzzXwYosty0gPePdzR8/F19HByGrjmq5
8Pw8DUrnZzgfWngBxLSSVuQKcR0mh3QgjOZnNquOlGX8CjMf6DuTbD+6mAJPilwf1F6CoG5zXusr
MooY4wuGKzqkGowRnYd1avCypfEdcd+dO/FP0FjUAM1yfyoelJdpi1+Ocel01t1nqrKZBR1iwaNw
9rDh7CvpZwKeFF0mFmkX49KZDbQmOwgsOhD676deNLFjTclf8AS4E7WZEYnkQfh4a7o+3YSs68GK
rtKTjGoZoZc5nlRclnyRbIccYbslgMjReaCyet1cJR7HAxq89VSD4esjHLtHqHDo00VkDw1kgp9y
Hgx4kpaUyNQu/pWqUxlfSs08zgm67+fowpo9gmoRTjOM5qt5MuVzx3aKOu1Ei6t+JDe+bWVIILo0
6VNPOjMfWaK+Nc7radz5tjeC56eBnuJGaivft7yZ056mMtmn9+xonZEH9l9UmQxZkG96iU6RbG0q
ZbUWOBy9llLMWOeagOIa2Eb1MPjT8FTRoKU511sCnmh9pqjXwDUZbNx2UqnCYqU9FZ4YhMo8fMa7
W02SNU+1dgYRcJnQwGHysbnXlhAURzy4Co1qo1ZgIDJ6aKSMfa7JKdMXwwMZXMQatdBotHkCfj//
Ek0oAfDHI0xbuVrkRaVwF05VB0b57/m40fKhVvDVZV1DjZQoq0DqlV0vsrLjVDLm7mexcSBLgBr6
/icedv0u9sPV3IXoWJUIpjZnxKf9EUS4bVIVwu6z87ByJZV5XB1VRAW/mABSGOduvdeNEuUEdIlP
r9vMI9OFDzJ3GGrREXCUC/T7QaHU5YpIVNUPZuZ/ypXoZGEgZVc8qPXmBHFN2dm5howgIPe5JKoh
WzBxlLnAMLSxLh1N9ELcp6Mo4tmADAp69jQTy8hzLhH2b+e7VYUV+XJuSQTnR6ZNk2pyAuRpLlEJ
GANYaCaQcDGTJe4jpyirWSujJILIq+Aw/lZBmwp/zFPxT8xjAkNn7+7BX6FsBsRzoBeveZ8akivY
DVSSg6Zw8VANKa85pGUDNqexasdxqsg9d/RZAfoIoT9/CQbTHx4Gt4QzhdBaUolAJz6SsiHxv6hm
dDAslGYgb5azhLyixgH0B2FH7P+Lz3tjvw8wgeGOl8X1RQ+sRNppBKerNaKlTY7rq9SEUOn9VKPG
0qlVde6VEF633f+uK+Yn0xuKiocAA/B0eNPG+xTkSBDls5TaMYtq7uBTQi3oGYWLljy/5v9ONy2C
GdzaS2cCc+QvXvVW9bDb5Yhi6d8+pbLCdE8Jzj9UJhlbQEimy/OjlzjiJXl3Ioqw9FeJXGgCu9WG
gsPJE/B9C7aElwXPVGUxtwf/0TQnru12SqiM57DbZ0zeoxU880VvFX83pZg3Uo5ME0BA01JJYj8B
QGEeCj9W0ccOi0B/WZG0dbYRDrxo9O3RNBIMO3UD48/xy1yOM0lljzxkbjvu9RGvTw6dMAXJjSDt
ECB/tSTaG9F8vhCar3WB7chBMlv/lpC5zj1PHuAGAnnKL9jow3A3gjFQTGqBTVP06R/7bXhH4QoV
aZVyJ2vrc67lX3gJymTSXdOei/9+fnx7iSkV+dnDQQ2YyEW/YZpKChoHotjp1shU9RSowlDTrlof
PzRY2lVjlbgGwlXXfeQ6/dnwjvXcSFaXidt0RQYkn0EjIi+qsmz2BvKCl2fHAa3M1+JNKczB7Vrh
0AWX/VlWzBvpAHNsWGxje5cLibNKw6+o90I3cHFiALrC1lEqwu2h4OupW94CSV30apBGw7LnfAyz
vaIeyrsO3PlIJceZvv+uqzQ+dzrNZ4YgvkVR+1dLhJr5L6fEy/QSE/MSQjAVNo3qp8ZpyLoJUReu
iObeDQi3j6Wau9cO2nRQFgRAfmpwEqIwnVOq/9C3K10KisI6Yw00rVKXtFYBOv6kgR4IbXz71/p1
pTz9sE/Sz97S5Hv37Ow8Mbs4PaG+VtP9WTzzLkN2XY8H7wS8E5rX2+cVNvt8TpUpz6uM47S5sB+1
feG9/Yl2HIfRQvVhIMHr6JFmNUCxhC2p/LScTmF+aTZWzjxmkci6byqkB9ksKkfHVV2qqPerHLmq
u3q1zQVU3T/8LS5i1dvOzRKdEQNmD4kBrqpCAsZqdpXS16lrxu0aXBgtgNbAOS14Be/7YyvJaxLW
52MIZFfYENEX4TDAy5HehXKXg6wWVYlPNmURFPEorikWR3yfpI+xcitYln8cgyEU9NF2yBW4e4JH
l3V0vuujSJxvmm6jDEX1Ouk5mOnV8RiZgv97ftGmbUQZTWuvrjn382v8x897kn8AyTmo/j14JEf1
Bkdf+A1U3Nx5u+qZDinyC5ZCFiTISb9/V3L6/BoFd9Y9DJqP8PKt2S0I+ZK7TKHwNhDEJyOCp4bf
Ww4bMARxT4J/7kRaj6J6PsbqPqtoptQY9Aild+eovI0Ckm0ISVLBAvC3R89UlVz0jD+UR0eQrudV
ZN1IfCA5ZtTdqPmHlrvfZTUb1Xytguzc1zM4cKLWpr8oBGo/+rvuS83nnB6wnS+85vsPCCMyrTEM
Fv62ii22nJfa68IrGn8x7ZT+TpMS5QRC2UmBvTv1cRtSbFHWMKocQM7gwVByk8MFNEZn1D1BuA+Q
5zeLo5lotHsBoM7cEr0Hg1zzbZ22WJvcyMtHVApQs1SOzyhfHeMaO9jwtb8OD44MKYyY2E2MC9BF
sAjcljpc45SlRZyx1Ur6TCxDQ9vqvC0/LvEHkiohPelC+UEhCqCeMrV4Lta0IfPD3QarOsRYEEHD
bwNzWWUGLyV784hM4BgUAjKefOkADA7WRwJHX3Tm2LEponTwqa0rAUdzs70771+4JnXPIPYmGQ/g
S13qC2fVy3kMrHvJ8VLput4wkzkQzfwk6o1Ipw7C126XaaOAadqomD8kbkIy/qlOr1iBflCngp7N
F5lChmlX+yILlw4073QoWLHecwiV34u4/TXJDn3ByrqZDVOwguVch4q8Qb0AfFfZLZptdyR5Ygys
YlHR9466qG9V5zOdbrmJ1JkcbkOhaNZw40N46vW7o+/+cQSwVTRlrf4of4ISafRXWmWqGHVcCnnC
lsI/hSfPnuBRs556WpZIxiHecymrO0VyiNEZV+KeWbzNUKEHgtELVk3HYLQb2aSC/iIY7IHaTmhf
tMPjXM4gAwUuBi3Ql9aoDpHuculi9/0Dvk7qa9cXuTGx41MnvjnaaUlfuCgsSIDSSVM1AZTd4fEc
2ol+/4dr0e1WgUUJPiN4mqRarp8YHKLHvYNDeaer/1d/JtKmowyOUu1p2vv0RKqU/NmlVXVIani2
MQLM1C0DlkZqJdou+KgJLjrEY2XWkWY4TzuW2IzhlsFP28LU07cCkB93KYhvyRVuVHVU7cZiEwII
iSYGQWP+Ef6xlUTM7Do5mTivXO5HnlGeYm4PFJl+N4M42TCA49pi5cQOQ8CixlJT9/agBja8Aa+P
Dh9uFKKmSZoT7EnCK+qCxzEGGkIo9gifcpB2vtRJOJTfiFFh/fOL/DMkjgefREtdtTmTk9W4KJAp
/eQQ2Oa+5/PENa4XS8hfiXsDk1pDnBPWCdKH4VK/S24/pwGuQfoPHSBqNy41TOB5SaLo4+nX5gcF
wNdLbCM+/j2tx+Vk2ZZAXtgYKtr2xeudh9OSl4s6ZBXIvdKlATO0YGnOKnofNPMwS9XXAIEHumjB
pBqKbsgc4XLWLN6lZ9gjn/6PT4bdCwC9S9vLuFXaUOQlSSwhTTFThg2T9ecQHgKIfWsQvub1O6zB
KWRnjp8ZlEaEw8MMFWuUoabV4phoKLagmqpvNMfNKYn151CgBXxH0Co4AWrz2oLErYFfi8PiVjRo
GnltgkPBLS7x6cLVEpQywAxcgyrQxfaNe0qpSAhitGHwTzKYCs/7qMPAMDENltncUxHF6KzeeiEP
RukRPKNl+qOUQV3sMdCIWHZy6I7hJ/q5XuQPWRQNlx19iEH8oMMkU3XnNxub6UVzofdLQC3WxQ0Q
GYO58ulrKXT2FgKHXxM0sjeTRDA2NjqOO3LmhV5/xg+LLuJ35anS3gnoraR/Uyx+yMu8W2kr7TzW
+gE/JNP2IOitwVqT/CaaVG32cDWpHN2pUwWfh0FtQ3o4rdlk4KHo8bxsdIchv+4ArZbqt+GjPTnQ
B85T8sNppXKH8QLiBV8fewyWpP5jUS53pLEN/gwyueMhyGExvZrrJau4XzkDA3gZ3gzilpLB9CNL
UQCycVOYlPGLg8oZGENyt78pXzZg1ITObsvR37tDrEKVnftUavUzaxsRoL8v6fR9f3rsbSPfVhwF
ITwMMa3AY2tDIc5KFFg+wVvNCz08emPPcUqScEQKx38+8Gvzf4SWRIZHm+RToGCZHZoLUNOxZOaU
h5katMA8Skv4FipNckUupgJa2LiT6ULZ8stlGGlmXMTu2YuzN+D0dxgZYEcepBK921YJgMqO/BgS
nC6mpJGCm8hzJqLzx38qBGOa9XufPqu3QS9EeWObKTDxUNyyHkTOMZUqkhy+u5nY8IbCcILEUk8v
1nhEMCNuQrwIX4QNO3N6iw8dGMC3+6XBQQfP7BVsbw0NEA5HT3mR4pR99vLUxkj81gnAi6jnVCPg
TrkEzlVeuJLoHA+rrFjWzxlU51nwb4rcIeK1Z9NkJtbdpXPyPEOq9dCrwF3573ZfIAdDn7ulVzG+
1WNQpAxTgeNpzTGsXx9QY3KLSsWjLK08aFFsIi8j/pG9XPIhG9Hb0FuETlDQuRIcarxdh6EZhabW
pfyBOBDdWC3Ea0YMeMqsm9O5+fil+s+rHda/XJk8L4OxjHc0XG/m0rohW7xO+MB2sD7ROzYYbYmm
eMuyN6z+O3c1ICuRjGVeAZkV+Wszi+z2H1HKFf/4C1LUaGEaqU3HBYtQKVRBJgRa2ZVVl6fgPnVq
wBOUg/Isi2QAh2heRaLknN1jESxk26ikvCPVnnUBgu4NjYCUUQzQ0zbqGfU2150KconMrRzzLIoL
z6lQOJaYyHg47w7k/xkxhUUKFLhGus5h2mL/7/L4483HeCqe+ur9q/wxKAt2+mzmmfiU3vkd6au1
vGavmfFiYKp4n4PnhS80O3zVBYwQ1o4yjYrF+05SjmCfMkQBP+dhYJ1cTe7qBzIZIBhwylCb/9V2
c3zamPRDGtWf0bbK3iezPAitSX33aiRkwOZ4SZQ7jJocX/mxAHjmjctk1wr5QUxifsopNdPRtPtw
4xEr6zSrxLAngJYL0ixIuOpgbG8UpzpEltiJfXkQEK+kxTvVAdZ0bea2yVOXeb+icOmbcjkZ70fn
viDF4nhL6j284hbfdDNT0pQ4RNf9JLraHUVMc+PJvMJDyXVuLHIZ9Aerc8krCh+Vo2DbcSEZ8YH7
TGzafXy2Mi/fmbUBr5atDnMrQRRlkgm+qMPiqQ/QXj1aPCiXX04WADBom+5m0r8Bn6m3MDleF3Qc
/hcSBAlDQnaN+g+mZojYy2379yagWhmp+FN4VTcPxiQm5DWIfh9OxHxz2Gj3HUOsc0F2rCQU51l/
7QnQa9fK1tpITTg4sGR5lp5utvvey3kRU/Rqu+0JApcyE4NwmOPvYlfUOy5FvVWO+GE6Nch5gXmG
KseFbyPXq6OAyfG6A1AcejosjRty7efyzr0amuRnbyIEOCvl8KvaBK8xKtc34iOSrsrKNnZgzcbf
FmiqQX/l1I4kE4Gr5z8vO2ZiI/6O0cG0jKN3+FpreCdATvS9xCcOjAmWrAwMajWAm//4BVDCTFLB
peCpIePFvc7YxHse70fk3GJ+BCP3F//ziXdWhHy2v3/sh890Xcl9K/wAvSDkYwtv4X7+oUIuiXTV
lxTuJe5GROeDrqJk/RPYXFulDjC5sog4UgayijrBNMlESzaf1N3La3DSK4DgFqr8HjXOVdGRcoDV
FX8YcG73IrUFZRi2smWtPXwYbFNTXCf/5L/pnS3oy46LjZ74koH6+VQRnXGGDprjOJVoQGBzDUSB
UMx6ycaQN0rnfaNFiJllEjbH9ncHxirDttChT8kck2Bp3x+MT+ZjdlBofY/3CYNaDVTlITNiHELW
UKkpr/v0zFFYWEFbbto5fwLXFTxxaEoZ8Buqh4AuTZbGmDNcb66XoLnhatG0VEYGzkVwC3R2uYn+
0laGKNb3VhJSZ24tkx4hsT6kMmEHUJFY1arNko32+3EPHxwE9bY28W4bb8Os+z/LO1ISCPS4+RNu
yzDf+ca+JikfUcgf9MbqGGodbnjGNe5CUswQX5o7cGZbb0Wqyvl+0J9jcSDg1Aj1lwZ19VpmPIWk
17AKIX3OBbk2TuRIss0JjkT6/SFQJqMGifQaPuNVUH9wst5RcTNqtBq2/HMIU24O0x5YqeO0FPIN
QudTURtVOtcsBzooGE+/sK2JISEFXhrqi0d7Wegbn7/BKngtO+Oy8YZ8347miZ77qvvrfVq9xJlS
2zp2dqG+U5iC1sHeFqJFYtB9DeR+/QEmRJkFSFYF5HYTT5Dip1+4D7JgDmqEBFFBYR2VnYfeKZPu
1qXkK7KMaI1urwnH2cK8OKY/hr4DdgbQT/bM8ppMqLxtRF3YmYHyBeX6bgEcwd67CgxrOBDOZQBb
VdW647653IiK+IGYxkpnpiMWrjtkK2ydYZpzRpXyJVGfmqxmmxBy006Kvk8yPgGZH4hV2zXh0jcX
DzU592tFocYMz5w579UPKodTVJCtJtyziM/ZEPSPC6yGnl4tsaXBghypiT0VBrkWSfWsMjNhwZwM
5cJiQmhwqShPlVXptM3GVD9iyKNhAPG/y74iQArZZxmRAVKWvyswwk7uXC26KQHAoU6eBnVeKilJ
3DsATJZtfqpBbO9bh9jUcRKeO7A5KRjwd/K7+9OyQwQonolViqiRfaD5Dd9JAMA7GfSG+djPepK6
pvqwsU0W74eIUXjXcKL7Pp/3QL7+pofKm+3S9kmxGrfUBixJ3zd4fF88sUfJSAiL6WW6tzCxM5ko
Q1fN8bIXAwblCcaPCwQCI7knh1/ySYS5KhrF29iJaNF+LGbsVeHVEXVhd5AmnJMMFV6szEykc4Cr
gP3X+0FrputMj4Qr9JL5GMeSf/W0JouS88rlHqfoMeP8sxA+Nibv3YegfIIl7dXzn+M12/XdfEjY
jrQDDk6IHUB9OiUDfhJ6M0gFFtO1xIe1XzJuDyDQs0j9xmaGPeUQKMqCm2wIL5JGG0nrT4+diefY
DNu3HSIZKe9FxuL9A8PoEi0OEpqUe4RHowf+TC5XAqGf525/bx9sxClI4BpcLxBzR86eGi2EuRPa
Jol/nBFYS2xalw5iV2eufhoV09sQvUHTwaHgzgmmjmTJXC8BUDDbR3HHboGFB/SIQQW3JRq+KXzU
YrkOFCFwroXIyE3xPgH0gDaZBcDlTTDKkVI5WxDMR7EyExiSjQ69rg14tRGnJ5VKT1QG7V3XwC9x
TTIxC7rXvfAqaXFly9LU2b6X7C7g/vk3A6SSJ/CdgL4BwoM3H6mtpBxoV8oQXZRUOuk5hTLJN0kX
fTHA7wKx3Mz2Yd9Szr/h4tGGOTEyUid5RleAD+kfy49oQDjbWkKL7aT+0AdPkf+r+bgy68huUzgL
J0zzaSyF2SoZbINf6uuJ8zdtKlrtSy0osDLqc9Qyt1iDziG9+2AJNrsMxd+pJDrMHQJoyxwBP9Jc
kr6xo6noW1ZoQP1a6tjZyoD+SFZIsZvUcNym/E4kAHTZuGmJhiAUy7MV6hOhmRddLYb3T3m4VwRE
VYnbV0dm5ehHVF+A82QUkjMNpWBfoOUYf952H8BZItAYwUXRJjcOttAP0hdqXF2ddYmM5t2oTeG0
bVJxlU0vXnSkB5ybbNCf+1ahiFRHU8vT6g3MHGafphHdlTo7WDglKAVYsCuq2/WoY77NBhxmSz0r
VE8IonMBbBvV33z4ie9fqmyJcwnG2hKJBwZURtMMJZPRVyL6MNIQZjOWLqia1yc1fgTg/OwoMNtq
A4Vry/mwdTYs19PEgDJsrIDTSh5nN0Ws6TvEIv8tWt8oTXhQ5yXbzyfysGqF6YH5Nb+WF+KNRd1U
V4DYhgllV1svZIBLD3tKqqi5MOWJrHRwayEny99pHDjxu9Y5ltVWsgIsa31tpsnvSYE84A4oYErs
RGZ6a3BIqJ3zaig1Dhxn8GuKNb4rZMi9+vgiFqPH1/wU8EdRp4VKtflJpMly/8PvvUwJNdOvQp1w
X/9jd0sG82yXXuxfEMqOFIpT2YdoVGXuHwwEtVNzSMjJIcvsPJW0Cs6Sp6mw1Pc0+J16wnVNY3ci
yUp2rb4gZZRwmNW2OHEjIK9sD21VTKySSiUsXDUqsQYky0aonPQNpveIuDz965qVvIWVb2Vz/KWl
B7Y5/uLJqFwCs4RSUbw/HEWjYkum0v0RDqnCTvEztAtfv3Xtc3A34D+tSY8YhV2d96nFvIAOUf9i
wvdSlktEUTvOf3ZBSVQXRc7Vxz1DVlS6lGhGGrIX16lFJ6jqakWJ50MoscWgny19Ubefyjoe68fr
qkiE+V4jM+9FfCwFyKL7MwJkjYiJuib5W6P0+HafitCkYczpRmfqxLU4koVGnrvie7kcohr5qwlJ
PY/f9o9R15d8nffOOgSWHsUcFyjeFGKIEljiwPjTk1p12lQJEoDG/6IG7cw1zXTmZVeNcMUPOGhv
xuv5zcdAPpNMnH2hRWORdUQwsKmQtsPRixeoyYRyAJlHkIxIGPWhm9L+D+pC2K9Af5QVcV4Nh2Gw
d84UCvdUXa/dJ4SdqAlnEspi3PZk6PgUBEIi5hXm2r5Up673PXi0wdznYhvWrZNRfQI/YLFUg4KT
JolinzZNKe4/lVvUNeZ9E1/88di9qln+njWq6g2upO28LMLn3eb3kYbGuWY6BQmowTUsdCavVP1F
oX+dHSZY42ESOUJtOcrcV/55ors3y7ftdLzrjwqto194kYaAUmbOCByC816OOLDdH3KFXmmiFM47
gKdJS7vQMZ4zN+4knlfLY8b2WqH1e5vJia7bI0uhDsUtNn7tUWFnmkdTzSkikz90hZUZpO12r2j7
GfOIWqvidziDGgtzNEgn/EpdcnF6MvheLsS9KSNr+gJj6fbHNp+n9KJdfatM4BO3YGnQvYGwLyfc
UNn9sCYk/KS1pdUzKKzZD0ORrsfuGfKjMhunD4O45TTtfkMjL63ZknMHOCdoMoR7zhnp/kFe3hEv
/KMk5+6cwZclTgcCDoFPXycg/RiORbfuQJ+HjdVr5jL5TikOl6/eBLGCrTzzRw+yNm17S8kjzx22
5xcJu1ZMvyiHuJJEcaP4f5p1MidXsSGfBT7VK/9MlF0Qoh/RH5q6fEdYitGegUxFmS92x+e5WNzQ
0QcPUCiaw7WUFivYzgOYVNtiCeTV5p8NIwTnUEW0piHxVWqAgIG+lTH06TS1XKvzrOtsHIY4bFpn
4iW/Drogrmd+uZvJPI0PgwXryDMbL2ZUeD1AHPL/eS6KkpUKXwn7369VveRNJOQeUsJPVfFCr79V
6agZnF9WeVknh8Q/2pwDHtiPPRQ1xd6A2LV/oXZTOUqZZhBaPkmye/9hRmYb1zCDkESFvL9QDbgZ
RMgBYNBc85CIdKR1Bw0nVtFBuf40XO3Vju/SElNTGTYFpNwnsf5BYue3AgRduL4lSx6ltjVccrkI
O2bLmDKq+RH4bT84ZYSQSCfQKmGDCbGfgGC63j/TjixXuzHL8LyBPVUn6Cfz6G8niyv2TXmpO2Ta
RvUd3I6PE4rJ0j4Mb/88DlgO4/nUMauvJ3a4p93qgWI6NvXa9NCROJSrZEuEIZL9mDG8k1npBv5B
0ploKv3GS0XJfmIjJ2cO1iBdsBzVe9UuRm/f0hwv6D+eAD9YDCJUQykEc/2RvigB48GP7oAIpCzA
iA5IKEZFYA9ESpV3m0cUfqoNoQ5rzpbE80J2kanoURi9HJkcGnGRd7MpBk7T/0A5netUp2jQE6Cw
jzHcz6w0BdXkh2adlwwLaA7dMK2/7JvypFGwz6JmFzE/7fqQ9NsCZXSsQG7fcaIWhDzC0sZf9ZWC
8qqrGCzxGQQ0rR+nK3Y9S/3F0RX7o4GyctI75plH/L07BJ29xCp4kHm+OJ1BaoCe5PwuUE48H/Ww
R/F9xvG3vtJ2z49SZu+LPVGxE1ZcvdTLvyPmkZJZeQ/GNmSfWhSwN87Fft+sOmZfhfXSJgBm9TKi
XNIKVTYSVhVSObJb0rkmAIfEmVeIA+3ZtVohwk/ijdWde/o5b0tXcozpH0Isu7u4sB2S/E+RkpYa
sOaerE1lEEh9dZue2vxIGJSj3p4R78mITeKm9K+mYGTlq1zp2kyiiRaXw3o1joBH8TEg+cXdmVTV
1ZrwNvE4XDvhFRrkSqvIPhpZpNT5z9B4CpNq1Bo698RDZVTMVoBlkYbSWbJIBydcD5M6OSWz1oHN
8SzF45aFbUy8VQhSk7He8r6mpQXcsQwoelHisR+LrwAuUEqBZCaXZrJH5/Yz5JUsC4Gch3CGHUBa
CqMgG7vMHgsN+LiUPZ+lNivRpt+jbApsxXKz+RLFWuOiPEVTGHvZ9E0PNUmPK8yBlTELrs8KNG0i
NDfWinsfrgBIRNYkj6T19fyt/KZ5jYGwH7Koi0Q/mVPlJnLsUiOF05OIJAMXS1D+BFAOJ+dLvXUQ
P/JKATqMwC5bi9WB6YlUVRs24AIwlrsTSvf3kUIIRN4bV2PJCrGIBXJDYGujbSOAf5L4+WWU0/aa
Vj9hbHPxo/FmomAIxbtwJ87uwHl9z8JP90EjlAs3IYEW5+Xf8Iu9b8yNy8o5L9ctfRb3p3QWAJ2Q
O49h/vuUy06qHipk2djMQI4dU/w31p+cH/deMt0Ku+fgfCZeIwws4MnyMnwktr9C+XvfAgVwCeiD
nPlbl2XPokD7kUa5PlbJRhEm2HQYMcqJ4SkTgVCbGOcOnWvPIh3wtTnkpGlc+lSifO8RCXXNrcip
LkMssqtZEdiRRtd/bSLoNhDr2YllYAL6JCZuZ81DxxNbNWtZ1gWUeoPFoFMwUrbBjAAXeSwpEXX9
3dsV4JacN0Bd6ItQkiDzTsA4C/yS1qJ7+qNdIC404W7KaB3ZfEam2WNCJ7iKLzprOlH4TLfK189G
lGrjj8ifEEgI6uBBl7QissIPUztfopVcaLf5GlxK8wAdS0uqe2LeUBrXHVuewJr/X1R0sJpYQ/2r
tUJeDxWIu2idF6+7J+UnzD1EA/fT18iZff9dmwQ9S8buheFjxHwm7abibTTb4r5XoUUZiesC6t5P
nfZ66hm81md2061UCaMFP2vgLRDMU99rVNEgZCdYsy5tCLCBtipc9gDnyTtnBqW7Fmiz99kqeWBw
qHzJAjAa4K1PLnIUDNdyH68TyQ+fZmwP2UOFI05x7OU9t3cB4WCfxgygIb3JBtDVXsug+TlSo7Ne
xb33wPkosuZebIrvuvBBgvDHCWsJDTgNqUnTfoXR8Ia+8JzU7nm3JWEfjFVUbDvQpXrSu4l1jBqk
j3fNKF2jWYExil+6EvYBD8g+ku3Hq0hmWQ9X971IYNQFWUFT2YgMQcwTliW41KSsn/HxAcSCT3pX
CdRdPlna7xzKJoRUc/uoWD74daaEmL/Wf345hoq06MCEYP67birfhKnxpK2q2KucyqMW4BoIduaB
vez4LR4HPddGslTc8rhkhE/sFFJygVAJKIjh8SMvQZevj3kXEEvbo6Pu/lV5H5U4EDr9J28fvykZ
AKJYYpgtzBxjLxilsfiLLfjRAAE7NxlTx2CixVmLXv8yxBr15nPnt8ysOUm8shbnmRSzUgBvbDe3
35eCuJnKXTc8+9c2KiJlg3Az+aIzpBKm9EpHn42Hsznb2HYJ8FSPM5HLGfaoNWmnNINB+2e4OEpS
tHufkJN7cGnEJRvoOnc6sXfU/HemNSDZ6ujXfg2VI+jpQevXUwp/2h8Avsl3998ewI8xsXU9S7/o
M39dJTs2MluFRFvHq0fRT49fOCyh4w0gLc5lvFiR/36W4rW7Unpp6WpwF8xtlAzxh7XD5Fv6hdil
0Vzc/sdlHewfxnZYnh8C/ylgQjInEbJfiQWGUnwVyDu2pgv2wyD6O9hEpGtttNJrX2OzeYoL+V+P
s0x65kRQgQh2rJvyzgRe51SrX77MvtgBoMxAXrXGr5OS7V1wJBWhCSjSJ8YbtwVaxXGDYwXscQGy
mPiUAVQUyopTN9lD4TIYnWrXw3wIN8EDlFZ7WaEIdiPdG3yyv4s8cIbPRD3bxq3sh3EJNY2xinj4
29AdXa33dKpv9j4erXsTHu2VgdPyT/3rAHbkQPRbeusMtVrM1v4Qepr7VuJVhjerJMw56nDkXkeC
KwZoqDT7tJhPH+dCqilo47kx+354A4/pc164rujuDgPxyYKFVKY5qt7CYqH57lckwW6Fi+k5bn6a
EmO7PmhMWauKC+GOcfzgcZxBdkIgojsWYmWyKraQyYihIqhm94RT1pUQ+jTnRbd6XCmEItMcQ3E3
9Ifq2vUrACvfr0E41YSExxKxdmlf7zDEkeC918WqLooWHsNXM/P/AbJ6ILKYNrP5AouACOCLImyH
F3VquuSvn9jnmI2Y1/DBctdPxeMaqjMoRZ+sItc6xOS+LT+fAsprvsZ4A2GckFIi372ad7WuPyjT
qjdGNnheggd4I9lWT1538B1Wu8Sr9CMPtDjT6hs6rNjHeYKMnq9R//mv4evDNZjRVTKL22+XIpUT
wUMlzotRHYmr5JGl2BI9EdYJJ4s6l5SxB/HBUNmP7UvKKFzADh7rWpS3bTNCSB9AtvFasfzemXI6
oWLr6qfeFwGUPcfaBhjAfP5qTlNxK7z6LBlP15sDNiZ4F30/CLAcEeSNOHz5FuArc2vSAVlEp8ct
uDe3OEnFaYKJ6dBVQ4ZekEbU73xFPpau0XJdZAs2WWqfLG7X4tQUoIhkm4zmF8hqkUUEISWON+Oj
L5nQUvySG7y1UOLOlEELRLE1G4+9Jxrn5kbvPER55VivHpKWWmjlC1ohTiagbEbQCyZUryvsYJrb
WP+LNj6Ais1e2tKWYAwEiIT2GLicjS5mCpQG6BUnNKjJZVn3QiuN+1u9ouGGEgwzWAWDwveufjag
tSVq7Rf716m0AEDsJfpXYdDOIH4VzZSPH+t2MiQCyKZ5qAf4D0VO1BdtJcNunjd1xf59slhdA8Wq
8/OZzy7PZajGR6QldTQiq2afY+ykWcXTHhFcn5TS5lbMLoaNk/KIdcTUEhfE+R7ABAa0/3cMJN3Q
1s6i541Ym80b0m9AuiVChCCA+BfALdfCQct4fxYwdhfJ3LyjjT8H9RBUwHlDVzBdGTowQsIRDkhR
k2/Fd1dALc+R/A2UYL51KEiIYhB3vgRAw4WMQL+09EL0XvkiNE7OeUQqmDQODliUGPVytPi/KCCO
4zMBmPC7B28E1ep9D0A3vRmI5Ep6mdf1YpnttmCxCe4mGrUfiQxkwR9xOHRfOnrm9FHH5LI92WOJ
1CRlfk9GKLODpdfzzERxQ1HfZcrm2Pnub35uJesMR0TLY20U6eQ862iC/qaTfQsMKWQAzRDuHMat
DohvwPIgioDW/RUOMkBUsoAaVHJu9hJgM1NMBPHPCt1mJ96tIrXbD76zdlEio/+B8jU8Jx4q6ryK
5/H9DSGxtYJ8l61tgGNF7gJq94XJubzXhsrbljq105jcp4ktcqNawtCu8aDTW2ACwBFVe5s+kFsD
7YocjhGmBi6iERTGOvdH0vZKThloDkC3J+QAf0DOGUt21xr+IScJElBTFrkg9CmwntI7+Nns6hEA
T2EyImTCMEHwPeSbytn1EmFrfbbMwDnxEI/3N/QpQiilkNZ0IAi6d3TKYxxAmmeGXbKbgGUvblpZ
cfFMg63RSm+rcLBfbuxkRAhQRcrwmCXXm3k23Egs3Q/xJExJ9UnAdpjHJk4IjASIEo4eHsjtHO7h
afY5Z8+ClPFupHrzU/0Ju3Sk7QNLjE1A7J5zCTFCSBk6qw+fbwh+8ePu7w/J53HECJ7mppjDU8ri
uAwPXfrX4jqx7B++1u5CW8JYfBkEW9ct5x76rEqJ6VFvTq7Vup0i4BC/jX4Dsf9tbMkZx/JgPlGm
2Xl0mAT2J6cYAAgJ6NwSJsx7E2NpuF3tZ4yjq5pEh1j5psyLyD4kxbo/5QxSY9NYF8qfE5X2nGTR
QYZjVQhsrVEzF/ztDbPkpPhUrhCbWPIYqYlwBBAL1MMvc4/u/a05Mi4O1pziLvjRLhnrRQo4kfnw
SdzFhrEcXrJM/dTYxvcYcELpOySybN0+m1rDs2nx8FpsrqJ+/Qo/bIZwcViROvwaohN7SYOkhIKd
1EgCtvvAqSOKdu2U0yriUSe3OHyHbLt5F17Xim1V6YJ36YSsXuWgkNy2HyRAI9BYpdB394oD5WTS
mG6OOWC6WOHeHgSJI+kUVf8CeKhBRVTcPTpgyN5SCdg2livD7IX4UiVnl5hUnsDKJ83k3yp3Bbvd
/aohddeL6jbs7mEeHpOi43jDdzNKvyYL2NegQG2sy7pgZv4p1VCeBK5k4TuOQnCRdhgvClVcIoI8
NnvXGRK6NUB49MRu2u1WjfsXx0aAGGnqOqiHGOBlLkR+dM4kjxLwpEXygpImIkOX0BFSpERQGF7c
6WpCr+1T3HheIGUWtPVCodA2y9Pph4pI0s0ICT4CrwcPGtbRzPNRYOmDisitRp5P4FWm69r7wc7o
MLKZJUAV9YBwTCvhq/5AaOkQvAZM9hoLk/4fmgHt7KoEs1t7HF0TTh5AAg5lvXpStbx2MrX7+4RO
2FHap73PNLQRE4FJ2cB1JbA+Ja3PU4pFcovPBeahjm+sBB4uHFaUNY++WfObEVGrFzvrfh8xYCyC
hSVHHmBHXfv3+Jdfe6p+aVUmkg6v4bgOTjuj6JJZUWVveJw4+qSbv92d8lX5mpWoYlnyXiwLefyi
rRQfSuXV0Y82mEhk5OG0OHq68uRTYdO9Fcht/4c0Nx5xpyJ/8gS1oEdeiOUikM9Y2Q8jrPsreqpi
LwKQjr6PxBErj6EgFdguF+ABb+qYDaO3yBsmS0TlWDx0s/a8BAQE8fVOVdhUGZvSx86QuzhJJWdb
e1zciVhyv4aKd5lerW1aGKYe7Ek/pP9F53dzyH8kw7X6kaIduWUuJN0DNk9VUEXUTsyax9DxmU9r
NGRaipjSjsLXj8yRl2Qu0I85OMJHoDZQlsKENpEiWBljwFB6u/lmXIzip43039PGFJhYsWakEu9z
mBmsSzqeIArqSrPcCgw7JAQAemTbSeEQW/0N22mIdkqdsCO3tTqq40M4t5M8T8TI5ZYKgPmke3Vr
StUlXhWCMqCtKJWdF0HgOKdZ2eWG7L0lCdvrc5cVwuFoq5qJ6TZL21EtXBnJmimTcai+EjtaVue/
+gPfY+J9I215ZNZtCXR53+Fe4yVbOGPds0lNY5a5+Z8g3hb24x/aEFhW+hTyQGPdIwOdF5xoNdcE
OqCm1sBSJ8p1O6mI9x592Yp90Pxu3iPPCQE22INPBOKjZSGv1nLGk1OEpFUXURV0r2y4mI1ydBbi
KRZRdbHY4ybDkYdNQjimco6D9gjyPGKdWLaAXDfJ3QkK28yx3ulupx/kdstam2Ujnrk4GfERzPlv
KOX2AtgMCiHJcduNFUqc/MqrLNz26EPNXPwDQeBtnE097JVDv2AF7tijYreSvKOoJ808wCsVCs7T
LpKQe09P7NeGaBUUNeh2moIJxqHTJty17/TfjzA6qcJApejqU5eB9moVYUqxCODR3Fk7RmbVCxnu
/v+w7BGAl0kRXdzu3fGviOYR+LkfyaSYybKpkD0peYceWLUFNI+ojH8IP2hN0ddpT7xnZXoF0ScL
mz+Wsdr0Q+cQcsYDcWR4gungWS+wYkxdwGxUljZaHMJvjxEVGnKWo5vM8MSrKWRMoQdgdoIzm41R
4cV1r91FrDmt7BWtx0iSoHohySMJufpFdAkBVzq/zjrm00PbBaNmgxlH0lDjWp0UzZTFgHI+Y29J
anHCDmC4locw0HefE3RtwE6+H1jdgyYPMI5hBA/9WwTRYgpbREd6qUyupH/TyBuStmakNhhtaUS7
dlqIktsf2bh0UwaFg/NDIHpy01XwKqgK+fs3j3gCS2l1nw3SOFfhkO8ntXeeK6dVCiE9VRt6ZKp7
UvRPrCKi4TdyFPxoI7TGj3aZrLIgTynzNWG/2W/KI9OQWXLRBN129+hkUEFiAa96tXpI/8DmHjhC
VSytrynzJ0/uzLt6tGa0KI+9oB8kjbrzhS4ZUEZswya09hq1+m/diN5RuE4XucsT8Z43kiFddnKo
PylUiQLPWiYRvmBDcGilHRMjvIitC2XbMKqMiDs5li+zCD25AtSz5JJ50NOXM5YFESRUutypDpXz
yhzjp5UoMMW4OWxcvjwpMVfPhTj6JXJuKeCtkEeA6YGDXipElM2CqOx09GBb7NDF4rB0wlOT1V/Y
6+M5sf2gcGzXVAG/SmOzMYgUmb05sT5jPpDBx7wv3aDz3KgGBVCM9lhLCOZ4x8c3pvpzwBy3K6BP
XIRdUfq6/8Vc/CwqPRzUMYvo9RoDg+f2IwVg8oOwdeh1TnbRWhxypxUMmoq0klrL4TsaHzY1C1IK
ov5mKRvLZzSVMW3F3fRl7IYS6/v9WfSULwofZWO+3QESof70nW4uNSbXsL6xtFGEsht0oNpzPfM7
mb0UnIxeL2sjB+i09A/WfJx7CukJdLOQoQj7sD60WhdUakAswUDmcNktAk+uVcdgMkL55wq6w4Ph
qKjMfVIWAvXKFWiSQ/uiLPexPVl98UxRpNAu2RHzvaO9EqhKctLkDslZni1I71sn8VFnkrYmtdUt
J0nHjCqIY4fhcsOiKkagZg3ZaNl3R59De+xrC6kxzDtphqQv+Loc9Adp5o//aKna+Y2O24M5D7px
hyvhH/CEO0yecc+Ew3UaULDtg8AISoTmunDpBgamwzxSPPvY2lSbPlo+3Hp0gZVlTSnNUzo8gkF0
UY0ayszg/W40MdG98ssr50COTw8ysOr/4eQ7FKhoG4cGM0k9tzL4/JuKk7z1lPl+nOSwnTPgNwGl
wpfIp7xX6AG8N7MPFNpBAJfEHC2OQQkoafxT0ZyQxFAh7c1OzUafReVOXqsHnWpB0Wnz2SfZ25JN
oreNQURhPa3BwFriev+5t2R7JVHSAqg99f50r8eR6hWhHc7dqUXQPWL5IullM8+MOyM927ABNwvG
twhQUWhCUfv1FeNYEVIIVEk2EsbPQNKUHGPqM0lTNx8+6r0UADlWO0xl5Kb3406fYjfY0zrrblHL
zDNPfPOPBb0++G63C3juuB0PPiKNbWXMM2swNP+BgRjHrkQXLX5br9lqTD32DLKrUM+lsmvGtXcT
2GF22YXWC2w8hx0EL+X5ZNbpeuCpZ20ZAG8cIpirdeCvJSqG/cW0aw/FEgZVfZ9E56IJ5c/RWhIV
4Lfdx1pWaXNdU8aPy+T9oCQuHJuVCTaB2CNg056srNxOWbE8+9u3vkdC8ngJ7yxMt8LNTCo1zBrQ
IrlzzgtNozoTQS4dneO7kiC0YomR1jcIibrPGLGT6wSt8grSABmtw74rchr1B+6SDJUAnu/PRkQn
Nfr6tf5gTTlxz2/m8I5C9lrPbSrFoUpXjYxVXCy3fAhd5uvjC5hMyk2YZTwgWAoXvLBOIfT8c4Vi
69bBUUhyy1nK7GTdpZViKaXvgdwX0uqItL2N75Rpbhs/VUkG84duKSNEz/H9tTsBrvW1Ww6zhvaE
CP3WoPPrjxU1D6u04ZAS1TKUz0iGujrW3pXLP5S1RwQ9rDTuWmUdNGyK3OfUFJ5s4KIoEQWUkTOV
WXewgeBWclEhAhzebmg7Gv0dAI2rPq88Zf6Lni/LdBFkPRub+kwl6XVyKj0TgS5NyMrolzBPfhVm
IxKFoqb9WPwHWAxsz7vawbyA0nUgo1gFL8XYZLHPZC0WHh0Ps9MIMJ/4Jj5elPqqJ+PYCDCEmSSr
njxjCEXPLSQZd1rb6WeG1nC0zsgR7LH7RGo/skw9nqnH+ZPEOgZLc5zM5aynNRw/ZH2uJS2Gzqw0
CzkhrskMqR7+239+90kKgtng8oYBVQGUU25ko8MRp7FI1ud3zOEBYZaKUxgXZNiW2kHO+2V0+bVh
r+6KqKSk0sZL7B3+e/bQ7WWcnN0XQSFL6ecFKpJAgiju73KZSaeTpeGCB4+IThFQ+otpEYMQuDbG
gK+UIAgQnfpz80lhtGvo06x5KT4YSrC1zef9TSVm4tJTvnwdEHAqpURin7xZ7PTfLuwXGN5RsIzR
W06PHXlM6s3fkxhk2XCmtPjl7b/VcNiORhcgnoM2dqAffFlMoOATk/SIl5Fu7sfcc+R33+pr2AaH
/f+hTGW3FKxIZWtbTEvndfaJg+h0URJ1oorJtBvijyaCc94MieTyld+78Z5zKbGJUnPXXef9RSPz
u1p0w164cheMcZk2pRLoRpnr50kGRfGywMoh2DmhvJ6oCVKhlciOxImeFfE1mX+1kALiMeMll5bB
+GTrCPQB5Gjz/OM/6WdAK+iHfiuc9zAdnFr5OTsWxBuBoMs0IRxIJ7d3aRC9o5tFVwd7G/fyCdze
JzzRWo+dRAWBuMVn3Z09a1mbCLgE6WXnbmCGUE14b/g8LBvDiyxVhSdCP3RIEchi4Pk9z0xNHTaP
rtv9zzGR9KydXP6zlsl3TnWMsDWdbhr+h6lXjikYHLB14mxLssfqEH5a2nmk70fxivRHqchKBJoT
FvnnVSOHw4bM/120AQ6X19SlgzPBZZbKOp4kthWzG2bpa/MTVwxuGfqHyz08PjshQ+SkOKW3Cbpr
37G2e4WmKFjwoyR30KtabaT9AKDskLAtq3qHM6svZplb8GGenv90g3t2Tj7LMvvm64F74FaP3lCP
kpgplvUEDHIVqcSmvSJzKDTLCeqUjidFqhDL83ncYZkEW0GceOpFe51sd+76idRFLtTjcEoVuMnj
v905D6xs/HxGBZ1klaoYeozHKXydQxDdjw86pH1aXdGFMCHrVR2vXwfhPI7vABDnzcgjxqCvIuJH
VjHdndJis+9us8w6OixkvNR9WRgdqrm7Cg0vRmRX76GwnpS09CtBgzsEwCLBKwfhd4ooMIFaFXmU
iQmkgFslTsgHxDszRHI3a42NA/UEmZ4+g/N58iT3UD2WbQYeUWDheAjr+9QxfyxxL1V8rsALk7Q5
NK/1hY55xNO+MW0vxzdd/JHKfol3iJpOKh9xqclopZW1DenYlV5a1SwAiHqjnB5rQks4HceOW94L
P79ouqwEM4Jo1Pi7x2vRLIuA1mrLMiI0MSurfss6v9eRZx+GX20aixcEi2k+tW7I320xgQf5Pq6B
csQGDguCyS4/ba8Epl6mJOutuUreBbJwpghIVOfe1T1llqf9VQU2N8SIgcweHaa46cHaZajJC6Ul
aQjrljVvGXn7+9Ay24zE2vrHYUlsMLrsOG8VHU1oeT4SickWLs9CfdzcZ7AJlckRkj+Hgmnx/bjj
x/ACpzOoclQjQ5nsI9iyXRYUV0V5hpDKeXM/u/igz/uiNtcZlAXtVsFMqmwUsdD+0JfCA2wIPQQ6
QkVyKIrj3uWo7l1KEktbB846nwlXyh+RbEI+2FdP2E3iqIQFTYyoWCZG4loJZCnd5EeAncJOx1Yb
PBrzz0CYK8a9ee+k+KfzcuBi7pCc3Q8O4OhkSLGScMr1qAFU/m/JtVsCmP3SVAFORXTihImQhhXa
Gnd41t6g9F5we8AhP36xF+ELICn9j8ctAi32+uouLKUNN/4bb1rdnf8Gr/F+XKFZ/s6ovdFxUzs/
+cS/M16+EgJzTfc/vj0j/vWUGa+TJNlG08FK+eX0gcuXpi1m+Kqvn4evdYulpg2BAoU19oA8lEZs
naqflRDXkZkh83fF1Sd19jWEhoS0lkEZ/BvqyS1IRakYWe8iOq1ae0ly52vNCqz+4rjQHPWtu/25
pxmZfL/12mw0nkk9jeMfyTCgZUYxBe3XFQW4VRyZ9qlh0k1p8VDB2P/9BvbiwdcnDDKm52dMdpfp
iGFDKptkM64VtJxM0nnyUUh+RG8SM9FCiU9XgPJ1IzhYxRmDCA9s6Dg8Mnc6mvrZJnQk/q3SAanR
4rZweIR0Fp6T4J6S+sTfPxekP/PkUZIv7SVzd+UDq6o2jB7mgUo4wLWe5vzfTfoXVB8Bzh+rPXtV
K9BExoUCoL72VDTo6AJsJkUorvkR+aWLei0be2WxeodfMGD0IT4l52zYiUe2GKGNfiFkeFBDwa2A
l+bQa0m5x0ujAJn2sHK50eQZLvSXotENNFumDNWDaePSNndLVj6ovZbJoJQHfUDiUwFolL2m0RPS
rJIZOILylOXgqoZNVzzYsOhuRyLDQcgVIyR5qzu5PHskekg+QrR3rOXIqd6g8v/Dpy5YSb5Sr1s8
18kKsGkTtO/R/5PyFyGYhNIfvGLCD+H8RXTfC443cJB2lHByDiR8mElxEj6j8JQFYJ5rfZ9fDHl9
n0qkLF8Es1JAL4j0mfriqAreNg6WvplneC3ZH5HYD8Xu97Rn7faJ5oqblNFTu7k1o0eSRUqR2wxg
mDE26PlSy3UxcAkKjY8jBZ6sPTdAs8cOZtS+MLzh3PBeFVc/gRHQ+VUMp29tOZ2HJ9j4YK6ZK5lK
gi6gqOhxsOtlrM8h7io7L6m6c0tWkzkZJWaCENR0SVHV8DoX4QGocuqvMdrZ4fqrHt7l0n+Wjqzo
twa7kBlABd9sPOuJuCYmPYxBYMEksQU5oAf66yhFM03BN+Yr44whzQGlFRhfm4o/YLN7LOyurf2b
62ib2nmEpxGI4/bLV4/Gm6ReTo/dFD/0PTflk206zoOUxeyqijiEQFyPpuJtScvmN2+6Z+DEVwh3
pOp6OMzkmI+NGM97+P7uaBAtdsEhVrESq+hIqrelpJtb3XzqWirqdyfCv3zNmbu5CIRJz8GgjZsH
KSXobtVY2tcCMiqEwmftIPVRBnXn4xqjEZHzEGkzwbctNn2wHCW293w6UQNAgC12Ilo1hY4Iz1KA
2g0qe/FXG15uFzl/RprqtTcC1TWtom1qK1Dv5Hb+Wad+Nh7GVN7MOo+MwLTEbm4PhIKt9OLwjHFY
ppdsM3dSo8/NftM2aKzuXKWETPu58YlrbINXICfpEEx2+X24oRYGKFqBw/dBVLxKPxBCk2/sLYh3
uCmRiZEOLFGdgofa7BL0m0JXsn+l2CebPj23OQcCGI0YXIAaCarfXbQoxqK7ZuXMcWBETphfHYWo
laG6XkLVyY7KDSAKCbIFRCtb+NXNrJFRqQQGI9ZquEeH3UMbOsoIa1bEYIL+iBEUDRO3BXMBIiyQ
+S2KSqLeAsxwclQE6z9wqRafObVIoS/oWEd8jRVPgWX0Gy7oNikoSP/ICV1Te27gGc1IWF/LFzTv
i0te4jXRV+ypNdINR+ANR/Ku3RHlXmUiJamVY0gWJu4MBGxK5e2a8Wr1KkJjCjIZSFuqCNckncBM
N73BZGSNOCZTvUb5FVhJXc5dD5dZkVEyDHqaJPp+85oRlnOfIxEzClOTMRgA4vFw7piOV6iMjhYi
x0RwUDhgFnV4Vdhi8yz8+Cjgg5HNTDRnWeRrhxEJkFIMF1D8v5rZ1bNKaX+PkH0PsAV8FdbX/sEA
1G0xymJnNP9UBQMtILkhNWtUuVjw6R50Bh4DmHnzskV1ymCfhtGuAUYuq8HkoFaxJUtnRFXX067j
/6CRV7xWFmJLCdoTYi01OGKP6uBDIq0P1zgOcK2wCQuoKxpgZHU+AAprXoCMSfPh/mAMV2+m4TVn
t26Vl81eLkEhHGCE7J5MK0J45CNAqFANMXtmizlDVHf88XVfOqe+YRJngWXMsYMNxv+o4goiplua
04AgpaYxD7Suv4lIIkmRuxzHv20/G66TucF6WVyNuG/2Od91Q+O5Sbbx9E+5R0EKUTFbJfQcs5r/
51K1bWWcfvbVrYWw85kdRhqY5Dy0UzJS47vM5epq7YzrQi1pB+sFss2T4KsVkm0PH8SU6ei+qauy
W/rFCyjk5yG9tXfKaKRBam9zWg1SeMRF7PrG6Ls8LeGbUmjLCO8/0L2HpmR4mXc2um2ks1MdChK9
XdJKypE/5H52Steh9e4WTfDBtN6HiqtH4NcKw4QUikUDoZ0OzsoZJAJDMeucjbJHWMch4+zKfcra
9kpqn+0qCX8CxfjaBai/wrbqIH4dz2sKQrNSBgmovbznfFbBb7XW3VfC3+ZylpkoVMeiSYNHk/OX
p/5Oj+th4RtqjZ7/qR7txpe161IufB6Q9GYCoPeSP/tUb18YvTN2zrzsKntPc1vdR9qA8MmbX5de
TeqjH9RQdIGGlpeEP5zrnbRjGoShmHZU7SeMZHjQZPjpA/FZ4MqD6s2WhxAMpYcKx8TN1naxNzkO
ql6za3U/11Y8ElXqCDOobNORNtRe7OwY3Y2XJGRwtT3kSxqUEFgPJ3CvN41MybLE9mZw0amx3Jui
sFZoWG+snyn4HZMWgzTrUwamx4Gi4lOC77ABt2sMVEdOsMzrb7Z+60V3TMx08rrZCnCvz4lDLvK0
6WSa8ghm4KClgchnp857dm2nZlfR+Er2AcNXId2Wx5lR7sVY9jm0mItuCZqrBKYC4fDDosV5/TpC
u3PWXgm0frNQTfuZ9vSmQLwdL2mtNnk7WyUOeHL0RTaoBN/+/0Hv75DuJQgfbxdXM5r0iWB90bV1
K/c5XZSoYGExIaV5HyaCCsugudPTS6UsS9wtidIk/gaVkXMvK99SPVrXJiuArI4QzH4Osh/i3xr4
1IWYKNFsvSk9cb0uvmll+3A9iHeDaRqiSXVV2H8Gw0T/UiAv7hyttZB8AqEhtM3Sgs06UllZV8ru
Yu5tg+bXZGByQR843m4Ts5bKVmR32lrrYdl98bobgCSY2rWI0PKe57B5jEtpZ1s4wOhbC0Mi6Kxv
V6kgb5wV4vYE4o8j19/X9BVvNHy254bBfUXmrCxYK3m5MMn0I2O8DckBlE8AwzZOPW963ozf7WK8
wBJZMLj2oxIwYWwBSuq86+gynsT425T7wpHd2UxUBjRXpfsH7FvEDpfo+shWwNb5dxNAoaauZVaC
VRCzXkGm4xzkKgbueRyv0/zvPWPHnfQCD74sB2VUZrxZ6r2OyCv4ptVgb14xQDXsGpY4xAL+vwPC
Bdo6hXHEx9rPqkcphD9uEeOiQDFW3qjWc8pQxg11oayDv/HKXKCyBj7lX+GQ3fDU5F4VVIab+YKK
E1iY58zxXSExR8HTiHRtBbu24obqM2kiJNmfns7gzQuBztm1bmvm98bdk41axttj+gcfJpCoRwbu
WQb7qTuRaQDR5XXPI0O/V4ThzF0Fg0X1MzUAWc989U6jkt8mqJN1s8K8sEHZJsbFS4fV4L1GOAMY
5zhG99o01IPQxpB1vD6fIyDu5q4LNOYJsJuBioqtocDmZvt2/2a3gN+u2k+85ljZnwZtun2UFnqW
IWTlnmyPP75Cr825YdUf1Vi1UdAdk4MHo/yVEHlbKV5T1b00K3ToGsVP8F0J00ZtoNalGhs+cgCY
3e3mrXPf8b9dbqPEvob5z85hbLvmOsabhOjLlq6dwxX/yBUGyxaRGG1HAVtSLgtgtrHTbmWrd5M4
T+fUz5mRSNkdmnvlZHPc5s9MdKrxQegZ/bwg1NRq2qFDrsp7l8cmdWrIOGkAZJM7mFFFra0ToHyA
1K0J7mIFafjk80XTXflBU51KISgNMb1aPi//gSRjI41d1Bs8CM30D9qP9EKt7Vprs+G5PcfN2Nds
WfXnJpckUn/GKcB6gdy5FNHjEFDlZ+KuLxcVmWjYZos3J4Su+ZKAWzC/qCGIgw5pFv0b3uWVVlRq
Muo0DIqlbrhh9mOji76tqqOTNncWG+onx5heoHtvbkwECvM7KVL/frdyrbnAHgOfgu7PNbW5pqKz
SUKn/eYRk+2giwOWG1PS7IGOdEgGHLY5vttUB0bc3q0sMGnhQ3bYHg8ztGvozo5rCXUjWVkl4yPu
Ff+LqmD4L9cc6h+YWDe67fVF693B8lmKXgrQE9OYUMSx0oo2L4w7KMEu9dOL9ghiYWKVLondkF2V
C4dCcwPgUTwMUOJMB9cPbtwhwIFqHyBrYVOcUK7aiq5kdCJLHbCkBDLPD8yJZijQCOhodC0f38OR
YgvrsbqnFs6IhmUrWlMKVr2VD924+SxvnCcLXHK3lY25+Llpd9OWEA/nBgX75T4Aq1UZeFBW+lOM
iauXsktR2DOIDS/TQMy9l1S9lqvSJvhZQLlL00DVOTz7hSeizVQbIV2gsruH6+PSxsGJBHvTlwpq
jBoC4VMLZFLW7g3WHiH+QgkbyLU0GMqd8ppk8bDulk+cGyALWwstnEXrRe6WHxJlhiL43L7lC/5v
zKo6sWsoPzXfu2P1tntj4Fp+2OXSC+jMjDHmZcDJbRu8uxVvOxbKp3G2MNfjEhBsv0RjNue3Nqdo
zE+ijVGu8nRKxrC5aW8SYZgK9LPPVujeQ56dHHcdfYtmk55Kf/0DXnDy0Y0hHMMQL9F1iAgd2vhW
s1VlnKB0GqRrrE4Q2lUdzu42Wy9fLvdcotMVc3NLxUR8O3vApoGxacLf7pWf3h5ZwZ41mt2ntXZw
sy/4nMXLHckB6FoxsfEIKwXxqQmrMJncQ34TlOdiaagB8zYUaSo8NU6ttZsPBW2PJnWPJiJdrCsl
vWEQ7/JaKtAQB2PdLAZYUCnFdIB0ofXQbsPXNPRlssRCWcQ94ro2/m821zO9XeNufQ12PqRTvjLb
SUwT08gIBd3BUzkfkCnTTm/OLvgds+9WNvGUw8UbZMBc4cxVOhWtrD5Ieq11SfefZf/l+5BrQ+PO
f2dBp5kLCrrIffaI4JIks6sw4LfsN6F9sxGGUOUepWDnfnFQ9hzDgApcE0ySyREP8yE80zZTje1w
fYVbHXfcw22z9z9ZKvx7qwSwnGVPqRsF9E5bG2wyjNx9V31urFmADi2xSHy5rIlCDEvG4Mhy5Cbu
Ae0o2skNqCTrVNJooXzAeWBVi8fDeGyxs9+rRm6o1W3rGGofJIuAhMCdFX8jATyO4x3iQEMENScy
6KBvW70VQfCOFArpH9fLpig2l40fCc9uQO1xMmzL3jS85S9+ho07M05y8JRsmnZQJH0/VZdS+iuY
aqUGM33+hID1feDYX62LMcQH+hGQlueuTLeLyGPIzIfBejXt/rnft8d3jxlVtXIG/r/ft2lB2rUI
C363l3NKufOdhV2vfEJ2Q2N81KLZjuIh1+0B/vpcY+1WvFhncE8hqfbR2PjvWqoa1AmlPeNreHuy
On/bAmFyrKMYapNA4B5NKbf9oncMlQ3k9CwZ1/S7xpfgnFjmHTZYX+m9q3rDrF4slBcjPjE74JZA
9A+sY4IRB7/85f02/Fx7eDKhncd1AGrcddZLGDrxidkg8jN0kduSFCY2Ge+5UucMHIGtwQHm6GOf
ykMmPhWM1VNPx6m+jpEJHFcnYE0A6j9yF4X/mX04zchLR4hUTTjh2tLBbqcvGkgN0kjqtR5S9tWI
D+8p0Z2qSKL/lXtVmHbftAEDUAjjwUWSEzqNehNvmP0mg0cj2g==
`protect end_protected
