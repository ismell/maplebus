`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Oo6legxa5riKkzLaa6v9AxgXpzPdVy7DbK1zivQAeLXG1Fttpk/BC+kBkutYNQ96cArsLFGRKy+f
lNdLtBZMjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pt9l/fS86YC8+G6uB9p7TAEWsdsbsITIzUXMPvVy6c20p13HRN4q16CJNyoA9U687ujlRA5TOhoY
pXMvIkEy4wGje/UiiaUg3izpfPqKjgvoQC5w+UhMxstlRhYvyexzQRchmrOoyISI956gvAyAWBx/
1/TjlrIzRE1PkJfE+xM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FLM1Tm4wDYDKJm8855F4CZnEQkv0da+2NnEyN/Tk9Tc0Xp3e8M8G2SttTQ4RoiAFSq4X2isFlJBs
XJOtDw1AABs42dP1uM8iQgRs8qzUkNCA5eTfJeIWFaHj+vLlxRDsk3XoxHIx8HZnhgsUVMxG5Ymt
LNa4QpRVP7qp597+u3E9ZrUzjiE7HxZ7KtuKBdQvJE4/zfuoHzHZ5WuOLo/Thua6u/SFUVxqy8V0
BRo+k86EKX1wfG9JEGCgmtpGiy+yOyWVKMhhyvukQ6fBadtzuEVjNCIfdilL8BYA+bNoNqHkLPQ9
wC81L0ke0VJn6vR99a4eMOfhoysg9bEBM7dgmQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KR3So1UW4ADGWGHrH51Xe2+e4VSGYNjqCydaCP4bzcY4ysX1nL/TXaMOBvP8d+BTJGyDSfBE/Z3t
0+aMMCVli2tWAHOdswB0edNJiHfSLLfTnJ+oE0xjRXCjsA6/O+aTAVniLXss2dX7gkQ8NpJy8xXH
3Zu4JKCGhfi6N2dF0o0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TNpAUsZaknNx9bYChQaeGaGpqeKRElLovPpCA6eMwCmSisaYIjaJBebdhrKR1npSX/c4bGfTWNLm
9R9d3vPVkKF4tENTnkxqccFOxu4JG33mfheEixBwY73bw77ieJrtGE8i5RelNXZHdnz09I1N8w41
o5Qd4u8QDnUJpHcSxRk/zYGt0C11aowDcnRYIBQzXuSxVWugWBjpdbi3hPTkYGj+2Tdh9lZHAj1S
0kSSe7FglDzE0ETzsmFiLnthVr4Kbrj5KNsYWOCmIMk7bPddHlW3NC9OHVlDw2VgGwXMnTiUj39T
wkJIL1h4eMQUCbmFloYkIbUXsf+lfnCV2Ae3RQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7296)
`protect data_block
Z+xz6hsYlTlBzutzG97j/bhi+lhkon24NIfynQt/N0qU/gpcJgGZWwvbVeWpcVRgz79/Dvb335yc
pEg9xwaUNVyV5QSM7YMldHsRcZhLTiBVTKixPCSWsh3O2p5wPjyy4gUfhjErpT741zNY/PLI+OGC
O+N0YLAF2lpqhPNE+PAU3dixB/9yiJ4/TFmo69ygreRuMseQcJcnPCTwKlguYgGhSkPioKSfdr5H
6aFp/u9Lh7BCLGih31YsR28F49LXe/Rqz8lQWmMrHA6O5kRBshfUCj5G4LOf29OQb+neVD/Ovj6n
UpdvUBUfTUTR9ILrUVWNEKJcNLMffyxJWRyavzz6G51dy1tgJsRtt8ICmYmDoJrbCxiDvev/AM0q
9JDX7mlqzpcPLY8TsHam+DxWmscyFNrjyr1LpjXe3n2RcmIP9syf8MVtiAlA+ibf6aEfQkKL0les
uOtb5KjV37J2ch40SNeTR0Tvaq7sD93oPa8ma1yfKN32AkMbmEYKdAU6fcdd4cHGFyUwktltWSxD
nCI+Qc3VQDa4h9FeZIoijZ1bbQNTsabokVaHBBklJ4XWdA47luJiKBpPnpk2eecLDBaqq6WMcxzv
k5gwEnS5o4TspNcLA3d//ari5SYzSsQJxKIat+taBW6VpnDT3sr26zsNlPwFHF5+WDJK3yiYwVCZ
Q6TUWcsu8492EBOGgS62s3tGAl2DUEjgwisUZ4cMPfAuExpjmx0FKJBGqR4rCTRqbcafRO7BzG2R
EQkfTj2LoTlw0d8TAWmOiLgZ6YY0JvVKhJhFFkPhIlIdIvUWx/6/Rxq4ISj8PTnJqFDiQkcimU+2
oQ0kK5lCNWIH9IZI5Cx0JUlbNsnaBGc6xJZwF7J0uIH4rzhwIA+Athfy/M9T9Tk5ZZiMh1NDHzIo
JNWVcS+YfrlfoEp7muHptcv6pyBqynO42jAwdAMS1+kvg+69zLf6DvuamHt6rJson4oUt8W7ILU7
nX1ScCDAMAzK8CXC/dSkhIDog9uWCgohydkBgjXyoBDgtb5mCX/B10RovYGxyZh9WRdbacGzTpIo
n0Zi3AtP5IJqjNBHssAByW1sGOfQgNDt/GdJj5y2CwBVRq6DKo+TItPlMloz2p5cYzGBbYDKW4l3
0hEteVYXdtC4GMoDnnO6/ES3g/dVFg/UCOrjb7Z7OiP9hMq5Q1/lf08zHYLm/yEj/eEIosdbGYfr
jKbi+eARfN32glUdiwirqSeqGIgCoQEU0BJfcLs93V/USPli4Ffr9VeJo6/4pPL6+Gye5ou2ekcl
vU9E4hk3VjrPlK6PVL6jovpqiVqhyHv56H5yrWjB5SiNX1LSnx+QvSV7bmmlPhvOFaBBoQwvuTwP
r9End//rVPa+0S518h+xwvSv91tP3qnpyiXrZMQ7Sr24Q+Q/TJOQZuQSgzwGPr4x9PpVR5tkNNhV
B1Zzs3a1NZQZ/OlUFCZvXPn/NMNnnWLBi3oFC7S7ybdv1F8DSqtA07vlOpBr1oTbiaZqcmcRNL4O
aSCkl6P6CnKut1LNI24J0yoajb6NbrvEi8enKbKkbjela6V+edcQj/2wvWGXeveeCptWfd87WPQL
7PHCgte1Ur6ibSeJybJFYIo57NnyuaY89qBNB6lQ0QBsSca9KND8LQcNbqUJlfrsuInooMeALdZ9
C80RLFXOAc5Ozf/W2KAJpmn6pe03Z4nNs3aQLTcNOtGfMGRJ350QecXJ7e6d/+tprp1+W2ZVTN15
2rQIubDFGPgnBT5jtubRjr3Zr5ir3bee3uO2zfjIWBhInpA9x8s1VhGr+aaRdigR1n/wB3TfZYHn
SRHFWZiaL37z4yZq/2FOuCb4h0L2oTyTPr7Nbgv4rupDvswlg4spSrvawN8iIFWl9JMt4k5NcWwE
7m6vFcubpypffKt2XMQzxO4USwFyV1EIyAeL2XrAtU10nLUgYFIRx83V1fnvK/2fXxQQo9dSjnae
mYMmf9qMbbtYnDx6pKhv3iZqbNSUSisBIniznIqZrSOi98kZeW0BZcKomACYlaPOB/ZRluyq+OH9
jgjKTybEjH/aM36NRvO6KiaS+0PZKXvJgNKbvI4k7LbG0nBNt4RXS9fQFG7XpqqxnQGrCp6FeE3m
mi5KoZhGYa854VF8RCeMZgLB2pBdXttooS0GXTVe7UHvWWTYlu+6LMC+vOBbgkz/MGQns707un+K
HkBIcN3Sfsf2g3dKsMXggXCAqAWFk0RUin/FZtX406N9VcNi/LFyrTwBE64NgWt6wUhcvhcDyJ2X
gsn+BEzTvxbwlZ1jeMhxgEDhlPVJ44EXhyZTRYAvtzOnezNWiUHZCgzlKONXI0QJdpSq75uQGPGU
2hp9jLFahVIgOeMXM1/8MIapWsQL0WbIFxFwpmYfyFNWKfJMo5xQPooFMp3KIJ+t7GL5DiNdHCmi
UZpjn9sRtMVzRuYsozFyzRSsJBC6Hy+RZDFaXb8oUVZvX4NszAQ6NLWohga+rtEnP55yOy8R5JE5
X4sO7kZy2hQoJLGfuOmZxP7sPSFJUtHrsQ6iBHSeE0w+UjdHmBIKATDietZhEDDPpqv7i48hvyFu
KdmAHkTepJc46tyGHm4TWWt+gfyq2r/2R0fESenOkMjBkM8LBnNCFpoYg6EZA9M6gvqidbbP5Cmf
voAeKAtYYbtR/Uu1eRQrXByKpjASxD22tL/9IoPmHrE+UykVAdquOZg3LDosLOE7y+LtRSGNAOim
xcYE1vmXlub5VcI+fY2fdoh2kGag3yIzvdZRTejzKNTCrcC9JbHMwHBVJSgRmUVMPDOHjrUz8s+j
dUjLC8nDX2zJHPyJnujvmbQFBf32l/yRrE4qcFu0Ekq1DVdBTjEjQS0T+ux546N0OOdS4Caj6kEr
MMbXmNirSnA6T3Kolgd8Rjb/msdTIH0ZTA8dFLNO86DKhclMRGbBPS1tZqAIVzCwgHqeo9pCy+x0
xsJGbT55R9txN+O2iVwXgvmzcyLPaH7ZI8f/oAx4zjRrOGKNRzFHT1zoANdTEVMVpQlbdgH6BCh3
zpdTRhhc3u/4RToFQWNF5Yv03VszFn31mr3MtVbadqvtJlWQCXRaLquvRx7oY5rapF6Ym8vaXhRZ
qhJTYA8/hqE9869xR6BbzZA7n/2NvuwGPfSLfoYAAW8yOHTJ5YtD2PCiRup6eXhp1gTKnG+gwmtE
Gp8LDv7WOvJUZOKEs/ukCf8z8UAsW0YfVi1RaSOv+Yt1/6OG1y7XCr1qtt69yeht1JzrTUv5VcdX
MxpBihvm9rGQGkOAOX9mqmQBDQ8BFFUPOQUbT6+4GPIDp4MuOMNeannSPz90t0yKVfurg0qWq8bF
8fOeeJc8AzfIIPfH1Q4Yr/IItlOp/9S5dTcGYT3VqMjLggXOebT4Le/Cm593C/LGeDkztY6wK5yt
XNh1BAeEl210DX+2mSstqSfjoSoJ4Ip7jBLT1MGp3nm0+TvUT68AU6eSj+hDNI0tw1y1zYl5yjhr
nmInCJg1wGvnu3/rYJrOP5STZUe+xEaWFfUUjrN8kSIfj2T8IsPRbABRMmq88TX7D2ciNto1bTOZ
jRkI3Y7alB+covBmvIhYl88LRlx9kB4LEchNlm71dp+qtMkI+SZS5zV6VQt/0IsTkGGNWCKh/JRh
2NjSwFYwfDI+doBRq6EWi+9KXR0ekf9+bT+vPydmkcAyonc6kIyOqElmovif6KsUhrlnIkIBQACg
hycvLzYNRmb0O9UC85tVxlGXN1Kr4ImwoeCBz0yi8lAUNeNTQfULpFmQEH713nmP7vdbBT7w4IEA
Z/r7BtSKgWj0IXNdHrqTw0tbvuMUq+kCVz8HxJdMuq/Yu430WUBaIL9C9EJTjj+sam+TnHk7Gi5s
YWPldqr1sHmp2qJLnJpUuXfDo1EMPFvVot1uCbciMbVYk+JDFbvyyty6JvbHBpegqoDEHTJYEGq3
H4LgBPKooEbB6GItlVWiUnhPokAdmJcnLZZYeXaDPQJzqg+mZ9kPp/QY+KML2dxnEXNzfLJn3k95
DpUGGX0Mu88Cq58dZBg3Q3LJu7LXHmamb6abPn1JOiKnEmpfS7H24RCkTLtiC/R5TU91Lbw8blm8
hZpiL24fjstmwmR/fZDiWcfChyj1bPiNv7UxKc42WJG/gcOBfUREUCBJQsoiUEJnwWX4Y1ZlIcs+
zw56o7JAGg+3yRNJjnvN8TpY44q0o7bRMBMi9Y4TsjFVGOR+yPvh26magDkl1m6ft11rpSrVEBzZ
BFsVhMOGpr0ZarWFWqe2bUgL5q7Cb4DmCSQTgjefZcdreseulS30Ppe+Xo1DfLDjWMr57iivVg6Q
nDOWPLC80J0eiPyCTDEH1ZjjDLwusTt30m6wKqUxFcoLwGhDK/0FaDgxV22rcUNTvGScxDrjgbQZ
Kv71HKrU2JhN67bCkhfpwjxQ0UWd7vIKkyjVbE+aysH6TfviK5FH2rNuIZoL4eJnKXwbwQnst98N
OXlZbuB7zw0jXnoBNwL6nLVLENpAXAMVzUjQlokoyt3pXKb+mtDHmVBcIZgCHvwaSkovI4q5FbSC
nNWKtliL3xW2N4QGWQuc2cGkWqYmix5ItemroqOh4dYHPpJ/fxXOh7GPe1IlmTnLjPpwkvHUd7YX
dXk6SreVmPZ5tQrQHNSO4I7r9hhD8mBrl2noZahv8QYwGhy118XbH12Gmwj5NqsqxNaitUplV90n
hHzK30IMbQX8RcXtQfVcd0HFJYeZx8rJPGpvbOkA5zpJljyYVeeJAslQ0G2bAwxOfnOJ4CTct/ea
qkt7TisPwc9iQmrdMdQ8I9fkVxwPC/qNqoTNQXB80tSMfZlpCW9WJ60trIu0O+eXzLCuiabohkn+
WAHNJJMus/Sbrab38YAkixdPaLlXTuLDJcfhtqIRUovtpVpkiXrUN4T1jestuywYhLfMtkuyMZzR
tgsSCT9GhaW19c3nwDK9dBAGZFMGcycaWdwmhpxzRom+vSxYEfpKH5hawvluHoYsX3EGcFlaMi+0
L7YmV04BcG6GWf9qEgG2jIJbNeh1RTSThe/57qSlutXPXWieWYXE7WCexs+S+UrbnXcuA4JJauSk
mX832fb1wz7vJTHBbdqBHqEThvNgdgmfRQ1IZWlN08nZUaQs2jGa+wu5ANVap//3iGoinnQeYuSw
2RUDBjhh1zZlxbKr1x6X/eYy1uvZJy/2UBjzTbfxyX1fOiMvd4RV+aPhBB3fA5vJc3iw9Sfp1odU
IlJ6WjRJQkqWaTVYHyPviv4uDD1mEWEeh/3BWT5dMJujEnB0JIEMZ5Z0yiGMTQmsaHXV92s5Q5ft
ELSSdkjBYSZp+5foEr0wFBrvJFg+0cFdYfDe779uBB28R5hvwrUGLe7E3pFzmKfB30/wx5GSYjpO
ZfvYJDzAgV37nfHA9evvQo1cWlQPeNq50t868sZkFNRPVAi5YjqsJauuoqTIgqwaX3fhbHciGq7u
+CuUvHFOjKRlTRXb2hKt2SRYXJhLjQqaCCwPFfRlpr1LvNpOtNKoPFssBzuJV+yqmmcstTH0LMw8
oB7hYnNMD7bTWMHj0e4iYPVmUwjhJxWJvpyVc/PHPY142NfGbLgNxe/EGpCBhuWmC1WscraQsvd9
45qE7NCpZxQY+6VUOigX47bZZJtVy6zDMwkUHOaBuLI6DsKeSqsmRj2C5jzeYQXQ15jtV+4LC8vR
OBpWnjxx3gUuqJiWIUNxzUM7FGljvVJS7PZiZJKgjc7RSj5ygdKOTLvALdRL3wXl1oistH0tigFZ
uPBtdKqzMv2q8nk7b4ksQU4ThIL4lYjTdlGOUCUoBfnGL7G8L2YNS/azvcyhEwXQm3EspbL/lO51
N5BbNOarCegEizao5/EfHK9OGRXtPo8d41RnuC5+ygXdTfyGEGh8MIIjpMRVWXhRh87+wvOxnCle
q6ZctARiGzB7/0xwE2TsPNay0ZiI8f3YJ1HBEg7pieKHOAOQfIFBJiDZqaasBuIxGMVE4W6abShw
13CbQzcw1kuQrlWY+4SQznZpa+WZMY+95HN7I+xWWEsisqfxTFLhM+kwhpnCZJ1srB9eRIikGCJW
ropb5Rc+ewSl+5OwTGyG29b9+MmqSY90lzHYDIM7T4nLWRIkvidKCxfyEdwdnkq1nuZeg2ObqaFu
/qi8Vor+pfcW7369LgqazSJdalGxGm3UK5xIW2ygyr2RAcfZUwHfSvpzl62S0FrkAmLW7dEdZqSG
vQTG+wD+DnbSjw7KnnFpAg57D+iujArRbOLk1lJCgiPiz+EAE0Vd7kyfEgmS0AZsNXdGCbdIV4i1
FywOW4PEEyicJ5BmBeEpO9oKmtsjpEkuXGAHs0rQiH2cgQqSDmBerHTb86ApSuMlicWUEPDyG7Wq
ORP0J4+uEG/hy8Dr/rj+f3Lp2Dyc2klzxOwQjbk61nVWUgfE9tsJSUm4bz5ycZm67tbNqWdkIEt4
NXtJD7xGVEJEdobvXKuLbqy/kIEHv+f0+m4bFfIpFLQvFTZ5fOOcV9T1U43DBqzCpL1xJzJPwTiZ
O3uVQ6zKe2vy8L1zIQ7RYFC7zSAsYt/aM85/ohK+kpMy3ekjrULshXf7qogh25EqlmzyrOYrBv4G
10aGzqGEZfexXPUOm7SUzhMnh/oIy2qau6x1GU0inaS9IQgAPivBE73Tt7SMjq6ahUWzJA+6MKDE
s/9dMy/L/NdgQtY2dDN7nR95WBTUI9ibgCMdgoDqGFYgcr82An9R6LlrgmJJKd7lWZDMAjjO8Ol6
uUF03TLciNwPAQP9PU5bmKRH3/FVawzoi985dtMnsMEwuhkT5PGz/uDEQIy/8K9wM9Yu0cG5Wjqk
EWy66xGBdEnw/wspz2+Lx2B4RclAJq32SGT4gtjjVlVIwHo9PsYFEUoGzrlPrV3jTbHlwNCRDNE8
ZhYsWfA5q4EDfB8FZcBBbbEvQnLFZunkCc+j9KtmdCPb9d9uIm3KPd4xKZYPmMywV5wttwCjJ4HN
EkcDCxohB/k5ZPoD8fXSpUu7ktMlyqchhlYr/DkRQtZ6M6vN7WBu0JjyqLeaAPKk+KF2/isO4Xfx
JV58sxeK+L0OnSM2A3RcxGS8UkhjK1JTzt0FXT+IvHSeyHkYz2kgTVKwL4MBkISSy1N283+g+Kuz
6O/FG/7tpUPKiJ+ZFwEdwQq2x/baYyieQ/FobnfvXSsI2pvauSqRuNrzr8rzglAuMmH3IqFcDhl5
9HDrujeNj5SXYP+m7j3hWfPlSEK5TiGv0PmBBXGMNaY8rZ+8UhW38Cso0c/nQjhRNa/W6sTHnESK
8So6LpdMtr+V9VE4Mjn0Ogd6LPZkvEpp8FOs6uZggudCmPy/YqBmayPklRfRAKlgekOE+do6qNSm
yVWjCxUOAArYrPMiOsFOafFo93cH2NonHRgpcjCS2pvvmnLDnTmU8Fzc6dejAHRUtp1GIkyr+Fu+
X5jl03PnSWCBtCPLO1UI+TLXHcj4cUSCsC56TNyQ43VOQDdEP7sSl2hIvKD8aIM1NYrpLtZC9eNG
vwK0/6x9OnIXhqIIR20QQ0+o98Y4xU+f4a/FwQVQ0qg8H8H1QV0bkN+pI629oAlqkE8NDoYu7P0w
xYwpMIwPt5Jcq8vzRUVM656ea5ZqlZqqeOY264Zv7XBbUilkPcTaHhtjGwCil3lITJyTyhH7xMGr
WCE3D5gPbtIEA2zDLotv3cdq11owqvUPWB4XNcF1UrBOtZUtW+KG8nOW7aKbaRbmFQdKI5VZzAAB
wpngfcPYxmF120rsZ9cPY6rRFzjh/uaE5ScJNI//HN81FojufvUpPeOfYT7P8dfGc0DKfE0cCg0W
wL0EsrJ2oGxs+V6r2VmOfFyLjfSgH1u9Ejlkd7+0zhacgdjkm2gnMyeV8Jm9/wdmrpp/2RGiInqh
C6JfKazgJuPN4h/IQr+9qkIb+kxFW00dwsMJzsuyMCUJHPjnSxA0I7OA8BU1hwZQM9DLzLujAU+L
p0p0bvb/lQykk/2aoVzUPdsxEnRqP2FImWQXGbNHmnl5iqiccOMLd0LUI4xcyJRyQRhc3figNZGZ
oMs7aG7n1kYRh1N8Hv5H4FaSPN11tRjt5+hpDbiK3J93RWLyxW8EUQHohVKSc44g4DSRu675G2iW
r5jhl0B2j1/rsHGyDc+3IBzpK9VXR8YOzWmXuSGy7fv6sfOxpiMLwPiKV27Sc9fVRzOSb9xj+mcS
7DwLbfQ10k9S1YOP9N58p7XlHBhwisB1KE7QE3LWzRHbLRaNynS3pqoZLyItF0bylamEp4eXxUyU
auT2/GlLrzMrikuIhn2uajMM3kpLp5eAzQT45kTHWERwVJrdltAfledelGj30qNbpcMuchR2fN+G
MfvQF3T8hbm00Uu8tJaSnQbd/40DIcEMrPHJ58RqwDq+0a9HD/5ipEcRZ0Fs58GBRjEZWwOP8yQb
NAiXmoTYc/IG3Mb1tjk2RZZk4zhFZgp5q7o1rWE78Cjwj7hUbhIfAZuk+rMg71Nn1brQzWGvwLTb
gCatssXfsEVnkhz4fa92e/OP9ti7K6RzaUnBrG9ZIRVbKW9AN0QNrvMmsns/LqoMZA4XixZUZGtD
LFkBv31zXosXXzL3vuPp60hb9r2a9AIxbbYbFosehaCG6MKMUepmuGZsS5E/HIgY89hEpwX9gtl7
2DK/iK7mhfqzvn/TNZ06vUvF+CgYSRCft8psRKceTCH98aISyyByFPT+UMGqmcF3RtWNt/ufl2my
IT4uBoRo+vpBuMGnE/IX5YgG2aZCLnmvZi9pT6QbWJHZj7AMSOu0PzaJDRKx/i0LD02cDaPagim5
ef3wKQJhLuaSSuLrw5ecuYn1448qYcAaDZlKGitfBF+4DEMk/ijyugWVX3u6hz6sdcVy2TXDKIcO
VksWVJS3AHbcZgXzRf6+39KZ3JedwDBTRytysJs3Lz7cXyKDqsh8xe69Pb34c9tPnoZ/NyRxCTI8
szhyi0njqacJUEEIHmrj7w8jPhcGWbaVMY7oFf53S8saQlkYkykD4sQpF0ekY5SwtnuKyH10Qmre
ZqSq0FtWw26BZOiOEG7X1/xx1NWNie4s0SqCxlwW9K5JLvFBFMWR0daU6aopK6FPcz9Bkm1Rb1OQ
p45y+MIZm5x5vW30gKqRXGsU7oDhC2X8dYISzKux77aQuU74p6n/Wz9bBbVgHElj+uBGE9iykaAU
qt99biq8wtXoSzvkvXKg81QZG36za7y4fqNDBBFbGuhNvktnt4mBr9sYo/ZaRVLLkXjTOgl921eZ
050NBRw5J0PccEHFbM1qdt7YSetsCVBDNHzMYQ0uIlucm/Hb9/oUhxu7aT9CNXb1Qgg0jURYtH28
N/xNvmteu0vy0bsjMfY8F/oYoBoeETO472yiK9Eo9oc0S5Kg40vuJzmDaMj2Q6zbj9cFg459tBzz
zkUQsD6UeHxmXUO30Ok3v50mtoSYFaCV3rFIpbeYPAxVHtogJLK0IZQpemPo8LqmdC2RpGozU60K
WD0nyTt+twS2XnbEBKengPcAteTPFPl3wHiDo0Khvi36FqN2Q6XCJ7xwpZmTebAP39znWRLbnvrH
4SckVatSoTytMbrqDmgb8O4mp8Uty5yr4MfH8It3XfrPKFKTL7Es6xMmeBkjQNiJsGfltlE/kPr4
VEfBUIQA+6nymEBmbtLHMuaL26dQYtf9cte+jmYJeWRDqf2ptn2o/m+WvRY/LFK4ZeplqE3+Rnm7
`protect end_protected
