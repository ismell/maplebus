`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j988rQGPJkSc3p//+LZwMCu3Wy2jaN5CprVWWNza1QWYGjKyfmaXOFjwEt/qwbjuzHbjjAfjGbw6
Tql7AHe/og==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j2uDSRzUbf/Lv3j4SMAzi4tR9lklbNWs5SLm2h3shtrZo60pOO2klDsHaE5bKeyJ6bUnYWcnHoHZ
FCxbv2P4AP3MdSC/np1f+WsjY64QkepPYJwjmJsmBY5lgcjdRkYUfgCYW4e1yOpog/eI+krhAT3U
Z9oy4o2E/NIU5n/cW1w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eksap/1cFJeLg4uPEMslnAPBTHpLZq1N8tuPwR/Hcf838RQ2Sx/f5Hb7ZWTJUpMd55t45TKqiupC
KIjq2EIDO7qRI6rygjFDjUDidh8QtXdfBTa/SPQ/tS/P9R/tMb3v8eiiwti34bQN4gtExHd7SjuQ
u6xXMrNLbI/fqTssUaDunpYLPgACrPKIKpfMTc0H5WnAgi29xvwoUNvUV6NIBO9pRj5BSBpf3KjU
BM7eE9xKo4/XsY9t900HT3ZxttDYJDvGTN0BB4MX2AdlfGRKwCEn7LJ3GsVFa+EN3m/m+aDZAL1l
WF+MxJdqGEVMTFJrgwCJG6iTFRUhTLsGVMIMMA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UIjIqhUqlKP93ALs3sqYQNb4DqeDY0JMxPMrnLsjpprLA9IggvJuqLiuHT8RD366ieAgCIQ2Ooxr
h3wIIuw/rp9Isrpqag4fDBcX/QOuJ+T6N36CUjG6m7zngqRqA0oQ9Iw5aRYOYiYlUiVaSdL77JZ3
QIWZgPkky035XImNqzs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zb3mEJvC1D5ZW7MTHXbwlIgCtA466qg5KcnOUvdWJrwOWBj24wG4gVt9yUNrd/uvHMTVvwkb4LAn
Ksdx8TXZNSQ919tg7lRcg+Nl4/va6jkqNPhYBEcpDv4Jiq2w3Y3wDmfIwSQF0ZJ2y7CGjaGyRM3U
CQhLre/ksPLlXyuUj3WuCXaKVHQL5eRVPNBVfKr8vFWroq6mtH57slhC9ezuRch94hSqyXnWl5Gu
inAv3QO1bOKRqrEZ1p0EoGeSHvVGq56emiutlfcePugNZPHZoZm5cGX+UqNB06dg4/c1SKsdNNcz
r7HevA+DkGwWrbS5G1ByJEVaKdncb0RaUKS9/g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35376)
`protect data_block
+8y3FDYQ0e7z+wyjs7wy353MdJYtQqaOm67yVCovEUTYCDfjLWhNtrBdttiPM3sDWfHo3nikMnhR
NKOvwPzfpBpuovE653Lk+DaRj+FYMd2riZxL9zwu1orFI2Y0zSNfOAdqM8tEukOb2UikUpPoGfsI
wqXWQwUwJAwwvTT/iiEKUBYxk/YhtbA2N+T6lr3ZJUalraBofB/+rYIohQ+07WoYt9JNpm8LXVrT
JDFo1ggubqtcGgCYlT3V1WjH/0LAruiwTFoANqpDCidRGufXrLHyYXdrO/hmfi2IBu5F5tjcKy2k
zjsGHW8pdPaIzAG2KwK0vVZpMleu70R2Up3J4th3xsZjCv29wl9KT3Oei+1pval1cqibUIL7y/AP
YyfYCNo2jNDdbWcV6XmP07sr+teE4fmqnEzDotAAiDC+pix/VR+adIxM0ywcjznt1D8fx6m17lMS
MNMH/q5KevPqC3PTMiYEHSIevVpUFVa1T+2fZ3EuCyyqdXeThuN/3uXcdR5DmpDoDN9LvsOQ9GCU
+6USCKtsnZQj6dWcx5ltrlir4/qvMFVLIEjor1+DajMk/e8Dr/3RJIm42zrRCwtaDCPLRBndVaIS
x/QG/HQGq6lPjZxRnHqYDI6xACWY0BWoDqk27/GEPdo/zHv1h46DczNvXGfZUFZylBOorsmgdXp9
UIIJES+nvRSQTOkSJ3c4gg2gf5LnnbAVGyPwBco1z9A3weVcqi8jSJq4YrsWsOQZE/rsh7QebFw4
U2NGwFG/Hzq93+vazU4N+1DNiA3IjiMgTYAFR1U9O0kX4bGABKdw2Gdgr7es7sVgXLPhO8LJQkw7
FQcafu4bMOGgXZodnA+OG7umoHaiZnW2JeC/LgSDpuUBcf2v4TOwhYFrYlHeER7WMWocKLzIF4jQ
iBPuK7xcjRA1Oyv4UOx+aNqpZaKOpQNwOTeKBaOoqQshBf/JM2zlN43OtMh8Ty1fHGIG4lx58g9h
cAUHGmtaAh0CaISqInNEk3Xzrh+nDkt7qVEwL0k4hmxJCW/lTaUdLjK4QtV/H1lYOqD9DbMkEN55
DoF4z7Xr5r9YVl50Eo14cc3MO13HAHuykwQLlZwaw3E9LO9B2qkNVZQzu2EEw4BxiwlZNjazAy0a
ChRNDQwxPesHhVWvxZfb632ZzwlV7T22HobqgMEzPXcxRJHLkiKQoj6GvLzfbRbykxkey0r2b/eR
bPI9Jah2o6jCN/QUAj0zzqPqes5IX4vKTgbKa6GJ6ddgclhZl6JNwQlmQysumbVg1AzmJyCgre8E
t7aKA3GsTUhJV5QgmikV9KNX3PiGwor/LV0PwTDLqGPV3lylS/7ltvGyK36TylNE/8XW16Q9ogHq
iw2km65v3v/+Pcrhp1/dfCgppdwQyVBq+aigyg9H+/v9y5LtGAWAJeUe9sYewzNAhNskFHK0Iycf
iOSuPMoBrSBtQBvnlNPSkSbdkSb517Idx95EHBn6nHnK0E9x1K0BRnk5COoEpN6bZnDoae4H5/A8
XmMIOOv/UYn7bVIaSOh0Cc0JZt+yBKqKV/K23HgivUucVWEVFe4cwHtFxNuUpaqknmmvdgHG5ems
5GB6+Qh5uu9d3u4QuRGsqHp49Y4p42t2TK+hy57GkEsUjhucYGBMvZgEhPK5ng1/3aUc3R3SPrFR
QWeb4OMLFA42Ve0bZbaREC34rPQRu/BYn1aMxgh/mE0PTl5PiTZpkpViP0xUx1sqiIS2isRpzHAk
ZSmoJw+1aY+sWj5ZtVc9TDSnShh5HusEEmSCuvmub/zRjMgGuqYbUkMs1yu4Dmhln6C7AvLv656J
y+vpBj1FpsEHEhxCmL9alPoPTmEOEjssDE83eg+lkn49hB1hkIxctsaMNNC6VPi6zMpRUClstAgf
sitXR7FVNPVcJCUxKgr6cHmWCejg3eC1AYreJB7i782TW1VQl0C0W+D2IXAA14ugDFHlzERp7KM0
8rxLlZNPrIBppeESm62cv92VSmDhi8Zz5FgxMNpGDOMLRHKNLBdX/MFcj/dbKI915SWvSH8A7Os7
CxUo9r3vbO7vcMm5ih5NGsSRLGKfiXaa2bgmPYnCAh+7gtda9tqgEBsMhvF1DSxJTZEOlqJBkS8M
6V5vwcC1gTcOLIjxOxx5p6OAZ1hwKNIqozdsI0VBpCwDHgHHBDYBXB/4gV5LYYO9SSLcBy3NdMd/
Yps+HlKj4FW92R6mWYh1n7biS7oZL9Dy268woA+PXinrABaFBjXZv/xns6mfdFmPRsgxsFp7+c71
jYygTrofUx8EgOiX4JDTGAeIPLOH0UiO5kI9mfJsG+P81yFzrcZOHlkUQujaqmXDo7w9OjPFR8NU
ZV9jj33XzivacATI5k9wi9CR+NDO7rhxHq5g9dqdD2/URCmzp35BjLZ0KHh/KRluTc6uJM1LyNo1
UvQE2KAQF2B/Jx4IuVUk3meeUTlcoTA8Tg9dAptO/NnfGAAl2mA+aoj8oPgrw52nRRvZGNLz3Oul
rcifEKjbNzdgafPWzhv+zrJLItge8R21aGYkta5eIX0jN2uJxac2yMYU6QQpG+yjDO9oSndT3xL9
rGQbOOKkmI4VEM9vZKjEetOW/ryWPCvlQIQ4MAvkaTPIQQPAZn4hTWxWJndpVFm2musWeO3/R2ed
L0HsGybfi95f5TQEtslZ2di6dRKeIh79q4vIuNuMnFMeTKBU8JtTrcBf21ucYkowik0jMaoNSVJg
HIJNx/dXVp9i5a2vMxtNz/vOObBH+6nYpx+e1KRLun8UT8NmagbqF3Q41tMFe3fpOkS0Y1MEkchG
xp0qHNPHCsFHblTdeRdl0pbx55HzkEKEz+Z41qAYTn2yg6R+LOQyfxdhfw5YGkxrvMUj+8dlobOO
QTCyxbLZQZEe0120CyS+2H1k2qrSmLyPP6EbtXjAlPMCw96SUbmfk93LQ+3oOrKQlaZLX2oix7N+
BEDMgsu7Jc/E4LIyWZ/XzwkxuRQbtMmOQsnItz+JaM6ULSVugwssuP6frvA5RQzpz8DJIg/MmJJS
W9+qKC82aTiPsjpjwWq8DoddiSUWSeUreSqxrOfT14b2NI6Ou2NBuJ85OJ9V0Fho1chUGbDYSxPE
NI3W3YW8GfjBmUWStkFrIQnGLwP56jldlhypQQhyTHEcYUWVJZgKVN2F0tIYWQp5ZQt1VOa0KJer
x2reCRuUC5XhyqGW2sGWzbTW6dCwM5Frdsn0qHhA+R7HCpMRmGGbv5mMMsRcdTCFYYI6EJH5lMki
M+l1krL/KIEa4U2liXX9187BPhE8icdp/tSXB/JhjYGAZVtVWp86zC3ZLUFLwpSFvWjkcRqdLQWe
xZqG8SUwgXbp4+fT/gFCtm4OfTdXSfzAosRSMaK9CEir1TmiHZsK9f6LxD22xGy23XM4u3a6Pmbf
CEz7eKvN8oJhAPKSsmv31p6LihMrxNGff63lEmnWUee/LNcrlLF4KuainuEydclu3vY13V0XJHOj
zFi5fx8rJNYG4abx2ImhPw25fnkAeDpm8+d0w4fCzO+MqbTcMnMQGoip2mIiDBvqOWJ2siQHeE6Q
dyWk/zXnO4WE5+TPjbXplkqgyqU1cEeXvfMY7wvClvkLTSry2K97YEiehqmsi7Iq/Zf9+ChRiCzu
DvAPF24a1dsn+AyPbawJMJeffBqARWOReHW8mRHZB2mzVFiPWUW2d3nwy4yihhb4PVYaUHjuiN6M
rELzEt3CK34+gXsyk+oKaPU4JSrR/EH5F6BRtmVwHK/vcggbITt/ehLuMCNknC7zWvFGT4UWDQXW
8QeH8s3qEIjF4L/UzDGBJMz2OqC83liCrmwXkvlVi3Yc7uixK2MgAupbX+qlI2TEFXiYJbHbh0jG
7zs8Z3sqk2K2SJfpfktG9qiTsNBp4QeOy5zrtraSs16foCKq6N7AW3eAGo+wMxrLyXmGtjwuTV2E
G/EBlLGPJeBba3I7unqecTKDXIC96uo+8mM//ba7OrEC6LJmhscpYYNr6Bs13+Frr38/JEw3JkYi
LKURJTKWE3X1BTQHOPxC3bBQuWtqJeukg5fZbEPSuYcK4Pja027PLrwB0Fiprdcq3XhB7rggbVWA
DvG2LSSQId2kPAk3C54rKBqRF+Y/HwQpL1vnutdQN/4G30Ro294iGnGVIINHkDwSrAuK+QefzIF7
ayskj4PEFglq7bK8h4xRmNSUnj97uyS7n1yqZf2Kf5/55inZpf1DHM5oB6vSRcF+vgFB8tVdAgTk
npFWp13vu0bOTZW3JjOkcmsCfCu65ZZMuDSo8jEKLQdb3ciSOZ8RSPi3riZULEv/bdMFYpkykCQ9
vL1vm5HKXu4byffgDR7Zp261P0KlOAvN6tZVCFXoNA3UV86sEI5nqaN+zZaM4+7wNjybvse0j0cE
ZI/xyydDTOwtkxrEJqlNk3ZYIbTx3rtgRBboJrmyUakMajNL19pvg/Ig/TzmkJxRhAN0kgrmIZ0U
3o7gWNJaGofWNA4wO+R3lMG6giyP2X0nkIvIBXPZsnNdBcHKtSitwBaMI+JPWaCIMsk8Az7Wjp2q
a8YyxVE/ZR/glLxPJKM5i4U/0kRFMhEUQxRIuAHbji+N0zkPt6J684yjWIyVYpUCrR+NtKM07nDu
Hhtc1gOe4knMTmp09Ld3YfwHJUqpNmUygvEjwhZAE2/46U6jy+yDhQWZuT5HC02l+upKLa2YpLcn
lKjRJ+NEh64FqMKlUUy2cszlWe9wor09hEc3DRCiD/qji7WM/mKIvJfrXvpuh4/DlqNOVrPQD/dA
WSQWZEV+3IGKVeuExak4AgTMhme628ca00RBDlkL2/dGiIlTYIA1/iIJTcw9QZdtUg6Pcp9o8dEQ
A3wyFw0r5WI/Ct72mpUCiSoGno7NttXFuJ8QqvyRcmK748gyrYvyIarA6Fn5Cvo+1RWt/EDLNY+5
QF+r3GbTLI3Y1SoA60vWpsGKJIhEDDWuKWUVfdeUxjSu1kXLnsur6TDHCKRr8phn0JfQd2lv3+tK
rLHyKEkNdOeFgladgIHQgD4ze5Zr7LJ/Ef//ihptgLr610Q+sOcAnFFX9UGdGjiM9fc9iwWVqwmu
Wzf2Z6RuIERAbV6BXaebelqRnyrS2F4hrueUAUgMJ+RIuU62FpCwJKhUPnzSS/dwM4/ogz37e+1m
KkpTsHql57x5xIT7Y0MKgB3BrAB376Em5Fnv5Ocxvt/S7+d/CxcOyTK7yYUyjZZlNqYdKkqXgYCo
B9P30FVZgN3OdA/qNuP8btQk9U0x8sgSkHc8NN37V5rP+OW7EhwfDRyUJYAjabQLYMoBAOmtDYTQ
IubY/9xX1Zf5YXcmJdXPL6pgnkCM205jLuR4a54YfLHm1OwUaXuGXX1w5YKeFc8SAMAhTyCJ80mK
fmmjdKx9pWyhiE+s7DKUUaiZ5Wb3zEmx1aqaMiLC4dkzhXaVLBjFeklJSzr57myGpXjFXCzpoeuE
1crUUMT/R3B9RoLUyixl2p10xG0Zcol55siukQXdST60ZkPKVDFWgB57AoAW7ExIWSTZoOo4ronE
Bk2+4GNQrk+HQPKIpuJ6RlHVLwNFxUcPjnGTn6i21LAN/CbtCDvnsjRhrAtYGFSTl2Xd0CNeIPBJ
ajuHrq4x0VpP7eeFMQhYUdfED3foxhSaIGtzUWTDDQSWU3xYsdQyJAP+55pyhF/YSumZbuFU4PoK
98u7pEfbSvxRrYOXVLCQBVPIFucFKlyI2bN9wCW5Ds2Jld6rB+zCeGUM2jep3ITSNrb+UQbPe+52
wmGsGdnyvMuYAChLgCVZYZz8HD9Vzw16rOmt1H51m4cyKBFWZ8XD76RB7dkKdoxGuLbj3BJncJOp
FtgCGGYlzqr4M4td7v6+Uip+0Xv7Ynhl78n0OkpsV6PMWtSCb7tr4Kh9+SvCOWJ2IRYaueV696zg
9t4vyHlvXNtNcEtn5XMK6mLXVyYI9qcXX3EvJwdmihDMzqB9wweFIkilaPmvjFp+L0j8i/GhwTz/
ZbS77/2QluvIHiZlR6BbjJLbXRa9UMT+ezEiFamNeJUxSdGfyVlI9RCjMZutvMrl+vqENFcvWYLM
Ib4wcMdwOtMZ7igNOv5qsPnJBy1ZEWQVuaORLpjfJw1DMoL1QWj/eo94izHPc8lzUmz434hrgOFR
199irJ8b58bKpDm3B1qx1oRwnPz19cZwnXJTD/RBlEdrUwt0z9BDY3LglK1h7NZhi8pMPGSmePIl
Jbj9BX9BXSdJMfGxEO2S6T4A8cj7kKGLkMxsutcdGbvrj0lQS2nX4TXnN2lXcK7m3YSJNtb9pb44
sDu/JzU+vvPj0GLiu+M986DZO/wB+ah2vffnkVP0oX2yFYDHhmGDLIdgYq6/5KFHcPgP9X6SBuyq
SaJwtx1/J1xSA40CgRty6beEHUPKPA5E72XQB6IQWpIBrQ5xbiEKWj8fXSUNev0KnswQxqZ8YcdD
pCRsHLojW+3UWpZfoc3GvkLVesfF209LkLwy8qlTkPTqG6TuQ7D34JVHOJDguAbsJACH+NF01TV9
7cPf92yG1gvv0Qkxt7dONwyR4U0VmoTyuXRkr5e13f+PoE6NBzoSr4aUdvZ4tCg9PRc544e4Jp14
szchIDd4dW+xyTquPu1Bc21usOcMINNlPBYuH/JWs28UEekunMIYOz64Jocims6yxxjeBYBKJm4R
zacIw30W/AZtw6O9XrV0RamMvSxhvhjrOqwRcYB+ESe9iNmelwXp40+xs/7S8HBYjRdjSwit75iT
EM2qLvpCcN5rkhSbiYKad6mhaLof+BN/4EsGP40deWyFScXjDAdbOX8xV/FXFmuoUtA0Khc6nmok
x89FAJ0EYqpAKmZpMd1qDau3w96jCSy6CfsgtZEwc0YLlD2bZEYQ3VDSrCOfttBo9OYQp5Qzdf/9
2gDfQzwFTAUZlSCzdfWFh69W+jTVvdqtigOHLn7kdL4CDAK5AxesW/n70zQ5c5HpmrRkU5xcf7P+
H5IH3fHMqyrZxCUslfifUbFD/9labNPgRFJ3tnU/XL/1U8URkth6h8Wp3hNWtVDXl2IvHwVKx9y3
XYs417caPYL5Gul6ZoE7rRnWTsdy4w9KjNGBfFKD7XzJFn0TOXloN6uPsdk5/lQdnfx0NQH4uKQT
eXyn1Tg3uN2loApU22cxsfqxaXcm/25sgrOStWbp0mTLHDQ8/WNyXzZCvgs7p/3xduJAa1QdH+vV
5eXYCzkISp5AENXPq7x7h/hn5++DwcnTUcsJA1MHAo1cvgWsDGY7ZjA84v3fCR6Ck90aonYkm6CQ
TMcP1KZsU8z1z3nDXoEtGcsejm5bAVYpD2hHXw+EtrYja3trPNn3xKHNJJtVQIoGR1xQFB5Dfvmx
SzCY93FZlfKC0AWoIz/kqEAJUq8CW0tSCqr5hqfC15RjDqLBvnYPh99YTGYi/vVjQY77yADICHgV
vFhAL0ImEeQ7C+aFtq/1n3dMWazWR8dK9AObM260nbSgZ4RcXUQxDSJ/cS1iw29n2nvNY+DgiJo9
qrpFrn6YQA67w6esmGVg0BVxov9v+syh0SlPq1qhEW670camga/+VkeKFNVsqctJhs+Mcu/QB1Lp
RYlYg0YCEmj3i5c3/q9kGJl6AMgNlhQmAwEcTMpkniJb3oCDm+Du0nH7qfECJ1YLANQBEvWppYVe
6Qf1x6uq5XBm3jt9zrth4hezQZHheQx6ZEHbE/UwvfyBbRnFWG73UWpH8rHRaZhX0UX9epygOMmc
qou+HIy3AaDIwDUtLVm3oe8Y9k5n4mwgXPJO3vQolBawZkPijqo6vSnseHEO81zM1SKMDvHC1/0b
5+vDnqSTccOs9PeLfvaAI+2MQYWMKWQh4b+o2VujcqOMBNVO3tV32pVq8miTk3W/kQVpjWh0hobz
EGAOal43eo0kpWS5SHTS3vdCE6pDTt06eMo5YTz5pUF4RYXI/VZ9jaObVPM4JCUqQYI1P1MKPd6A
FPHA5huSaeXNaUh6UDNA5uVDENKb3lhosTgVn6OeJEUozpWtE3+FkvO8K9fEEQjeOiGGie5zOzc2
7yAUqX3hDSj04Yq6TTb+ifTJ5zMLDPO1iWfXZ5uWML7szwfn24cItSrdGFbjnn8WnFfc8nV+WL4S
KA4HWt8C1AKbTDHKn3bkBfSLob7QHubhywQ+QMzCYNUZqpPPwQA2ijC+me7ZXUDTiYbMVFGbH33f
q9r60PGK4Ex3KizEE/RfIfZawApUD4DYwoSY9VLIWoY4YeZGSBS/+9/QfqoGfFDMPu2jxwjTq2u4
ShH+Y2nncDSwLQ4IqCaSzxpfaHBKp9PDO8naCk6FweuM7XHpwh2lKWnZ5tkNjgeBfuFpkUYPRptL
reN/NV7mjbyKiWsyKtzsCEqZ+O9h9YqhzjVqLE6mFr5AQjcOI26fN+BVB9pTUl+enlO8GdUPdG2O
/WCgfCZdRuRriKkP6YvKNOA7yJ8lhA5lTRzrp4BFBy/WjubmOrgIEGV6XQ/ptG4zdwml80iXCEzz
jioeJthCmdpGva5B/ZUtipHy8F2cffX1WEx5mAIuZ54/cBk9TfOqIQVmp1Vs9Rs7OzB/TmEzm1r6
l+/dckfRxv3JGfCrNe92KH2dhdRZ/B4npYYcVx1qYfL0IASvukzNsXh8VKl+YhiWrqMER1TVcFyO
V+BK/8AMyxJP3D/bW3Kx7olH0oHuAMtxiqSBdmTTsFiI34om8TdVVCcK1hlLGQsJrncrMFVyZa2s
JfjoSfhQ9IVkQyW1A40GSleEERKqXjDpbon0CWiDPBOnlVUhsOCXxeeRMInlh4hkSmwDK/Gdgxow
H6CoVP7QZCPj7VAyy/BDbFrWylLdZbHGVEDfUQmffZzWKWmdWz4BPpkHoYyraqXRG7e17PzZRHpp
0jj8JTwZTgffsFS2Nha/bdUxM/DZ9QnIUAhnW/kIMfrrc2XSfhyY+GtVa6HIUOwqfmM1GlGQcZ//
zIRBhzcOOiF61MEWZW2Rw6qMJwd6Ej8i+xQSiQSaOzcPrUdqTwOe3qBIIJRPTzmrFaDOgTeckrlx
fvN1rDZ1IBzRBfdu7BPX56Om0jJspTcFgjZs4ysHBn5T6EvyFXmhCUBSuoASwG0TZdJFbZuczQPw
BGWAf+QqAC/r9+GORDLYVFR0TQav+h31iH+E7RZXTcjqQc5kr+NhSCGwT5bKC/zfXS2UOlfue0n4
+3ilwdO+eU4GEwuam+Es2WxRNwNdkvtSWc7rCpQxCGfxJpkfMORyRIyEccAxfvJVmaNMtYlvRmo3
5Nz9JG7w17Li+9y1gqFs1ajiSe1Uc6tnXbnJ/p9sOSXTB4QPHKa5r/iL89dLQV0jyar7uZgBDEhc
dkQMwC2sOPgEFueq+BfRGMpahlGCeFhk42UT6CvplN5ZJAT4psZwlm3rpCACt7c/HRNDNRgli6tt
3wgEHABlqX/jtM5hMsFdmXxC7hGVcm3PFg34d8ano+TFE4RJJzuU1TUcKUP2zEJheWd0+nlrTWxA
o+lnar6ZtT5wFGIEgjSVDDhiPakytCaKZKTbggeAlpqSm5RlpXppElmvVlpeFQlioTArhK/Tnh+q
ff3Y9aBHlobetEaKWmMSSf+LTJeieqg37zkj1BMhF0QFuowTt0EatS+QxG6saxsquTxZIKsbkUat
LKDRk4VWC6kyVFdQzXEyE/INYQnTW92Y0lnx6lSl5HihOWCpAoZXinCw/lx6GqmRwacmfwvHgkz/
xyueIKm66yWInNrn2xi9933+sF0jsTBXjtRTLalutvk7Q5924B5hnJ4MnFEghuy/aYuDaPhsGIq0
AVFACflDQF/SaKHYbU7XPjon9GKjirljGtd4vOyUVAzBIi7E8TkYOJEUmyGuFxKjdPYPHSgwwLY4
94xOyYpKXJcIEu5bzv3l998bJJzZAv6PtFk7cLYe8MYBUwwjLvsrGyE22pJzrJd+usLvJ4NSjNoa
a1xBT1E6hhaPUhUz7+aPt0PqWUi9pAQWlXoFTm9XZJs2Qz2Cx5KAwDbhCz81DVEdoWkdo5GojCuj
fk31MsPgsmDnJaqFB8xm98+HfDDRK7dynaj66znGhgECTRVZ5AKPi9zRS/ZkUTZrZAw5UTXWfGxr
8a0xviopagB1SkSicOu+a+sRBCN1DxM+IdEcCw600k7hXIrDCw+up1swCNRd33AK5FmW9KxYa99n
5Z7w7wIGHHZyB2chIpTHiB8VvnoO7USzTeNlB+g3PNBGFXwaL1rRM++n/yGd5RiHIaEQrAGPmfdp
QyH3Ywq/1vz2N/pG4iwnezpdS4BXRDk90mEcjVycT3HLv3p+TX86SDVzkt5yySn04csIgi9CvIzl
mtsvLIkLnIl5PKPmzsbfg3Zqt9m3IkxyxKgGN409PieKxZxUMgLKW+zdeZ1yBY3AdYCSJnu3u4gL
CowEA+5G8SoMHP67XsawQoJ4wRrKXNm+FR7t0WU3FfDPBb48L/GAZiFrlfpBBYo9R5MHHuf+koA3
wDi+0z6vseZHhQ4DGapIbHNYk/OqzSTNYUc7beqnM7Jvt68k3keqA+EkBK0Zq5STqLxV2m8vwgFD
QeJjojrr3BucqcdRfgx++6WTVSFlBqJmHiVTFv9GTjfT4TTNjPty7mjd79ffuV63uGr5beDoIyFI
QISbOTjN2cODpUEDEntAoCmQNQi/9gc28JJAcJGqlY9CqJ1weu0zYl7gP/GXCOWejFNCgmijqe02
d2jaP1JJ9rsLczlaYjaPezO1/TdhpT2GjmoEvElykilhXfZz7FUK5qg+jBqZj/B85oqIGtfQU8mq
yf2hcgQ/r5u+KORUUzQHypQ+opuZU3jTj+rbVqMeESN+w6m6lhA0U0YM+wY5FeMfqlfHDr4kOkfs
2CtyT8usAybUQ+u8ZbrHyt2BdDYPsAzQkJn8Lq7IhlUZNAnc+lM2IGpnRuJFQcg3FXDGJFeqU7uD
LFv1O0C/8LoY775lS8zBjKDoHWEMLEE7rPGIIOgjiDaf4P8s0csqNCoGn4ioVfSEApcpo3o1kpe4
yTLtHb/fBN2VJpe8uPbXbiNHMBsEVDTxKIuyTARh51EDvGTPOmB2TMjE1Jl5Je9FhCHk3zZka+3z
6+R6XDVbn4u2ZP83GOXHsaAWsdGOg6vTf0YG9qpLeNeYiGTLh+r9b2hoqd4z3nA903/IOVlnCG38
YmNkpIqwtY9EvtAR6RYYc90qTx8Vu+jOqBIvfmlz4GAygQjVt6IIqQT6NuSM94YCizR7N99ocFGf
52KwpujatwVhNrxqyfw1lJsExy+3AFCxerHJ3tNWMHu2Sl9zVJB2zHIc75v1dybJAVeqLn0e0jCe
VOM5in9nmwYVMLTvKm5OY3tf3wtad0xT+OlQOICxcH3DUlSyTZ2JAH2J6TOHqIsxj+cdsHV+gkRX
eVh6qtImZOty2KrFT/dd0fgTHErVdA4r96BT19aDMvoWIKbeDlEDbXl1Em9pUV6DwcKRl2vMSMfm
fctVS4qGXVzTV0ndeukSMCwXsH11f/jnb6rGqZvVEHaXPh9EOZcvyF5FsvlEiSFQA4kaZg8GqFMM
koPtYnwxoA4hxa+1KGFPnHbmvMN3x+UXacx5T0k1PAyau4fTlhnaTDZ+M6pLvXGzM8nhHhLV4fHn
Phrou1nabEN64U3Hk7QgHYOkalrf7Bv96NeJ051DWych0/NCiAS7fZ9uDX3xf0gDmwD/hBLXlLs3
6V3+g9a7TprygqKIzfJsMHCo53tuwfrbRkYjHb6/q3445CccM8Mm23xLewXV5sbTWWfru1DQuVRz
RVvSO7aT2by2pdpJSrEIQfAHzKtN4R56eJLhdkID0KgNWYmI7lN2nbg5Z/ynJyI9sIZZ3t4eNRUo
nEr7iNDDwS8KoLtSNKLOQde9DwYDX6pvat/aoAPYNQglyWhcQT53H1STWlfx9d/3+b5PffeksoqU
iehaH8EovxcWg/jX6dBWgUXpbMRImdLg1VSxL2rmctTvx2B3fXKmAjo9OBcxxWOmfytxhHGhwuIE
Z5vu2wUZnC2aXdKyD8qUdodSO66ZAapj5XNlGvHOidUBQSRL9kR9zkH7g5uU8QN3xgoNLjxfTfhE
OLca76Op0QrO8gyDqJ8ppRdGgHjBab3xG6DeGbgb2hgI39wwerxA/7ZL2e9ej6FbFBeaVQbU3FX6
kK3bLLTXzSI/ONXrWhU34YhsHdC/M92uq75NxRjJ6Fy7UykkZ4RIl0zGS6ESjOXyV7OoG5aJNmQl
BGU64GzTO0BQN3Yw/4e5YQr4ELYHWApM6BKxqkfmTIu9M04s8437z2Sa/x3o3oJQOPEJfsFSwmx0
enIAaxdXRwRsGyid21jGHIH5Z+MVoH5xe+XJ0KVCU503tSx/NP/tjcrcN3zHcRnuGV01MY0cRRs5
B+LHMRYrgAqkdsvWiWu0WxhAox9XJWuPIbt+A+yZLJmnSREskdr0uPBWWAVNaoKJW9hHXyIpK9mU
Wa+j9gtQt3cefQO5Zw0TVedcYUHCqxlauIKbhB/8D6Gp9NrNcVU2jqz4y7mTmKyZ28L4tufHoqTn
nqaKu1IeX9HXK3ZoHakKbavnz1/XzWrgthY1LvdOJ+5CvW/QMqyvcOB2nrNVdX5vir0kdoy3bmBA
qsjx7NujSCxL81RGzlsu6Y4X8Co2zagTvxwyIqKRn2mBNEl6SPHiSwmpcEyHO6oiu9YmdV4kOYHV
F0uhGDbBt0twNV6MfokhERaxtSDqY/8t+PlnPQ2jXW5bKhenv5bKorSmljgnlScNLAAQ1uKW039U
mGEz1YA3/sHVoDWMAmPsxt0Zl83KvHxDGKiMhQ83+ICbw0X+p+2JUg0y7E2pX5ByR/umrEgZJYCm
cwMvRatAXO8KD44H5xtwf5SAHidObiqy7MwnNDAJ0WJ5TDP1pS8UKL3wR/Y36rmgTbS9mI7L3ai8
l4ubcmoEhq3NuaqzfnBgaXUtLohO1ZiUV00Yn4jfgxMT1CYVEN8hEImoHA5nXoypm7oLvuB68VAr
gOuEyP6PZTXQyFTZPapoKU8SRlG8k7hDt/Upud+MWEdwNfZTXb9w6qFgKUbGfrApgWMPWAVYgeYy
Mb4/xExivBpkxNyvOOGcH9Bgyf6YUWZ6pKzLE0kXnBsxXmNAhHS9b/jbyn9lo8/1Ofjx5WfUXumm
jZ+BSq7dp4HR+ZSrZGv4ylzd0aCpmollVW6Q5cgxSIxa+cW0p03zeOKvSGZAxUGBuetZKbJfQggN
+dW/JELmaFRTiWiZz7OmNwus/2qSZwRgv5hnYmMYuRM25EYBJPvJu8yzDT7ZDBn6DTmk5A/I+9uM
6V2ehnYxJUXZlYudM1eNVshrvUczFX7r36wD9l1j22nkFlMm3TE0oBCJWJCnFgevxCJyPqX8tk8n
bPrGhVC7MpqnAFFgqLtQPISCvsPab4u19eS2BUvgWOhyUIYGZ8GRqiwwdmcjkyUU3Zori0k8IVwQ
FwLIRRdLWMQ3Soe1+rcMkr2kDAiIefThawqrq6ZeM0NESIXMNV0P5F4HI8Zv/CmstPtWUxD2qMuG
F9zRacJ1uMHi4aewS5TGM34/T0vtCUICL30vjx1TwWQXLANdyYsjbJY+VNxIj8jv2IhXm1DQA2TC
xynSahvwWxmeDLDg0zTj0JSVYAiJMjaZzxZ3Yd7fq0JmgtWD932lpigyyAXe9LVlsCJ57aca3/i5
aVSRGxIiXWHOSbQyOKAOeWckv9lS3OUXUgsOMCZXK5LndMFoTEaKbMf3arIPCMtl4+9of1AVP61c
7gMhxVsaRyYm8Qn8cwU6AGkv/4hrBe1/9GAWV8h1xr64zCxfdlYYi+knEBDVKpxTU5oN3NlyRFRS
r8wH6hYVD0P0AUmDRYL6jMZEQho97RYsYBPdjq3e3YU+ej9jfyinPxRcs/tSI6dUxwsz9sWz8JU8
3ZOQatmHCq3iHc9qpyGtUYUZ1yUHV+3QR6T+dJCjQgg0eXmokhmqPZlW3J/iGy78dR06WC3RjBfT
2mkPchBjb26daLyikTBht6wNWfiWRdZ97amaWNy56WuEr8OKfwdDtGOLXDxC7NBtfTKqt9gw6q01
eXsefahFXKXRbIoVYhSuv+aRJA2eBzqMLzP343ad+BrYrr/Ci2b6vwo4oruPX9NBuyH4NlDBXmQI
VWionE2cXsg2oG4v5VwNoubXwClxkbinwn6Wr73jeSzDfDAfre5pb48th3pAKq/YW9oDyXlXNfQR
0Co19DswHomfmogjm6xlcgxDU50vxDgsJ3nymMDVTlXfNk7X6yGCdm/CLSkV3nEkGQpulx3zbdWJ
YUjbq9I/rn/XGomY4/pSPV8a99mwnBE/pYwdxdVG9w6EbFlS6ZuiYcBMyuQQbKz1oyIUJtDpEtD5
NBnQQPUVubriGxNMDGDN1MHGCBXVWujZhbew8wOMmHv6P3nGV43QjlvzJ1Iu84nIknjX2VOhNYUy
TVvfgEyOzP//4t4sLPm92fYZ1qx9l13Ws5RpvghjZwgPCuy0Pdy2ELyunpLM1MQDCbCh1wMOSysS
8MaZNpl3OUMaG7eIlsJoydAHfcqIA6XjPBMoYBPhMSaDX23Gy8mNounA9R+YxB7JlDTxfQqjXyeO
O+6OGsdZaJ7lrOqhL2PhpJgIUUj6N2G1itOLcBmgSaMbECSt+b/lgVGp4ngc3qcJ0ccuRMIdfrQv
lGUtIWa7GLydSld8YZ/iYcEJBzMEFBqupthhA4rIB5Rg+Lc8JLrndgnZfVshvmaal1U7QV8WidCa
6poI0eQy4I34jN0LK2rbb0oeBLSb4ApEIw1+3/i5tmFKZDERp22f4q/7uqQjiHUUJ5/rVtdRxKKF
0Gduebz5BCF2GmlBB+Bvl82hd6oCdG1SkUfx98T5D7m9tmyQ2hVokBgFeDWoJgYYr7NV1/9SSKLZ
t+NCDVBlkpv6rBz2S01ASOM69jXx0wexQoD3nY34uBW5Ihqhx0+vUQO6u70tafC2vTjxy5vJVu+j
5DuTQHTVdhKwXZWoOg8gZnc+Hz1BzncB6QPL+xAfer0EyLAM+5f8rbWS6ql9uCUTCxV5bWgn+1A4
ESpRt58MvKq3UHqQCW29nks38y1syh9uBPXr4u4kfsnwwj4LGgDf5sg9sTfd/9X4KluSdNEL3bAC
VCJCpRZpi7sixm1EX7Equ+UF/XB+B+RV6mYLIqwQJPXAmqcLcRxKEwFKbUPZwof6ykY2OBK+uC/S
v/ee+YjlxmFryE+u9yIsEL+M5MccbvwAmIhJFd1d4DD1qfdiiG2ZCulI/dCkpjjjQAj6EjMcQH1u
MEF3YYuf6wgPjerqsGEl+i6r0cF9E/0S04ao3wMsGPIJTcyslZskHRPdCFlGyEKdMp7FTkaRVSlS
N/7O8aWkhIuXm/XFJHFEwdd8GKVVVDelVkTBq60hBfccKBGMJEcVQo6km+Bpssf3VikDgsl0xFN1
KetQncf9a8phi3k8TWbPtNW6D7bObFhpODkZrU1YYvmlvTV/OwZaSPm878OJpvGWLB3CultzS+ag
MtYmn/1s4K+zenJH+o90968UmmmZajfXmKz1DuuWVTJQbP906Figx0SWr3X3aCUT/taxLEhtvbEA
BClNApzEwqvGULtgE/VOdE0FYdqb5+v/aFJI0RhHyOHYrh3snGvd+erkLvlyi12vCGK0WBt8qw8u
lTwSrpNSS8hRMxSZu4x14nLYwovzXQ+TPVTONLMLaS60rcEbNtMj9EaB7FSgNBcoHQ4ZRR4xA68q
7C9kYUTZLGEW8Y0DcIM+cmgFdoPYgyO7W0tn3xPd4EZyP8zRIdof67WSbx451C+oFKWOTvOHRUZD
1ANqdcnvuWTVpvjNekkly9o6ZPWTBjVQ5nwJyQdmXaAdNQhyPt+Mry845RATpszQdeO2HoBtuQjx
E4DQ08YsYzS5rzu3EYyZprLWriJ1E7HHUNsgDK9Ajx1w7S/KDHFuqfVdSBsO62wzeyNgdwoVgSAY
pk43ZcFwXW7c2Zo9e9Zesa8ZLUMhi9pncgTBFtBHkkIMSgvwK68imKq9oIxz74+vgTcverVthdiD
tEIiKumIKMnWmGB4PTq2kOQCn8Qhrc2LLH8e7j9HjhaiQQ7RLR2W1/iqg7MwQaoBbdf1u8zuQd9O
aINdGrvKLzVh6Gn4dFaWRrIa1D5VwP6e3ro0y+ZAf3dJ11xOiE2vUc144Qw5HqgtYel8bcxhwUkq
wndgI3aFYZAEL0hnzrM0aY2nnIX3yGSawaf0mQzj+JRmoxTkztov/xAbzK17MTByrbykO48NQ+b7
roAMPfry+srqASrb2vVRfxYHLyhbf2p3eAX9M3Le8YVnovDyZDSwE+0X5smLjaS7skITuJ/VUeuv
I/hLVivL82p39vrt6VllFVoXaHFXwITQNol2eeIIdi9F5FUFK1OomzOByXCDeJWPF0gbp+8Axh2o
zSFUSEOKR/lFf7xaK1X+sfcCOgAbApLJmxT0gd1yL3yXrUGL06lVrhc2gsFZrkVMMFY1AApAuIkw
8WmohfRIdmDQWgrJKEU1lCIfV/jRMNreiXqPu2pJGY5iVjyniKD5D8zu7vo4KjR9iznFSbFclq+E
GX8jH93ntrUXo+2zuIrc7NhlYdkVVk2cUUqA1LwlegVTcsiV9sNjDAXT+5Wg0suqwrv8SmXl8gJR
02pBB8AyEqn32R/BvjXQckPPb/K9x2A15h/nMFMJrZyQ575gHt78hBIkRVvcmqN6EjWcTDPRTwek
OluSVYcCRawyMOQoCoh76Cren99LhmsXN00ePb0KU6RBuDhG4rld2E06uV4vM1FsPr0rCEGES4B3
Xxd8QoxWlUk34ARc5wDyy666FB/DrRGE/wSLHo7MozymJwx/oMIVYMuC0xATxIsc3r3/+dPjW+OD
AeSyXXLPznXJIlhqKNrqxDycCJyuTx1ykbGv325Nwt8zFZO7Dhy/K3hhFe4/hCIdJnavV8sBVeSC
39+FGQcUvlmZRVztVq53PBbeVCd5UqLPconBU94To6kuFVk+ntD976+22GWt7rb30IU/75VtfE2y
hko4vSQRcpo6xaVcqQtMU3I5L7D9g/5fW09NLqO9qHVjjWuLoID22AIFKxbRWzoZjGM0WqX3OH1e
OS3MBR7cVdyN9lrG8wZNgPhGk0ZQciMP4TmE06ahTyZgMtTKCWCgCNXHEO7p3L9b4SzABt1iR/fl
yhx9camWjZlOiBunRD8e76qprWZWv+7BbLlTRHmmEX0RCmDUSyCJLjSYfaSewGN8h+pflp0ZrzQ5
x/KjorZ3iHStJJTjuizXi1vPpjqd+/KcneCQGqAsiw99ICNChVt9bRbxS1KeKBNiFzKjJl76NQIv
jKZCLvMyoxXfhBk8dje09gNKUE8Mm394lfdnZkQgKYjKn8Ru92O7wuravmSackvgQ8PsDqJeIH03
ewzeqRv7gmwhpYJT/AuylkPeQHgkz7GKHYjDLPKCTOteSX1vwVguvs50QwnZgWGdVAjy8N1o5KGH
FapG7RwlAKWKpjRFR+gq5D0GMM3fsm21s57EHVzPidZLRKjlGynhc5tWk7mEtm2c64fsIDXKWDTY
xk/QV6MkepojQrO3m/a8Wbb61HFb746vLmpbq6cR481FQQfiWryZwL9jf585fe3dThpOsu9ezn2X
dtcNJqazrl7lhajDrguvxV7rJWAeUnKg5IIAIKOoWZVIMaP2hw4Q6jk7Bb9fX3SImZwznMA8Hx0U
TbEFnODxnH6sCtccrF0EA3y8ILqHN2uUocrkyS6qYdqXlswErDgHgA7ZxtuzYgyayN4FXd/5Dsba
Gqy6OKkdZWL83pedC6rPZraVf2doN58Lk9SeNtfguudM8PNMTmuVRTFA/83sheQgQfAQ4g0Mly48
xERuAm35tlgvhaVcJK609iFJhvrYd9ee2Uvz/VKvMUk7Rl6N2SY2TdSOybezoL1GsUff8iMJF9fu
2VsGVWKFMlgDtJfZjMJmUocHHxIUbYSIPw3AIaLanyvc0jujy9v2eqsCRhvwGh/Zm9Gjwl4j8CJW
6a78VNBbArcUHr0wLjbwvx1/Hc1eeNnenoak9LqMX6d1tWE8jrEKqoVsqNyd220a3VeArTfYjV7X
5jQJqV84LLwAntRzD3xqPbNSHj1/wWUqDcoBt7yN2+cRi+clSUKhGWHQKiqRfqTMxcV6sbnz5qey
YRKNypBJTL3Hz4GbJCEzURCMS+nEbzvk9mPxk7Pdqac2wF4IrPmuSxsuMKbs5OnO2hp3MN81cnak
K5GN9xamLtAmh3e+GXb9HZIyEGwoaPTp62atnfIaCfIxJ+4rUhi0FKHIVxr8vCHaphGgZkHKXec1
InlfLjxlSYya+04+S1vXgrtRoagvrlHpqgWgsq+ENy3XMV7Fx6XVWXuC4WWQuPKicHFM8gABSP48
OSKpsAnddvrHIvudwsTDXV60FNGoT74bre2vztVF5bqgQZ0YsuT40GjhsmhrMKz1HBQXdKnDEdAy
lGgDWUNaqWnX1CxMvuBud9tynu3U/X+6+oCmY/fxSMsf5wTK+/PPxkRWOgxBAfvUO+wbBT+Qz/Et
7GkpQWAkOipJQGaLXd4judtRLTRvNv9vp0Wzi9b+Z5Jyezy94IclYENC1Bq/bgEOFV7OVvZ8WA9A
mMiKGNF3ysij8ugDa3tnFSVN7cI70dJ2ENXSK2gAg6LVTy/FXRQsX28LQgDYlbDfNot1RJKceXP5
VL/6v5NgOJUBUfRe8jPzQoGvex5vnO++kMYIqw4S+H52ZzIzYHFDh81XCh9l5hqF/cSqZuJ9ZO+Y
1KGngrX7n26Zv1P3g2NUs4nav2IS+tq7MJ33XcQDZ2H4lAatj3wPajxSAMPwRlB28pGF1tmX1+oM
8iSeOjq0hfNOmR6TfK6BKYrX1hsjpz7Tej1fqJFuQzGND+yLjE16ZSmjPLmIAeyQqvXTaTc/7FzU
KYH6L6D+Er3P32QuUe5TiP8bkCx6K4O7AH07oEB9rLtCQaHKsoTGRhqJTlM/u4KJ2bTMVoOs03+p
kaL0gzLwlVvtyXDZ+3mOB2uGtBhBZNgEyX8SVxCnYWO9PK04FV5BSjajyGLPQQJc7HpulPAWwZlB
edxL9JRELoLK+/uOAo2qOaZySXEkpqrlQH+lVdrnDZuk07OZuVfb+HoNijiMNOSDuwg6nFKvloCY
HIDNwBWmg5zYeAdUV0tOHrtBdj3NdklPk/Pu4zh95FOppqyHXcfcCAmyVuOmUS/bbf1H5Y7IlQCu
CUja+oMjiw17so/fID447K1oXtO/B6VqM5G2VxXvBr8+Z+VJ5SsaYB4D46SH2BMvL+OfpeloTYT0
MHT8F64AmJiWUyj0Wy4aGyygdveBhkWyt/wbG6CsY8jjV1malL1V07RQ9J92VGKX2eIw2/wipzaB
YajtX9D/rHC/ksZWuBh0iIeDZOIhGrNDa3ESvq94o6A9tRRUjuINFeD39kY/Bkvr6joTttiJ8l7g
xX9bn5rTgHfX5wqiJiD/7EUNc8+6d+FEFRKxkR2tDNFFUl/NlYEEEaJIyQoRXYCpuC3Y/iPbktkG
heQDs4/z6c6naP9Wz/ARmSrG839+QqjPofeZ5UaIVXKm6bubWwQ4/YC0Qxa4zNtFdImeDbNqArSa
F4grwuFMpo1iDTNzZzNEnjMlkNrhyGR/eKZLg+t0Ttbpp4/D5w0gqDQJmj9OH7H+gQV+OwOKOn/5
dnOtF4JhaUDo4j7pIVtSjLXBv5ZzDmO6coboc28Vbd2H1v/+iERxCqgSC04hXCviARstD0lgwwtv
ATSiVtRa3nAUb9n4I9z5AZQraS4+MvJ32uLuLj16+zM+BXDBhwEr4Wz+QZeJsIF4KCdwk2UV/puj
yorwKdYzFHBLZeRyaGT7fvBqZR5i4tFlX54L2k7E1TpHPmGF7I3Cg2appXvKLI1ireZeXL3b02Ut
4s187p3AuQtWcOSr/IdpTkjxGxv0Oa5TgGALkGHYZUczGjS7kV4ztBiLdQL8D/TwqpHb4SC5ws+2
ZCbMN0TvDxVo7KEouKxp5egUZebEMNWevHTTdJVEeA99Ri1pv0zTQo/1cI88pi3B2rCTIOvA9qH7
k7RR1t8vqgo2WnCLcvENk5RRekZM/jBHRQQA9VDRfCpUoRRosi9c5vNonLtVG2pupJeni762IoQl
nsetbAhv0ure59Pao+N6t6fL0spB+0AattG6y2Dlg/DmOe3Fqdx++QpTUsyNyxMGfmgBEZMOrWpr
IbZmTDmzJJKBb3LL0cMXQwrFdWJaZ1HqhvCIVq9M4CkI9k2i/NP+NYhqydxfWWAtm/T6Ufcu1ZmQ
cJd5Lsu5hTApvqwZI0IjAwM9uDr0t40FtYNsDPVhAjmip6jKHHoDwMd61nJJodVBCbg3MKWxNK9H
WsMY+r8ia6Yn1CpHSU0UTwJtEngRALH5xI0Tc9azmQA0IJwg/CFWnWVAnhpDqQk8DltMGwAV4njS
jjLk9+vH/dxuhy41fTZl04kL2V7qfv4djhseNIpDLoc8YzC/Q97Tvd/7VwdTM0QVbENBIcu4GJqK
V4rw188mb2O+FhsuQZc+r4DUV3iTHur95O1T1iWMHLZKNeREQtPLwVrEJq993qTHHS9oaqrJLwzy
bX0dOZOZ0tr0qPJ025jbBJMGQFp+LW5lg5ePf1frr881KOdxyhK0ScHSalFoNviwsv0UCWH6mVhe
aaooqv4wSvTg9BK52Y/fGd6LY6ZGjr6Mu7eexkHJVdEQ6z6KrFqym9cI7swNj2bdzR24ocDaSqaj
/9i8a6cohcWKZZMeF11sTacOfK8kb/O9I+7YCMI12BWb/oiWasT8whXz3WphFjPgN5u1bgLzrXwc
eMN2HgAabEhMfOvGElAL3JS2yhO+tjLceKE64tvPOyPv9bOH36lkBZ5h9ubxF4p6R6eFu90POxp/
UzpVhYdmbussbpuVxrZ+ll5E4ghA3+ObHjuJaXxUwVAn411xm2gTtUH/gWzpeG2u5XxApRbOYbpf
7D5RhGhgkfbVOfb3WpeJLeLJVHIbaygBthV1Q4LTA15ehZnIlm79qBDk9e15uSh8gByKi9hOY4/B
AFUInT1dVLdIOgI3PPetl4wAqYOLHpBZqIKhfIoSuwBprMVM2PaZdYiFyQIknWqvQ5+xX9gYfRcX
VaeGkewzi5DNWVsW0eXFOW+NDMTJp3+uys0GVjbIvsR3sUtHcV+hrzlVr8d3X8xq35gbDw93j8EX
yxUlS7oJmL4UlrEdXPMPxB/3fDk8ortUGJefoaNDgk/Jf0ZQVj7yJ1Zlg1tQzUkcUqtbmiBGyY/o
T5QGm0V83osq1cbIxBUh0h8AaA+0BCjbngdwsJY5PdNTVDWH5HHVyeKUKO37R7xzbBlCJ/RYlgQV
BZze8HtV9m2a2yOqfjyw8CaA/rJikrBqMRWLotoAU17OlOiQpcXEuOqyt8f7/zhMW20GL6xmVAUj
sYWV6VImtCGIkMjNnBzzLrUC3fbOzGpjosegdhQ4AsunacJLrYsIf8xk5nK0SeewXCUwq4f3rmII
PPQqNuPw0UYW8apQQ4XOU2iidFICHgMCm4LzIxO78mTZX9BPD2c6XbJH8ujE/8IpVp7bZRhckMZW
gPqTiikj6Ulrtzzrr8zYGrlY7ywRdS4q0qH+j2PDXPv9619lrcxjX3O+h81WgG5K7TvGnmdMv4Um
gPEmzWb7w2tDUU7fKoTZtqEJPaEFfeAhYefWjkmqfC+eeX+CwOZs0s2vgZtF+oPJpLrHF5k5wRCX
txBLP4XqrkacPljd/k0EpgJ7uDDg5LOJJXDXAm5z1aqNTeOhAj89+EgPdtGAyEcDr5wes9tqpWak
+Tj3wm023+g4oGIkjjw+c8d/ACIzlFsTBBQYTHroU9MYDMiY7kael6ROePbrq8TtibT1oXBqb/52
KERz7AAG8OgvtLiu6cvVLHSRAquBnIVicoYnVbN4vsWX8LeHerbN7r7rmj1q08ffrkXheOR7zH25
OmVNFv/KUOzqcInpxnxgNqm2J6hAL65VircWYBuemVMvsThuCpMUOgVAKT4rIUPhfIQ++mFd9vQF
q7Jy+u8lHeOWvCDoQKxS+2KvzFNXho0RcLD2uOdUfrP9PB35KjzjfWT8Q+e109xCZNYsMsDFGsgp
SwyLb2qJANFU54R+hl6X2z/bQ8CKowqgej3Pr1v7KsIzGYbkoIw0NQmDFDpBcFgUJmaZGG+POEag
gtZTUKJhTm9Eiugc+gGXxj4pYqJkkuQ6giJIL0TCKed7WMUUrmhdYmA7LKgu+A9E49q/x86fjiYg
9JxtAsyas8VkLoLjBmk+Lvkm9tsgFTI2zvJHnCpC372viY4LQjeQpzaP5CtXgff0dFBx93jqdgwt
SSqEydgQRCzQoV6Fk3UWU2dMpAm8c+yUkOMVJ0Nse0ybkmKt6MpwMcOnmNo1goshekeybXX2pxll
N7G3O+uUSo/qjMvTC1FhXPSYqAEud5BRraERYQZmHGGvYawe0z9gyeLSEJO9xgwZRpI9Qd4FgjXg
EPDW6XdkchxXvsYsTwxAlUdohS7PuF+x5Jd9n+smoNtQrocvzmYY/G5FAQ2m9g6tb3sZj5hLdz7r
I18qFxo+M1Tn1Jw3DQNH1r+SDr0Ji3jrhF9fQhtHYst0Xma7tdjAUUew0wnwOuLgIcIQVcIn73nX
HhP8FjUkVA1p9ez/nYiLAxZtZDruot+9s+B8poKAOz5OdsKigb2F0eKCYm+2x0RjgL2FfuMTj5+l
D1OXQeDmTpGIj3qd2gECEbZc5Zd5+FHECL1Ab2CxnZqLKr2lK++1gvzffm8L25LkRX7DSsNa4TlZ
XoF6ondCD+ePR1FGW/Y3HwhSj89Tf4YLCwqG5qKBoNZV7/lrVZsUHpRlJRqIlypxZWnrtn18e79C
ExfkRG7B8xEK5AfGe1OAGaElXxdF6r/qZJGjp9cWsqGy483YnlU8sPxWnRR2pzhAeQQAAYWaPHQs
4dEr1h8ya+8m6mGeMstawQyQ1Ujf64nwj8Ph4AMGH9zvhDHO4gxAkPvJ4CS2N0ImyPvNi4uR2/AL
DUd03z7KQ23/HxIboL+/8P8YgYS4Lk8UM6uexgPKOYsYwY7LLA9IPvVaOD6A6qxo4Gw9KWZXAPGS
tUqGJR1HSH7bblncr6Ca8svCE5hWUeQSGaJ9hx4YdobR9ZEyzUF9SSxSIhbquMFFFnqOEJ6NW5L5
ewqEcaK8pXa0yIEn3AljedZyHDKGf0PsiC0/lxqpcoLFrZUlPSTTI3s+C2Kz1XGd0wX8XXDj7igC
Ct2m9otA/urLSzJe/3aNcvkToCD/4D146HEAfOVNYTORNZDEcHP75PM7kYGYrVEyQ8n2wqgkmZXA
QI31qBcMHg4VucygdZdlKpq6Oes/Jcrth1A63PuFgCR1LnhNMUHaZQOAbMQO7kKdFAya/EG2eT/N
O7mHQ/5MYh9fCzTkikaxNuFrXbMKE/B3k6cDwd92PVSmk3EVQjHyU6OH4bfJKp7xhGqkO8NogBpN
QcZx61/imSAlJU3jhx3pXG6fQqQMmEVGNo2ey8ICqSlx8UbymOEoi77w+i1EDeQxB273dLAgq2Qo
LixtJ2zuouSDEyOKY8tzSdlq7MHEXnV+TNbGkLz8hq93aV6E4rnJU9VLnPJKXqAHrN60uKEypQap
e3a/serGit2ZsAh4DCqTmIqZIHC/ryMYdqDl5XzKOFi2WZxHpP1XGVQrt7Z+dCvp1CSuUzadKyoU
EQ1X7m/ZK7cb8vi+PO+FZSsIEDmrwfzOeGR12f9IKj4Rn7+JvR/hJeODsote26Bc+1Jx36b3rd/A
mJvWAxKZ8aGaCvafuhzmArGfACQ4Za0Dhx0m+GUT8SEsLX23zFzuYOP1HHrUtDdFWBmSzVtULN5R
6TwQ8jM1E+7vf+zTwP92clMRTRZkMsuo3RzOGbQNR8r2815NakIf6Vrh016y9xbHCVtiNDvkxNjI
URacnq9at4ceyUyiMAiNZYJNZyyn+JWyg1a2BMlf/ZDf1R0XebNCsb0ON0C4s3MyxxESubLX+Kvy
lH6YujQkDnZhmWFodqzZwfEnRZ/z5ubyMIrwQKo1vIcoEeh6VCtBZiLcFP2V6S0DzOlQobeLqwCZ
fRS7kntWcLAeAyJj+YpAc9Xve1VaWCdCLXAsZ6MaDn931/PTAKzgXvp51/uCFiAXzROZQ8bqrGJ/
wJj8t0f+lkEmIx4hrZzuugr+KguuzqcNSud3k6WNEC4CwX280JZoR5c4yuBMA477VHmwCxpERMQi
yIrt8LCRNEhXomUFqxkssl7Dci9yS2907hf8SPQdcB8GPKTgbsBP2xLkT0Uml97GZoQpAgq+O4i1
h+XQ0En1iwhZ3Jdel8l+6ejnNLCAZApOc3xhPEncCesWYqNagnd8l5aRLF1pe4ZGQyrcLQTLJZVs
fXIUOO8ElDAGG42Ske/yQhGnyDDkk2BZRQe5j664WkPfd/WMjT/uhll4xVx0khazMdlt4oX/bF+6
LB5gbxD5PXhVYucNdsply1Q1ojvaYcnTRGeRBh66cGBtMhFgYKLfCnzJpBg7B/ZTbJtWcjeTUIdV
NvLPcPaHFbQNPG5GJs14n2z1+2ADy3eHte8cRm8Oxdrx2lCuDp2x+08iWe5hbmJ+dY1IbzUaVbZG
M/B6GcUR1BmezxwOm/EiHEwgeo64WdnR7KjKXiW9GBe5othaXztiPhEdpr7wIFYzCIapsdZRhM8S
2Ok81MVxJ4rIvGWJ8FQ7dqTY7VtojdS+5nSOmdFNUKjqdhtMCkfjFzt2L1BJ5FVNvViM9mRoXUIe
nmuk3Dp0ERy1OYgoMD0igX+CuXQQQASFB1+1zFYx68ZY9GeA6FhtJe/D1fAr8FbVWf+UozLDHbUL
HqD2Y/r8csQt9H8LBL3U1ZeD6l1us7L+hN2mgkEz4ghrDXFG83eQ2qQvG7UkOO7mj4gThIikk/Ar
blEc5KvqSiCR51kRsn6qB/4v7lwrIHhcrv6anNsLSPg0xYKp9p/X20xvWGrlTEuRRtG9j/WIb6/G
iHmpAild8iVOy3HvlQYrlDVYRc8RrmY1lLvMajL8YJ/GoMa5Ys/LUD8uy/LFVS0uSXGDyoJJuUeH
CAOh9pz4viZCwsxp5y9Lt2pjzemQ3hdJVXaURW/l7QhSOcIrdTmF7zkv0088An4lcYJVAmealElX
1lwXuwW4sa3S0/UiCu/yTK/S9Wt4RMls8p9zss8KG2WS1NWd88/DpoSUfrEITFps6T8G0lmf4QMn
Sd+4TP5eXg/XTRrLe8FG2zzuZcYeYIzVOCLUF3RF8zH8psBe2GfnnSohf1jwfCiKF7IIbpA6kmJe
dNK49FUGbow3cTlbqfqyFv8bH0YcTtTTJWHYzCPfwUD4rymGvJOv0mT3aoxid4nOlJ/VmrkpPUQr
aaXZy1UKDrNachWmPmnD11zXKfB07BFvtk9T4EXBubSA3u/shnE2xES42wu40VXMjBW4WyW1SEjG
iI1mo94ETeu2ybxniMHMQRsOBowigX4vzv+fxinp36egIAj7tPUp1mUG12ZC89OIioXsVZrPUgtx
DGMRiYV1+BeiZPtKSTnbid9qt8Xx4ZLrUrxpvorKgTZciriSX/zDGdroxxApkfbC1+8q+Yd3pjEY
oahLKL5gbrw0lgbVzyzIcUc0HVDQEw2LPk68BWJbQ9RJomgT+fvqd7YFqpyIYOoZlvqHGtIeL/J1
UPW6ZpKF0trO6xYQxnryWImLwzF97e+zQGUPYGRQwo5+H3n5g0kLGOzQCaiXdC2Kh7jgCloY2BR5
vQZfpFJIwn8wX+MpXrycgCcuROm0gD1d04SpwBcmEjopARA3qi9bFfgD1OD+0OQ5gy5M74eFqMg6
14ofuH/0bKRpSMsPXEBpTPxI2m/qWREbIY8eyUSQfiINoHHIfMISC2+gsR3wkCngbjCPO4zVRFZ8
YDCjdJfmYa2NEIzPurCupMmMQf9OTPCDGmUr466mjdwK2Byzt+DlL0hhz3lVtMlqxSUsnBM6mXiT
kr7I1VVfA0hI1KEMIYEOdwhqrWThkuQ7SUfq33BlDTqXTuDD1GM7I6jF1z8r6uT4iuy8B7emhsaU
nwIXCHr5Y+wKfgLhfuk6a4SHX5FawYSPQ8EB4vq+mTJGNr6nhmVT4eAZevosikFEbWyjsVKLyKGt
8NouBLk84dLjOaBndvkXv01TPJbgROVUTHng4B+OjdyquE9m9g9XPcSj0yFczZyPkd/9z6Yj5MlS
hleZNTWLwl29S8oxvTHmfyvzxbWZfkKxDQAVSznTTDOtGqstz4UfUOPauKIRtsWc5d8lbM8SXRIp
JNr1MdLBrp2VFHd3APYgB9uu5s98NqPUZ9i8tSP69kEeuiF3Y6fFpee66wL5fD1gfqDONPG72U5P
a4iRgYANUDK8EuMKF5wA/qLtiHwuM9Kf+Gb74cM14wpYaxpjfwgmMb8YKyEe+Pz33vApTsgIqpOH
v7oQabu0RM5L02wZyu7Ouxr6k7M8qDvuXsg5IUDOAXMauRu8upccvNAPTvFYGzBWxHy5djXMSlVy
L0FHD6o4eTvZOQc3IfPn9sNB7lKFxL638j7HztiitWlyFelPWbPq0sc4Pm2EZQ9nVTgp4ZL13JOW
J1+ubz7/nAuz9NQkG0g5JIYSrXRo0M086VQKCG7EVxtnUBMQT9ArNnCZaWjiwP/HEZB8MujoW5GN
sGaSpT/w6nJ8mB2E3dNPXlQSoiaMu0OGurM6+glZc/qabP0jd5ad2bvxuN7qTJ67NEOoa/UJAbg/
7wXLJBtBRLB40B6IWZOuAmNE307qN2PKkWdEHtIYhAWBIU1GZXsbdU+k0fJU0vpsgyHoJUxKkcXm
kq4MobdWHBvnKVHn7Xub31OO3O0hiMyCiAm98e1UQESt1IKZ1CWI5tK12QjUFi6S4dVaEGy6CC7e
3hokQbvaLQ01w+V4cPLO8GAavnGrpwLK9fElxKrR0ACsGgsnwA1LzHmxNmiVKsKfx6ho6Ev7Wa+Y
u9OewP99FJKTsAdMAaA9Z9E6/L/XbeUqYQVAXTiSQ31l+TrKmeuDbLw/jRo/53nDlk1ulkDAOqB6
i09kxL/CegY5Z7GRNXh71aGTLL+iNJAaGa++Evr09246M7EtemgSs2MfUL3st/qisFX6xBjwy/Wv
Qg87pDSyebRZEPXVSkP2+1fEnkFzX6vi/Cnbr5PRnMyFoV2DM9835kgKA17zBJiT15YaIG+gWt1B
nuF2fa77k6L1J68mYvdIcBApxfchgHui1FEhg1TeaXSMQnuLhUS88HcjoHRSgxZwB5iN3LwmX0zB
R9n3R2uJHQhJcnREoG7RUIoEOH7Yol+W06ZyEgVsKvnTbbul54zC7E/U82BHrx3unr2MCPaoQdQQ
swB9XOXNVX78kkXVxjhpgZqtR3GSs6yikWyPzHQt7n7iYFVzKAOosytGTxkCbjerarFKbnIhKNL5
BV5Xxl4SA2zbqbS4NFiuYQYy7KwwG+wfX9x3SSYvRejDIPbpj35OublWq5QFDiguhm2gpwzmwD69
klMfaZ9F/hYWBLtot5+95ikTt+5Z2Ax/R1i6IcfVw5Y3Oo6JSXM039n66rx9iswpgpI/1TgbEhpm
3fFR2uC6UVGSYXH8NWJQD2D2UQ1eU8adRQMNQbPAcyW2Nrr04A0dqKTZUWT40RhyXVGi/pHTKbY0
vkkf45CShoQ8sSh2HA7oSCjDOpJj2MVFEUJEXIZaBPbjSPS1nwois7yRRtFkQm8rKoxAMBPftYN7
DMbV1q6qFOhMozf8C32dbMA9blZOGIMlNGBZ3nFuiCLSb2kgqJG3kzJT0ySRjWouqLdvE9FpBjfz
hkbZzQ/V2oHAZ8AKTGGbdafC2LRGqBW2rqVGewY4GrlURCEggL05ZfNr+8R2oeSOBO/7mgR2YwOi
owb6fk8nj1in1o4v/qQ8gOPxGl+jlOY9ecTHhy3wLCg/e8zcEqWIRL0vC8YMMQlHeFScWYstUzAT
OCU0lAeb6jJBCe2MJa7emguC4fAKiAZTL0bUXdBp/UT2VHyT8zlnGx+QuPR7NsyM0kLlhI2LPCAS
pXclyVP/7FpZm2Pe0oQEIhAh8mLvAafGrr7ke0bEuLxW0dbRh+1wM1UXGOTNk9OZqnByNNgMNoCL
1y8ti6BUy33ntIPSQ8Qvckb6DPVJdHKxRn5NDImxp5JfePNUedKRxtXCspuCnE70xyOqXzyL2VIq
a6ZO3G04EfgoQ5gL8Kt5YyxdOVDSQP0ZZ16077ILuo9vLJSk9gQTTz4+H7DFc06//BRU5FQpNJrv
7DdhVpoO9dEUxZ57qqxaWb9roze33UT56K57SEBT4bmf4r4QZJ+yWNQNLRZUcMrvJM9sx2DOPScY
cU6vkYWXdaiPP5WmRo0qAZaJelQ4YEQ98I3rd21hbD6XfvJPe+NRcix4o1Lc721/ekjVNt7ukyF2
1n+6KVJd0qnhDP8pTU1T/iskstGU3+eVl0ns3PQlxzGjLHuqNvP1aR+65N144nKLHgf+FAMsJUDW
/RBEF02UYQgupWtx8oCXyo4TrDWSAYQKKl9m6vS3v0d97yTtYtEqeu4A11qjdYLWyNnkqxbbNgqz
9pD9X01DSbsaBfiso6T+5Dr/PdFXSDU2GonFJ/G4MCseFG78Xsx/x1Kr/VEgCViVKpf1CuF2XKJO
jVP1EPWn4D6T+LNUYT+dy8aB833jy+/vaqxPNnqaO/63xdngogb2IBKIzcT54SxfCfkofhjHXZIB
p2sjqMrzr54P4dS/nNzRGuDGo2iSaXpsw1lsg28aa86wif4Wx9V+VzwKZNCK+Af8LE4f+42Un2dj
ZNvbiG69P+VzBPmwqd/r6nq6lcVwXeLfr8qadYgHrmHrM9IeVxq7bYGzrIBI4gAjvSGMrRAU1elk
g24PY/73U16ib+TcjaPkY3VxfUw2xNXHi/5J04tNqz7VaGrgANZ+LTVk+wQAHloiMwgQA2Aekuf2
zevHKnQEpmmnzqAKLd3AQJat93rEWLCCt1/NyUuDqoZ6IJgNX+J0YGqGvEhVBo2j4bdKqFtDEI6l
lkhyFc2xmZKsvM3KSLXv/2M6OH2FKUKxZEkVkxrJlfJDEpBmyueOxyyLv3xS/+Q+CCbJbYz39/Oe
giVvRZsVi2IkAPn0+KlOm1V3+XfgFakVPgmZI99OWH8rix55/253zfUsLgxFedode/8cM9JMI82+
/M0CmRl3fHIkHpf2C3PKehLE+K2lx8Bk+HMCBR7ThY2TTdfl6qvDoQQx0YJHeuQMqNk2zIczZvJU
3Q54Q2SX//cj5qSUk5irQd0Dn72Op5j5CK9hyOLLRo9+H79Muv25nAcAk58mOeVrJQMZQ5/DZyKD
aTRAbqqUZSmALqsZcTPy4gMOXI8JWlG7VOzY2pPnZV2E7U9g4ciJVMAtOAvcAISfLIOUJ00Wt1u1
R0eAQF0Vz5XXaGDdDl8m3b25Wj6+1ZbClG73vgewkX1HA07jQVHKa0O8dsjTapJy30XD84p8Xg03
7nMvOJDu5uLieaO1MVblZ70jOnIa15XACv74hKHi4uX9Qv2ddv5Z7XFLNMEjqOtmYbtAlGycUc+S
JYqv6EYRJP/wGdY3dIfOp+GW9iZ9SZgiEqzwmmJ8dzCNs88Qlh4tDGdeUUrLLHA3DEfIECdAkxG1
Cs0NHQxXuQ4cWFx6dgiB8eZt3qReO5ETLfYDowjQFSpfQl5MNEvmoFOAFOMD6y6WXQJhHHStxGkH
idnlTUxPDDRdnZNqX8gOARoLXgqvwvX+qp1ZvSwAPqJOtXQQDiG7FqYgoB9kOBoOuwtgIja/Cl2O
q8QXJ0cTQ56jhDPiGp5QkdiT6YmIbn40yjyp9De9PhzZ7j/CohfWJ6TbNyy9HsJtpw5F540c0OWP
bSFkV1bA5Nrx2LK6rtb3cqrTilW+Lvr4vQSErzWrsnsS0JjZmPw16uyaOckFPVAeNm72Q4iR9ZFR
/BOX/nQrcVqa4f5KzCegqzsb8+pXBix+qU2uULZjjdiT1HHLbt7jSr9GAd0/nVt0Qxl9xmoX9GDK
p4xuhaz81AkAXwNbMaECrz9GJ/XgX0ZpqvZQ3wx2bjxrLHbA2LKoYUn2thQnYb+spejUSH0at/IG
m5xVVOrvtP/5XG3LLPmANI0qt6RyVmFugqKrnx7Gzzs7ryx11G77dwP+ZUqOLMGX7vyrlJaXzv6T
Gcla1E14LgtHffaKP2M77kL2NK9mX1tl/LSYg+fsUSAni91SvQD2ry6EXVgAVIHClPFGFVKJwzXZ
fSqJnL2rFwoUOmz47bqg/0jW3osassk3xzuvGxu8u9+uDaoftGY9+TRbKLynw385ClUlhm4tq+yq
JLKAio/eftngUtnlwMYbpjmeh2yRzqUXQ4HiAQaX+l3YgVgHJJI1tJqh36+91uP8ruovYMSPIxrG
TzgymlJPsYtoYLAj1wADbHb9ZqYWuJELr0XSCr6iLwHIIuIgQl0UEMbjOpkkp9kk3itzO/ClfXsb
vCemSTE4n50dbjUk4S3ND5Rd1zWbnVJsqJVBPneF4GXDUscCwJ/807j8BtjlOYotOsAuL/l4WWm9
JaVNkpzHEDO7GY2NuUAjktvGvyt2TOjVRtsP+9oN0+X/LHg4FHAc+mAAfZVQUnfDpLmP543zn6MH
qTYrOHoZKjVrN2kpKdygU0vd9f7DASxfK0esZqC0STnmUbGpqoPNYobIL1loTVL3/BcySlll+3Mg
V1XRvGZh0CC7WktOrcjx301WJMXCt7sFAse4HGPjWr4dyA+A1NtxpiJU3GH8ePp5NNQNApTHcNj2
Py8rXw7UYnSlh89obW7Hf5JVJ+oF3IewjoFH8YUxrMp8tikWb1P8gISWe8yMbtO6zWE3s3G+vBbA
ydHnhGOF+5gqDV4FV5xO7u3BPF4dFK/Ara2uim0UpJuQ6J50/tKhwu0wmIqbvQesaQ30tnSheapJ
vgwNgdWjNWZv2RopVI22ujiJZe1KbhOAy3GYQHqIbtBXKXChCZpg86zBW6T0Ui0N2/UNVu/gFsbW
i5xGAktq58Z5bzyKD+41Y+izRAD10BptI/TY1KhfQ2dypIi210lyyjLRaKvs4BmRW5+6XK3etJMV
s+/6EIm/I62PORsYAoU7fVGTYTBlAQuMIDc6M4l1J7YCTBqZHoKKV3aw5Ta1ZORO+WYa8Avb0Tb2
kxtdvx+iR7y9tjQyVdDFkT2KuVG2Xs229XX+/p9/+n2J/jiH8jDNkKaLL+6Ljl0wL5V1AwXL5u/Q
AVJZ8DiS6RhF7UWPwPBdWYY7ayiixYh6xbYYCzmDbySxaLdUNiX62UCXxvT/mOC9M5oXkOlMBy/J
LB9zbgTqbq+JKxX2y2KRpkpcgka0Sz1rhs6CBnjH+nbtiOFW/M0lS2JKP/yguBTnJjERNcO4Ykdb
FgE83tx304+XNhUGf+yYRg6RC+o6VjanGpINet9cHRSSC4aWB+IfETAzIlv8R10SVFc7TtjuLf4/
bem8cLRTUYniDhIwTuwcJc34BiQXzD4rrx/9eYHuKPCASWJ3Al1VeU498AkG3TtxnZoSpo1cTIo2
w4/xIjBirXpy9ifYgfq8ZfzUHfcY5kh9wdxrTmhUzwXLA7xG7CMn7Ft9/SDgqLzBmxIdLbPS5AaQ
G7FtgHU9ax6M+56Z3H7iUyJSJ6/B1yEvRmPfA6I9L6jcZBc/fmqEQ0H00ODo2eL94HW/bnfAWQQ7
NvrCvkytRAxIGKjrL9uIeSQyY9N/3IDOTYdCutxIc3KTEgqSbQsq1H2uKEwL3zgLZ6AIrYEg+X3D
xkw8rnxCi1zTdNn820diuV73AgIsWz4p6r+hxmQJ6xYkQuq3oxQSaxXWY2VYT7iNRUSBW5iG91Fl
XDEukUtMJJtDieGcXvNVqjiFfq81qMV5YiX3AkxMq4S1AKESvZBLbbhaF3eNy3mRsoYjgpjDICya
LzFFdSLIRrEV8FpsDAGnMNe4nZtwiqZWxsMvGGVZZ/ZBwr5hfcnwU5JPpakvXEEg+WircJzPoTfb
SXWFWHoJXjuQP56aYgfyGpspUf1hxq7Om3JNfrgR9Qn5g7nI6aCYsiijLTq/j/4pFtYEZBNzydUq
RXw2K1EjgSx+nfpwqzBhTTq1GET20tF1z7ZjrYvxodUGwwDqFMQxl1otqoybREcVRXrq83iRaIit
DwpUWemvJyYcXN37miU82fL8jEYTaZXUBPjYaRUK/wifC4nCYHsyjv6zCuEmxB/skLY0W74TdFVY
Rat4uyaA/svGPPvk4BLQKXun99/m/P5HdTgsip4hvs5OW1fN5w0zIq5097mwhHXlVN4T/EuHsz+x
r3Wpe/j5Qbi+cB6jcTmsmMju8e9+kcYqeWLkx1Z1FDTQwye4xkv3PM5YbG9en7PhNIywQjGfuML+
YCl6X3ZtkaR0PdTumrPO/ULj12CMWJlo+a3KfMz+JpSKE665YJetGxTJqi/k3YKBPJxqehiK37WU
VZ7I/NmS5G8B/GzwN3nQhCr9VkKDWcbuTgeiLQDMpNs9IyyLHgD9sdrNb8raC9zhF6g3RvKfIsSO
BghS8RZCGlgYmchZJzWUmNlC9Rv41t8K/w+e9EF8Qxh+DcL7kwhOOtBajDf6/cARBDC0PoEtJhQI
lEwSX9ybu0+goBaLjEMSbdtok5ulYXGpfjKfM6TRDjvF4hPxBrVrl+XvKTiy+gMNAcL8iQJUQaug
bMzM9Iz+cbLnkTwMcF3PEp2fPRjYu36xAQdBrP2Bgg0wCYKV8rjwlILHSuoqPlKsF7aGldS+nAZ8
7p1vFIAEAIHfJHbzu4E/g8I2ZkL7vPOxLsIqdw8GBXhDL8rn8gixdSJoX49zEW+T8luqHeu/SGd5
FpS5/4Z9bWwiopes+y33SYdz+nL/UjcBLX0V49WkfKgHrqRVWtTiLBuaioBxuz4eQWM+9ezjQEiZ
fKNhxfnyIr5r/GenI+xDQqfLnv/c0Dum3lQSq1XkYmkJ4Kty4e/7uXktF+L4EhHysQaSAuCHzYyL
InduVVlUmQ3yj6/El7biq25gWtEgPsivwhQJS7UyYwppvFPiubSIs3dVNC+hAPO07ze2/2ZyJ+xb
6vhd6MMzJ9/fqk9iQ73X/Dd+t37v1Ulyn0sKb0YO5HXgc4opsNeoBU5M598vOYNqLDnr+nA6Qx5d
uGEwQntrKnxdscbM9/Vbgyn5BnY5QyAPg2pbNg8jGT+l1F5zGi9dBXFJyR1mxwtxErAmM7n5mGPS
IeuEsmVmEEeL2ALfatblNPGTz2wImEEQYk1rLHociVcCBuq6TmT35d/EjjDQEQ0IffMddQxq89fQ
lSxMHQV+nGtKh+NkkOqf5RtJ3YQs1YALKssQXkb9bhcNyH98kfMWzvELMwulWxcqTjowjgyLe4xQ
eOMud+kyFo5YsqhAS+ZKRI7BKRmh2ktiXJrcrhaLVExcjVnpdTS2TkzqRs56byBLpEjpnMCyzUDV
iNEDdCod60AgLOswTuWzmITh7GBShe9sRoMQbk16lU7MCR9+u77CXyrE3wjbqXYPg/LUIz1a1l58
+m/q8EUW/symbzbc1pM9gZHtaQoQhdvIwzB//kqOxyS367u6YiSnd9lH1/gg8z2ylEM8b8UZw79v
dTWV756B0De6Nu5Hkp2+3UFx6RAhwMmP373T8CuTXTkaK/umcQgmuLKK5cLHyu3F5dP4v9scX68t
OfC/XDYJZgFzzlLCOD5dw6XKeYvlc5QCQ8Gwow2RsxGlQoRHTdPTBHKYhQ49pXDYkaIrosXHPDJ7
BAekkxOOt+04j+aAWXFT5FxmEWDQgQmJ7x0l0al8B1PCDZo7o36veynb8c+7WPUiX7TnJ+fgDuZL
FzJjMOjTaoT7hWPFFFL9nEhN5/sgtUJu5bV81qHtIhK3zK7iXTWF2j9s08Eu2jAL6Ww6u3bzRO3h
AfCBSud6pLtrQ1Kt8t0YWEB8IZMaLrp7N6Wk9ezo3P2161wBu/FfkmgRXYprbMEpGow5+O8ugN/p
9rokPeEiy845f3x7n/l5RUpLgVl6jcHN43v2NukBrpAaoKuDeyFFYO/slLQHt92gRKqIlFIfcLXQ
WEANdYAybNVnrXqN3f8EV3kA2RcEWOtzzWavzY2ecfU/pUYnKVsip2qYOtIhAmzGUWn3jf3MKJZa
du0Qw++6Cs5HLr+Nz4fpQ726vOzMmVSrjjvlhpSBZwJwi3/YG3dgn0ewI4Z5HoCL32rDQyT0QJCL
esjZeNgpopO71CwYL6nsNykX3v4eBRrqtV+go8YjoecYlLjb3RnEBBUEYfJ8Psg8BOQvtsggR8Vt
0AC+U26AVSBgfSAIU+3hFYQ5b2Tn6BQ8d+D1JXfYdJAsqTV14PG7+oUntPVWIzpmz8CdePH2wN2F
qma34OdwN0UmtYW0x0nPPuX2DL8Zh/VaUXSAYytVGTCpERCylISabxEGq00i0YJv7K0unPXxVMKh
8IP4zXIb1hTwr8Qo7pnB46XFoQx7kN7zLLagYTpCAD+efuUx6mlYLfAnLnHs3rYHiXSQjOvOeKLE
2kRezlmg439Z+eJ4WDkaowexnWwbkLMXPRQ4q+fJVtxYSww9vM3LX8glkCY/6KImGOAisWcr79kq
iIz6FpZRIiIG4MTI8JzC2zRE/aPKd9IWSxOeVNyIF8+7ZU5UxKiOJg83QTL5nsKlH2ntV1A4jmDR
klq91li/d7NZ4uPKOUUQnDyG4Q605v8Vh4hJfW5O1tE6ITSewrSK+uabnADXQZBD4ldledh2kBSA
omYz9Ke5j/Zz3oHk6O74a3jNnqCAudKEYjAmKpUW+MiDbrDNjFhBiEWgyElVx9Sj0GcsVO8uk19r
WAsqrnLhOZDAWqy+OJFwYuBw3vW4TnhVDhPpi9Zg7NlOF5Zr1CLWhmpRhsV5lDHHtyIBee7tbGeI
UluSqv2ycON6rGFzbHJeb4kgZIUaM30Pu7XPrYuYGt2z6b03kM3WHqzGSC0od9OKxLnmsIZFGZBi
EV+dw8c4PO3YuVZf24kdUqQ2oKh8xiMJxpzZV31KLN4ghA58RXxiN0EyRQQk3xrnv1zsXhnvcvyU
umaG/zLy8xaA0bNBzV/omx8yB28Zilqtfh9Igp3LvxfpfF3y09pv2yN0chK1a8fnJz6S+lwax5C0
G8FW9s/kL3zYdlsvS94aHIwCvRkHXjl890fYJmYSFIbMQEOONt48yDdRK/lp5X08pwX+OycwiYWn
o5eISdX7B7LGs7VKU6BClm1p46kPcxgUeAUtUxV0pw6+GhqUeXz1NwqmgigOiWmP4ZqOf8TVK5uP
fWWXd4BFEMsEcT6PkzrUVsAhzdFlsMonlP2xKD93EcK3ek5Oojh4FNWRapNuWthjGU+Hk6WouTQU
pa+H8a+yWw8Ep4EhtFf6eYRrS79MdrAHm91DfkdVRzWYUcZZsUcjZWHG6OShIFnXpKA/L+VOO1NK
ZzBq0VGaYJ+pDJvtRiIF3y9U0aU3D1++UjAvDHOWuobA5X9+Hre9tN570JCv9JTjPwG1m6eu0iJ+
OQ1Nr2MwCk9CG/jvdALD7OWiOoUplf8Eiyrog+nhmOn0FnpY1lfjMIaqCxOufIW9Wg5mjNNirSFP
p3BMpKcCBwV4hxvpxeL784OkiigKQUDYJV3BiONk7KBajMk3E5AVPDkTpwqk0YZTmddLVCuwnVMG
fQABp9VNO5UbSY4cG8MBbxwfCA0yATE0DM1zqit75Fu85Cb2binw5fdEesKHbCu/O5aAZn2aeUY6
aii7wnnzfvOdLtHY7ulm/QDcTxuVO/5FPnYdiGgqwr9aGaKH/D1pcEh+i/idW42iEEoF6wVbzCyt
hHJYAMDa2XJo2pPimKuiq3DQJ1cuXiGLjHELzznHIYC2IS1caVk3yoQW54+4iLrNxHYoGbVRzhz3
dZEp8zcNGd7WvIgkQjRZXgFhp6gMR4FaA6WrCrTTaAT4u18PRG6LRtuhrnYICdap6kPnrTVodu2r
p7YLJH3O5uBH+kTEb02k4+olSED949scwJiKTv1pjgyXhKM3GgP/B26P0WQFMlRzrx2un/9Ym2K0
Z0ApgrpGOxMOD/ycJ0zMm/nxaIRhTPhtzu6I+uNNhnC9/ms5yGD47MPqn20sDEqBg/tdiEx3SXXB
0SkK/wYNiXrFxf/wOZ/towrsQqGHBiTuRiKnlu1cxfIWY52/ScPDkUKTuKQDiaMqxAKY2xBNnt0E
awDhCy7uXYxyAQb6jjM4Pso550uMfq4ZFZU1gHpyOPJAt3ZRyGpuSeT5Hz51uLSPQerzGEcbY4r8
4uo4bO1ovvBuYdNz7yz+Jwkh17uHYuTbLhkUZmStb0vXrGrqXwOm+AZI6wEZU48cp/5RDZ1W43JY
q3IdQju0HpInnCeQqh2d+76wE47U5ALe22r4MEGxYOyy+qLRzY14D6aIRPhZnTAnyeeHJ2jANKon
qleFmXoKMcR1Z6wUrjE9qlZT49V13uuIEHqNVO/ZeAam+jJvLGyOolQMjlowY4tDQu4IzV60fZ6W
8ZHq+Lsa0uaB8GztB4RC/DNFJKIzdCRdkn2cwTD2j2BTS7bvvAx9v+u0C4pXO/VwuSYNQ+nj/CT4
Jci1dhVcOR3fCXF5FI1rCgIA3FB/pVjaCNrNUK4QpnXDdZ44EQOWG4VosUOQRBLTPvmc0SuI+jjL
Sr6Sd5UCih8E+GSKWtwvTavBFaCU7Ug6VqUaeLnFyGc9omHbGhfE3sI7Zg9P+vTAN55qZBMGDbQA
cYzibP+0OYfXpnZU79EmfMGRM5t5RTZ8IYlQWFwQTPD/U5EgEqL/FCh9HM3vaGZgKUsaVXzJsUPV
Qqx54wccIb7mfrxxmCS/P2453hTKSRWUX0pGEocRS2Ktk4GVGv0yU9RkOrk/07AgAzDuJaJp6N0Z
3tbI9Cb3nVC5FSDAMB7lFIGZfzj9xjFULcxRxt3Xqktb5Vdd8V4JAhyKJAppJMyYhzryAPgLIq3d
5SSsKAwsupePLcoJg0PijulVuRR2bNk9fhAJGLmPKGv4M07GnkTVPbhe3nOdxO8IF4ofJJUVCisW
LZ8SmHVAm0RQm62zmX64OcM5JM2oK/gESVwq/O3bkrKsvph5k+zdT4oeJnSf5GHsy5qWwxVK46Sc
XP6EkEcihrBqDe0YLErCsxaT7Ms9lqk6yQiaRUR7NkQOHOEHsUKRvJLh6qypPfJDjla195/0Ov24
mVsnASuGfWiucCgN/E79vqA3nzm3rVVpGmoQU3mmb/AfbinhgYtHgjVNqsu2KLydk1APxZ+9Uiw6
o641ry5ihPiqi51WDNzJY6U/kNaHY6Oi1Ii53NolHqL+DumZJmpnwBepcmVsggYOvYZuQCsX4BwS
vk+VezlRZnbTxGOLqGtrISvag4RFl/T8tld3sKTADNGBH+mHHHugZQBAUr2M4cG5vkEGrdkFnWhV
+gQ5moUWZJSUSs1VQgWc8BD1yAT3KHs+pZQphEnfdG1zGgiuv9jqNvI+twDqwrmPbLV0rvxd7S7P
xzskszR4FoJHwhVho2Sa7f25sJGiL2wUht4eEtSLJs6OOM1hTO0eLr4gpL0ezV5c8vS5lJQydbgp
db7jXczerIPQMR34/eOepzjuGz1CamewS04FB6A3vnjKsE+wiDTE+nbWw4RCHe193YpRh56NKUso
Vvsk5UL2zSmlUOANnnk3dxRUAKF3L45X16+EBDDGYxq796QaqnMH20S8DwuLpZi65nrfnkoBtX69
HlTxkEEvq5aD1r5y47VbgTtMCxOnOmwNbasaWTv+CYSCmtKyneZavLoVeQnQpfHLpw8ZIV/yVpKI
b71D0E1HFo8vdOVsVcjhgSE0wPFbukSd9j3zhQid76z3lOfBE6gy7xR3WRACL5ljs5C7QdZ/wxyv
gy+MwuROINkRkPe/jRBpezCM4Mjw5i5882C3KnmvUIPFxLE+/ul4kE8KHRc/nJOpeZKB7RpwbOAJ
65Z30AmbgFQ4FiTgGkYxFQWfc0otnKgevzEM7g+sKNrz+pqdXqlFRYpmWNKLO0MU6mtBRlf/r04Y
XF2/LFFhJYwtqHkpKOHtWDFdYnIk1uAxRHS9FktfcsRJQfHqN0daNDPi8uQW6ljScL9WHKqnoAzL
yko7hJJKg8TRgXfLPrYX3lolb5Blw8wq03+4toqXxPd5Zqpql2NZylv6uP9dYZgj+OlrVpQgGAZg
/fOLmOYS0HUaLA+7Kta+TDrfsMPcgY9TJNUZlQ4+rdqoaZIlsJc53jS7QHA6nTAa05q42Ij4m5Ub
lpErqkccwvaCf1qqLBefNdct6g9qygERxUSlsd85o3pBaOdp8SDOE/MAXGKs8lmmyym+nImQRWGU
cg17E13YIAZrFq7VFoHGWvG31kEOPayfW+ERscNJOtFIaIxdR4DkoQ1FIf4M0xds1hp2rBIB7YB5
olf8f4lOKpIxEehMN5kWSnos1sLilhvmkUCnLzwNBYeTVsUIkZEQN3T+LKt1/mEpDQkxbtT1VH5K
TfNI4xWvZWCFRxgwnS7CAvriu9Y8jBFUcnnfNea7imVKDSZ5tzHeiKMMO9giS44f2zQ87uKYmBUm
KUbPUJbPfIc+1o4ZCuXKn/NPp98W+inlSQ6TmcDZ7fn9tT4wscO3UOET2PZOs3DemGUi+JC2GC0h
Yk/m1xF/ROlBUu1HRKDFvKKb7juihaK1inr/jQ+zgnmfJt47ZZVbYNjn215PY1FHByP7b9BgL9tb
IBhkUyNEk1rg/lYppJBmUaoDn93iDsnVbFpvLfOzBp+DgdwJUpY7Rgrwny06RJUYtBnevlVwLOCI
gn6l/9vAtHNVIFWM+MKXzSxDHd7/vr60Qlpi4IbXw1XC943hm07NREw8nHuJAyeyis6vnmaW6+4Y
DLsoDfRiysvjHszjIdMC5GBPChpsf43XtLRame22iL6j4/ilRRMNf0YUc2AjFbYwEDYMH+cm9x/D
7ekTCpvhC6/DDAuaDfVrEKZGvVFAnu9o3TPb47MUcnkKJaJprMGKpp3lydNzF7XOz/cOoFGLA3Nd
A9ExuHJdxLBQ8dIxOlfdGa/6gvWr0oviEZHRoAUHJ0arUQ5vvkHZj0Uek6LUjOI/7TnDhyX6lGme
g1KnKe7wS3kDKd/+puN9sWxl1c8UXE6LYuATs70IUOindV3RGjnWQM4Prxlva/yLuFk4afEGaboG
S5+veQiI4ZRsrGoKWxlTK4gCpamftRvtd0pWHzAHeQxiTVotl3BGUKHpDCnf69RO3yukkBY+7OUQ
ZiZlZkQnQaS2T9q1VczZjw7FI3T74Fzi6kKVtVptKCZm++rmWuqVIwh+NWBE4I7YuxHNA0/DphZL
vUf4BcDatF0NZaiZOGzlv7dw2VsY15XDPui947c5yZRiCPH/ax15PsB5JHYsjP1QtOM2NU6Xq8S1
J8MknbeoyPo8pitW7lWTKgzPZknnMtAHlHf2nvKyqfeKkgkxWJVnH51wyCnVqQDf5c/Z8EA33477
RLzoPqUqOQsVLpEoHjTjKzg4D5ndHHcRHTuoV0IZoZDWFdhk8zbbfWFrwp5fqjoZtP9kuhJZT/K4
R0amlpynq9vGcO/CKMC4G9zdhrHpj64e14L7xFFh7Z6/nILY7D58uH3I8E7KOBRyg0N6gbG/HQwl
CPyzcmCy7Z2iiU05hF5w1Jv8CpIB47jBeDZwcPchHRzqjOqMk2+Zvn51bIesstSRsdsGKlOp+Wiq
iabaW2g0yKDBmNhi+Ep2OWP11BJD+ypgBQ5rntisygBV4JUrODlGfhNKxyPdW6XLgdOtAtvRaOP6
IZRvNjhdH/ayQbrs1QzsAUSEpWZTGElGUThVsuAG5txtCooY81nDLYdGO+DLYbqAahtUcKPkvzdR
6hWc+SjEiszxr9khjOdJx/+a0TapCfz0xCPSlGjwUfyPTGBqx0RWjR9tUk7an7ppHKMIp64wue5q
FNzHzrH7JHJ1IGksKz0ivMIKhnpRyCMGCjoIgbZBEKdVu/Hp/jhT0ksTehNtgw/6CV+SVmFktPt2
w4haD723G14HsohSVlEHBSa0d9Su6cqu4tdg9zTIKZKrrQS7IyRctzilwh80IHgc8JdpoYxoXe2Z
I3zUx30a4E3B6Ad+1jGa40TIXZVC4GYgERamAX3A7wMAEhKCzmjYF4/K/EPbAR/uIORf7X6V/NU0
ZHakLCXVw1a2xrk9CzTI6agfTPPjkGTYVzXb/y0LV2UNdbdl6K2mRPKqxxAnKm+wvW9SqSSJEUrq
7dr1Hx+rb8VMqCXFMmLPAN9vkppSoyftIWHS8iwSt6GGByRvEkHo5MfxShP9EBq/rvcCPrvsq1Hn
ThsY16l7etz8hvDFfU/iHrdz3XNCGDmzz/ovwFLRXTIzmF0WnUpgakVn3PqVNAwGnImBS7vLK87y
p34kS2kRaXPBf79qKe4W4wyF4rshIviOCAFdHGaVi1ui1aVD6t10Ky4atcFrufS6HTQgYwBlOjlQ
HJMqavLf6LduETBGmHQO+Hz2HdDEPHc9kYzUwXntQg/FNfCwOHXFBs47ovPt8z/Wk6FrDsnhT65p
c4eOOIVig+U6ZfMQmlfed9Wej545Ha2sm7rSGZrAlWfnFNU5HjJ4jsBNDitTBkSu3VRuvJPOk4YB
LGqI4FT5SbuHlFHR4sFZBuOKYbAQk2UziF2pYTZ922zmUNyIrPlrHSqlcdGGn1D/CO4J3UyFhSjb
pyOY+kCejZvSDuUyfExsLcIvBN7rWaSgonrzwnN1yuI6dz4tic0SZQvg0G6bilVkPIe2qdnSySah
NaYrPR9eEThRwpRjULAx054fjYzc5Zjdp10xGE32Y00CGDxq6Sv85euZ+QTy+HTTms4BNVjGMYka
wd1bWhJ2mP2MOBTRBAhtawg05WHSGCOHe8GyEL/9lzKfR2gRgk83alA4BgqIDuQCj07buEL7QeUu
FghCfeJnf3hVY17YSXD2GejktFSLrss/CqBKLzdU9XdHnFZixFGqmF6C6vHcMHS/VelfjdzN+Xus
cbjNgbyBLgPBIEj1giUf+6lmnpINV0wHT5REIX+PTzGQudH8ZId23piuL2Rc/71Y6w/q8ZOSTzI8
oFlmSAb4aO0Lp4nXovIiBTTZ6GZuTUvdWIGqFtLTDOzMG+ouD/AHHSlN8ZbTMDuTrbqRZVov2cVT
DcqUU1FvfnhiEzZOVLVYVehFZfpoDSGk+nkTFuE22sMFPjsimTZj9097KYfwzY+/2hrjsFXSe1Sl
Y1YIJKnN1ZzolxoJOdsRsmZmAz7S7iKp6m0zHfASvACyITwX1o33irnx+K/hRQKDfn3kTKFjSPfR
bqW2CHwwpL8+7gV/birjMGp/u4Affl1Vs/XIKvMbbj8/cf+prO6B2IfVLo0arsfk/DEDeBtNCvc2
68meA5Qi3VQHXRSo/DcMVtinMWpg8MGmEM4JmP9FTaFr0KL5rxdiDGU7aXlB1qTm9r80mio8+0hO
m1RsacII8Je/lmVPGO6fvssOFsF8pgdxH1oSRAV4ljrlu9iVqXxzaJBgwAK+297ZtkyXLxGh5C6j
WqcEyjdDee7fOGmdgwEsO5fGgPPJPsL5ZXc2EwBCrwWMnAtoDdZcWXXsh65uu2ZHzI0AQkXndAZ/
AUnLpc+FEyk/NGwojOKwVeJzhLcjoUT0SYiJ3L1BdABjEM98sQojlxuqPqkDLn8uIaN+pwSg3oUk
z8VPIZqj37pUGu33rO1M802CtDBmFrl5RrTORwddyvu58+QIjuttuXZ/AHVVPIZ3a4AYvlqhOHGa
yyJjWr0oT/dSdy9/PtL0tyxk0AThbfE0y3FjIbSTaYG1aXlOKs4hZyKvv+gjiLJ8IViEtYsxQ27I
SIi4vth2gshS+cOkUVfGDQJJPGUancGI/k3zuv+iCHNW/8bGSngrDOLsB0ASeEqh7/OjFJLsoT9F
HwdEhpQQmTofVY9smfMlo+ib5ioWuFJvgAApK2SCZBfNX8HowaHHfoo+CgFyFD3B3Tu+M8eeWD2p
EpSMhTdv2mgjmOanrV4DS5nR3+fj8lgLik5VREJ0NOZZj/JSQIwBxEVwtQo1HBethPtpO2s+eLle
lCwlszIvG9skiRS/xgAfzzfoIMmiXPpMamv2ZquBCo0KhHfTuxWPBgpiDJ8nJjbDXCU9BwqkWpbh
+yVZ3zGa9DcefDhVw7UCsT1VeS10l+1+YLEAkVJluZNJG2eMgnPNweaJ0lRXX3OcNJkgzXp3ODjt
m9O/THmqnChwopjKo6ET54S/P1hvol60Qqd9wP2EYS3WlRrP9XeqMf5t3HESJEkLiCCwII5oHJC+
fR+qL9rr9rOc6rWoUI19qFRUTOCEuSFfTou73geF2/d+f1Kv+qbt83hhZyrvQK6/+aO/D0yMeR40
+bw2ZwBO2WsTtWDOVLRS5fJx0qm43840CLDQgWT++I1jvSPqTLHW5KC1GbkibQbX81eWNwNusA3P
B36ga5C7W6Qpz4b+O39u4ju+m4Jr+zS/SXqkY6veQioCQMArK68Hmxvqvks+5bCd3U9qgPUw2M4A
DZbB+F63whkUuXhxUnv+NdycqMs9XVv6GIewJnM3VNOPoi+8Z/OnuJQ4nZF1WLgtjm/6ziTnnkju
TIw3MVxAIKiW+wI0vx0M6wl4MBmBUPBz0+d+HvxGGTF4WVwDFDDg394zR7R63p9VYNhDrbACKhS5
nL2ELGSMfem4MUr8luGISnkq3haY0NwPyGWefWMcYiG1vvMAhA8idLTuwnb0xG5AzaDiGoacCMXI
4D+q1gInHxpqySJ+6kbyO8il6n6bcM2DXxvdTDRSIKRW7kQYbl8Yghj84ZBMIduWxRLnRdxtysDT
KUTDquOq8xxk1JyPTYSZ8uI+39OHvSPhF/fBTafysjAGwMskWOssk5dizZvTiP/wDQwrJZBUduax
8MtRZnCw4oR/8Pt4emQ8u/Nrx1gHlHqI0o0RjTQhEZxRjGRjTVM8PqFg/Vuvap+1DAlonVSbLO05
gRh40TH30EfD2w9dC+I5ZD1kY4dtYPgVLKlL/VAGCg/Y58QUJ6kmf5txoWeOIkDBDt/Ybmyjojzo
Nbiz9M7kUhIqOA8RC3hHOE5IvY3fSdEEyIh2cVLRbF3zz2b53wRaglEX/jzZr1dSgLlKfX9iTWmS
P5UY1abC5CfcospYEH/uN9oW7URxLtFMV2t0FCH4/NcSKz/0tnA92JnLTI1bI6csRVegT9ZOtMVP
RFfCiexOYrYwVTj76GsFgslmjXaVRIYlANcHIE/ttpokJpmO5dIIlpD+TAP8y44hP0piKVGoZjJb
7ymDqA2V06mj6l6133mIVH5v1sDJVK71x9sQ9YTGoWfr1luQJ/yTUyAZkuDJN4Q2R5a5hMz5s467
DLS1zUxc5Z+cFOH8g/u0O7Pk5Q9KSH2OP+Mk/TJSrsaQ9RN8R/lg+4o7n4JQdZujOoBwyHUPcWd7
fPGrilnR6SfVFbuTJfP4yVilgf9R6M/3AK1m1lrxOeUmje+4vXo/yBh6J9YFyLIuvxRFkUsIRclq
ziIOXDFGGlmp5kjmPDAZMoYpIRpD6EuX/Qv/I5UAsgN9iolQ75ygsEul9n7h7CYoBXxJRKjXPg/x
LkUxYDouB8/WO0CNlUsDZ7aY1l1qb+oVT/ZeH11payTZqZNOSWxakKO4UaaKY/TlqXa7lm6cazf+
tXcQMZt2ViNgGRy/ejhaOFfXYYe0o3SJTpIipeOJpp5t/E84nHck+hSxBreubLcMn2giiFsBzpNb
c/2cyLRLunkabUl7FiZkRdyls/OQbbez5pTqUt6DOSzMADiBTX/k1ikLX3a6TeFjnfgmk6jLFZsm
vHgwJJKdO+LeK0lwqYCN/qEAn3MaZimKOxce1CGNqZ2EOXFRpXKPfzl2aZufhOckqmwtxccPCQnc
Fk9niC+jstybbyVyspW9Y1d2g4FPaz8c7rzHtWFSFAd0vQ0f43tYalzGePLa2wzq6Uf6ayf7Gwo7
Ca0mJSsaYTcez+XP6UwNWfqmBi5ZpvggSuVjVBkb6PA5fBUjfLrpl26kCnHSNiJCith4aYHxI1Iq
XU1UgBVfbDSN3ImEEpuBPfKTABGu3IpFOAxFW65HYbysfJs+O5q4xk1vQ49T/n32HL3D5U5oMIsB
rPm1G45G0rRcmTJTkH/67XIHG2mq0GPz5x9CAm0cf+gGXbVBmHqeVwK9atyNWQE/ZcCT8Ou4salr
pcquxTYwF/2TvYO8hsjZPJd+Ey98aahOSmFkdx6YGx7rjC1UQYzTVrLSOAtKn/N7mZD9rx849WUg
Jf9AA2ayDbiIbSqQKuRpOQ2MhfeWfYtvlDz1bM6Wrso5a9QZA6sZVKnOOyNJEOsqhYMxnMIogTt8
TWb905Ow/EdhJ03BERP1CV55Zhx36hXAwKq23DkOvFkVV6Y1L87ttyYFPR1zcQrGH9hlws+jP6+V
g2GrQUA4aJXI49JxuGNddIrAKjg5yHqDDhzhgh1rkADZ5oQkjIGnTRW2LD5yxwigRGDuNYVxcfls
6+UhXh53bcrWGqzwUwVObAFboxHvehN0LjifKh1Ml/kjCk7YAEQY0IyPt7ovz2eXuM9ygzczIvFW
dpPmr0a5txuz5puDLu/65IGhuRdYv/Q8CrCGR79UDKWoWArh15lVPAlqrkdV+G4RhRzyifntw8Ct
aa0MKm4c8lVkLJFDmZ9dOg3RvJ5F5/x89S6/t18YK0OyZ+SGn/t+TbYvHaKMW9z2Uq+cDoc0RTEV
ugH5CLyFAaJfPOYJ6bbRlRsvIeigf5Liwq2Y0PjNdsAc6kZzoEeirPiCWya2tsj5zqi9aSle1uFD
483gcSojVUZCMS2cFDIOdyhhmC5MgFXC4OcGEsjiacUPgXJ1qkiS+TG1LonYitjsa9RfFCGkShZt
ChZUfuPWxHrR1A6wzxEqZHWKjP913mfNwj/jraUjUUnuHv1PF2gZ0C1ULvwcy5qjWUVpgZuBsTcy
ks9P87YqOaj5oKzBazmO6oCjGMyRzr6QHrKtFgs9PPy3nVhMwRsNruMutwFIS9l21DPE5U/1tAtq
+e802lQkWz/hoPXDbtDS1Df2+jMjGzhhF4tBGtG1MFyucOzd/TcAUihVRrGwckZhXhmS3S/J3UoV
QR+PF+tbo2E/uFOz84Ip7RmtaQyG/ut+kcdSTMJtU8mEVBDW8bm/hPvOhk4f3V818poFJ1fD3bLG
+mifC9IYX6Ido6Y7vFw+55TaZQa26ix5J6YhBCZXhvrAoWJYA1BP5Dc57DAQ47y1BsnvFZqQgH7u
HleJ3IxIlefOamcf1s6FTbGU2+B3I41xcExcG8S/LVzT+157cBURQ1wqJ49JkIT6jZoyDfGd3WXL
MY5PO0E4dPzejLLo9qXIJymoD2dl0eWKGKt2DpIilzf6wggHcfllsgvO7f/sAQl4GpK0UjycwCi/
q5szWrDaZrSh3mBPrYmM32eq7Pf30cWRoQHRsXN2XX+e7rXZANJvgp7kscuSU0KBsZvQdou8Y11U
4N1k/Rk1Ao8NkRE7YeuKAW3GOd00BdtoooHJIrNAMxt6ZR0QJS7gm+LPipttXOn5z6ksH/RG2P7C
KPqW28ck47qQiJGcOYYjzMJnovmKiaUUfCAJXfA+mCzf3lSnrZvelFwo9vwNKxhdroTGXTpCDM08
Ps3yORhrZderDpIBTgB3EF9P3OrPMrPu/YkZnwOlIPHjpWpwQWSlSt31jiVhx5KV5P7XlbZqxGU7
l6PSfnnGAq475riweZyQIgipLtGpXH2Pytc2yhesT8Iphs/sC7g8pCEA3SE9oQ6fTdZkXvmnnZoE
JdqbytJX4Dvvw0FG8ToRmT6IhRHvlwFcf4NVHiFlXIXLqlO1CIJHGAbNDHGmLnNR3vuLLoV269c0
yYhPPVIDLNv6v9Mp2l6BOEctwDjKjATScAr1a6KLGox7sGaeb0NvR6RrmDzv1byp4/E2GuM/2TTS
ph4TYg5YznGQJgvwc/XdBEnFTgjzBTjBms/SUiAzQyAUEQOWM81VnnLQUJiarjZSZQUS9QhyuDTQ
2XwUtsw4R603MthWygXxDWQY+nnNcC7XUsCrHkxnbM7yxm079qbSt5cVe2Tb9zLf5gI0oYTWDB0l
nQvzltaC+D8hTvPLnimlqBtH3ikKYa7cyd5m+qeDzYtqBhpR4WynGvfmc+OpzucvBsE2cIKh/bDG
+Lzo6+U2v6hXRfbCaapzTjSF7muVR+/9u6qk2aytP4Vu9MQmBJ2zMtyRg5Nor6m+W98IPrreJHGv
vGlFrnJ+mFj/tHCT4q1UonmhEGqtl/WATH4JpJBCXdv1X0lhj+D6ywz/DB0y5PJJ1JeyGME1Mp4G
rjVMZPfT8TJR8SFI99WcFJhUm76QtfCGVMyFKrLajhtYrHt5xNVUOvUSBEJUOsM/1Ej0thrJ97U4
3aLeLuWSJR445dBvyReWMIbv8ruIexymdZf9nm8Z76srmQ3J0GVlZOjVQDKN+JvAZLQk2z9sTmbA
xvGKki0qC66oie29vWWj/dumJNrqbuxSk+Vgnffube9IeYwjBihhzhMzmCGOHMHzCJXitwwefA1u
hQ1Ja/RU7iYQ0zFf3/vFjCWs6ELKFzf9AsF7/MlfIm6gWCu7XISYmwaPKTbsmOCuB4YjUiGRriw4
ezs3VHeIFMGCqJoNufU8dBdoKSYW7cgUv/zS21jK+at/Ko6lNZIwOk9rA5LKdroYUct8L1Ywy4Kv
aqisl0n6RLUrbFtSKQykQLFccBTnGWSZj2V19qgHP+5n3TGr+ehB1hqzQoWLQSLId6iArsWj0Av3
FFqhg+LDWDsYyGAyoBapeDQRYcMysEOYlLPPyaBSvcSuFvCojDLlYhnTP3Rbq3H/g+RDsyPj00Cb
ChLyzPU2dbsLh7ICStDCFYMa9PsU/jnCY3CUnqz1ji/N7+oIk1B2IlDGVf0B03mQq6gENDFTQuub
73LMIEK6nnGqxwgkyUrTC6cZcRBveoHw7NRFnwELM/Zz4EkV4GS5SToAT1osuGDnIb9Lvkrxi2Wy
BCL7AroQ4GpncfILBG1TxO3mV5WdwpZlpe4zEwFaNUq2S0PCpc9e99kL2E75o1W63z/XaEQRMG3c
cVIPJsZzQp/e9aAtXOzDJg2L/5WjzfVcL2P/gRIcnOC8HB5WAOOVp4Jor/PPXTT+Yfu7u7Mh1Wfu
iDC/oL5PY4Fq04WZIeAQOdZDRKRTEJy2gsMnAwdIf9EIYN+D
`protect end_protected
