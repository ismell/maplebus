`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kB6UzV5k+LtqW00OSvpaAwP7y+LCUNGAOzLnWdLyxex+z48926XD+BW9XL9Esuzg8k33w+yAGcG/
w93YBcL0PQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ifDw3dJC4/zsZoXBaDP/Pb8AAskxDjXmoPqK9N1plPQeZMMSbQV3H2aPHmDW7kRjMVLXlu5Yps4T
d3QWLwsMRIvXDdkKidcLOcMP9rbPGIibksDSp2RbBjjE9j80HiwcyGVGFMGx8IslF9PyFpLNVqmC
JghFFYKIeNYh5c3c0II=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jznIu/8Wsmoo81jT1Gjx3flbIS2YkGja9FUSEZ0+v19YdaamX4bCjZ65bG/vMqdoH4ytVaJrUyqV
3t//grfKD9ZusYOwjjDvtp4txeEnHbj/Y20GNbJk7msYUWcYsG8hyzFyfOW9zDRZo9Ih4vvc5ng6
yw+bbkLHJ0FB/wnAQcOs7cEZLZ3Yuf22EBjT1DOgoGTsmcdJVtGquEXTa6frU57juOk3RU53j29/
+QY+Z4wztJG3hfErpJeflEgBfutHI+sHJaQrnEQUhpq6fJoYF9l+LE93lXhIR+tM5PgwYHP2kJAY
YfmSbLUW70QWVHAHLv6XvPXR5zeotxoylQn4/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kN9r8TSrO98SyZLp3TmcXeRr2jesha3b3QDiWPORlnCXyi10PBjoz+hvimDBVZJqepSQsyvhMfzn
yv5cfP7StdMG6cp/iTGTbm7KAcZcnNzA5l8KGU7m993ZxRJEQ9u6V75ZXTtrAxxeHxN7Y6NQUSFz
lavNOGQE4GH44Wg1L2s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Grg+O4AXq4r4IkSm4d7Mc/+CYiJGsA/ujVFABgoI7xamQZstiWwTO/GnBsLxwYFJ/RAkJjiNIpo4
YHCYDrDFLn1A2YGOud20bOH5jBVtY40cuibYst75hbZgisVa3uSP0O6PwpP2enr5e4xY1H4fzRyd
Q8xBCgB+B+WzSc/ijSu99CAsDAtI4bb263EoF4WCRqN+rLbvfPSfxd/rJ9W1lmrdA9wIypSYE/7b
5Kbo3Oo/U1iomD19yrdCz7mxsb2OuiPquHn1RayQ2dss+jYpBnsqR7CnXWFm+p71x79IUVbYoP0d
IT4ZRR3ysvKkASRXxGhNHANPvDdCfAXVDp5P7g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64848)
`protect data_block
XwEcTRZBLpb3vtXp+linfXbRnm3BBhR/+cSsFSs0WJuPG9G2K+naBjC3MarzimKxQDGPX3rJE2cy
G0PwIcP4CiKEY4zYQaBTJiJFN00dgJrmdMBI37mwPTy1wNptSox90ji71vjnecIt0sH2DMOmqEuE
sBQulnBN7felrtmMMVAviCPWzZ1N8y2AHk+HxQjlFhKudnnpfPa+BR5nmGPHdxbXLKTwbAOo8lui
GvoMLyiWlrfkV6qJ2ImdZE5HOv507BjMmd/CRCmCZh0VY+m5p1/y70eIoypvleiTamlymGiRiBPG
ta5gIYqUYcJiSyF6m5poaWH0EBp9R3pQGF9JuF5eXGkjBIlG+JcZBR86r5uioiVDfbhPLv4vB8zy
xO7LU37Hluwll5r4yPboZqZlWqN814S8F4rQU8zdGeErbJZc3/HKv41IIZ3/OxnYseHxALdHHSP+
EJx5joE9bevLIUCC36p/Upy37hmivQ4lHCpxpvbDsJmu/S0SVlTynSZug9MrE655VRq16UHBP3zl
2JGXn9Pp8sMRkToN7A0HbDf2XZyie4NCfXcegS8Ik0Hg65Ou/t+9cjh8SIqlBUa63iWUOYRuoMex
/49iwMzCN3CDyiOLXb+fJFPW+DVE2SZnY5zt7xgRe/TwOJPXEDxz4JquFQxSyn8Y7HRT8r4veA9d
KsyagiKnS8cEMVtKMaRoMXGnB49HTh+Yf74xxDy+iGCJWdeIpjuLyQNS6oghP9hJvHYbw4TPrnCK
k0Wxc7Nijz6esSEDW4/2bwYNeoel5GxFDicTDIbFfVvMbCeduYEym1Ai890CbWkj6zl5Kl+p2+OH
rnrZjfazOAAE4Ha8Gk3zkRvxpVn+xS4OC5XR/Rx9xqSKqEIApQK4AwDsflMhUj7TyeXsV4+X3SqB
muvv5ILTNeysNcjSlffbZ9oMBWVyOphOg/2kqXrQ9sEnjAmgj0tGcY21b3jg2ieDVJqQZOC75NCW
vTkyI8sjp8iJIIh0gC9q0vczcGuW9SEu/Lm4GmKoHaeOP0VRj+M6Mjoa3YIwueIiK4Uh7hoPr/4b
GkNxTXGNjBMRvhg5EwodjUzouv6tJLwHm1NyXyCSQkbfZFCkmT7B5db1BFegIIpuq9Xu/vbUUCCL
nXj41jWxeK7ltXsFYqRvdBBbA4ssqgTT0qFPxF3Z2CBU7k0m+S50r0pdTYhkrvu6QC4hXr4CLeSo
NqdrF5YsqucyR29hxnm2sNKo1GpXF9aRVnGWBEJy7ET+AJHy22Eat/u5/dNp4QlbOyke1CxBZ3yA
zMtjM9T+CNvzY+5vHxnXkOJUJI0ArPYHDFYikF3wYPj+Q/PrGHu+bMSzp1XyFfDLrD8Vs9vHQmqY
8EQz087YG5nWwY+UnIHfUC7NWvHR2++bx+O/ywTDwr8grANy5dnanlnG3aioiEDa96tSCM9pT3Tz
qyh9/H8sPAYwMQVQKkBQ3y0SFM1z4dl1/cKUqz4LYXC5yvmWGleul5hkTy12PrBP0GGXqMMbs2qB
zUsDWYN7fL0aMpvwdBkLQrErnve7BGbxKAgvZHeABLRBTm9au+yl3t0q5RgFYe3jkXnf/yTczR3Q
p+ZlzLhu6l25GS0AauasxSloiM1j9Hsx8RkKiNdVZX6kvPCbAPS7WKHDwiYB+j/DAZ+E0oRZZnJW
Stm7Tc147bMP3s/RAsWIOtHNSj/iDtJHX9AURQ6BYHKuSUBCN0B+p07UuqylPvof0FKO5zVNlE/6
cOquExZO9F5pg4pGPMSoywae9mwfZdl3osUV2iYEKue8qKhpRE3kxyClVUALl3ONOiox7vKT8PUX
7BINce1N53kRnr7AukilEKJxGfOWxOLYjqyTEBysQZf84fxhbYHgowOewkDgmMz7+bBuhy4HD4W9
Ic7FG6edmXjgT4giyqT0QJ6gTAB43IncC/agrRf6NZ68vm7xDULSfoXXbVHyDs3M1tl9qA/6R5A/
E9T3lRS6LBHA9L1VrnlMF1rq3JB2aEUApfepckgB2anQvMZNYzQhLwT1PkU9F9FxQHGMhAcAwX6D
WSj+1VlYQEWDr66Yu0Q3TuANiQOLhJarSDMXB1XuSh9HDx6Sikywpna8rcTiivg5NxAjl/PMYq2l
sKBuEX/nU9Fcwg3r2XQ8wpShhilR4U61iL3vBmWa1Ke8LeCp52BoMP3LGWnmih7kAPoCSShj6uXg
4MTzuF9Iq8TKYyZqD9KW0AzpZKh3T7Ik4rF3BeHvCqG68hMnG+4ig/jxrF7qMvK1pnZKZiINghTX
OlTxDmVQBTQ9JQ/aXJDLQAD1lGCj1OnmOiSr4/sg8VUyBw0btH4KFDWzDbRfW+0hq5O89QRSlPQa
WKRAB4gCDsWJEbS1Ly7VpXMrh/LXIzr4HjlXY8hzkID+LXh8T9+tHNI7XLuLNnmFj6pAoNudqmRz
b85BLKHQNfo7WLSSHhBKXglNWAv5OLvDG/weJixzKjstxmPYPwZOFmZtKPP8YIl80JMY3bGozEAA
CEzrPfmLmGwK1tLyUMLEKpHTigIgmYe1xtwITT8PSoW/xT/Ynb5meFZVCpmjRmcXBz8OdzUgLO6u
2ZbbRQAy3OCfoRxo9OFNcRaDKuE9BexmmM6PbWZsQN+J7P2A7kTMZ8xmxsmQl44RAlnxLKrOwhO2
D2hiAz66UTj6n2G1pC9jwme6mBng8+78IPVCIoLOIviVYTXwtzTIGX6n0VO0htrQDp8FuRl5etDb
7iJwf+65SNaD7EF4nUAcG8MIsO0hqp/l00DwKV8GyOi73POpkXWd8CnbOwf/DP4svf1FWTteEMI7
lhfXq+7tszIg7ZTUhAZbn55/VAQ6KGYCRHtZSK6zOvYV6AdYdCEuHolHbv1bToVkejWQbT+Z0edf
ZSM6k6bzkx9RXevsSX+N5V3NYz07djKyx/AmNuOvt/0ewTiWp34JPMqTTwQyU/cdaNJ0mIcXHxEc
/etruDCE8LUrzModub5rjwNcbcxg6Wm/WfmeIgZYlmagu0PdVWDNsX/h6dJwiQf/umPuSwXJPGRZ
3by/sUkJ5RZ7pl6eaQcnXC5i4ssQq2hvE8ZvJj6kYRu/GPznJoeOWNyHpDlFz+moe6xCMwkL+dD2
PztAUVccSpamc2gxO75jtGuZK6SO+tOhbYzSDDRRQgDpHWG7FwcheCNr07xrHipByUguqzor++Zy
vCMuGsJ/AT9TAZ+s1pKqeAetGsS5PyjH/BnKlJcAb7pqzIV45VPoEazwpTd0gODMU7qUZWnnAcGA
XLdI19UaYP5Y0E2ioChS7DJplnI3VXsm1judUb2ky+2eF9S1S4V8rPRmeTHM2BWq13CLI1fjvst7
hxEeYhW7kUzd3qd0RxIPGdLjxiXlRQdmqIRRKaKsJOlazbqZrbZ63Iqe5dNTQQaGWe5KpTiXA4Ss
MEDgUJUwqjWzevOGHcvwziKJ4zPNP6tJmdAsomhPXsgalqs0zKpnZfFXMyMp2HtpSU2PPPDAUgoG
8JdjwBqOrGu27giwtr/Js3LAVywBxht+P5dF87ASCFrLlXKAAfx9ckLQbJkbg1ODerO1JAOm/dPV
aMfvHMnkH3Fywk44sYzIFGnfh/TvIAI4VCklCb7Wh8nz2kIhGlmhvdgO0OYwIrbhGbOybQ2CQ7HN
U4V9ZTYPpNHJ87oZ8euwg5MwTNBGerxvLCXaP6qEKFRmC9SyQ+xhNOvpA5fGpqlH/SqD/URyx/yg
DZyGy4GNm95RGYjYYYsmoRRXGuFRF7xTp0WLp+UY+cSDCBE9NLybWFrPXjYLUqzZNDEBf/JfIspt
l1VOTFsjisanDOQ7rpD/hvkAUAMmT6lbfS4QxLRh4DVBxT7aaD5WFURndCZsjIN61QP3KpqoEA0+
QTNVTDKNwHfILG/LH7sRxxqXfA368+vRHvcLGbJA9SBywTaFU1PYMTsK6YjpyUx6GAjqnitE1TXm
oSq3Nw41WiK5CWKTWctrkR74A3EHOFx3EvQUA/zxEPimgAlpBk25TXhQKK4T16ukxJ4mpcy+rx9e
xyIwFORjUmePjONr6iCKzR2X+1x2y0raJ0ECDPdxD4VN2s2zcvfNFfZ6ujZpugwWYDHQEU9W/twi
L00KlXxS5gXUNgI/ZVQou3xcyoYY+spOD/Lbai/0xJJYqevlVLw2+qVsamMCZg+ckSMQt39B8NGP
Ampcb0Vwfwt7Goar6dZDZ+4BfvC0qow3I5O39cgAZgIaViiRVaFM3/4DO8yFabrqz7agfm5cFcT3
v5ZILbHhEJ4/+LRBOCo6TgUaXdMwy35nYleadG44/zxNtRvPadWgzGttIfHnrBFKcinrArdLadMJ
SLnDd81LSeI0ln+XrXRJvgaGLQOmR1vZPmbLUWXoYG3W2cp2RyQq5v1atECIFPG3Do2O7TeSbh8n
JzVoFX7ACwDvoq9jiGuZYehkKesvDHLCTBQ2h4bInHSB+aGGHFkCQeZ5iutg+cM5vtaFQvmN/PTe
1nDfec3xTF6ArrT7EiJsYNoLLhjYvJvR9zUbSFZRk2vuz/eXWsG6eKok5v5dqkBUeJj6b9eU2l69
S8RGKIjAkUsgvWBkFRyrt2BQXyC95ISIsS5NBmIWeJl5KGaireFjOkVf7fNBGceQfpNNPh7fqUO4
5pEC22Z35kR8qDrzc+A1HF/vUzLCju0PIuLdT2YRZD/veMH6gwaIhU7M8a1ihj8n7gNqDgcGNKHy
GhT1dUMwZmTQxvxDhTKq8rtMvepi3csR5TOZ6kxwH34ppg8ad9mu2af4+8wWvavXaHHHhmD064tF
93Pi3c00okbNs13DZr/Ih71iSV3QcUAGBISTLeFr5npObG++o+B+tbGpKKjZd4aF5x04i9pIcpoK
i5TSBZaw/dA52/DJumWVRMJnK5vMwBqmxhB1o+jjJ2cYlAIxq5jVoE/IaikPtH7Rb2YMyhArRCcM
dg0VVni7GqAX6FJHOGB5qlqIhnq+tvRrh525S5H1FvJK1IU9Z9JTP2FeqnSUXWZpyckAEElzg5M4
DvO6m/SWtRoJXyESlb9FNt5NwPbP2Wkqazy1K/yhmhatTt0sBHWxq61om89xs0oKF7DuOEvm4SUo
ltLf9cQJBtLf1xsY5vJhQgm0S/hEpBv4+0kt+e4Wm+6Kuz9bxKRxNJ4nzp8roUVJLWF2Ttr1HuSB
uI68QCKUnq6AJJLHRk6icOeCyjpdLh4AA8V11MBh/F+Knc+pY96/rlkEPPre/PTv9XLps8XCbofL
wwxjCIDwJtiQWDBOhPZG1m9qXG63LkGAM5ESrzWZWz7lsNtASBv/GDBhCZEkWphGIMWQssUPjkU+
0lPResoAuAEfQStjmpLwraRPnUE7pG6IUAXXYj8gcpzo0WTt4kWjSw5Xj3nntGL0QLYMFdIG5IoP
jjsTp5LmyqNjO8dWxniExbMRWKjceB0ubJmqbWdaXcbqwUyJU6bxNyLwme+WUdn4V69F/kB/tc+i
R5c3BsJi4u4evjgKw7lnnfVYobPcUlAIDB2T8atBqLMlWZhFQg3Y0dxN0656vBso6GAKexv1Q+Qs
SINdmvi3N95HBRjqBm2Wz5FY7tKeisDq8221nqDA4+3XkB5q6bBVzIr3wbme5HqmxMSpTk8LoLgc
8GRbH0soG9MglIWStRn+EMRGfVH2Ve83JJ+w3gbuaZpXX2LY/8/KzI5RIHrwCqRmyHIJ2tK/3Gcx
Vh8Zz3fH3brswPS3CpW3ZvhHKaAInTZAdn2d2siCL3RwmXkdEZwFctjsWVPiBLXYyLV4ib1Payrq
v3CJGveJLYoZhQ1v+Yn2DKd6kVsx1sA7liDLvfvviEsPIFlaQnMjOekhqR5AtlTKOG19j7JG/7d3
vci2oc+KoOm+5G8MXO6vZUcXWw+KalGLNu/fieC54G/KrxZfOBetAELsq8saPDovXq2zu/YJ7lAK
YIXMi9tlf/bB4TMWAtskrEdYh5/87ErNOlGtP6/glfC7k3LRUayxCjK0XcZPcIUoVMjfcLtmzTSu
HN6otebpHTsWvY55raItoafehkAQYj07dQA7YB4Be08rrd3AiPLObZjYPEBWt80s/mQdCzG5dilp
ae9GSECfhFxUKJ8nUSC5tM9oNGdwCOYmSRvSMLEyOpOgOtg/ZSJWdfWnvbVpFjnFqX+CQH4viIZ+
uDu8g24lUQakv3tfl5Wl42EE89QUGOzzlVzkteDdYfETdD2abLOeHJw31bpLJBdJSJLvP3mi3KOa
HXghcwtsrnm5U/TtjLJt0VmzU1NNZzg8MRfSRN15Pv90rKJ304PSdDe1k74dM/AYOyXb51TYueQu
tFqeKIK6Mfp4M5aCsXtj6KPkD0iYWZVxC7Mx78cysCOpzn3cE21h3L2r7b7gw1or3el7GfOsvBRK
8JZ/4Zi7Km0ZMEB5XVMn/F0WzkQJJDasYyWWTCCMbrfHvnarW4hGeRXxyAM5FwEQXahq9KNOs+Ma
MeoOPJbD46TUE4plDlDi/pa+ialjT3rE7aMYnQ1QZQbYRuFBaF3S1DPfdQB2svXuTC/E3KUXgN0C
C/BJELVdH82DSUZONcuEuUvtrFQ1789hwJHSRIL/Rxbn/8AIUoKWgMZ14n60ohYlMeZ+5vZU/AMw
xQrXfzA9Xl+5XNc3n54dY5kliojFmHIRPaZ+rtC1/YASQiSo7Q9wP0x7lukuN+IX+ydajiq/cZQs
gFlbOJZ9YUP4mqDX2p3bZSEM0TD48A+na8kWdNRHInAvyTiES1+L7K56McikUKquJ+0fnGlFBnJw
+6EnJj69WnmGgWDq12jMahgi9F9RKc951MT0n/5ULKbFaZppNUnONiWjm2kK2skwOIwJ7nDe/yiY
sXhc6Bnkm5khqsAXVAsfLpztygvvHRckbgC6/vlEE/KAt5M6r86MYnXBvb1tYWIMFAOm7eL03aoQ
iZifvIlvDFtdzcRqUSyM8TyAooyS9vptXwkw7SZtMd0vbBfzDES5mzGhTNnrwWmpl4qArH6njBHU
PlcGHNDQrWdyIEJonLgSRyJ9AkWLjMuROUnMjg5NTo6TI4YLzEUlnMyKcGM0iZ+eV1yB8nq66lrH
QusPDhjJ9Yt471XWY1BAmk0AswCQk8SP4DaV4eORlraYw6vzseyyeAJ+zouNrLrufChMXztWhQD4
TpX419iD45hkC1NoHaoR6RCF9t0Zh4pYDq1QkmwKKMmjeKJbfyGWc1HB3YTlndesBZzee5rJ4Y+F
YLLywbZdXHITi+dBsR3f2hdLLb84f5pNKzzylNN5qUvSRrLX8yafE15+PUrKIKXx+XjrnwEsfJR+
6HeXROvNj9wmrs5q9UX7vAGysVyGSAKE0CUvEUYr0C1AvrTMFXGbAcgGZBcazCiEJDJ2naWBrnxV
Eod3gLLTPyAwJxEVVJ2zkQrujZwds0urq+sZ6zJoFKz+/EBfDN6PwMlbJnnGiubzdgVO6ITH0keM
ojPhFIaCb9sOwI5p4QCYE04VT9WF9KivuwQJ98C6HO0rPplRKoQmp08uzhlMB0wGtrQ+CVUt7DHT
Rtscmei4i9LeoF1n4s7QZ8bxpUX/VVaiknnVdnjL/RViJSaL4DvF3xGO5IWc9oMJgNNbGbLqoRaP
b6mGdktdLbSpbvgJkZEiekZ3dsOlnYzUh2O+lR8HMYH2CRxVrPbGRaWFhqeXUUxVSB24LH8CpHX/
kUugPGLPkdEi2smUruclQ2u1F9O0PRcoWmAN7UqH95JwYcyT8V54fV+zmQez9B7WADX+cY+cEARl
8B3In068hLnRJ8T49RnkfOuxiYs+kgtZOZtkfMSVXNlns/1RO5xZ639O8Me1dLBtmnmtVKz7GV01
TaIRnV/1tbOD3E/4AYWYjkjbfddmNvSFwPbT/slHcLnexaQ/KQQx7L9csqCTgMpEkcvrAbfvKwOe
cISeS1FCjPdqjdiIvHSBtN+I2fM6caepRtgvD6o179lvvY8pSWmLRHBobWOCTLmfai84hk7oTGoA
7BUyd2gx6yqt4A+K0rTVwmBRtegLXBNGRB4a8bFbjtCIBQZZRSaG2TuPOcDUlwkDqb/fn7w49u5f
JSscIQC+YheqjKak98rYvVEb99xe48T80Ke+rC+IBotjBABipbCbFZ6vAr0YZX5jmROfV/1LD0Fm
cfio0899WZT3fJ+Ul0vavBke0dfSJvq/FS/frDwYpkr9oSJ9+stOZYZq//lulWiDV6mz02dn9ooj
RXHwbvy6pW+QYRiYaEIWqR1c8wPV5U6GfJtq80s69VIZz6WdZJkS5E+SyYFS2alVlyOeqNNK5nOc
qM2/ezg7fcAn4Nu9RJTMI3BJincUyHyzbDV/0eu9WjrG4ccXVfgumHewqdEHJxKVqjgAv4CbR1EH
R6U1xeYIE4I7lnspSR1inwGovIXkzec1aErsumLIYq3YSCqfjgvSX8/oEdaao8tCpIUfq6McC4S7
qid8aDOy1EUKAhjxJk0s6AH52xnvn0pLjCg0YHVEZJpNGX/Wcm0oU8vk/igsYTL3FsgiwAYKubOn
DDCQNw4XD9O+x50XpNPblDjuc1VRMmMv9Nz3+ugGft9fiNYpyJ4895HHnGto+DAIJrQjdhYDkJig
rFyd14cXi0gnwyq0QVvj2fqaKl1+alij6xtOB5CHTVM0o+9kZTTcbp/mG6SgkQguMan86ODKZwb1
Y5/9JWvlFLC3WBzxwAkvfekzgYrOimhSvmBGNhL6RWIOKnoHKgNBG2SRKqq0w/M8EvKVTWM1Valb
CUDhZ1UGsjwUFeBfNP9AkDeGUrIMUKV13eYNa8CdnA0r0h2Um++/2YRo3xYRWUjfdUKFPlSb2wog
kwQOeJm+gwyi3+Sy9JYE3VZN63tmGUi+hhLQcVqA++UVxtmW2LCgY7VJz7ncgG4GfG5+U8ZnECzH
G1dzucMHQMIGnsFnzva/QX+RZNSZLjHyQe3XHzNMXIlstpL/zX5sgGjEx6mS3lHsSWQQebkH3w6Z
XgkIO+u6Vs+DQN4VipcD0Ch09x/5yKQdStJ3aK66zuAFdHjRYIja1gDQmovKSzX+IxbjmdZFf4+y
lf6nyulgHId7FkKZeFx/F8Jh3r4/tlGXLr07Ls8lZJy0hRs98ik7KPBOk1aqES2g1S9bd0AagIuI
KhnPu+7cXPiDqZYyrrRgpIt3oJJt+uO1CmF3AYh3qOi3rqm1yoqN5bzP3S5rrtDomE8cHnN7PpNL
yqpGptNmk89CBvvJmMME6yOhIUmYQbujw5bsDCE+N6lLl9zleHRHsle1gvwplnpFaD6dtT/N+Hh0
dTP0v8CxCRXbB70tGlPK+V3U5OwtKCTtzpgKMaT8MWiRZO7NAjzzJnEwEjl2gpPH/ZFOxrmWWfQO
yQH+IyMR+ZQNyk4zq7wWwgv+JkM7ffzSTG2i63YPrtn2/88MsWVHAEIMRas8xezYCHJdYEjSvsWW
B3D1JJGZB5BAkABa4ArNdaoozTrCNTVQ+gBIQFetY6VtukNfXNG5/6qYZx63WWZZZfahx0IZQZ+f
wgir0v7QYSVMTeEobvmOae9tspyIMZQc3Vipmn4DW1BMCqocZJmqAkXy41ZJeZBbWrq4uw9k41JK
gl+wx48B5FkreKkABoh48bq1rEU6AltKH88olysu0St04jGK2K6WD9xuQCQAAilBmjwcaXnCbxG9
u2bxBBWDBrlAP/yjpsGxd9mEw2rW5vgifZwFgIodPmeXTk3Z8aUWL/LMGMPbC9FnwjoXee2r7fH/
48Qsy1g2dNeI/0D+1/syU8YLO3V6YnqVjUfayBshypnWTRUmofwwOoegCSEV2HXFOr8KRKGauKKa
MHzpkgCsxXq7Wtz1zqqz2ONVDwWu9fcGxL7QsRHhpmvj5/jC9UfNdSw6bNDvogpBPihMmROP/ffF
lAqjJgaPFDTvx1tMB3RC2dBvJFAh/9ZGbQhnOP1hVbwSokueVhpmFkacnbSFS/u5UABHh8mj5epQ
2cS0y1zBnTbI9e+N6iWXO8CprvJND0L/943SOGsRuvyUShhVsxmoSeOxv1NmljG4uYo503dnSF0h
2qZh4oPDryC+ecDI1WNu1VExO1h5zu4NBEMIs9k8Xr0B7E8CIihZVvW89YHptVfQksJRiazYVijM
Tpkh06gSxGLbe+JHKTIAaX/UEstjvmpTIYtAIBX6WOhRqM0gIqOTcQCp4ASdOMB5pEgQYafXs9KW
v2I1ih7zfE+KQCRF3zBsg6VNQRYundQqSd+Wd5noI5/mNxjj4uLZWNit7YU026ENdGtuaepGw4lk
haEpNzTWeqVHGFcpDeGgqwP2hDbV+sGgzzmtgH5yi3ZAJ4J9BY9kiFIFtQKw9Ou6d2w9WjbJZjeP
L89kd0wJME5cjWzXgIf5yVjabWhkDXFfvJRS3rRPoCrCx9IL2bjhonDgMGouDDkRu5L4BAnKRQOl
g35W212VXRua14bpKjCrBDl2aYBqdLt2xIXiE9Z80YxbAPusVZmYQA5iKSwXQ7JxUSj2BYK4sSD3
kKAUTtlbb9Y/2OoaiV7ELB/5DaZAFu4Bg2xsEFR7E28gUaFrOdF5ngytNWY1gB6J5qXSdLkTfQ6I
LiaIryxecFPI2xmw3YBRSs/sNH/0jiPcCn/vqDz7z1XYqVbVt5bFfSLN5UnCRpsC0YH4/tbUm++z
W0MjTKbbVOI/CYOKDB1Jt/EH5XbWxxsf5DEd2MvTVwV9jgHs/omiCfgEJjlJ2n2pl15udmgkRyKh
ZC0ZkmK2em0tmiC1GwU/1ZCiSwhEutVnRN34AwDAI+hHL4BQgTxre/1ZpSh2oo/P+MPnGMEar9B/
gS8Xf/dxaRZr6iHhU52oS95cBGV0RIS0cpOgRJHD3aOPfp6L/222ADxNaPG+2ZD5y8TRD1FhU6N0
hA45QZLl9cxy1kxIFIFI/k/57r7l1QdZy5jzsoTaO9xK/0tzrCp5fMSBbpb5JbU1g99ryRmwHvrm
eTfockAmzZIgz7W0aa6C6prcPlp99y+v6FTf7jMNzfU0PtK4WtX2S54wW35bmAgNA1m6QmHpXwDW
RHAzEiAcr2fiQe4mg2+1fe1E2GDMTJ9r3qvRkjgGf6+U8DPobpUF1Km+/rHz2pdq8P39ZUTVuROQ
6jSi3k4hueGjZvgKATzk+nEytuAeq4E8azpqbSSNIWyOPtFpoDNfRS45S5kn9RIs0SLELGvZtP+Q
nwX7JFfQbPzwPaKtWYkogb729G9BIyPtCBwbLjg5WrD4we2eSSb5GvIFNqLcyHWjLmvuil1rS8/7
P7nyWAf5qO0/Le341Mp+2jpn7y1Fx4QszmxvBe6X6Mw3g8lpMaBIgJI6Yss4AqatGJZxfc04YrKF
LXXMKcm9fNAyHDqgwLtldPA2vlBmP9QMbDVQS90Lio8LAj5GMsDBhcXJcyA4vCZm5UMsqUl+eWEJ
P6Ek12o+t/QwU4NTnky0TYc3mBuRjUE5ks3+rfnSv6WuFd6XbseV+kts4bys3FaPCaz0m3dM8EF7
XFHhZFXexIJjSsbd+P+NFIbpfNz0LE39iLdkg8InNAb9RToZvN0xOSrp+w0EK/TjHIASYD4T8Oqg
kGrlRwPoQ8EpO4TKCNo6VcrqjvNlWoEPa1ii9Y29NaROE5P5XhQ898j6NBSGrIz906FJiLipOHrb
OKciGIoOKXUi5kkcJTDsNL6LILexE5fUYAQxgEl34w4ZGu4tdNukSmWcGQGJLYCawQP7px9sXOyD
csDIYvDyk4MQ8FVkm4MeoBHHAysur+lkLefJ/U7R5TGRbsui/7jTmns0lKDD7HW18HoeE86AAuJt
F7R59yHk3Bph7WV0cSn0sK2kUpGR/AkYtzJbs7/ax+1lJJns6VyJoF9WB4thcnDIRFlibB/GN7RK
G46IGlzs0dX/K5IGHguQi750167nj9Z2CRnaRS8g0Xh2SZe7D0ldQx07DuiR0CuvO8ExulfVzlXR
0iPcDg7/oLwWN3yQiifCJlL7NFXiZ4JF7rZZgBpGfC7E7QYhKlLcl+0IxuA66Co+RfPk9GIzbRQH
oOUrmCvaXJF1xqMRcQjX+zMbNirYwXsAERqk0Tg+/EcIjPijRvQ6D73sDhVeIPC4t+bvRc02SrVn
+kDPEF1Zludp+SGfx0xHrzzYSx6/r2YGvYQixeHTxd6HVInNQY2ohH4vqjIQAmXL4HEtICeRVzJQ
fVx6wRcGhtNzrpnhsc3JJ7HvDshSRElWiyOcNiWobgDET/Vm9lBFOYwL4htYraohfCbbTHQ6swRH
gCvQ/oAaIBlkpwTeq6kC6RUC1AKsmAb+EnNLoqEqb+zge0nySAiSewuDcOgoumjvTpk459A32G8P
bZnOUj2PoPrvZw4gQ7KLRP+9ws+qzL5Nc6JqZYnF6ocGRrnYgg0TN0RvbYt4vUm9DGTebCTD7X3C
5Q+BjuxpEOuyoQTkVsa07mreq9D+/miFGbsmZGp3l+znOQ9c/OVJRn9ZD/mnPfJqqGwkJ0LvlKJM
qGcUzHMDU6RiNwfGX1zOjt2mLX1x+jKOgdPi4HoI3NnVkCAqIBHodCefFaza3PtQzUZulqI+DNf0
Hyy3AbcWZ7oV0FEUbI81xiCtlFulpYXCM9rqTa/3O7BOPEAmNqSiAq2UzQ/RgG/08xTWZ9yurP/n
E73xqnm5uFdgNmBR7g2q5Y959olxBUkAd5KfVmkazVj4WYT9d+LQSmxjDozGpzxFywUEGOPJmDEA
oNqddcKe4cF592yT84f3AJQmVusX0jWS2knxuRRnk4GaPoC9XkrqwAaPFEm+Y8M+zYxVL9l1wd4E
kq0N5b514IteRW0kBB4pJNpMPN0NalTRZIszibzwOEHA4SdqSqVfTiGrB/EhgIpAbH4cS/2dewwa
kmGzEHJx/hHlIg1vnAnlDXTw2mqusZSZMGu03IFg2kGIPp40TXSmiHNovOqwaTFGh+QpDJSlQ1Cm
9p2cpLYtd83x8+u/9K7wZCY0tqJTNiFVR5rTXeqt/eAMkOCPieVC7R1ET9YhF7Vu0wnonpHaQUQq
FREhtjiJHcLxSmWPcQWOhVi2W3yv0rfxOQhul7eCUUQ8NgPjokCEz6ads8KqCFbL9u3E/T4WdGV1
BwmJbYg66xYsiCPwlAabtAvWeIMe5Esl+CXbtyN7vCh4FYDNOCg29+MkozrUCMXx0t5ocNPC1otN
RZFA5OynHN5ms7zSGWX1eI++6zH0FUcud9Er3SUPknd0T5YTI/ccSHPU6XACG+oRvxMaJ6fba1Id
YzDW8VaDord/dMnmL8z+sJ7lECUYiNWOTPT4l+oVPYK9SESnlJCP9EWDxzAYvYmQZWlfIfNDio4R
6iTBei4JeuA5QfTPJsaiIISTyEDz9qquddwmF7wysgBnAp9wBK8+MEew+xDYWJfG5qMYU4cT2Xhr
4dvPYDP/YGZpTUoJIb58iL2uOZaEdhFAXD+Jn82AqZszWFQquSAJR8BqJAFTMHtLjDGKwZimHf65
IiO/nbRtHPifbVc6aVZE9UpAjTieGLlb/vUWgH9UsgE54egOYXUmx9jdZHFTq2LM88gi36guyA0G
hPcnAqH052YQ73Q9MOAvPkT7I+gzPsYUBtl5pM1xgfOuDoushA1El0l4Nx53XU1G1yYYXMzLzQlX
ZN+OrikD7jYaX/K9I39Wet061hcgjXczolby0wwTPd074zlQO0adCB4Txf1vYvjXXp4WmgSqLHxA
WDCueIhX0hPOhN5eFEbdbzKyJzDbOAdlFJNEp+eWqxSntrnqwHJpVkAIca0a+qL5SUiWTptIlTXk
CiWopOYJw/A+HfcjuArDcel4jVqCIsgDVD5oNpgqBJ3hTizgbw1mxu7hoXjksTdmNBN8ajvXYBDR
WKZb4sC8TdzwhDB8Tla5XdSbOpRvzeuHVvKFuW7ilOTJBccpTSC6FwGCpqnh5K0kpqXpidbQy/r2
zuCDKywHDYUh7PC00qBhgB96cUvWskMiita3591YixjStlhc1Vf5fGswS9xOBXoozswvwvybeKfP
CWyrJi3dTlt3NfV7KPlgvWFsP4wd3It8nhXJ91HoFH/IS96Q3Y42aGN8nCAQP+hpWgqkWxV+PQTU
F4YFA+L6NDEBtAjhm6pcXMc/minCewRdYNOx7EoFmv17iPwV/ObUwI4+GBwq/+ymVV2Kv5oOFQPl
PHrCu0h0eDSmSDTyb/e1+JO1sCMxVnF2gDF6xsqWl0b9tMTBwTcAYYX3rzQXrTw8libVTmq97KFR
gQDE19Caw8zMt/T0JlAcwt4EwoB/RnNFhWSrUrWZGpx+e0yD1vpPvsWtN6VEBU5tyv2g0QOOOZjh
TkbTrKieSam1465tqk3wnC04F4z5l6azEdW89eI3gpQkfdSmx9OUKosDuMQPkcYxJ6aZkDPyimJP
EK+xUdgmcRY9josKfL7VNtu3SmmkgjLwqLcVH5RwRyHdrs7hMMgyIPY5oxw0n2me++Qx3H1mvC1V
I+kLV26ZXXQKZ4igPQZ6ThCR60QpJeE8VwlnGUOJnfNSRSXXsakEYN50JCbk+wv9tAjvtn/uD4Xa
wqadppD7oi9FBsMjTqk0d5bbFS00e4ZcKqLDg+mbx24y8Ivylo75nHEiHKUozFd7SMotN4aB66db
Jj71+4W+PS7Gz9c0kCjwqj2DRYTB/gKE2/2ZLRG8r9VqLmXuHZefjc4qZWDB+AtHpWoO0SpxnWEN
T5I5bqe0TEokNP0eijIv22iDydppemu22YB9yikmK2YVzWR3cePJPOiyeT6shYk8xhPvR5JKpABP
cJ1UPbNmBDWMFzeQVvVgNSYQ/Qwrm0Dc0EQnBUzuDv4SMiKKhUgBuk5zGQVHFHYn4YzivdTrl3BU
aC8KSgGG0dnopugoEsRHDEXxFRI74FH3XGO6hEW4b/PTgHJlMQyG3H/oFad87h5jQ2ps3urUSu5s
lezTSXtrUAjPn/qIB7Rg2gwhGGHWHYD7rRaB40pwLRyE0pBY5R2czzNG5tYCAm660hpj7zPVAEv7
RazM0JZao+6h9pj9iO1A1rhGjHELgbzpwzsqtQq+6AcCReGtkMu3m7AVIjm43BRh0Qy0i0J7xUYx
zyIEI6E4fA8m5/M7O8VqrmIwLju0+q+kk7SxQ8Yk1PlVTK8j42KwjV7HsY2sXxY4igDs/9o7rXXB
qm6jBJbk+04fYBxv9NUTadxwIzf9DcBVXVHBoiLvhYKJ9uLhY/FvG8Z7hBoc2SEmyB6a8DkpxjdU
B+DsjTwHvjnecGjvSiXTBYSuNj2Lleo6+nAjBWtQOsl+uxm2mTucv5RQTVK2nLZoQ/3djPAiynCV
d54qXof7rc7qPb/2LMseHwIot9XLNjG6KUCVc44tNuXPilFMZgQfTbCJcAgRJlaJOOx9ysNW0JF+
RGjAoZkMkAFvEJJfxAMmC+XoN9peqmkM8HJdUw/L08N/JCs6Bchn0HG2o/Zrsiummk9mtIVVp/6h
jrBjW0kn+YuXmZUkteRrBvduTL/gcEGwXp6j4WJLjvQwQGwRn47bKZeGGGXXC2m5mqlaFgT+NHHJ
3gNqyzEN4N2rErV7Igu8P5fx7egXg7xuw37/jZbi/JREon0lColBc+9g5pNOkLAlbigWD/Cm/UPu
kks+19wGHZdJ7VyLyjRXFpqfxFfA+fUf5n8jAjlbNzwiNvw1HMY7k/6R0MgL5lfnrXRsCj2OcgLj
jJ9jwiZ+/m4V7ZW5+lbebdqcCqJSY9HrNVrt1JzO43Q3gqeOd+ahnSpBfR+UUQCM6dB+fQwpqiPh
a7uHTNPqbrunaDzjUMga+0ED7yLRDTae0wPudQKgPnYWtu5DKro2R84saBqM4TW2ImffZP1BuKxO
IKMhmXOopi0BGOvBp/c0SZZmmJPOIzwHfeIU+dAQx8VKBhoooKPqSBXNiORX55qqUCbchzHx8HvY
d97E1oxL1rM1BXQJVChP+1DiH94VnrzcvhyzQCEYqQnrCcnWz1hUj0F1Y2oVNhi+hGjn7JATUAIi
nDMpPRyt/mNMZUvIkiXEZwnUtyAtvNarNzXDbu8mb4PW8G0ueV6DJQ9XkvUVZ9kO4rVKd/ot1lz/
09FRVgiyiktAbRvsr6ElwQkzVc+gAkJspGIyFWAqUhqgu/YUXmDp2KW4rGwWTlpPlb5OQYgJ+/h6
lnAkmiaxKBI5b8hgAo2hh1U3snL/SHBR4pYjiFE38K9/Ke6qumotSMKbEZSgFrviLWSIrw5Lib7a
R/pUOLZ1zryr7nU4uG0bVjp/EkzcH0lXYX5VvCj1JSXzMyW8nzrOu2WXXpFlxGQyRBJAKLSR/SBa
N7NSLQDww+RPMXEU0FBZjRtT+CgSuzrtnX+P9IgZONTGoEXkOmu+qM5EEFNHjyrDcg9dnc+T9V/f
vPpG5heypZGRdVIS+o/dLPx9lBE4DjgXMEt52HxEyEQrKzF1DHhuSN4WaAYRgbqgXvgZlIvMBx2G
mTc9zWNGYnHEF59J/w0iEDuMKV07Y4/oFTEoqUetI1OO+lBPuLXdL2qXaZH0E4r+Y39Pb+WCxH1D
TesHyFBLOXojRdXiRqS/Z/nB0u5ILt3HLPMvLCzNt5XVYEAqXb3xpSbF6vQs+BT+VOMqd74yJ3fl
nIGAXqhhMCmYHfAPFrNEF8aHAbremX8M5OLebDhwoDLdHwD11hxX8m/v0SmnCbIN2ZIYYqjd4Z2i
lYwW1kGH2anyj3Tm5U+I3iNM8//iRFWWeojtnrqX72r7buhSYdq8n9PP5lrj3zV2EzYhef+5ALN4
DBmmE+Ci886tN9Os1K8o3y9lTS5AfEXasHQqC0swxtJzIZMei4MS9kfdk/Jf/IQJrkKmm9q4L5qq
QtV1o9kM7HyUvimEMolVs/1Uj990xsytcWVblj6kHOrqzH92aNZJ7Fn5fDjwNqPX+sNuvVLLKpO6
zIY4ZxsDG8au3eudP6YosaMmzwE7Yo0uBLW+Q2Lxto2QTEEXhDE2TGXeXFTqsu4/5drz3XZn+SUg
xSeY02d+tOrNz8FRRhasWmT8OhxOVpXC4sWFDhd1X5xwRc8n/nGsA+38a2BzP+msrAY5pYUCoy+C
qa/9gMVEGy7yIVnDmOtxV1bVq4O7CN7ULB5r4JH7szNb9ebz/hVXKPAyR7HYM697mR01O6wBHOVO
G4BwnrTFYqWuhOndICbuvWfvn/yQ3TLLW6zMvS+OJOQVAO+pM9siUigZccdEYZWBJHJUyJa2wrfC
jYRAXfiM0CgZJQgSIKusFoq+ziR/638f8MBUPERnEa9wHGGS2g+qI0eitjigB4nCMv4ao+6pPddk
2xX7m3nRaa/ktVs/oJunnMTTdmjxZoUL3wWF/aA+P58VairsXolHKKhxaJ0AbxfWwikiMh6DmW8v
sLOaxd3xqgQzzyZ0/3gyLVauaH8pGRknQ6SD5PRuQ5itKFtcGlk9vTjoGK+NL/LMEUVVLM6PGbOB
iaKl0Y2FS3kpZj57foNu9uyY3HKdY9ZRe/evBMoKm+PgfF8qo+MQoSJPPL8KUAvzlXfAmLqey0gv
LF9eLrAySMsMcJwO6ZdXfHEQpAXzGss05nliQUu9YFgcrO61FkWD4Blh/FK6+WnSWg6TnCxn6V49
7s3zaH4QqB8ZxvjVWYajtQKd2DZNxeuNnFXx4+4+W0Hyja5ezIyaAuKGVl2zceIBdaT9zuJp6xBS
adFuJDNyYR5nraub/T5z1b2m5lxdjHKwe36d9YiP0LUbGiuYJsO7VqiXdUi/cvmJe63A1HcsdiOL
2SCVwRquk4CRb/x3HHD6mKMX1SG0lQnV7//njY6UgBby5l7qPRNTtb1yHFbn2KCDRcoH/4a1TpPQ
zZR7RoiMpFfvu6WAx8qtLgjwNPgD1NdvP7Zmd8C2bnyO8cBLsv2PLbR6LoxcuV2h7kwsI2ReJHyX
9vwrns1ZQYg6DXkhp2lF99wm1E23tdSvQpTSEIeMjHcGJuCeYvXPTtasCCKtgL1SgKv+QwNov2F5
3aqb/WjgU3sQHQMPG5+2zig86yrLDiy8O3l9z7ts5UlcxYUbVw4NrSKgjwTKp1Og2HTCf9vw9385
J/pywKd9adrJuaDpIIa9Za1sNPY+4wjl5iGMet0A75NBb8iAjJEmCTVWPKww6ivktmI1k788oMyZ
yNSx6pV8hw+fsxsl3G56ObfyRrYl0uHOYuRpWh0lTpbfXTGbDhYUUABXB9bGH35FVwuP/CmLIfb1
JSPxZLDrPScgE0zaBZVSASNJZRqC7PPzKDj8M/SE6Eh9LpwcFYVNA9ISuVwXxtDvy62qO2xhbDOA
iV7pUYV5ewrZB6G+Eh3vw6y369UzLz2XJxVKCvDeDWViosV/twJNJUyHZfIEuwfySca0ppvfY/aj
CGVlunij8ZtCNUrzSD3+Q3RtVmVejwfWdVVwOCsLX7R7LAhJhcTJe2CuxzTmy42B3nLlIfVoUuOr
tWg+Ix1e9TSbIiL3g6udLEBEyxA4hyRFkoVQtxOE7+r/safIsAUhqbUpGxIlf7JUAK8szy2raKJ3
s6e1ktUl65Ll+B2ILOJsprpjoDKUNmdsBxzSv5bEX4rqfySXdtJb2P2ORIc9PojS7wVMQjT5HyWn
xjtA+p/MwZtbLIRjEB4akwIkXUejRN6juzsgqlb/LgWMse3sL9KJJMO/gNTUpnj4TOJFrO48zpXT
e/WuKY6tyZv6s7L6/+3sRJqm9WHS6yiggy/vQB20mFer2zXLl5mGzcAaChWrHL5bAa/UtFKi3YrV
iWKdaElwF7OErIV4Bdg077wbGFQc2aBjWN7zYrHZ4XsTJM6NbARlxP4orkEg6Po+Wr8JQi7icQeN
Rk+bG98ATiWOJ7mZ9usRbJ1pOjFvLYZVhVFk8/E4nkcApWerXFhNYapSh+VzlwM4YC3s+mdkkwq1
eOQG28a/6gtA6BtFGAjw5Rmts6ldH6WHFOpwhR7Rm632EjKcbX++2wMEWV9mYmkl2Snmqv5Wmz+q
SkQAWK+UBDSEIQ1ZTRezqlrg49traa1V9FvUMbvVYSCSybxt/hO4uRmpEVcWAG727k6ixcgklp61
bHqGmX1RiF9VnPFx6gIsdeQNBkulh/5TMZUXRPIlUSGTjsaCXUFSpMZ5uUKzMIvvJlM3OMJ+FOG/
BPWJId6nrlNLnQpusjPqBRdccof5j0elNOGZSjrLedZDUFT3q9s7cv0SjXnYKuU3bgioo+oeAs7M
EPYC8Qm3sDNCgqurXqNUMZOOPCoERzLl3jbWRXTX2AZv5/e3WIIl0w2Eckub7U8GtEYT6lKXuj4X
1LxgY2P755keDnOU6bsnrZVW1Soh9CspM9fRqztfDxat7hyhonqDDkESKz6wSoCTTCQ6A6WFzMgd
6homtL+jQRysC6QqH3nrstXtTCCtboS73cBfUeu7ontZuvJiGj9J4y/HnaC/fhHUCjbgbk45TU7/
XntMErv5xvzCKtx2T/KA1t9POQRcY7YqyOWc+MiHvKb5W1j+Hr/3CjQ3HXMXAyxlnbwEe5Q9FD0S
5VkYgocaJH8uVJlrzYrvnNh/7fAEEkXl8/3JOQeae2dl6uxj8n99PpwsWxfa5O5izfzP3oC1BoOh
YZKGW0VVrOwV8YIpevI3YJChGNELlfKMtZcuXVlChmdrm2q7DExUrke3nw2fT08XVER8g3mOaCzA
QIBP77pi6ytnev28HH79cYL0I5S4KwN905FujkZLi6qZXPZ40ZODbiazFHZin0YYgh5DWYvYKshD
2WQ2zIAZIeBGgWO12VMOuP8ZLenQl2m8dPLIw+afUSNFLDymqBr3VBVGXnerwbDAf+RUp6Eo4z2W
3a6lS9m0VlweqIboTbijPEOSasuAKDBRfHEFadrBtPlMwn4ZvbivyY/a0BNHlX7vvlObIfA53FoP
1pLujgf7Gu3tw1h47Ta1lFontrcINLl15kkl1rd5qVURwWOnxxlDHQbf900r6qaZ6Gwv4xXZvY5C
XjxOy8L4+c/9VxyX/jXhqMSn8mApwpjiQsZx9yn6p+EyYRg/r7HFlFG2TZfbl7X7iPTSZqGBebJk
yrQpopE8UwBsdP0cAaDR2SUVXIYsqGgDdt7j6/zs2SyWsixmP79Gudhep7crqx6GuBaeg9R428bS
m02MZOq1sdcVzQw3MD/2Hj6ssIMYIC0sBdigNmlu91YxZDf9D6N/r7QACxO7IgH5sKBZXsYLOzCQ
4XOzOGub6H53xW7T5CT9oGms0CKf8jt13GslipPGRhFfaN2A7KU2po7f4R4udisOM9CVa7bYvrlX
JS73jMhT2sa+nQyCiXIsnMaMcAr2+1uva6KVX7T5PO3I90wUAlYK6EVKthDroJtc7BA3kUEOnjKL
tHjnEjc4DGT+/a+B7g+zrpRNFC8AVltvJP2tEIf3Tea65QBYidvEh7RNdpMVUzrWP3v+SjKpYcFX
o4cW2HQT/SQ+unYRzwk7JdMlvhs/pi1hdexEsOY4+n7e8hEGZIG6kI5ZXu0L/TeebVdBaKPoYmmb
rzXrTn3S8aDhFuJiQe9KCDFktc2v2pvIbSYoAVC7VHxrR8a0rhpyy6j01VIUrnG4DJ1w7NRg6rHJ
DtmyaA3wMNJnojasoh2AMUo8WC9nPqf8mOG2hYfcwkwJdI+N21Ws/ksaDsolIlZ3fAGcL1pvcdED
xbiIPJ8/Pj+V74jVKV4nxyZYPbnMbk2PeFhkfHWJJO/u+6JQAAzUOVmL7Ih08Zv6WsXUu7L3nxUq
x0ThwwJvRzl7i1XSOXSX2Q/cvZaUNObg51wv8upclsxSIXxAlgTI9KI2BPZ8R13m8ciKJKl8BAcl
oQLIWq2L5jGcqT6z5CW1V8xbEcWSaDI9Zhp2qSr7IEhV/dbSTvr8Wv/Rg3O+DDWIeeSxeNVmePWb
4myA/ZHiPEIrBeJAgGqfQJVTqRVJe6eQH/khi5sGaJT6kivMss829fogS7cP68FO/pf1JmMgqR8f
Q6/eVf3obsOHQbO3OO3CvGtBRjam525iG3al02Y+XWkbVFKM4CUsqAOH9/ukIPAGai6ixE/0FgCG
3STKbV6JpaKwyDEjNFazO2H8hfrBCWMT4249rQhYTvzAXSVEm15mmdEMC18UGkJQqbniVc8oPLGO
LWi0V63yUJbeObKEW00/n52xmi3b3e3YCAoH2pQ9pk2CgAu8BADLFBHA2+3Q85BENvxPvjYOYVEt
tMj/agXXWMNaofNpF578ibuXUObBqB/FhKkNYlbJIrrX5ujUALs23/66vsYmvCI4gzsMyDeZUQpU
4iJC1wOck/I0XlScefA2OQXhmxUxlTgoML1zWY/N1sh8jwL1vpI1IaxqIVK1LahXQcAiA1OymWob
zBcfk9S7v/YJgtedUbim7J9hZnpgWB3XtaY3qNxMt5iaIqQiRKP3JPHM8WuYYUVUZNSEGmbsaCHj
+XDg1kFxZFALWP1zjiRkfyyvJXR9RvEAUUSDfroUWWIphw87x/l7bqfwDQ7wtBrmbxOwVFu/TX+2
St7dbr3+SjTu0TB/CekHSKrsx+RXvz6nTFAar4AC2Ve2jpLb8IXQuFhZff65b6leTTxYSb6qjtMh
SYmQcNaTn/WZfBbw/MZAHt6Zl6zRBcZyNNAM5XTAK+2qAi1dkVGhw2QETktAAgNekvLxuC3ijgfp
lEpRqwkPwZuiowMtAINhhg9mEcEJYHMQ7Bc9gRwdlgjGnW4CgaaVdXNl2voJU4x+FJrU9ypqDBnL
c+tDX63oc3CuWudKlXOduJqPIGRnrDJK3fftnh6fgVrdVqHPQfy3uUenw+m8uJLiDOhqidYMGQ3w
LK4AZQXggDcq8UTE8N/7zxdfPIMZ4MfqRnugudXKzFX3oe5HkoWdukK+yKx6vuZHVcSkzfDJJa+d
ajM1SFyXaHTabI8P5iYtW5GMP4NLBYQzIxofQAk/SsM5jfVUN+1oVB2dZ8jNRQap6Ljg3Nww+1qT
0fL37vq5tdfqmp4OZwY1d+MG/ILMgEPEbYZysvoBlPhg4tQQRvv92oUr7wYwBpXQEyfvl1k0kASP
/3fSLmFAVSYvHrAkG1bWAu4gU+1B/FaHb0S9/vB8cfy+rlP2PlGVvblLDsUjJaIad1uIh8wlpkYL
zFmlDc5X+Y1gl0yaLZ2pb/pEJBsWLxc6AI9RVS244U94oE1IjV/e/zLPEHMAEe5zvnmlC+mbY5Ig
/bM1z2Akv2wSLi/u2naIy1K4ipUtzoa5H7gmMx5Vj6SZEAUAfO6MR9gTXjECOYfU0syKaXQHBYqo
7AkD6BYKGkdOwWTpPV6i3D4f/c16sYPpYczkwSTrIhwRid38sTtz5Cb/BabFsv6JliMCQEdTA2zf
DrSTkqbzvcdVMvmuBr0gSKrYgW5ZfRfeRjxhlFDYcbqk/IENDmLy+WiEphDgClCmxSM8Z1C6oedO
gEzmUxSXHC6fOF+e+cO2ZByM7ezMa7D5KfsB6XJv7bZjLdo997xkkBpiKK89Vc1+6kodVIySmhnx
SXXXg13XchX0EOYzDwgZx7tGwkBZuboW79GWpNGc90uhIa2ZD7LKs9c+uq4CrnMGDveBv126MqRd
fK1bxez7MYXwW3YLxZ3ToYaWQl8Qo2l6TdUxu1b0gm9euP+CBEHjaEOjIqa37RpyZf1wp8qCMBgO
rNFKbCxbrRO4lzoInjHy4ZMmsciSA8IGcMTGdewotONuRrjERg4U9F2LLGl1UraOZE8tEIcwVZuO
qKa3l0xevoZCwuW+cT6NfIUc6nkR8dn5IxUyeEaClS1HIllOaXhWQ+LeHnKtoHR8CEydFgXQgyrE
LxsjfhF2A1M1rR4l/o6/IH6l1HlUrptJfUN8FSBHlcH5w4zzki3uTvLf7EDmgWw878yN6Qv6Q9Dk
bWE2/haPIm440EpJC6GjX/QuDdrx3DOr2o+3yD0084gV8087UEjxnMd6yVVE/84V/LMQgZRBXp2i
jDUU8Q7ihYZiCSt/mXf5JbMTw7hKXstTQs/nqup/rHm0J50awH0D1BsNsNxGrjG7452gmR+/hi5p
LIMVrbtreyeqJnXivI4NWrbDF2xNbuVoWxtE6AH+nTcpcAS9qMjNouQ82pFoCG2x15OkcY7TN/5z
TeRvQnUF5wWmsR1w+t8wEsAbpTXa58zr0jJh3G11W0KD9m5R/wu+TORVB03jwdSGEo+u7+yuU8pS
IzVee09OgYgC285buyz43Vw0nNuAC9v/jVPnJMGPT7NxTqq0DaAxJ+2pwofxxRW2lj2HHlzhwU0b
thxqmvqpbddw0cAEJL2HfPYyGN98OMkmNcmf0sUKa2vHPyWFaxzNPrtLlHn8s5Olk0PBMmExYMQE
Nj6s2ZUV8Po6PR1DZKEnCMNqAW4+ZR2mImWnZJyZB48ClzQD6Pc/pUZfJd81tuNrnCvEC1454tB0
8vTuFgw0xXtcpLCAH9VJLW7KNlbVRtekzfcrZmvWwXzpkHr2Po4bxRGbZs7rSTMjTHTdfLSVRJry
DPMD9oof0Eu8XAM6qzyDIzmDQaOKwF6ll91PqmEOxdwVrotkh8JKbxTETNsRsr1VyaqFNM2eWrlI
2gbNSpAR1lO9UXMmNbtdk5xsIKCXZjG0qiv0Egm9ACP9aEf5VOpbdft1jRd1xBaj/V/pzF1wJ3zP
L08Jx850k7S/8Uwl3FysebEwt4x7YkKS5SjdukXy5LEU2eq54g/73EF1UNusUVVxSKadadcZyC7h
QUf1kuwZvKw4Mc0DUb8MHO017pkPaKCaau3kuGB/6BtVxfjxoW1lYWwptXs9SUjI7Qd9mDjgxku9
KVmb+QhpwzGO3pnnkWjeXJG+lwkaob7j8HRGJz3mnlgRNSXf3gaRco2v9UaA1jGHrkyzFBi9BaZG
yYROGbdbpoKR8Z3ZWjCA8AzwJXHBV8mqkuCvT/6xL7qZwnRMWcz65lTmSLhVGj/tUt9xSCoZ3PQX
z1+FBatPRAIyT28gs32OQruUTDandelz3/34Zhc1Dopx3yMc2hbXukSU3tACYiNnqB5mW8/5nH4n
CPWcdmk1PcdB0FG5iMnEaOWwObyaDEupwffC1kgszeeK34O9MDdzvL4QdN3mCnohJfffr5iMNbZk
y708mHFIGQroZqUt/V+mBxiuj+ZC4Seug9Mwpm8W9zxI6xNHw227cT2gwl3OIOE+Z9Cc5jmC1iGX
2QSe4Yik01f+5b6jmcg/2vyPvFGmufZhOAGgOuz5gr6bkP+Z/dXvleyXK/nY1Qn02Io/XHEW+49k
xs9fM+MXxtY7WYDRDs5GWQcJNRowh7aF8Ahy35X/UVjHca/uWuO0HJ2KE2+XRC6ZxzPfhuuj+8IF
F86yUBa3r7Ya5e1mDI3v6m9bRC5I9HO5njvs8a4oKc8pAko1DKXlQA8LTrzX7AlosdnZvmd9jwUO
guF9adlNluTFcV9MCcbJtD95AsWJjCY7GUyCdtpiYb51HLDSDZ/cNU/VFR+Gitj9Bd6LOs08+NuB
j0CfLSB2oVl4zX5ir5/61ERx8Sz0KKuUCcioqDuFyu/6TmJBF2sz/HOu2iN/SJb7cdYNycaJWTu3
mHtm+yLkMM8DeFeQT8Wms9ZtpDg2cPP6V5cBdsAVc3qdPdHHXswbgyXx/1vcPuqWWTiEd5CfLqPZ
dSZ/VkE5fqUV7XYNF4iQteROdYA954+faEolOFcYDZJ4NgKCv5d7eWKfkJyc7Rc13Fb7rNuArXpB
4Q66BJ9anPASehH4v1IlJ07EUh751gw3FOB1aYTfFFeBJgeBGl3Mu1vNPMB4Sve5yQ4bjk2ZvMz8
EIOAAz8M72rCyx5+u3dqymF6kMpZKdV6r6gJ94EKN4JZYzZ3yZ3RG73gwjmBDGim3kxjLoIz/lZW
RoL9Li8h9GdgWd3CXaFfn9DhTYJ7E3QtCFoa/51c+tlxJxYXUXMWf2DSl7iUqMVya+K/VZsFU70y
mEYJSzslFvQX+nGn6b96hxUXPmOGtBxCeV+gRlXcMpLW3FbhCtThb0Jd6f5nFla8Ib7l1pChoz/P
AbpZJ0+yigEH8aiMgG1i16DK5VibOWBihzqLHp6YWcXHn5xyEFjjAYZub1j6e6bFzWtQx5tpRFqf
Rj/b24CUCXDV2O3fN1FB6Qlmjo9fWPFjTJU8KwfVeDmQAMK/93fNl/ahU5tpygm2ssNi2WSoRoKD
onJF24892t1D0RkdMHxoQ01DeoQlcK/NGV85vqmNDxpe3kjdALHa8bsM6MemlabKOZ1aE6nLJdnE
20nZsipuaEoHRrxxgTvH6Du+RwAr4M76oQVmaWPnrmfFValI1WtWrRppoQIn5GfqLlHdHSHOvdOw
MJ+ZC/6y7ms/zTRShYYkBhaGUFzbirhppuh2Vq4l0tf3BwhfRfaKgXqrv9e6jdBnfBRhEToxjXAJ
ObyiK8jfAu8ADMUXgS0cCVnwWwLgUmtjxz7mM7dU/DciTIzjoRsxJK14cFd+8ce78aaHEHDFGS6r
4lx9eZ8pVTpmWr2IQk5tMhgo2qx/L2ilNvJPRWyNM/dSJUXSE581Ocae7mHF4Bbt0SKTMhtwktVG
aeMyoCCFA5w0PPsoqtsO0jx2re0cKfUDkFQv9J0Einoqzeq5JwUhFdqnm4XuAmfqIGZbiw0cK8GP
+f/sPiUu2JfqG68prZEVo9VglaJY2QvMjbZOb/OBHh7IAjHoPXF+Jbxtc28vZP5xfBmaklUWKM91
/QCsbm/UR1Z6qwa8dbdBmEiBRf8rUM7vIiPNTDGDM89/Tdj3EKCW6xDEn6qBDic9Z4Zw7GutlgyF
1Fb/P2zmF0Bv2jwGxHkKod0U/+A8g/TVef7hgk4nRUIqna3A1DOQKKRzKt/pmTVLSr4dcf4B5yXD
NQe32TUDJtYhb+5U+oK4JKyqHbiXyeUJZyv8lFnwmScx/aR5VXEoZhH6zykFS+5MN9uvHFNL6w0H
qGH2Kqxd2Y5eKlpC+N79NhzAVj/YOE+NWVEfROByjcuzwOYkPfAlE3ja4HaIfcXCOeWZnnZyhKmB
y4JCIddT4DJjO8FijrDhJlwkboddfZJS0Pti97S5wIu0EeaKK+Ftbg6Q0OVO9h4kGawI/Ioc5h9W
n33ZFc4vzEtGlXGohdgQHjjt9+4PmUzEWoIvq0PwWr9gZl/iAtBwKvYl6G4nSIAk13Ms3WqONCpa
BL7Y21CSZJsWJueozgqpiJcztlsongzijEs5lV6LcTns7GP5xBU17CooXOnUSQmd5vefqzzVfw5E
zKhPHgMENjT89XxHPsBJmWVTZDYl2RAKMTGCjrAztSh+K9ObqrztkKIFHAykiLDicx25nGOc81o/
fT02eY8Pialyxb9jt2sD1VTGKfT0NLF5s5wWTutmgo//NnQ66eGA+sgguP4Sz1UF9TRI2hHK1ZAi
tGKtgl5TQpFK6NBb/p1GDVnlW2ayLJYVdpophTshioHDS7Lj3rZtKrubHIYIM73pRtqA+nB20fki
2fqNgDtzNTveHlRwDCr215BEhR8Ghy09g/NQ+RDaHh8FopfxsS7iFdH9LxOEAsyVVe2NHlf7hRi4
sy0Kt5p12UUaggHQEiD6S+grM72c7wqvIeeMo/9G60AYhW/qYQgFlyXFhx50fyyNzXqbzqvMdyXP
7lyfSrEc5UE7O60kBCG+DOQeSbh3NQCu8R05AsQ+f+ADuE1UUVm+fHw/wN2tenR72m3TLEEMtMgV
ys9/3bZ6rHOYKIqOVORYGgo3eJbObTfIddgetopG/KXO7ct6r2k/HbA+e8VlGJNGoquLYzXZCEas
A1nixL8aRHrt3ImiZEEuMWmXdSjfFuH53leeTzUEDVntGEXeWLBSIYVCyKJ3yhYxDq7/8cD+jrMe
uGupZd+KXeDRf/ilqY5GMog6Ibfhp5rOZ8rz+xZV5dRLGlqRIsGV6iv/qyZhmRNYulo85W3EVYFy
YiytremQtus1ydjGnOq6rNlwdnbPW94tGK4uh2Di+1D09vZJ5No7Mdv769f4+cyOl6ZpgTs2MNSW
WYJNWr3jXWh/Xa93zohBWXCFpNZ+lsjQgZ3ltzO9hYvBkrh9YH8IuE4OOSxMnepzq89ubSi/i6Qf
ZXfkeYW3zcqyPR9VU5dJcMLMghXl6tOblvB1G9TtaZEpUbHgPV631R9CT+mAKnNdBY0aZf4DswMp
VtMaqeX5QM6IXVIxH8mixeROiTTzsoTt+NsyaSZqnD9YbJh5jb6Znamgzmu47XjtPFkF77QW21z6
Dz2GL0McGWsL+ooezGxDoswr+I7dq0TnMNWIyZBQs2UbrgjU3S8OmscUp5dDRSQ53axrtJtG63kk
0PFZoPxjK5SIeHRHWWnmZV/UdOgV+1/ir67vQfg8h70EGV0oE/y4uyO44mgjeL//bbysGAjprCQk
I8sxH27kZzwvoSsBMOGFaYowVudyY4CFFsavU4B0GZOBbp8Y5Tggq8X73+q7/0Omshj0qqB2JpqT
EzZQOedBjCtm75YbRvKcoLWrq5vxYGvpBU9EVMjwFZ3/RsXklhUlZ9tNMVHUZBNpP/h0uYz0hDPN
T9i6Km//xkFegvgsO8iLe9kVMepsCv+QpsOG9enWNTXx+xE48Q8/l9t4DBGJsBxqDxqIOnkajuCh
9jsavs+pJ9r3IkRGGVdBgxa525ma0m9OXgQo7MOIedAHRBSiRgh8F2AkKN4OiQ1jhM5nk4yXGXBe
vVIvCV7CxuKjJX3HAvtbrRW6pwrIqq0qdjf/jkM2u4zoV8m4kxUhpktB/Ihw8LJwe2yxiw/UHabW
oN9/WJOqzZpSg27i7Ae1uL1uDOO6OIHy29WD46JShimeO/OoGH7dZRv4RCSu8Js5sxytGeVnPFWR
eCojpPfzhJibsSp1b4SZSDmQgtlsU3Pf0LdcJMsecAEMGIfN2xwrMwlr8BqzMfxP3wl5eAok58yV
Na5tTAYOLajB/MJ30z15OMeo8ho515fUUwAUImMHYliUTJHhpF9lbnUzDAQUPyBoUmO/Iv11iQDM
ZsccmA6xOkDexVDIbsO0099flb+X12SOzz2vPRdKwMB/+/yeo3m3zk080pEMJfVJ2c3Ho3IeWox2
+LorcjFF7TLWMGvP+/rT+npUlTLtmTochmR/rZJDWKbnBcK9WKTDNfnB3JJr1XPEma+HmsQDSvl8
8hTXB/Wpy4KtCS+bS70rU/kgs6ykGLHCA+InT+411L2aoQJqO3oorT60MzKjwQdbrxpJvij6XCVH
hoMmRek6kBZ+lBDOEN7fY+YDOKsuq6U1RICOGGCM0r0bDtEWNRbX1bF3NRyF7zAqpB17CRbQ12Qu
QlcYqLpuxhgyrm0KyXferoLLRa9+axvZu5rI66Pbpp3EnI6dezvlU8i8dcMkMfEJprt65PbL6F7G
h3yN4GI/dg9ngkaijOImfR9KI3Fl9Mod+88Ka3W86thyrA4GZLniTwKpfv9FcUzjfKtE2DYH/rbZ
b6kNmuJGIg5BriyonD9//IXwTDfV+Jd/0F5PiA1cgML3yd3uwCYKoBk/shg6KvE+d0vnmgVzGacf
6ih8MS4wO/c4BeHS8ZNaUFGOvcagtfVmACTTu08oR3dMhCBo0PEvlojxsvQdxQTAqI6afOmVA3WT
4yT6r/tQ/A0yzqE0oSHGUBfX785W09vP5YymnMTN73do0eqsv03DkIE/BMT8JD4nGOxBalL75cSP
E1N3ei4P3kVFszBnl7J4ZbItsmyKPR0ZtdajJbGIkanbSEAYOuj2e4O782h1j9IHi/4gwov3F6yy
YK7Ik589PQ8K3IXfVuEx/xG/zXdNglnnbpZDJ1NCXiaonqOScL027C/+oeAa5aByFXrXpGegDr9S
Z1pQ7szJsY8W81gfcOCoeNDWbP1rynKy8nMdOKiyXipNYXnbm72jEou0sMZc+MXlnhAy/hCymm+z
zhw3fqk6RBzQDH2NRba/bzZb3AYbGBODp62+hg2ydPJADUwpktGBZSAGkWaVwLOaJJz1ammUn5/M
lWjYSr8AjMsUmvzUQ10fmuzrlhzgq15WJhfn1Ytisu1qnBUimySN1YOwhhIMJt4ZSz5HDox6EE9X
on3kJLfQYbsj7FaqV89ocP6eM1MlY+gXy4+EWF9dI4TgPtN57TRmXKtqMcWqNX5VBOUVvj2+hIly
s/72dKxmjRYeDWUh+qym+Bhn/iQ3iBI8pkXcyH8SyrI8BhCVl05j59OyXRoCKvwGPY4zc9HcDg/1
L+SqlAlIo797TJer/wFq9x+zRL8tBFS4gBJeH1pmYzPQkH6a1tSDJTShi1sL0FlQaX8oHRH1oCGn
sTQjsVd1Ns3n1OipH62JxpyLvTMUXHf6SQXNZres8LGPDL02jKF24meai2f0BaX6iIKYlM+2UHV0
uj3/Nt0LuL6+HI1xPHYTMpKcOmdhMdnKzvvhxTAq9xP3/y8ZXfphxgm7z+55UUO+kfN98nzm8dER
j/GtOvGtwXmQlYTi2mmlij4fPqjnem8RNigMcikANfPzQT2g4uVraRD1/M9LcS/1PUpwL+mOcjNN
EF2NlN4O2kTwLpaFg5HGwuCXogoiCpkS/RhYSoQk6CTOITI/uAKHfx4YzZbK+yLxe8SAYYkoJQNO
gTqHLucwGXh1qa9X3cok7TQptFe/v3BHQHSoF3XQ1SysYsKeIQLmKONRAxfzLuDHJbgUMoLEE4gi
oh3VpZKndpMkIH8qAu8/BQ7+IuWU3MZNl7gNx4r3OyxImky7sjmTwdDCCab3r7VrVwoMA3JJkRfL
iJZgmhnZS7my/ZpknBDKcGfFI4tmyL4vdUuf+fSuzaeuTzH7YpQW0Oie3mq2tqgzDTgv6cBg/4SE
O4gPLZphOpS92Ueg6v/haXsG1HbMsq4Q1YymoVJo2rc8Sj0YzyMKUh+fS1MkcFwqZpIv/n518Qvr
EJK4GB1Ag7VWaiy9215gj2GWPtYEJyTUcaqlS3IYEEs2FeL77oJnMSfYxNr1waOUuWRsfX72b3Ue
vyBSRgwqVdb0+n+FLmrnrtL8EeyMlGsv/T5cmyaX9RrmpHEOldbWHftU0qkxcZO22dhKVgYa+AVe
HvIvhKir3Ll+1Gq0GlyCj2hKj49kchxcjX+IL3uk/CKe4NzCF26NCtaqWSoN6pMASWZlR2t7IpQI
CT/WtFQ1bEpUQ43X59fLpQdZZZ+gSxUvEFn9hgYNpttew73Y1mQJivwR2icchrZV1Kl6mWn3QX66
fhUlYQeoesnMQiEiPav/vTr7RKJhP0kHW0Qip3Agq48S3pBNdk0gQiG5K5XaiOtClgSy04+kLcR/
surkA6IbJzERekEotfOG5jJaEcvS5oTTCC5766dRxOGYkprFC06+n5RX64GBVZ2i6TxAafqDVyRd
71NiH/VcVtdX/DFQxxs74aZqXJVxjDhVzZCfqkWzjhBkkHlkD/ddHkrHda6Y1LG/5bKYjlQ774HS
2FyAFE4orpxKecMgi82wWFk1T9twZO8it2i/Z/XMCHhf0P6EvDwghOztvkqhbTtTc0CwQvGPmO5Q
kT/JdWi0nmkzgFREuujW83aJRvCrWbMaFs3bKjvUE6fLBZnrGn/hG9uhqSOhIuEVg7yARp1t0uhB
iW/JGwzJrE/+9LeZne0rSa5lb18zgrmVc+Y7iFcxF0fVHKY820ZDJt+KfYjrrdvnc3/pU8fIG5Rw
1df5K8ERZrEaCkki3TmnngyMObHb2WRsj5fb/t+whjnBqtAsmq8GJ4Mx0k182Baq6+rOBkaW6eny
YzLGMNIGNB7YzAZp8P8/pjbP4qLJeQ6AE8BUTiOeqXFg5Lc37PsebcnO6b46FOHyZJwcsGkxNevL
BsEzVOj7z4NqMHL7lDi8r0ghgZ40TB/87+K3ianbR6ZwEYUZjGDybh97uP+J1k6v+4FfSkvNmpi7
l5pMcwd49lPcqW6mDdl+qAtiCu5IB5SZfKSKVDF0bU/IcGCo72VFbuD0mvBiwcsa7hDLCnn7ymSj
g21nD9A83gbCowHx9ZIQP9Vo7NTwdk0877kOOhjl6QFBPuJCZbf8FBWfM0XEeMdEFfoTrDTy9Qys
NS1QSp5Nq54GnCgl883wYCJq/MN9bqmGw0l+Y9GMixw4CXYe9CbvgePfBzHHTrpWWiBZJDLb4zGV
a6pPZUaTQRDnKWgon36JgQQIggP0cHe+EEDPwgWXircvAYbqJj5JpKjeL2qgpuaCHmwLjQUekYYL
55Y1QRFSb4ppMonZF/Ao0L5/O8VUHq0JF8ruTtiHBJyVAHS/hCBCAUAsD3/MXKorcmNW5aCZJnJl
7BWWLXYYbPorl5yeTZRB9ty4aCAp5436seSvMtE81Bm0GoDse9vuZUHz4nCNuDkEd/g17lYB3k90
Xo5Y4Ayqjo/l1a2y2emv8kZ+ArBwqF01aczPztG3ETm/cBcZgEiKAdwqXKOvXW+FHuNOeixwTQF7
L/EmSWLCzet2NAUTqHvaWwvRP8vTqbDEFzRqBzOIuP4JUpFUEKdTtv3eJNpMyz0th+9ta7s+mWAI
w6eUQy/5iBQF9LYtrdX/eloQ2C56ubpq4ViCYrNaufFIOrMs88q24YuQpi8daMxUuQy3YSS0mErI
olKjzVZZFOLui7NjVGV86MpIBWTgNRwloicLzDrHJJ4BfeHmy1yFSAzV+Ws9gHOjzZLfDsaZcYKM
yiq2OgNj1N81XFBW345hFZqdiKaiZypOruY1gQm6X7vYKjIgPMaNn8DPY1w1+y3qWWkgIWnnmwoC
6vqtFScQ7+MRJSpO9Fmc3GQMwjzr/xADZeMIsBhcYCeoCcz7SLlWwIA7j6D0VFHrLQQfAvnuHAxV
5DI7jIplS0Xi1px59EVDJ3sIc0/5ndRdys+adfiG+2Gokr0FchyTlBekCxOYWoKKqX+LBImaLBZZ
GPh7Pla4X1rAF762yNxYus3y8D/2Y8dWZ9SzZTfJnkDY+0xIqqfrBPaBOEFp0Zh2c6LDpOJhDY5N
yzYAh5P2GdK0Zf6CjQjx1BVqIYXB5plai1KU/P71FAZB+tdW9M0M2B4t6U9lB+xHemOIuxkp/OyA
hcOxD6+6HmPXuowPE3Nh58pKizN0DGaji65r1hCpyvLsfzotY1dC5Mt1Ll16eemftlmZFIzJoMt6
Z+WWo6ojEg9RYwj1w9kybtIb6XTEu5t9S0dJQVXvCsw6mc4NfrmUuqt2DjpfGW0W84Mr35L0nKx1
hjUD3Zlhl0EKxVN3oA1UyH1l8ppPM7YDsabQD5LTrPNDKF6mtmJozN+dkRIvR/hzBJjmRX7nATXd
ZECt731AHZDRkKATuZbQJr9IM4y2yvOtZE+k7Hm0+C3b6MloEkn8+0mZfJ1H/7h754aLFcYcNdso
Rk6rLCAgzhFpN+aA/o+7SQ/JBjW+JXDLK/z+YC2yaAyo5AHZDI9EmGb3ntz8crkXhKuSfbhev7V1
PLrrGnaNPHZkVeeI7uN3DzqECNhOe5DAclT9wsdobTEKTvqOe3ff3oyrG/cCvdRQzM33niJETxtF
v12/f3fE/+McfY0cetBIzFeG89YgEXE6IUnXob/lZHqUz1zJ1CEbXkNCS1tPY6fOcl/KCoMU329Q
SiB3rx04DBdrn3BhP49zV/5pwHP0jJs/Ucqv8s0ViYAtWtSdMXG5aZQ1CY6ZiseVAs8ISz54tWZW
SEA6+B+SQXoszGzoJXOSraBbuDXFnqn0DUEUmTx0MzE9jL1ewmJIyh5XorwcHEr7KzfiJ7ziUxQY
UH0topvJOVAx8qy4OsXWRXbc+oTB3uSH7EUOslAzJ93SiA36CWAqwYRCqnez+I93HQ4S6Xwf93Gf
hEGLbW8t1Y4W1KZ58wBTE51BxgsF9oqaN4rMYDq1HZB1LNbxPH1xaXCYFVsnfe3OSj4HIu04iabp
BXBvLvAGWaYjI8Cc3dEf7vLoXcU5Hwhcx1CtrU4Oufh+EqiQ8YLdGrmLCPRYRCTZIRcwcxJJOQ/Y
JQdT2pWaKBaOjxrQ+PzNlgQVV+raAV06oo2Y1jcZQB1ZfKjIe8Zb4fIq1cN7o8Uzf1sCh/2iuiAS
VlJc5avvmgKXKAqt+KOcsdVkruDQMQ3bl5GAxX8i+9IA5A9HzQZc+kCQypJKFd5fi3uGEF1f7ZEL
uZRi5hqb7z83UHaYkyihzdRNT70b4up+VKbCIzeI6nHwehMKsyPnojyGoNbWVvSXlYtEOBtCa3dd
/CKcAfDFM1xWwNingf482wV72JbJFLm/i6BWCOP9nlmFvnU60TrJvfzBoG2/x32KMa+h6FzNZ2gH
HFRDsqaGnAwVmbG/eu4tlYYlWOEwAiRHtBIW4jnN6nxiHVdXPFWzVDsgUMsR0w7pxFOXPaiIhcGB
r5aCag/waNrK11SlwDQY15OCl2u5RyfmWrZJHrEZUVxLUSutYjNgLFhBNO+0gOhBTEDl3LzRINhl
ZTYYv6E3itFaBUfaSBmJf9+ZY7+/cNhMDMvuFITWuhj2V2sLa5xkgmnnQv57LradJvKiPPZcSnwV
ecIUoq7/7afxJLSPDozntsYRDvdMaMv2zcIfpRdLob3s36xtWSPeNlaelgcszXYceZtEQ83KNjmc
MDJbVifdGt+RhUbPYxYFkJrwF1qD6gVUXRVmqbuTQHFGHjUCjjQK/zW3mkIKyQHa8+O1ERocBGIB
JWD/YnsNqi69z3xB7z/KYC4gDaBmF4cghIclSBXpPJDWt6ial0db4UKAWL2VaHvuNWSFZqlDVTXh
5OsfCbCKOXGrr4zVnqxe8n9XDlSKmQtGzMuO1yoKN5rDrmpAIjQqpLD5MN/wOyWMXwhwglEu/PKy
dJQ2kWuuxLnAEJfS6RUJFe1c1azZm1oYHycK9Ai6rBdVFdy0W9Vwi5QQ+gv4DaKmHscqUFiyoEqI
Nyxn8hUlwmuvHTCMZ3/X6wZMsNZ5K/UkbRa5J/qxGhGBEn3hC6OPSx6k+5HkHuvzFrTfcgwI0IiU
cfz2dQplOsQ048doQfjBTw6k3nJsJAuC9S90XdG0jYshJrco4Ys/mb6CvodVbzUITkiCcyERZTop
tLoLQqot9FgkeYGUbEn2qBKEO3IcpSShfCLaJqy7O5qcFfSRTkm4fah8CQu4yJghUESk6yKrg2k2
Kc83hy9l9MMIcu3H6WRc9gfINQuY12b5n5+d89p52Ky2fy6v0Pg4w2zZrJdqrfwXMywYd5oXdwCT
CaLiniWefDr76N+E6oSOW3XU75NYk7LORNJdHgebGnRNeETmkrF5AeWmoBgHGAMzU9NCl54MIW/o
7dlRDtVtC0f+iey94U2quF+xdgvbhkeFsjNZc32W8FKXmocp/aLa4zx/WLHVAPxN9E0U726rmVAP
/UpUTFgk5rMAjahSmGDMeedwn4fcNwnrJ3PpmWrsUtrUCePTZnyGkECWQTSatgmSoZvtPzy0KiiU
PaqUw56K2B1S6iUfAdzF73b01vFuotZBWQl/pGZq+pcl2Ic+1wmUQs84f8ac3cJm1MyPhsOcJm36
/9ynhCmBlTHJL3VNe4dv8TDudW+vW+cCMlngxTYRwRiZvw6QKyGbfXYoHgQEoyghW7BmVr0t085U
5Qe1qW1Et/ey1eblcdJyXHYaY8Ak4RMS82MMK5teek6Auj4PPKLdna24DWY25AgIJxEvvQUiPrwd
8JysRhdgO1G4m4OY0Gubx2Gr3jkcE9y8hvwmrq7aYipsHYjLrgTC82mm97S2InTpG7/msUURoYok
DM2lanSOvQJhmOcmNKkAboFv8hrmUnIHkxZ661EjhHQSCFi1FZwgaIFJIb4EGHWsHeiqhLfy41Be
SDI9xjF9oGC5/ESLciA0GLUUiWmg68nAFIbuWTTADt14tFaegltYhrqp1ZrPJV4q/RB1rXoldLbE
IcDD/S0DMMgQfOLPekTjPx318jtvrJjBDNBphqgiGCFfyGQkkxlGlM7927dzYUpq3VA4J14kEpr/
qsIsklfekEgN5IdrNmYLHqZVyIk1OEpGeXtKaUbRwHNTafQnjj7w+GTpQziR5jYqJAXxU2PpRT/X
N0lC5FKRlzrOqWNRXm/oXd9KTkak+uFyuONn0ndmOoyQ5dM7eIi4qSiVCk9EvrEjSpyIg9748Cd4
6/xxlPlhmMpNmMwlLbwSxsQLJr0Oe71dWy2Sd1wsNIvvdkArBFcD/X0g+g4Iy+GiKzaXbyU2irqg
9Y+QfVYhjw9o6u+1zYq7D1X+NJ9C+OBISkaGJ8DIUCoK8QQ24QlaXUO2sAJvS0POIVmvF8MJNUEW
SyGMfjYoVlbAWFtLgBg7aFjk9WQw7KHrZo9kKZU3xSWx2AqpHzj3M5/PgikGvxyoF6LfgB89WeRA
280UNuX3rmP2MneZPUaQKw6ej52/Zsu0QwuNZWTzSxsXYw290ScFYnUC0y0ob47avPw3UwejVywu
E8xuRKzxViF+ctYV7pr6MxCm2kx2lkWwfUIVUeZJ/nOGCLn5+/Wiw1PG3OdmDY2ksgrNwULCiF/w
0uNixSxVQcnJUT1o35BfoT5PHu2blkos93j8rUWXALZHaEMS7lmWFH5bB+oyp/yMZs5Ek70R9uH/
ESGBoE0dfn+Tc9OJPc45mfT4KoN8GB9xIrCASAPedRnLxYP5NPgJFVsVGhZtI6n7CwSPkRki36pc
QeXlGKwiQ8OF0El2JVF+H2OzaqCdyIbNqMhd1/jwGR1OR2D/CS/Aww/WxL2hS2f0LP29owkSVPHL
ovwFc0tsD0UP4S4dor0R4dmDvs/sg5UZc+seFm8OZhIp9J4MUQLp2tbF9yINAnh+267aDJwmDJzp
3oq/A8imDLt2Kq7KFVlog7k47HbnrTlxQ0XR+TvdUPPBUHT1bobYyInRFwzSIj7vzHZOwioQJ5Zm
3Hymu1rFJFH9Z6QJSxSGLuxbvIjmMIyZXoRNcAji+adJz2DgZDUc78cXNWFg2K7OURWWHFxz14Is
C/rwyP4gCT62+FvPFOK1pE6Jjgo6i2liwG8+gD1UrfrMmEV25UzElsFS3X6OULc2KQFV86IboiGc
gu87GVEXje6lv5VqUM38BbPcirJFY6FQeQDjoCh9ifWX3Nr4gt/ue4KDjIstCcpzqqA3Hxhasaf3
PmUiRZuQ53ptclrrEQCMroKn+xJCmh1UIu4j6L0ouykfnavHj/i+vjzpA2/Qktx/fdJn2LNKKc1j
1/N4/NUmKQIdjulkHK3chkTi1XaioGPRANNlaUaRsLR/5hpkXqRDck78iXYM6lsZg6Y08wJ/EWqs
xzGrr14MQ+upT1QinJfz9Ob/zPiEbDkEXsINo8rzfPcdp0b3dFMOdm794WnI9Y/qxctLXQyyW1aj
iYrW8xOTwZCxBTzfIWlcmQWW8azgdsb3xWf/sws/Nj/0zngwKGKvDm4/Dz57HOFzTnNmMHt4bMMY
2G3vHPxYd6I+r12MNMoU9Oz+9fTdnrgQb5d3tvyPgPv4wLwcnR1r/DUqYxuifH2bcGqjrPDsBg9G
/3KMAxvxjTDai9eHawlywflv1pZ9eUdsYW4jojR2spqNIl/Xambcqs8yVb/4PlQn3UTOh2LdObsW
nmhNrnWiZQV1jGIUIQaKxHfx6qD9VKiLt1+PLxZT6cg+/7XEMuwQnRNx4LtQXHHmL7LAQWYwG+09
6DSg3TW16fCKLd2YzFOxz9J6WWTdU0jWEyNFZf0YOc54LVBm7U1wHzKctJfFf+XnTvOb8zDC4MWI
qVPb5ryM4R8g4TYcZ+Wn5bjw664Bm5d5u1Xis27hO0T0cNGbbIocwlnjB9lwEyPGehl4+ftYUiJp
KGgG7wUdqfXkmnIUfdHuY0PFBvrD3QviCVAz0cmw1v7SSWj9eVdLbDoF0wpmc+E9vkJ+A5K7TLA5
kddpXjb8PfvYRvdBFSz6P7FPdQeI5N6PqkzuF3QJRCMRtEzuvAf8YS360Dt9n+Uk888kf8i0wFk3
5E127hXf61aETcDm8x9T5kM+U8JGaAi6zj3dlRcPKZUc3eu52t3o072QwO+KY2EoDjdzIRLTFrVL
7qQyvkw4Wf9q804Oq7E/8/ISvS9J2N2zemOwQi15wHzOg1W5mmP60ttSnS42KovowvrLDc6ysqfl
ahLKNw5EAKj6FVNqnTtLzQuus0amAkpnA1mMqXpmiaOzhx8+5YLVMqoVa9t5KWj7/jO44hg1e4rf
MKWSE9KzJAYDLh5CxlZx+Xu1LiEtcvBCqSywKGlclQ10/xlUecZekMnjhjOPKbfyq0/PxboALRV6
DgRQj2Y/nRX1AoO8dytmXD8nmZFPAEEBlvTNKr/nE2316NbqfkHVKqMkkpS/BpqZNj1ogh2peb6/
8vw+mDL4VX8M3u2WA4ChLtEB+tJQoZjsYQfh/UML9RsI4Ke5vN96ajhL0ONyAd0uBuWmnAWDHty0
xh/nzKFOOkKjG8+zZo3twqGWb8YzdLE66UYoWmvCNS6Qsg2XRQPfe0/yVkyWopjgBKehXv9b1VLS
3f3+g1imtvf2ORiTUKMaH1JP772AeM1+mq5BcT4UrbyyBvghTHTSbSbPRgP8AFymm9sKXrptERQM
4fFaCXFYVuByTBQx8pVzBmrAxBqwm+HcJgV3mFOECDKrl6s7B8FmryTfI/a3Sw3e+DWgD9MZsm1K
oXLFN5bqQb+Ya3Nyo+jfwZAbl8DVGiX6/dopFiBZ91hlRhjaYLp0sOGhuwEtt857aCkI00LHaxsc
6Xln2BfRd5cjAOBsqWMGWT0pzDYYdg2sjnERZ7AWYYF6VcivkT7Lftm/WjmOqKtBjV/fsrf+4tln
PHuS4iyZL4Z/EROoOQg+N8sOe9vqWk6P1RFbgfD2SSRh/FAqsbZLE+GDTRqMpLOqmOaPnoU3uYuY
a/DB1L1Z4YuEPxShUDT6TYPmnPbiwFBEefpFU4tzDXnmgQQ4FppJfm9n8q9GuzjuvnrFzJtkWW/2
GO3NvZyo5iKAUot/4f/y/fInzvQm6CtViCFK1yMOtAWIcdQh9icNReKWYsPJp0bWNxcTMAvTxqjq
rf0lDVbgvtja+doD/C+lRPMmOzbLUloxk6wJUaKKQEM69/BwtLkDdjwoVeoweVLHlZiTRDC4797S
gCZeOBDLBO6mk+UaWw28HDgq3xcLHF42VglJPAxRXlHslqvzCtrkWUtuWzUyhFea/GNLhTR0zsxX
ZU3gKShenPFSiiY2jzLx8NDtd9u52SkACgzuO5fF52OWgL2/7PoQrX5VZxvxYM67Qh6Qb8oFgNhS
baKropm+Tzlsc1yuPUHxrZAlUrDlNSO5WYs2WwDjX3jFl6A3FDVE3vo8TJzTmGWF/xTcDiwL/lDd
TvUuQ7Vw3GxVeTA2wZnMOepIExBfuRpQFMxEFVB+6eFHia9SPYTNT+0f4fyXG32Hoz1oK8TAbSrT
R3alyjZQNLGiEeWKIwL+fmNBPGvJj6yM9/fv9qO3apAcU2oLmI/kutrGIt8LYrZSjwnbhlxvvYsU
urqILOVz/qKLGzM8yl4pAPnCC2lblDbw//xje+zLXeP+cdg9n1AO+2OP4LaN8R9UoXvSTY8dAlrI
phsnour9WlUdTWi+i4EkjqPtkbNxaBYl+IyEYhcNJ1q2HOh00Y6ayljaxaA1S3Yxq6C/iNxyWS2z
A+mIucKB0iN4+qRzlL1iy1rSPOnPXhixt4MkJQCrtDc1+IVgvxw+aKoQX+WNB8T1zXXGgLYysr+s
gM8ufOYbS2ivWK2NnCOS1nfX+zrBNu6hfkWUgGAvoC9J0AAz+24zOtY7tROYisTDL7Q7WlwYYZDa
luwgqmUfB2XAOgIsCAbMZ/7eAgfFSUiVYDhY+Xg9aqIf5p+kG95wL+UPI7+DcprMvaVOhWRUzCLy
dsue53dWp7wsxjP1P01DkZXCiTyl5r5t2cmDxHBslWilH307ovG6uvv7UKcgpLIsx61lduH2zcsC
5KF3p4wQeJmdZoFJxV4GG6XUgAfLQoOLelNa/SGKNzSGYtqg9Gx3qGVHqWXXb+RWuifWXVBy8ZAz
3JOwmGRn/fCswxFpFZBTAhjXdgeYc17B394Ui4VLGkPbBbqB/GPbz8oZCSSTl4Lk15gKfYCrYLlB
mZjcOn7vUpn9EyPrQ2OBbqOtGTDc7uphAwLithZHtHp6zOfVMTQP2JDilhrQS/tLvxEd8glqs5tS
pWQJY09xug8CS4kcf7bnjmKUwS+CRQUrLbShm/Nfs5CCwg6cje492EtzE0jFxgEeoPZBs9RsFQ2I
M+3RNDLI6Aep4Hc4bJ/Tavtb9shxfuIHOkyVPl+X7kKFTMy014PXNIhvmoGwU7xPSREdSYbPjnSn
2c6vw054JcpOysc6X3sPFcniyGru7x2SlVD2RkbuceB5SzRkH4XRRVyQ4Kf6/JEZs47y+Q3ovib8
Yueu8xeggMUZXQyUktnNwP2kZ48cgiNwdNhAx50pIZhAimx9tTa44yLGEjJDq05DEUIAcilq6PTR
uR3vkpmC+WGifO/B2RUIbWfs4nH2TFtOpk0rMm73HAj/Dou1/gF+T766lI9clrZRTCg7365cWcJ6
pRQpZGgXXLFUvKmYKZzbw3eJrkWrE5NQra227OXoiUskkxVDaq7rJgmY6aGxu+KqhE42UkHLSfak
YUqUFALG/mwz+OootEx0JWV3cMWfpn74GMUoMg95Btg6Rs3Q4uVJo+Zo0HcFSd4pF4FWFuN+HNzI
8aioXQQu/6XamNSoJNLLN0E199ye9AgYDIe5pO969O+rScC2uVavDM7bqehTPLJISTSdDCtZdAYH
KhwjagbQLaezrm0o+BR0tph2X2WurXMoeSz+rajGrovun3Aqwm+QhhilVNXJITsLduViFxawQocI
LBKZHT+r/BNhx+TNaidjeUj3v+/cho0RFvL10FTOAtQb2tDGGVLcxmHZnACvfi51viDOWQGqpM2x
0JuMCpF1aty0CwAqGfx9HjrVHIfHtiIWTZ5s1O4GqhdsKVMUerXXOrm0VwcT7yLb0OMcZj0ao3qm
WysB/uQ8gYLxUM4wNksI5edqTyoE+4ecphI67RgwxDDRFaRhcGITFaO8yM/MMX42NLQmQRprsV/0
GQFgnp6GFzL0fNpNu+5zLDmSzWAEEKJ59V5wBgekAmRNKA7h8LfWeGOJzfn0PDVgTHVge6o7cV9r
soOUjhnrDd4YPmoFB5yLpdcwOOab9tbeIt4/HbatQGOqrzodx9fIZGKjqM3CNxEUT4XdRaUaESw2
l5VUx2iecZf3iHB2r4JbJ3jIh/NlgqrVz/5PYSfc9rm/ZhgWcTLt7XGrLGB1KAkYu73xpgGsAk+4
S1B3m6YC3IrjH5Yh4pUZr4+oLlhHAMyPnuO6MZnF1GzWj9HlMUc0ga9vfIXRX7NezEUpCwVIoAvl
RvwOBcXD6T61ltw86xU9CgKmIjotdOtu0rfLPBvoEuMYBaeDOi9HaC9D21b4kBA8rbk9f9BtM2yT
JS2Nmg3qux73bLP23OvOIb4hdZOMHFiVgDhZvTiXsjZBU8UiGZXebKXKu+mNRIh+4led0HiuyO7v
/LvMxY3nnhZG5uaU028HFD5neeAHGpK4lKJp8Hlc1bFYPTQAYiom6X1IHW2SV4ZupAazGkWMWRJi
wFSW6WRQsp519JHjVIASevJ6SEwGpTWLDeS3TD1PKoowxPIua6a9nV0qsfYOD0Oul1WOoIQwKhaN
rvxwGqCH6ySvDJongoRzCojObFC9MZEffzPa3ke8sZdgO8YjG+iN3ChemZ2eKJpYOAtesPZQ8TnJ
Zx1OSPseQMkIedl6W+8sUPyWTRAGQXfhVBN63GBpYCTck1JerOHnmaTGWnQRSVee30v3127GbdFw
sXPt43/NQQtJ+0JenLCsZyNvomML17kdPC8BSmT09ZSvsoJkswBq2TOw8MSPAph/7AEG7GbZ5+wi
JPzn5v7Yx4h9f2QSCVL+f9kR/zMxcyrjam7N1tFch0U+2Qk+RsB0L2PwKIq4/3XRR23GC/faQxaW
qPNX3a3aJcafCXxjk77XC1VlcAk4RL66+bhj86le5C39e4PACL8P/yNdU+encE/xX0z7j41WAt1M
7myLJPzZ10mVuzIP6/w5B54UAcgv3Q3bPbuu5PkpsLgFSvQaAJCa/flPcED7s04WhtakkWZm8WaH
/M9AI0RUQ11uvWzpDp1yXp9DDJ2Cp3jXzL+UHEh//ZUtbBNO6+bnzj/XY+AD8lMwjXYc41TPP0YC
kh6PEVJ0UgPw6iRqXVUYEQ9pgoKCPyWzusEKOP5Sr6WBnF5HoZJi61Cuko0c3+li3SSRU0qglwWo
5vldj6BB4LgTfwc4YJPtGSJsYR2I6WOdeLH4/gyXILzMBziFXVX8/t5JZl7vO3rUWSUYAl5v0KIk
ebTUNDX/Vaeq4wKGvDQhEgScLkW0OkCyy/SYYD+ASBu1tZtt6AV6eYRRQEx+rWyxGR0pEqGAyfE+
uZZQqQfsWFbHPF37oeYmUpFG8Egc00pE+14oYdOYv1sZVRHdOz6fhULQ2KJKPR+zLPYzDybyr6Y1
r/yedRwxb37qwfFvge0pfIQGfXloQRlNo4cwL4xw5oZz72YDG75+1nNtkIVTXbJJwB3siZjhgIXu
1BtrIZ61fzHn2Wr4USw4DxOsA40LB7MCNMUAmpJwCOEC4HQUpgjCq1kMJ8byyvRNeo1sEsuxUrOI
mUGbidWB1LcvVaZKjkGsfxHtAe8KFdGHMDZEKIFEjBXjBcoVVojOaWHgAzbQzDPRkhYPRlDkU8U5
iDjzGF1L74rR5c0T78MNTQ/Twk+FEzQxYizjFGE4bT1zwHUDuToHz34Mv2Jb6VVzzPaiA5zAqnLD
XIvU4/Xu34dhafctSBwU7Ac+gmAPU+1FQsmILYDVbX5hE0DcZ3XcpLT8nK7cos+kW5E0iC4wsSa9
6TqvDELZi7YuKVqA402OWBNaip2zS7cyQU7zbtD5F6vDj49mevu8MEN9iKi7fEwJmwzTW1q0FrIk
XoSWF/4Eo3k6ha1y262QkcUzDQn+1c1CwQqM1Urj53twgRnYR+72G8El6j7cgM3orHV+5cZl64WE
pPLLR5kgyi3ialBQg22zMDfc84yFEkAxA9MAB8qIkICImz8oyUg1Cr9qKmCwT7YPc8/cQQ4pDwJ3
zIa97FfxvEPDXpiHp1rT2LIpaKa07RLEh1WgZRR3YqcpuFSsitXywBFZxLV1vDMaFP9Tw14oWzgS
hL/kONvAfJUcsoXwi+HTF5qoDB+dRFog5w1eU8yHdfPJXTF3rxgyr83BNEsMnW0XMxcCmKvKsoMO
keBVpHEl8P9zRcUB9P2F7rTp00rW5rbyWSPk7tHIdjOpIrCio7J/vCVBmwHwZLSmh9ZTopslw11r
fPDbA1bE1PgeuiHsCmj8SLWdHZqD0RbyXOBf7Cl34KAN7wh/rjiuagi3zOf5REhLT9aKI/1YoIOh
7zHaZz8s3Pj8f57G0rAwZpkPVlxcc7m9Vp8FWJcpKE3eiSKDfUq3xk6Sf8z8sNIuLI0u3ftoQzPi
JVU+nJ2Y0Fqptoog0ahDdr3neOVe5h9CTQ4bvaw5qhTu+UjALk9GPOsgUjFdbldZjpkFyjlbaGx5
Q68VLjtd7wIddUhC4Ht4pYn4ywTUcCOI9DERlGxknbAM6rhwn9D/iK0+/7bk/021cpY2x3Wk8R7w
BoXMVbcVu1ba+eb/qgDGJ7mMnPS//7Oho+p+2qqPyJM0pi9psNxE1raJkbV/0jcWUqqWacbTiwJ0
LwEh0xO3n7DAXt05ao/FRVe7PGXrs1UrjRobCZAzR/+gW/zkDEt3bhIw6/piC9ta1Z8UupwrJADj
xG+zxo2POc4ufR0la+0gVmBu/30+2jxuqKVDsiSRUSNhANK7LU3xlOH4zcZCbYocngZQMuFrh5f/
NrcE8Zz1IVuDjbZEErnG3i2xGnwWXtBjv+aAIlEv3FJ14SEEHy5S4SwT+V1iaMdzoX+YwmaCDrCa
X7eBt4+qlmPIEsNy4Qgn2P0kCRKFOrcamiGYwq9l8kT1/EWpgnapUFJAZfULTZMBCtJtzDmpdId/
9WTBDyWYgbBVBuCjbiMii78RkOSVieh4RkGerRUXElfwGUQiLZxuU9UoaUv8Qi2ZyJVVKf55EeSB
+IRW1jCtZ1reLtVi0mYg1yH0/d6NxHypnD7aFbFb4txxY7aLuXb9X23r2FQp4pztNDvhuCD5utmD
SDqkU3PVcfItn278WFN6ZDET9YypfmS2EzkA7cXNZfXcLICSv+2v7OFN2HdTlUPmC2NOSfMmD2c7
14S1neTix1JNX/j9p8SBMWf2nM4CjhJfQ6VIscD1TFx7h7XVC1IbmvcbazQKxZvHJsfCfDm4qEWy
y9da7y5HvT57swIR3C4wn6bG/5PYMnkJ/gJX00oT42NrmmU86vzb8chE3ugAHRtNis1izcWjD8Xp
G4lhSynTPt2nD6YXgLrm2zQN+hdjuVARzIZDvwDgp3Fp9WsBsv4Czwn3O1suS3QGm98bnSIiunTN
mbuf5ynyYYiaksmSQzDbz1P94JwHIv+AGi7D0bccVw3tSPrIwiOA+h4V8ycZ051iZS0N6JYyLxu7
hplL77V3JzG7beddeQpaqQrPTsT0nfG28FjW398jEVsu9dnYngymiVHLEPE1Avj/nf7fVYDdhwdl
tgvGNsYbNqSGHIHRGoQC5mhR0G9Fd0KieXxTKNRtId+FqVtTHBBH0zrMolrlMHKl13mgu80OkO7G
zuPh4MsbjzZ+l0RlYLuRJkqS731rjs0dTzPdRwTsi1d+W0Cv9OO7DmTJFGm+vT+LAn1mvVMXxC+P
j9C4Vr32sgg2eek7Nww4Ojl3plGXDmQ1DpoOrJol5zReaSjU0BupmM7XBby4sPo8d56NNWMCKSzJ
OCLcKXU5z0MDYGOS0b414uIWmSfFtY+1P09uUtCLXDTCPDZ8mmVoDm/8bwMxp3eCz/7uWlG4shMP
Kqprtwm2XvpqYxS8kR2tsdyeAYUsHWEks+F/tLC/j2YLUltUnWlSrZLQnChIw5zNpUXRjrphahuG
H9U1Quoh+V8dproMFlCU5g+nL7KiAnLtOzChyaZCdSRToFZlhiURxc2YXm3/9RiMYClfGaEilGCw
8rf8PeikSrW7RqRIN6Si5B5FVYCj/LzxxrpEgTzl0T2OLvok/WWJGWuSkGjRPJtzQkARUHgrx1EY
we4znnpPFDlWmKUNPLi1IZEMIR+zYg3k0GhIDfHEbqZSAK8i5Au3kpAXY3eut6I9Dj+jM0otYv2Q
ybACPrLCJLXvp4FgLbDqI+YMIz4t1O7ScEkwTTwylw5dSSdknOc30e+4i9l4k01/ZL2rznL72M2q
9aPdu2Hu7r+VInW+59Ft6cPVEvY/NF/1w+sSRoZf23lGmba30makH0holB4V8BYojKvDGXxB+GVK
33HWs4Np4TONHS1mRNrBXr/qRnfjFp7ffx2hutFPDGOGeSOxMi6QwIArKQu4S7M6jGXPWu6imNMm
mJGMY+jv4j7e0/iIkYAGhFFJ+6g6LdaXRl5qf47GGh+5L6zzdoXbLGpf0NydI7eYZDcwjvJ8EBNb
/e4WhkfsAY4d1tlqpelfQlsF9Pxblk3Gh9ykHzA3woNIvI0Nd1Qk+XPDG7CTX4gcsuYfh0nHx2nA
rZNQjaJEYTnR6eF2AmudeidchOR40b2kjBUW6nOQfDklBBKN+VrM26ryp4FuQNhIjrhLvSkKPlep
R/1V9JjVm8dLd4Tb9e6vBPIbEmoUoDhG68yGBp59R0S9ESO4eA0mrXfdAiF7By7oNE9EtIJRrtnb
p7gVYXNO9f34f7VdfG2x+dZVX5ItGIXC7mSfGbfLVmvUOeYxl84ie9OJzXS9M8hu7R/VNpWYbb+z
O8Y+hbyXIwVACblVdYhFSvexXn1WbmKtbh6uXb6dpgQyMihNsvfxzFbplYY7OGK5tWpl+zV6xjxY
jVTazT+wZgWHqBq5UXRIAsc2M27HLDPZBWdkcFY9tmrZCt2KM3DBr3zRJuJxAzCDVTmEFhEBvEIX
JdUmaenOqDF3T4xRRp2AYwu3FIl03eR91c8+lbol6biYfakSxSmLNB/mAD/fk2hF5nTf2IwvAlsv
WcBzN5UEmcVgw9J7dq6zRryuPVsX8D32lD6kkHhBjr8XLS9UzdfgQJJ8XyQzkotbhu7bFx6FszsW
9aZwf2GWeDLJHZsXmHI4SVK1ASLtCIS0eiDmBBP1WyCMKsSDUz/Kbmsn7tZLxSt6/tUgCWSzViMt
dd58RI8mR2dl8SLufLtX22RtaBWhlSh6UyZE85RIAubtsgvTX/qWmfEEWErxRrGqurZEags/lNV6
EkaHW9fsif0noGgCzzpSKglnLTa0yED776N0WrnQZN1/u1LF4nDTGjAmAYRyxj4HVlFghYfAp9lb
d+CZyjyTRJm7p8qXa8eIY62gLh9bPyVqFBNZr1MaAo4whBZUtTLTytpv4Iv3bVQnO8iSBeZoDpqw
MVH8tBTozAKzx2AFRYYnnnFw836UqLFEWQi1sX2t85nOsi2GgN1gtwAAeMne3XhTtCPVpZ9u0GyB
rc+bH+GBx3EpoG4H1t18jc7ElnkncxOd019E81q/eAthpktTLjuj6WPMGEocL5/yVtTGWBzPSdI5
nQ2WgGJ7dJ1x19EbR/gH9B/tOh0uXw0QRfDMTNUST8NYiPui8+S/yDI47mDfFbstbZfQFCI4W+XI
FU9IbWDAFptzzIxK8WCdUS5LTIt48IwoeKSdAfiZv0p09gktggFpK9f6LsyKUH7/ypW+X7jhJ8DZ
IrcP1bHHsEja6PL16QTfZ2PcrR9hA3Hy2OAGLepLKWefNiVtnEFZfqxomY+vMQbkDj27//mL0Lqp
mAaTLQ4B1kastCGr+rb9V8VDKnSXapsJWxKdo0fMVdDIMJjlhp4I1jxyTlFVspKQ6vhLGze1fV/k
NudxixMfYUGTOAC2bwl2Yw5RWdPTM4B5MvwiNT7JCApGrV7uOwh9mftr3OdwhTN04LoS1vJUAoNr
1RPIeS15TxEtqfypWMgVvqRzoIVOpvE2TToA7TyXV6y2oDDw33D5ONB6yuYzoFpDe7zOkQ0MPXpY
RRXd4ysvqN4q3YTjPRDsEXGrc5R4/Zq3ARGpDvSusQB30L9TBn94RXL61MXESwHbq0nSR8qEx08O
WFCVVVlxvUVS4o+4H8cgy3ZOukBSyKRmNCwHSRGrGaiR8On0VZxYdoT1Bkk8RPODSeRREP/wCDhe
75YxGpd7GUNr5PT9UidfjJL+cifGf875U9EDHOgjR/aroyteTmz3FdnNbl/ayIaywR2sc2tSE/bS
baO0wjozJjy4+FYmeUqcp0yK1yFQGR83UIQ33dBmTUlgMARoUd5ln6aAzaqFEolrPZhIOgrST3Xn
IIdGxHvuEI0ZA4cCxAE/8cC8VWV8WupWaeIjRs4RilLQNDSmfpNaHF+jOIcTPkWtpDOleXV5109N
tbdSvkkTBfxncLsNfqp6HLh+1gvnSSLnvkawgMoF7wu+IEd3vMvfwl2jYNL70VifVdPVhTvQwLU3
iwDD+baBB+gP6LbgfuYpcRifEUk2skaJ5h3sHd9EBZEmdN9uIeDEix5CmBqFgzdNiPyv/L6r/GrG
ZwViALq7lhj3TTT8P+lWY01rHOylGC8xIN3R8xtZ+IFx8U9+P6/afLVBRu2FvDaiSKldPklAztL7
cRL+FVsG28CPGuUV9kPFefzxMrAf4dn7+x7kTCvyuNkLv2X0QTcfhGcnEZ8ta27ckSwTg9Kkd0Ob
4Ks4iGVH83KxVFTWtV3zV8P2g5ws19cd0K5kv6ioHDh8tvOzfhIpKz65lMzubAiDsgraKFmfMiBN
v7G6xE865sOfPQOfu3Q1P0rnMphEcSRrO+Fj/UM9D9BoK0/AU1WmJ5kEvKAw3IykQdQGbpY6iOll
mTULDCZvH4u1YM02BI+S1udN8AHj6lTIw4tVcZvKN3bUx/hH1x8RI1GeXyAahqo9kFlNL+OT7439
eRv2ux7+QvT9Tynl2SilFmzYOj7slZqcXWBpS5c/bidHxdnZ00Kgm1lnZb7GlC1mQWt/IaG4O024
x3VXnikGvDK/Qp2cMYee7I3d3kymuDQQ4kt7a0wI7Ot/RWFuxlJVYKh0xXGjoZX7Tf5iPgNs+olA
XxddCept3nEeyZbqL4xRL24V4GAlal4zPRR/eP3y2xcvvtE3wmw6Rio2yhjTUpUGNSl9psTZMz4D
L2Fj1WErK7zmhGxE+VTPyDt8WH3wVNhDh2YZdqmprdjIt3xDTGQnM65SRSYDs4QClBxeEd5OoZa3
7GLNJ2bP4HPuVD8V+n7DV/PWucRGcR1xg32Ixn6PuXHVi0RaPsyi6uZ+zKGkcz1VdQdYMaak6l5z
w4TCMeoWYoKTiLGfOpFZk3D2CFLISt1p4vRF2R13SLvuyu5wzDwLAgTyGy1A+eXKYtaleVDK+LEx
UvthdGUj6fAJvvncweOa9mloRtVJLC18QKIuMtDA84waGxTz4WGaSxsexluW6LlwTCrWbJh46zzj
zDssUBLd8k/lhR5byKmOqTMTvL/y0+wrjbPJGEyImmp8kHlXu7rZwEvr3esTTKEZHmIRweL5Lngw
f7OJAIo2EW7G+SFEgzkmvgpb6BOq+n6cgopLp5jJL6PSMc055UbaH+Z8H1k0yjGEZ7h6PIVk2V0i
jNLTLMqyK1crY5KGDluah/duCUbhbbaYs86bXsCKY33sH8Lm31S55iU6f+8koq3hKg+Xu73RRq1a
OeXKxSUW0wb4MRlAB/nbGwtp43nkDJkhqqahqkrbAwhsCyyE32IZeXbsBwIAZrgph/+noC3WkAzk
MnWVB/Pp74VNYtD1492Fe7IxH09NxxVgHhH+hNW86CsWMpaFb4uPgrBv7henLnqQDCP2lecKpRRz
qfcwC7cuJhUeZ3/oWM2MvUOvs7Lfq8oEmi3ZMW6p+T22ZO3jxkLOJE09OIF+mAfLjbi65clEaW25
ya8wLthBwLlqliOCqYH6u4Q8q7shVoybaJsiMjBpp217WhowUo+vtdoeVB0SsDP7J6B51aZ81xyM
BPlbW69EACBGBwwu7M8QonAYUMTDxezcmNAN1GQalufWNZTNZIDVq/On/csCTjtv4cuafePpgLQh
cEYSV8UFZoDn8eqb5w2X50rkd5Unh/LHetalJJ69jSQCjqU7v42Vru04C7Emfio8LKSeq0fcMJzF
MNMEy0hfg5dAvg6HWH1ENeObyv4W934jghI68AFW2b5ZC337GvuqMsn9878k7NHJMy8HwL4ioItQ
MbUrvpEEu63LeA9I5pRBY2OrYyf0ENNP7Z6t8XcNTsbIpc7geavRbQ9nIHvZbjyZvhKVFFDZ0Mn6
WmxxbwO+w8FSObGn/h6stzPbZxTBpUjlq2Atb8SKXqnXZZ9wGGLnfBI5gmWrPU/RkvN8be3HFCxl
u5NLfJ4U7tFLSj/AiUJbDU0M8QUXLROA+fxQJJiYRwBrgyoAGXvsimsIVYG4x9uom+FDvHJvhKYe
RgotL1S2kXiS6rbgZSIPeWMllG48Dfl6qCSJ4LSLavOyaR5ChxVqTl70UIYDVX/lvglU078pnvNq
gHHTjQDOxb3n5pBq2k5ON6OSJw6vWU9qKQsaJ6fnIGRD27+3DnSxiVBhANdw23ubT3s8HglvWS7T
HUgBcky6zirICbhgS9Y9soGU9OzDDMeMJm86bgK88xhdk0DmP+rkFXP1x4WknLU3vnfa9D5aeUKR
NPOyXsvqcGGeHohzAOyAoCZvmnbhIzTCPiCssdy22uG6qdxjXuFa+Y3pjglTFnGHxcohScyHPfIK
ieERySk17KcG+ng3oZbecOaSg+yefPvUI/551EA/rXch+YYAMwkoR/5zwAbvp2+RMC0oQs503cre
aBzZHaoX/2ZxCLk4+/jPqvIj8zBgWvZWa5mi89UTBl2o+/09YoADeMyCmJYz2nFYnfYS3yjh1n2B
fgJsaaQBqY69q53aUgsvwKdEGb/3URTC8LMsC9us5O8gFpPc/9lK51PYgjve0yzgDu5e10zlclNq
GlnehJsECH8FU5r291XgNVhZDr1fpNbhH02bu9aWLrcXPNcfmedEAZL0AuUYUi2XU5POsUjR3gja
oSHbXE72xwWVbaPvUXCmHsY5Knd92ItkqoP3ngObJ3+C3dV78f3vZovgJdAYmHf16nQvuZDPNQYI
IgUKmrdKj64i0NJUdfnqnAj+RQvz5xafjc2tL3wlQAafKIrRlqtF21dqGg5RgqY4DPre7PsFyHkB
s0PCw73XC8xTrW0ASoEpfz+ZfOKeadoZ5XTphbA06QN64xcJ+jCmjGw5O/4aXZLoMrbFSVPn8uD+
LGpmE1yt8xnL3vUx/eDwwMOGk6V4VyZDMbD35qnBp8Q+n7/yRL6ZdTGtWbbA8D/lAdTgbEwS1/nY
BK0c2KZoIbvcT+c1Ll94lN2531KwGsVI9DCSnm96xzFWAWxSv6Wfnr6iZABkzhFjGs2EuC4ZMjLd
2Y0ZM9WajIMS+lhsxufGb0tFpUIggJZKeTLKmjbf+iPK1Yziytx2R4mmYwOlUXgfarCP5nOP5iYT
VOFhpdSWQ7dayvYU6IH6D0VEmOPHp/KExHeHWqOd7MDMfz5nRpJClNZDGNLG5FZw9TkCwn2dlVYd
kMIL4P2L5i7fZHy/hKdt0/Gq2khjY9mbBk1MWvlTpeHDlcaetJ9jUyJKjpfaOs69skHTKvTBrTNk
+XSek2Z5iSimzwqFSd9Rc430fN5RwznVOWKMUcVxFfT+2XOHLnXPlXTwdnH9ZkeXNEad6sOO9xmX
P6WsX2I9Ko9BrrwhjnnyHsM7vPRZ7HWB/Z5kEb/WZlR2cvFqxeDi5Uwo7ClOL777EHW1dPwk9UOV
RvjY29F1FM25VI6RnU4jTMRvqVK619EM4UpEQuMNRFTNwckP3AuVoZ2ytCUGjKyULIpTnmf9ZCqv
y/BAV3eumVb5dkrDdEdePagyoYWlYx5qSTIxFMzR+Wv7EjjdzRKr/LzhEI3XLqMWA2WmJcIbL3F6
kHz7yk2ol5VPr8tQuuvpfPK3Pu4qWTXLFdwY4JvQ9EI+AS33zOfJoL6OvS0f5EpQoKJpvhMVTJUG
XBT/m7bTP+CS5Z6mI3TrQLP7TypRlPR4cqU95k0YIoZwxPHNQz5G1rS+cKMzkJGJuLWx8Bgf8nyo
Fm2bH3+fmeC2WhkjpbDSJ/WklCqcssrn3KS4wt2S0aPhs+UwoN/wNvsAzdOCWq2ANsEPflyd+xmd
/a6R9Vhg4tBDfusoV63EIFynt/skJ39bjTeMAxEIRQtiIAjPPFoUfOY01NST6pUwstmr96zfcQTr
r5ObID3nklzY3KijmCgjCQ4udRRKD5KDkpHMuFgqWtAW0SjMzsb5YUG2BRyoOtEyQpZQonkcBZ7k
SuBUKQSBU8ZxRKo2xgKGguQOTYef/DAl3knqqHZ/1pViihWLhzYX5CxCM/QqYTvLt6Im4kLIvNTN
d5l3N9QbgmByJ+I/1vp223GOz0AH2bFoPwLMC/yhslr2LOblG7LGP9ibLR7PQB79X0NYYgPP+Hzk
9xvnujeXQjKmhIps2PmGLVC1YBymsuxE0MsGEwwvOECwK2vGZ6yuKwmdgbCYyZAL1b1PhTapeD3+
YTNdGHraneVcMkKHME3mH8lYajS9i/tlSZALE593C8fpuUU7bIVdK8iOhIFsFLbdK7dCeW5BKfQy
KUwD6i5+TfgNZb6D3gsjaIhdwYMAPEVxkDhykaBhWmgTpv+rR0nt00ftLipFCa5cH3tH4JiQbgEs
U+sM0ztQ//66JgowYGZCFGWOcwDnqMo1b3ErWMuxW1U76GSEfeP9JC91cz4Xr7m6XJqXYxS/7Yx1
7h1FvNwPMxNtE3M/1UoHEU7AHTuI9d+nRldtBDNIZVbzYPHMqs5wyhqDwpGF/WZRFJrFmYTwiRiN
FUmquEqQUf112Ape8qLG9T6tCokyXyk0u/oR/ACCjE9R9vSTD25+84TqOUbUoCKnS12duVutvO/n
cUe378Er0QFyBR5K6UXOX2Igj14ymSNbweD0tGYMEOoDlj0CLSBbFWuBDKzK5lw7c4oJIn06P8w9
dStIb6CyjZky3VurxXSvhLeFBJ/Da+1AyuppjaSPiKwLfXLd8PSVLdN7qNcfMs56ytfrwoLjfclG
v59xrLEgZYPWJhf0EYk2P4ZBdiCIGTkMsAAQOM6cR7TS0y0dZ09xWBUk9eDun2jIFnQXlbz0nYmA
E+3kUbZt/7g78W10/CHa9+gUmNrwspmLNomCUz4fN55FaF04mcJDY91GjUKCB8S3DGwMB1eTtCfD
BSokrFIVHj72TkbkuuTOfkMBJOLP4iM7JiTOlWP/faY84U1ynTa2gv3n1qVMZgj8S8kalVFsMe+/
XrFMtsRI+sl6w3mQiSu8ufh0Mxk5Z2jtIYBzdIzlHhdShakDlOnlJQ680preOIq89D29uG1QKmJQ
5aWEl1GVkX9q5BvqO18qU+WUxSsBB/IyDaBso/3yPzWBBkB5+cHI+Pwp0pvkDk4W36lCohTy2rav
2K7Am1FUXdJ1eTl2JGLygBPRet1GoQ6FVtLx/wfP23DFIMZ/AvkJ1+9DnmcEicXLAtIEVBgkXCDh
cfgEIwMv/WmsxcOcitbzfkRV5spAGuE9ktuxtRxB2fVtKNrfoWeDQQyRrfIuHqr1iR4d+tdYR1pI
szZAhNSbVcrw4U9wnP4+UyAzp6JVDdzU2sdyzhx8cMBiRgtzPm6ZhpMYjiDAvWeo/0INTHYkCiMl
A5z6IwuRqog3Z3ymgFxRK+dQo2LvgiYjhD0k4MSNrhl3jXMYNrs0WBYA40FC7731+daR8NKgpb5N
oHIIgETnjk2dczyZuejfrU7MVU4W6lbY4JPvqFfiZox5PWSNPMtmtWKML9fYdc8PHuW+SKeZZ11e
w5DXkHfMIKyZgf9DusoXDKkatJPlblyBkh45zqpSOs4Wynnm7KjkGEI7jnU2vyKTfPcQO8f+WKsa
K8ljVIIG/TcOJc9f6BtuI8sK1Nhz/tjEbV4MFzHAEATMxRSCza8cGCGHHrkG4HzYCw6hh5rmrgbj
skfaUHKULO6vDx28WDe6Ureepa5O2yKe9KRcO1hUJ5qxk/xNQ+rjpSlUOBXyCfqwJ9ZAIVu8foms
I1LelxF5YHzAtS1UQqIVx3SpuhcWZ9nVhqXHcoM2oHPcNNRxacseIDtFgbIPxoSOf44ddBWbssCJ
MaD+uVVg0Op059p3engXWn9ZO0XaepbjcFxpCg1dl5KxNIhvEGeSRBGIwRVP0h540B2RX40HFvzo
10PrP+idk5lU7NRBxChkYQ5TgfcCo7Ggws9SvpOT2Pvk9Ej/BcJKBVCui/c17w22wb8F1+lS4RCK
jIjK2rsAEABOawEzD99HCr+qolGg5hmNYHXOij5CGfdYV9gjSln4Fq2AQMcQPlBuITqPG4T1u38Z
ZmMjyudSkB5z69FqLxlg1APsBsUvJ0eOHmgftPbXAWDUEMjGQsDByWfKYycQ2mP9egCkzAa38SpC
FPVWzXCE7syUsNCdw2jO/8cJ8c/jqPecujlBC6d/AaZG6o0lLDze0VogCn2bkJA0/pPvKyrKCsp3
aWe6+oGMqYf55iI7KEapKuOrCMVQ2hs9mUD0BPhsthKl359Tg+7g+NCMYAFZugT+zdgVemI/1BAh
CwSrNb2a+SN4YZS1Wa3c4T+1haGPwUmBBqODmqUEW7Hg70WkaPPX+fKsonS/RLsH+nCHrqvqikJn
X2fXK71kIMwLbFnxToOMz0NxiC2IvH2b+qv0NzE4gXTLiWRVu7Y1Bul0B1u/TisdERwH0Dq7QqVN
CWXuxIz71PhAKtd3LR2D+LvQkJBwM5nJp9lfrQ1sz3QCeJ8VF5+/a4Wf2vi9HR1vtBhBsJuCJXCw
Z89jZumO+Bv/DwgJ6g9G9CaBd3ekU3rIMuUt8o/MOLXr5oAYGFf8evkI4p1wU2TmxihQ/TduBNWe
ldHbZ0vXafjNwVrrVnlDTbJPZMykL12snUg/y5jY18jBpH9sEnARX99pydqkIWrVuL5fufJKHpqq
zN1OVTa/4FmPEJr3kFcZkq3bY1duwdlHSvTZ9zEcH12WgfAM6nfFqLa5AP+pQiR3IvMcG+qv7/wF
2p3HUcHjbqSIjaKNUGlIBTZhW7EKKRr3kNSi+Myu/cdSgFrgQ8HLn27UOVZH+pwPFJe7kUBT/2Yh
0E4db7qZHB4wa+45Xxw3Vv25iTyndLVoadqvJvtUCXDckAdkgfNb7scWbHaJE9Ji1sgkytrKHL6m
iBIjX1eOiRwKDcijzu9sX1G5V+4iBfkODAdS9Z6ayYrMAeggaKDwM1CW9XBT8fkRRoCHu9E7K4rx
XQ57jLOJX6t64j9NWcO+0fTVEmPYIHn64nIrxo36vSMl6+2OSSuad9d7KagYG1GFizlcBp5fn+ct
In7tJbWdyhAHiaK9+mziuoUjHnOLCkIimJqvgt/Dj4oazjVDEnfDZohB9VKzLQJF0kAWk3yI7qoR
5fH5mkVKtusMHba+EiraU0sTuaXJLI6j3K0M9kMtEEh2DKmboOLOaZyJo/d3mSYZrunb03atdpIS
Xe6DeRuH121NdrIctaOR4nts39+28V6pHxcWieGOo9Damum3R7q8TFlnzGFzEP2vsixGqxwP0qml
garULht+wpi0OuJ099JxZKflwIqGb0G7r1IDG8mpdLFOhF0cVsQPePYQZHM+OanpSv7YtPzuW1Kx
IO4+lsga1N/MYftrsRR0VSzArdMygV0/R/PhV0Z/DQCY8ddBvvAAe+6KK6+HdnIOESSp/1J+rYiR
pYRBmw4QXjyIUuP1lPja6VLqEoJgilwQPjL42H3auNC5+o7iIrgdQW+DUuX8gO14rRwpwuwu9Yh5
cibXwbgowzApLY5VxRxWjQUX8WnQk2tJPAra9oVXDYaCnWO6AsODZFCOojqLuchfK8aiwe+xutQX
TsWapt00JO7+jMvrMDhtDI4h9RcOc0ZhqTFgqztMC8cLqtDYjSUPOR0VbStBuwtMsm1vR0b4xEaI
s36YNcJGCSo+5SvENVCFHHkITWpE3zhpzxWrp1iWGgQ8YOzU1y/SpscSIddx+nYyfie7VC77EHbm
Rt4CFzIiVKbJ0h6OrCSKQ0CEyEuqcfWdBcYuF1+tu6VHNHHNXX9YpEu8GQnUU28HfD1kFFN5t3FK
Qo+nlu2cZLqMh16qHFtMFmoKy1F+VRTYDRFEksyf12Fcd47u0Cn/XXuJyk08dL5vurbiNA6sGWGs
C88AMttD5cktZXU4UlZQmVxBZPrnBg9tMEL8XQDEZW7fppP9xfMcvcdJ5DlxaqZhq3/A7S8zgCZf
JsPXepuax9hWKH2zHmSuo+7JQk1qeShFnJVIf4wINJecsaO7kESxHTZwk/a6CVnOV6Sh4fONWoty
m9VBPjJYNWMR4rymh2JjRL1+Fpp1J5SANX5ldbCLZSu2MDaZepqP1nBof+Uc0h72zNjrg0pRYgvL
oA05TFkujFZalbkOpb3Hn4jDZP1aqlchxSC1xd8tOwtqFCcuqtahoBS+40PA/3FXcg0GT7VBIjbe
c1WH05c3lteVu/PVG0dBmaQWEeHxtbvyGJpeTgzx6H/SqyPBR6rj0DdxwCYbZ3H6/fDLLRnsNl5h
BTmM+EPoKZHkf26NjM728RdPfz6V8nbENjUem+bfb526omQ4ThBnKMRtcEnVVPcvEVmNvPLhj49n
EiPsg0V1Hpidr4FGyyJlkal5Rs9Ksco2GPu6SS8Ab2LNY05+Y6fD4d6EraON6IkLRZwuRx7LWoQl
UtFFE6lurtUFP4wQ3coqfxXZk5+Q8E7MOTYAPVOZz3q9mc9AlJ0h0NW9JrCb23Bnil5Nmp8JQNCP
Z6famBwSO8OWvu45OFx5Pp3bPpFF6HtF7giG0GatnwBN1Jz619fQbj+FpNnRtWbYavA4DzRUvzkm
HuFvsxSgazVVKNmgubKCVhnidD5XI6t7IpkvY0/1Z/4v7BcpoV5WLLHWdZOvdr5TUcENSSca/24F
oqa3VnaCE+ielErWXlVRi1MCK2myLe1LW6psLcKgJtkdUMgSDiDhzcAPo4QU17sRg4e7lmY2Um6S
CYTgE90ZvyGp2XjiZATeLyyDXNYpfzHQUUrIz8LCCn3pzydHrYirw4VJIgvi5DPodDPHJDFCZqsA
RbCuF62TXJ8ygYtryYZTLM/7ynZIboCh3f++6R0rlmHqQabcjczFF3EGzBsXYojvTZqN3dNNtXJI
/IgiaBE5d7vaoB8AMv3COXZcSgcVt0W6kLLGSPv9hTnSTz+yzKOIt2GHMK4pk6tBL4FJTaheej6m
CykuzeNkFyDNfDiN0bhzvP1QvmzRgiXTh2IrVfj9LVuJhLU5XjdiQvc7fgtE3vlRuRbf9aizd5SM
L+0X20gNgVysjkaLBPJZCt2YtDobhSfxrzdNFPazCJb5roPH7feKA4/kBdXbS++byfVE86rd0hP9
IcIaySRX29RzH65WuOFI+Q2hvA2e7IR8CQkyfdf5nExvH0x7qF+mVV5JdIOEr2Eg38u0MVuY6OTl
xU022NOF7S0A3Zbw/XO+CuwBRV3hFVu4yQkAB530mXOggeZ1n/jjUE0shKDBygf2/yC1sCfJb/DY
eGf9tH8ebcg1U2WjUQcViy3+onyczqfDyJ9OlFgNrCZCwOdbSI37jlIPAjTSllngEok+7ro7kkJZ
JpASvxYskKcZTHYKCuaGeB655jyY6xqrlytLi2sVk4mMq/2uzDdBofzmXf5dzG83utxw00GlJTOc
s/tSPibg8K5qzDuhStd0cFDPsOJBSamaFk7jK85rXYJw8ObpY4NBHoaqwS2pAjnFImZZGIDI/Sx0
gITFQWEhqun38+C3K3pZvapCtiTZ65kdfSXX+5TwbNFrWlkOC3Goiqo5zE6fJZyp/zy/UPvMOmPQ
3z5gfPzU+HEY5fV0kRmypYxxZtqvFjmLpMlp/fQk7Q+hDX8voWQdd0hNAxo/innOrmexN/Tl1t4c
xjc9y4yqnQvfiL+xd27nqo8BOZFJLffbSOp+vM8UPQO9YZV/QSn+peQiTAJb6cjP3wzUuL9vRu8N
LvhbLMY3g+zbKZiEmL7bdQac6xfx3J7ZeW2hlUlIs40H1ADx/6VufNOXrXueIq/m7/lSWe8fAt3Q
vGSivDqqdIiZSlSIFPshqgOjYB/KcvMFPISALzci6WHWMsQMZytvxsG/F+H6SOvS7NOf1sEewifA
pVm1BKLkpxaLjQyB8k7HazXIa1/FUL9WYWNeTV5msMMAznLsrW6nBJN/FfLtmaahyOpk9eeYkb8x
MfiUIyZ+egPtsoB1lzZa4LVk65niQTAh98003xo1u2PRMJFIIdVZuztGvfbNHt0kvLS9DXG2dM/q
P4vFwyHK5K0gIj4gOBN+VH/rb7p6xPzHM605hUXNjSNfVrNelwi/LGlrOkWxczKhGDZSq1uUmG33
NyQd+tu8VA0nk9aQT1BuSdXpGidDfaIO0WLtzHiACySK8VIigRFdEZxJbuxpY0BQPt4nVBZai0ba
AsKZ8Ik7Ym/etSCykIVRT58hM/KQQ2goZDfF5zD6HPaa3wA3efYy0FH/1xEZL4JtwBjm1RnvyF1O
z2yia6du+D46ft61soZz60fLNEqaHxgoZlQzvF18lXbnm1KfyJh8ke+Ia23VMBz6Qi33NHFn8nA7
8LylTMyb9Oy1cgBqQplv4WKQmIowl2wSFR62Lj9gVV134eA8OKRZQc9QrQf5gJFXvyeHW1lniCaH
Ge6Ml1KV8xTcozZtifNlsaUWpAlAiUfE1+P1YCajxWQ/016beAAm1uTdIp5SyTgzAEJ08D4Ld9Wv
5xd8KXDwVTSPp2IgkBSreMpKRFc64eRYnOELz4sogxlg/a8FRTS/7CYZptc/eWWM68rZH+QUra6s
+ocOEAnPBbzBh1RjiNqqLgFMqE89xFxegKZm/p3A35NWxBmu3EIYjp8IuzwacpGAkLjnVLPjm5uL
BY/Ta37UYI3uIQhv4TVPRPawaoss5n8aDZKntSwS+lfJI0jhISCbOpvZrZ9zrRF7ee4ISB2o6Y08
13DuxUoKOceFb2Rni4RXYt6k+wpDApGtizRid6Jc9n4Nyngq8+8Iu+WTtAcRjHoCwtV5chZ2eweg
upUohCW1X8lr82+RXZQheSZflBE3sfzGijm8kIHizRrlHM5sN7cWFSyWwhIyRGP0ObB6JqTBK5Ds
1tTuzqQu3FmGPa2LoJrxIGgoJuUL+wWeOc5U1um1teQ9if4GiwZpJw5oXRVlCD+CeC1iAnHm4yb4
hBhHyf7MPRBMzz8QsMRHlu8obBVxB4m+c3EbxNGHhgW5i+LsddzqJMy3UovLhSisyFhOL1wgOs+n
S9eqO71OrkCjR5f73i9/CXf7qYNIYEV/06/dMoepIu97S7ukjZ2F5qWiafIP/KOK8cVZ5uax1zkq
jdFkh22wWN460xPQfYp7pbZShwqBvC03LdCJiqnQLotxJutGJQJi5//EqQW0GSg6VyRAOPYnKr1q
XJ2BmKnJfmDhl9u5KMPxLz7ppqMEopgUmeteAOh80koLI0voUcLdboTxB4oePHld6a/kSXgZEIDD
24dtycQgbqgoLzYrLJ7ywN4vzTD2BGJtBq6sD2/o1FQF60HEEXX/gEJitKYMtbXeony+EkeiJIEr
xFlS4umjozYY6VA4JDLVNIzMvpQYGH3hCHaswXWciB6uiE3V10o5XVkxDT73tuODbyNh1TzQ+d/R
lCgImZsxwMRAWFJLW193D5494dofpmCt2+PQxVo92fOysTGWO5TOA+hedVxVbQ3VsyWqtjRn9xV+
56xGMYkyuNPvfpkYafa1nHLDWp7tSMGazuRkoNfAh0kSn3TfNfON6rBiWDYy/WMffHQRcaThaxe5
iqfe+offlTM29F8YdYVp8Jbs39lrm/qQr6+hzz/n9wX34lntZK41TM3C9Wk+e7Turhoaj0eTn++V
rxBt7OIYcvnhl4OUkAyhXuLFDi3qYq0JREEDLWg6oEkebfjD10V8RCSOml1wdgVk1cinlo7FdiuY
jTEcBrHyE4KTPUetqMx3sdsYC7/ImurplEHT1+86ZOMGwbh05gPTv+bv6diI9o/ZwlToJ7tk9DbT
Lx2syeE22e/sS1AIuD9U9CTZERUMDVnYshBCSq56PuVuwGtyv565TE34ogaI8zb7EYLU2IOn/K7L
Mki5BhbhrLu67HwEF9OXDZnRtQZCkUAa0/WwLnGJQd6heZ6+Mg/Y+1lOeB5KzL7HFxorrYQXjVOY
9BJyRvIo+N6hoabiV5j3Ukw8Sd3atpKg6btwGQiqPeZBf2jrsS52L+M9wBPfU6dpNHd+PbUbUgWC
wr559cUmu5Bj1maGx2PuC3hZEqsq0U4YjxTMKOUNPFIbOUJ9k0IrhqdtKjHIahWw+aSywZI//Uu6
F0oAiyPsdlm5gHDzH+cz5u2qJODkkCsNvZ+YNisy2vbGU+cp//8Jx0dytcUk7WsJwHZWykjBLQw2
9gaSUEKdEBQmz7Jez75Z2pAOiuRj/H8pgjNPvqHUHCayxPL8D4d5k0qZXQMluQ7gQsd6S+qzOvdm
JH76x0dnvyfcIXeCd+i+izYAlepruu3Ash+vVT8+ULwh8BXz3fINVaEuxE5qMVIgeROwset3JCIZ
xzGIY7HmEGr6JhRIFdxL0QK+2Omov11+xTFm1CaAblHvL+mSl/5h/YFnlwlXgxRuG9qXujVOtUD7
s1Uk9+kS2m1+UaFKplgu/s+o8oOq/wspjKYIo5M7tMgVEuiDJq7+ZRluFlyfrxy7A2Cj+ZTWUldM
hyCw9H1OairWmF1Om3H3xZRCQvhCkunJkFfDbe0fId9U+PwmcRX6k/JUh8/C3AI3N7Itnrfv8oyv
y3fy2a0k9mTeOq/ESsw7PK3j7pB1ckF26bmGJ8oBCMfy/HcEmu2a2BHuvuBMfrJfdDeV3v6tN/ig
iF8S/X88APVGsoiJETspVaTEoRK+1D6mGZ5a1SH8WSC7ZPLwX+WTYGqKoHBQ2fxZc4Zm+T4ugtSt
sQMxGMXoihvr7exjF+UXs8qXpfmieW4/Lc8yOql5mlXb3eA4U4Gd5uijd1bO4d+TNK5VZ1Q2aYLw
vDBwWTSyI94ldzTqVLds+mMbd4IIJ98khfuNIKeGm+PVfzRtkqoi1njmRhmONmwSyJrodjPz5OGM
LH1MrKLcToP3Av6TQKBxaFwJQ6ZRfmADYjvQeXIZ+R+EAJ44yp4fAZ0QLE8riTQVzd/Ogzs3ZA7Y
ekkxr21oPQ3lrgak9h60S6zF82aKRJIcxL5kRzt5x7U1x0DL/uYy4GCVuLuA+aJEqyQk4jEGlB0y
JIsHXF7r0ogPylRf7P1OFmkdaOA+ZgUNxZqM5utBX6/nb2dU1+gIPrx1UUDh8zIfNZp5StpROWAd
4CCVu5nTs4xaDUCAZ8EACOXV6U0Opwas5NgLjuLXxV/IdQ/QOGntCA0vLupxvs2aggb1FN+2y0yV
LiJfy88/EMi/cPeXueWU7b8nDVjYMfVSEW9RLFkVIyA9AgrxnHxDqXIf7iSGswz9qLN2cWDdWw/d
xrdtwR1DDTxFgRHHond7AbY/3iXBhmK8eGcjufjVr4FLlUPY0Mjvw0AcLhmceBwyXyFyUMoQOP2G
k/PcdXpdF0l67yBgz4SZt/rKoRGwhPFPvY/C3v+yhM6aVdaiha3BdXR6P6CP6NjBeQ5p6YR2MCgy
aMERZiRLsnKAArm4ytj2zgkuOwLgv+vfI0ZsyM+xbqlAo7AqWvh0Cl5NjjrXGMuQ19G6iRiZFzd4
/l9HObHDz/3mWtD9Lw9QDhdig7xtwTvmIfEV0b7ofcDS7cTd4RxDgZ+SgYLXFHufoRHHmboyHC/u
ScQWH9XLxgCjMfV8zk7yayGcg7h5OoeiPVKBRgQHeLZd9vEua+fHwvDHndkhDA8o1IlF35zqh9PO
WqEpbkMsJ1LGtsE72u3RQSo5RpvAKF5HKEV/29R3HhiV5XE2HigcD2raf1z8G1wuops/QKVNmuRh
LANsyBks9QVCJnI17eSCY7Hpn4vq62mEtfviCCDe20+UFWknOZjRxgcSQdn/0gj+MNlz8cGgpSfF
VyAb7QVw4wSXRz01k+hX8lZ9eRVb5Rkk+o9UOxblLqGoCMBkD8/+tnn4O11fmv4CTQxBq3ErOKj0
mRtXIJcS3WFr0Oblzuw6ekaippU/Ccbm6EN9cWb53U63SFemyq4mJGwpDyoLGNlgtv7uOXfJ0G+l
aSQ+h/IVmFhPW1TFjepGvJDdq0fQxAkGOtsjAukAgluGbVBH9sg1H/IJ1rvIO1ydtllH0Z1zl0by
vtN4j8Z+cxu8DkFe1Ttix9w7KnasYDIIlFLKx/6r/cDnL4w9KwyXQZm+wfqF7NNoAdUDDC7cEVv5
UH7lHSm5WQL5Yg5blq3Iu1v4NCKzqGJoOnRN0T3yi+5WXoIHqtGq0nr+3LtMKpxxJDO3FSFATR0Z
KSF/uNnOl8q4TF3jOQy1jcfzNQDrbpZB4GfRHm6lT31/4fN/tBzWfK8Hc0pFajqz+l9ohzxNgfAL
bJf8C+fz4FTeKBfHSdzGwWuwZfriuRUsLfQ62pewwvcciQkbZillRILr7NjdPPe6PdssZiFqg5if
56wxvBLEtu+xswW9gPYuSX+wHAXYy0PPBZVFGwCEJ7ZEUfMsxZGZi5POFb3bjKATmm27x+V1+/2E
MellylpS6M8WXQyNgDzmLT5izfcMixX5PxI7bZ4Pdv4OL07eZM/sf4gP7ZVlA0Q4NQ0JsxeUP/oB
s3Mg7xNvBVPALIt/N5HdQfXIjBte678YXdNwnkve48IgfbLBfsTMq2rGpmWO7ABfAmmaFKd+ttdR
jbkkTcgbUk/8rYl60LY6rJkowrLTH4VbRffQS96MwB8GGEDIpAMQAuvwhkzZSrkaHY0SHhIRNuYb
Kd/GJbEbR240hM5+wY9GnMNci2ekn6TX5f89Vlz/DFiDp0D4dmAZTcv/Bq7acS1AYzrdyMPABBHV
2S4N+AgQqn0BXY4G6HVwnvS3hVjqdaQNFxN/5EvKwEh1QAB4WHzB1L6c3/aHIZYSzolV2xFaZIMy
dDckz/v2nglYp/cwXgBs3kn/V3gdjAilyDwUXkWIev7tDLhcbsCYjETMndm3rH9Tger2q1zYdeZf
tzShwdYjL5PveUPJRuPvwiJD/JP/5YDpRL1QRKxQTxG4ObdhJU68kP+7Z9bpws+zy0yXPLg2WjrO
dJ8c0XOEmgGK5HiLdTLDketp2YGW7sl0UYMKlcTrVawoidm9Md+XWr+8Eozirkos3MsDzIaCWicn
fVdU/GJt/CWuWDAaBY+kHQie5ClmNV3Ztf3hT/JwrHZ1bawgnjmCG3mebAdJdL9hjYAZdQbqqqGu
aURPWOiNy5vGv3I44x0r0WRYkzIUYxbmVeQ9oZgcCGm914b98hS49J335/JFli2OA+9px2avf8SF
oVpYlQ3E3b64F//tfB4Y65g4A1Qg2xjLds5MND2bQggWTc8McKeiiTeywLAxt7ctEECvE5tVxR/b
q83BAmUrqNOhKi/WCtDi9rFMJp4INwlytgPWUu8xucpy1TS5NXirgKt+ZrhJNQHnzU73+avEcaHF
mB0xzggkgu5/Kkw2esOMJATsbndDyuUmz2JHQnYrLnzYaz7q4n1WjEPqA2VWK78KlBRKsYN7WoTV
5ENGdOBmwQBzdhqfaN9JtmwFiwnRDyJREjsyyzLztczigSB7h2W7UKiWPOHr0O5OM3T4/b87FqTL
+j6PJnkqbhcOeJ/eFDSJv/QzwUu9bD83QbhQCgHmobAiU1FZVr1GxzSV6yRjBfA5KvtEUy7/PhOb
utza8CtWhb8fkESMIrT22xkNkqTtFwUSz2dieP0q+d2LxUagA4jsYkpSgCtl5+De3vOqPunR2EbW
e4yxEsJoHd7Lam7x47dyqr43NWwWE3YIJ8IAOEu0DkynSPFU9DLNWIqz5HTbhVWppdz+qSc52MUX
aVQvLJzJOy8+44jfGIbrM5yhaXa+9r+d3SEfzKv/04GHX1QnN1ZZVQS+TmOOI82vtPe2dZgPwK4k
TaIpFxetG+sbVRcPfviLFUGPeuwGtzC9/Y8a9eU4zWm738PtyFYVfj4SJm74WH+tZkPRh9Xs5z2s
vZmXkAgh37HS9kxA+GyHJoci7LigetLlxMFy59ZvrOqsT64d1LJTL3uWqD46CpG7OeLQWE1HW+AQ
dsrKTy4e5k12tkGV7mZmBXA8+gIJzkanjlLmGk9bTXaFYR7f7diBo/4cFqokVbd/ljDkUTnEck7G
rIdOagq+c1OQVKo7Nt8jSWBMGetRWNdYUtP7gVkgOMUO4hGl9LCokvzK5521ObEItrMM+HosFwI+
ej4J7+BiZxPneojDQZmtjCt5CXxl44qv9STm8TDvA8kf9CyM7e5c1EP8bHRlvHDqBuxVURxNvmjm
ihkOgyzbLb0mRcgFE8sdIipDy8Yes9j0KNAM/QOg/9du9ah5sZgxq7c/w3CjE07XTxbmPYMpyCDS
CrAFfS8X8BhPEw01b+boB0iaJqQk7+CoE7rmxsYMGgUaWEi1O2SFUDSBRSBlPSbKphHcJ0gdqOsB
tK3zqXX48LwCbGk1QKUzgaefE5oArnKr3c+cu6ZdAEWN/hAmNvy5t9AnE9ILOY7AD7xa9SphQPfN
2m9s8HsX3N3g+i5blrHOu1UNecjeflj/h0MUTa4LdgFNaQ/1BlSJ7t62rL8IpZRIfN5SYGSwLAEf
UNfaszOutw8n3yUy1ZhKKo9L6Sw+YRSXAv1WNSlFVA7dbbuRjI94OhOxJg4jkp8KHVEFOGwqjSLW
qItUihCZE3bw/YCpfowVgcn02IO8hRxR+QHXrNqrWPGlrwyxXsntnlf2UmzRlzbdI93AvV9WBbwX
Hl60zBNPTaawpyI1FA2PJmcBvuoxaqE6HTypZo1rgJZv+rzykvTJRNswDOEB4+84/r7DLbAZ2j8r
FPg66VOO0JfoJycnpM8ez6szFBFcJsa3htFJajhtnVqPQtSyJTovD0yEfHLBzBUyaMuMQP6JM+ZK
yxk0Xpmi/JCvFJzvcuc92OnN5e8hbXxtURFIzYU9e7RRB4QxK0X97t3qopxWA2IShXIBfMXC9lPJ
iWFeG2weUbyGWA6efyeEJXSebzc6Fr/MJ/PQtAN5eBEQnBoxE6JJe74B2nFqdzHzFfOPZXWsmnp1
7RqNmEY6+pPYdzdOJiPwO7eyC7vPa0wkyxELdzulnJ8T13PF7fBBBOHdjZzTOrPa5VoZNA+f7B38
di3I2MPeSaUjArhyyiWbX1i2LRLeQOxOd41h0W3TrCerZWJtJjD/trQ6Ekk51wCDSEBgolFPUHNL
16YrGe+iTgRVW+qepn3PXxkW163pBLtzWOVy2R/Z6kgg69jGbQJZ4pRaow4FpJ2bbMyuenVzhDIq
rllzbRNr15lZD2ncQ3lFqXHog3Q9vrC8pKBo71zWe4iQN43cHpcp0bUUkzmWelaXe16q9jUTaCeT
KwilOmwLzxwRlryBxAorogaTnijCthPraLmTFWiuMtZsiMG4UHgj2vOb6VNB95ZR7GY7++H2mUyX
EdGKskG9PY2Dz9BXOMavN7sMp50cxZI1snP8klebc2DwDmeIv58Zngoii0cF+EN4i0HLc1JDIVfd
6t8HG0NUhf0lfGCgwnjCtZThr5XBhGTdJEPLcMJJ2m68IROj3+Fu+Ajev7Y0G/nDND3t6/7XGBVm
v+V3BInUF6OAfk4NNm/rmuo2G4CRYdBAmVYw1F9WlwuV8np00eQ/riNPd+Y/3YeJ3i9HI/aQvgM9
vpUy/wLwNImtfgRdMtTvVF/rMJSP05Ix39MXo9psFGzPE//vp/SDyjsxX639Fs0K3LOuIX+PHSjT
U3MLgrmWtevxHlespa94znOYnNAOuoo84cOqsTOC6bjABjKXjbWjzYjv1z/L2l07KuGHFJjXDu/I
Djskjwk3DgGrGepUDaU251HbAEjtR3LCnw6SdkQnlF3TxBiA/8n7FA/Sk718WfqB2MYBjALTqyxy
x4y5L+MbRahMSTibSVXdIckAgpHz13cVMyJclMzAhICfR+9GiyOJogmVCuR9l8HP4rVfSppSt6hG
D6B5Up4kUfvUzlJIcjatg/+uF36apQrg/pzcdpxLxaAn592N1pbKrRsZLBkp8nc826UhQBT0EY4M
WwXSu+FL1KHQTxtI/CcMGvnqurE1e0TkoK2N1Vu7aRACHMQjxSDK8UWUoG/f3WaibvILb9w/Bu+b
R3SS7xs3hcY4kLmo9QoXiBoIIzH6bZeCpFDLptQghG5cB8KT9GO+gVq8sblm1Ys6m9JzGUy9/gIG
0Q2Ce2T0rpvuGCWxTiWLccuGQ/77jSyZrYadqUYgOD79mFcD95RKd5ANchPkiIDmf4PyeeeyJkuk
8L1Mp/uZxJ6ViByvbvAd3XpWFvoHWzK5ll5EpcfKQHWZ4B16Ydkz8ogoEdtJ0aCuZuItrEPJ6uwj
YjGeaufgWoj90pbW89dRpDZXrvxJfn0e77VTKfwTlYXcovAwV8FS5pnfGdZE+L6ujC+0B0g12t50
fNlWAiup1QS9rTmmNDcHIjsp34cs8uGucnCwTFHBZnM43QEDvfds82G2Rg08RiIvdX1FwSHtHTf6
T3e50m7VmFptqHF6E139RQEaLSnAGD6+5pAcMS6TWKyvduoMKblWdLVDXQBhhXNEdDULReI8+j9E
GAkvMC+gtZGMf1z41QeUhLBIM24YnAH4M5bzZafF1AupIwVkGxr+umKwDzZwk8dPAmCFFnJePuGx
GApxRfOHKYv/Azeq56PSQD0e5bql9zJkLxbwqj3PihOjURc4WPQdKnOMFT7n89aUAWF5G09YwVop
vu4JMS4MYIA2YGUb/lvvZZ6VICIlAscl/hnIvRkyLfCHlnGn/kcf/kldoiMMFkedgo1yG5o8cecS
UXSVA24P3vTDBOlEGkBWOiWTg7aZoyCwHDz6hIDcw2HlSf032aeXQ1XkxQ9jYOYrmY6kO+ioqsZc
yphmkKXRhlQBeP9zckYwZCLEapFwL2UJ0me/ep+Mpb53TRv+vm/BXQasJbX275kRRVj8iIKletsL
rwh8ZH8zV/Ue/kSaa+XLwmI0jzsxX/F+bEAdhdZ2iOnEfEbmz1Gcx6nUuNSuC+13TQY6xEBGKL+Y
WUEgrhFrRaCqvNxEwjYy7NDZiIs0Y6zqEDXtpqUdInq5GL97c9hIrDxrF4VQYrIJ5PM9MGCCrIoL
VXJX6NFzIrc9mjQCzacg8bziqzWR1W3muotMogFhM98lquliaNnZa4V4jnijfKIZxt/zrRCdxXil
gMkl7puvL2QVkF6s0ji+R9WUuj+iaBisN2GhlInxCW1RdYzszHsgLEugV2+yLikHq6buEvl5adwl
fus6A1mfhvnFx9IoAF8wqUTVXQGbHAHg0rndmGGzhlOc1CBnBVVWqyGLR6ztH3M0+52eHwAtSmvi
XBgmraeBIKXvVPOSIbh7bxM0Io9k8GZ2ZroApDL0VVMB96/jm7cVAje5QGWfC8FYVlcJ/3Pz3DmX
EcbA5nNNC+7zYWRIVtjj6g0NpnD3fDKjkh5ydfTfxwvLWst/YnjDJkUoSU4PA88KMIRIztUBydgJ
jVDEhqx2H3GkzAVr8CLV5CxsaytDadPJxU9SpvmbbW6zwfN2TDyH7jjNagmEi4bNYmPb+mLYpd0e
G4e+evX+Atzt+szpKbICCQEbcJIaNyL4mtWJqFIdAOwe1Ujx/2cZ06+tZKVg/F10iTjaxAM422C0
eynK9NdCjRTnjDsPq1CUlwb1yrKBqegvaVNXf1RzF/joNdyPNUPub71hlJjCQJqZJbC7R1ndu7V3
YGKAa2AsFVlSJrtBJNpjWb2NOwuKeL322nRXeI2aMnXMNcOr7cV1eikjJyY9g89KX2BGK5iWr8Mt
7yiFR+j+PWuATDSVlyb2MVfdHOm+VDKr8dogN9xwo9TOvJ9Oy7LZ4GhwSyEs5i21gn/x4kIQQOLY
WsfzDYN6J+t89JOncQqysZkbjGG6bEtb3QqsQ0khh/mE9raqFlbzdzFcUuuLAO201xg1zaoLORnE
sm7PK9C1cjnWhvQTDDUN/MUmOKLCbouyjw97yVXzd9b2N9SwE0RrZ/PSnndwqIPTpEPnEk2BKm75
SPdCxWgbwikW0wgUZnHkJ46Y3zJmspIoDj+6vvoEn6+jowsEQyl5g4xQIz/FsXKVR+7XDKX2KoCG
O8OccYYmLcrf2c4I/kRq0RznY0RZnL2G0sPB6Z8AYtVDKIZCGBfQVn77gFHwnmIANrzfZUE86rNK
EhSUXKPeKuj12nSe5rM27N+2IJ67Gf1sEVotl0eusy2qqLhcJMbl+I5wKEw3gb6dh0GzLSkajqYw
sPgrrTWaz/vPXfNf0BEaPcJusrN4A4XF+KJ+kqd38p80m9gsWbMGrhtcg36Ctb5On6d23isoWWEC
ppSg5PpTUznVey4qpvpk6oC8zLuEp8hImqRqRRA5yhtNESOcgTOZNAaXlkv73uOOy94ilXp1snl0
AkA3bxK+ot0SJiXVSAL9zPNcGTU8XLM1V+XbqqvBFEKRGTslURzysGWVdn7OJpSwU+ek32lOQa8U
VTCblnXCvpr+szkeRWdd8quPDAzfwiklgJa4E56eFtKjFGAPy0/E7eRAf4ltIdwgpAkGha7xon+P
IelPtdpIHliLspTsAzNrMs5WhPtwluoRvCQJiaLNknwPsdGyzdkCR7hv83eZLdN4V+zDG2xEjwC9
uhvLkxFzJ3zvsB5XJSZioMdfkvCWzYHYkVQrtYhBIfdArdrnfS7wtTQbIVTVscTVSY/sPS1gYXa5
bt+kuD6lbso8cCmO86wAEyPV5YcygFW/NqbBiSbvd8Ne8aBlHRJGFBMtyD2xVJ56z9WEc0724tI2
YepwdnUQy4mngWpFHxAkKIqqvTz4auj3MTNhuKcUnQPOlj1Kvt6ZHGd8BMH6YTnTNlp+HyJlr5Jl
ggcuU+MeZ4tIjQcG3793oB1KSMkqcxKDsgGwi3nMmRUzY00TKMsd+hXGU7l6OBUm0pmtpw//2i49
RS2/6Jfys57i6JuTxzILxKYv4RObEd6riqBWt+JMTObxuUwU7mT+gaalpqrABsvVYGje8qNKHMyO
IxNQR+khCAjYz9hOOTrsiqEo6GgZAPDpwxxQu7SJxdZXvheHUsTbqS0tHBK5NC8+DdeD6jFi6SkA
IsiZhmfIdB3s86DOZpzmwmtQMwTUV1FJWJccdalBLxefLeSPn4TaINs3KLqCmVVDMnZI3N0jL7Wx
0QzkGi7n0Btedzj1Hr4qDfNuI6hlRaSzmVUhXto53sbLdUzNNZcZ1epBchnupKejA771M6HPBSns
8PiedTCxwmhYVd6h43aJg8BEfuPfYSOpociVFYePVFZalprdmZdg5nXIeQhC5GGO3sxkO7bzBCQu
qnE0tGDKdUea3gSMh0K6z6BCX2ueBHwLCXkTXSTI5H9dARXvbKn5x+/U9A9Usjya2FyTHzCp2R64
2ZE7+rDNCNWRfK8KrT6XrLGpaFV1dYu+3JzWzPK3akqjW0TJb78od/TQ3ZPucHoyxTTTayKi3eN7
adq8D2iQzPGbVhttpxFLRFhkMXfcYgyR1NvNesbCikvuF78eEon6qRnn2s7P9jww6l1PUM1e0PRj
yPUWU9mfTa//F2VRyz2uQ+5LCHpoGlc8rfnFzBQ8JukvlAJzoX8rPTz/PVJjwQREvR7xnDtouZu+
AqRXahXX/yGMM8JZ9WkW65QoHZ0GXbDHYh6hQY0iO1hH7bvv5Orn0gLLk5zICVRlH7ynwxe/ihPT
APJR+lu7a5eiEDnKG59slFUaah/dVk4Kf9MbiumvBnyP85v1SlcN5dj9kxmfD5/o5cUaWQxHGE4k
ZD+bEZjoXucZXjP3esFefYNyddGGtcrFjjNY5N7uT+z9WvAPExX+LDhFFKbm7RQlti1KHhhk1Ebr
rcQ2kUVeuD7ZQVzN/a3dAp5GpbZ+SQrkO4reV9RPClEt/267sE3YGgyZQxFArh+kJvlRDw+KSPUG
fOfi+oHMspgXEYpApWmV0d09flXTkpjCOqkfvTYNw31iy7HEVf3h5hw+TD+MqxGzGWURGQv+pRw0
Zf30O9q+6a495eVofX77O3m04n6VDjash3HbDaXbUJAXb3nC0Zywc1xjmWz86J2FHcOU4BVu/euV
TqlZpGQeZ5RYI0PzJNMZleOECyK4oL4JmMaMfgIOsliJ4eESk28mVkUifmHvuyzdzhKmRLYTN35f
OT77+bQeJDGv05+dkCUn0wMt0OWqfFQ/JTbUdAsKkp3o6ufJcu1xFLKkCrmP/qwYEUxwF5pFknrG
qAIO2qdbXYXQZxoxoo4n90fC8zfLoDaUr2R0EU0Z0/R9RUaIKf2rQCS6Xv8uk+IlegJuynAUIvQ/
qM/P9wEshS5D5GMfH7/6Xs5mWuQaCCsm4PkaVw2BFyOW/nbqBsJMFwxH+dZcn81U0A/iLjz8DHxj
RJiq+hKXojYtYu1Be55MVZTW06D0+TwQaQYYYwczrnfihKI8yzp/7aQHPpFxFlX21jmzfItzudyP
fiL5EgwiDz/pEKAoPpHmOkz0TEAy8Ysldc3oAiCwFcVqbgC638Vyrk250ebfXM4tARj6+L8qxwQY
QVuGP609MoPfUI4k/41VitrwNVZoMXDyLOi96lwDd/fIGTdMXOIJaSqN4qSzKQl9tYaMsC6bBW7/
XNeZ9wxUa78u76oDnRdpTRQSFBeYSIpH2guDwZYVqLPQm1Xix4jploljVSgyN1XBid8clckwV/fS
dTtygi9q96QkY0ACRoMIPsqci3nRLj1FOrdO0tldPqYclJY3eaFers0TWGub6Qldwo3XfdXN3Uor
6fM8eZF3UZFhEJnWc7e+5H53WqTZTmsEWBKPixDrIWOu9BC85R6BNiYb/ZpMKSjFzvkXMNS8jFoS
xdcVF+TNB5yT5554quwaIJRO4y97nE2HNQRelAI3+8RkQ675/4m8MAckkd/I3oxoGofeQxGuFBR8
+XeFhFOIJIVZ39LJNHNwLbJU63l8KhUiTbj74Il48PxL5TZVbVmpWJGwOaEB3/nMqrj9cmBNKV9P
nIJR8fEr/jHoHo26sWe0M+LW+rzdKsfuWMlDimkdXOqurStBR5HKpU3CUXbkR3AkBneTlHqtp2yt
FWYd+QqIILdFkHBdXFqy7ZyQIbhDEmaIkClhuUA2UO9kqIP6hultFIskMZc4o8BNn9JheiuP1e0O
PSvNxHdpfbdFSmgt6Knrh03ypjKhsah3AQHnmGcY3t0plq7+hWiDpMKUOWtaQ+Rh+oB/faQisNGs
WnyzHkIHJI0RMhcqPbqcuM/N7D+8glDRthCORwOdHNjVJ+2QRpsbjxx1EFobsjLLKkoa7OdTmWDI
pkv4fm6T2A4OjXWv5eyDNXO/MET/NYqpb0y1RsaUmqQCF8VHYVrxniTvWI/DyksCIhU7YzxFbfKb
qUvdMwrAMaXaj+Y5lfV11qCbzqSJqX4j5c2O8O8YaDd5c0kIFLe4CbI+ZMRa19YYghbi9l+rwiOp
X+Sz1uldtSOV1SKCgNyfxPandHQWeh78h++jK+Mj20mBC9V1wMRgpYs5u/LCIZjerxQke92DEOr1
XNpCwHy86qolWEsofWjxn3htED5oqDraHW2qBCGJzlnN1eKHOad9b4td/1aEm2PfWPh7962E3FHw
vas4aiScmLUZ94RE6CAH+6k9AMI5hC6shy8XVhzKOSY5SJKPvEDMzlAtg3qSBzcle7XjOmB5RuHw
1kaPFkC2TrNETatcbuJTTMLxz/3UiVO0B6V7CX47t0gI11ahlO0SENDptHoblSE0iXAqzHtNxRoh
bGBLYllDtpOyT8yx+LaHaIcBqaSGG0IZJPyxv5P7iBilhPQ9dB/V3V15rJUIIba30H+SSGHDPd/l
TxjDq0MvnkgdgsNq3QeCRDtQc7FGMzQEEJ87vgVd5RmxAANFoTk8v/isPB1HOjcPD6rwjMbX8kwi
ePFZHReFgLD+HFr62UUtJeEhewze4o1rTO3slH40Qk1Bzta8ntPW6bslmv5sLCXUrRHgRH2IT74o
vyhqKD0PNo5KdkLtZZuK//PBChDhKSC/yubbMZxUuvt3VF15lDPBbz+XRQ+iuftM8t1Nu6/8LI/k
HEbTPBBSdVSEELkW6zA5WgzBuwjS9UYWQMXWaElE3qXW1MdR4X7X8m/QXzE+dsBapGAdcomt8DhY
UlU32ZlY5LrARuQrpunkm9SzbjEk+3NFSj6bah7UOzzyJdUzxrIwYe7nQh/pI8VbBReMRXnpGLFG
dugLSPBmndPzBFAmh7fX7eZDv0/XeeDBk+CTJj/mvt9Fc2Fp/J0jvJ4G+PCHVxgVC89uYipvBPgS
QW3JVnYaYnoeUVTPwQBL3rIChQpNg/opidauZ2w4QAcgUb4Neg85LC2SDWo+Fo3sIEV8mDYhdnYp
ZXehmZNIbam9nyccBdvoZpV3iNRBIxftrzWDI+fYm4D/UlRvYOFfxBh23rZ8MuESr/m1fSwYm/4m
2fYK1NDL7iSrvzpcewsUrXAsg7NwGqLghtP5rfxH8FwHepHtYVNx1HndDrq8zMtLtPuY5l42THnr
FhRv3eV8BeCKdcHJBPZtBp1bJ9+tieO77WqIpjTP9SKhx75QS+VGorXJ2dnzcVYqtrJsK21WhTVP
rKBECmqUawdbAjclaNfRvV/cmFSk3N+o/xTRSv4MQyaR3euHE/TMtFSdDX0YNmv+H3//cEMR8vmW
VtWASggNUI9fevaH2M9j7agyMwEmSIBtqxYb8JPrEg8kOUFXM9vspgRD3CQl2Vx/S1eqRKwQqgd5
pxU/yXsetm2FM65qmPPGFQ2XG7DdCqAABA+2au916Ajiq999T2OgsFOI1Rs66SBm5lM8O1xVehX0
QsQxC/fslzz5v4G8nlghpMmoN5DwniBVTWFQFKyLOH9kxmKV7BwGkweja08U7wKYX1Mr7kbT7W4T
QJb/rB57jKlDIceJ6oHrCo5XfEljz/NyujFO8oA4800aJsFM01HqX3qwiv6FCLODNYZizQ3rp1N/
7sOnjsQcdUiK47nezR7LSZM/mQMINy1CRG/ffggwHpYfN8IwA1uvTahyYWU8n6EU/zhP8qI7zF0G
EEgvFyPSIjxC6RCrWrxpkKE27EhedBwq9iYFdVBVjvoQl7G2h+HXIEptbYUAU6UsXq3kZn35MmJL
GyIzrIp3gsVJ3flhMxpsCAtH0xfC0V+JuqtkJGM3vTu74w7m4G6gXpVfxhU2eg4iy1fWDmZB8m9b
EkX/SI4zV9F/G9C60vlFuzCzAj0PaqFSPg6BPK0m6DpCN2rgINmx0i9Gxll/wK36QNTyVqSYqkV5
8ZveRahtlWX+hDC6wAQEEiQF3lwdr9SV/PhZJMRERx/buvdshvNZ9n06SAkReYv6wTuJaweeCjOu
amh7tdaLZmkDoLZR7ThN6gVqOe5IpFUFtVOFQ7dG9OLdPSlwcUo3npaagxs5aUL+ykmq72Qszr1w
pVUnS42k+8ANN7lxkjZ6Ox6FE9EpTZqHP1NHujNO6eK/CRKLOxSWt7Cd9UXkR/zNmejIhIapTrt0
rH6XzkYeH/8mm+UkhKtFTEE7bfQN44Q3rAynGimKdUxJNhC9OuVDIlA/PXqjGP7OI5TX0yeLQTYP
PdE5ZT23i7TMGiZ17H4xcFW1uJG0BKPv9MWcY6VTcv+pdkEmRG34OrH0197DvxXtm49Gx+8Ui9F9
ip+OhaLvgBa/u39mkb7UzhfpFs3pZuil/3tBb/Rmlckqdb/GbuceoJeEPXGL2itNAy/1k3l7uB9V
ySLcbabFeCgcX9F3YgVD3dunUT9oTH4e5vGt0yi0TSQeTBqaDUPyzZlfJovYYxw7PsGIgkJNXRjK
9oCyOto0z2n8XNJ7+7FhLYQI80BcimSqw0kYKlY+LCjsJnq1E+fkv2pBq1uVN15YtojnJN3ybesJ
/VuIbkBFcd6e0t63snzWJivZM+2+9OMy9UJ5qnpnVyZrmsZQT2CenR6n2ZMmE2xiEeknldTX9UbI
PETktNPDjgeiYXmH2m2OcUWHyh5FdTcHm9CKzTwKiE5AQ86xrukY1XkfC+6ULjWKCMVcSY8p9dM7
BCuUZmE7qldEAtttXPr4MHhH+6paH8hdpZmimIJ/eQzrxUkxFZiW//CcD8iXy4q+jxrOUp8c0/pY
DIwrPPlC/B9eo0PKXal9SJ90ZrOf6NQz3uK9IdhrlMi0fVQ1zuwCRvwEPb/811qL1XqmN1WW0PLR
5SCbQH3zKMh822MS8qs78+r5P+Dp1fdtoo79HOHYWp7WsvVaZKwYZEydDXE1rLGhNMCLnRCCcJDs
5haOlgNNvFJWysOLCe4jLTNHaGkM1oYWXbHl330eXMDLfz7On4j+MRM/RuFFLyolbxeB8c5FDuUp
udTPKJY+8EoJHfkWYJhniAEOSJGLtih7ef4fYIpjhONvMP2jZOcNlgukDDQCjOERgmi1UiVGPPZB
gdeHFf+uS0TM6kzVOeelOpGNMQLJJ6viPic2NMAfMeF5S4zk+C0RUWNd2YHwsh7fbtOCKJTbyEWt
armnaNtY5d6h1ysLtc1cKzhzd6NN68XquE66lcMHdLe2m8WkDQTv03E5GrKUpsR88J2izMdPSW7M
OkXnvUWGhuQKdlcBBlZECqOhFwbURJE01op/L1xlUq7bm6FSGGUqZ/ED3He4qHURzbtKg/2bGjF/
FW6cdxuZDQi+JJTmI8paYCeDhzHejBxiH6HH8PwkSFGuL76eKz/xIsvvy5HKEUevDK8OCB5D2sCy
JYkdw/5XIFbc10TEToawhmWthRwjg9uBvmbwmoUB0lsgZd2Hci0w0kJ5K50h19t1CGgp4c8AXTSC
gjvNtdNkY0w15y9akCbpDmHiIbIgGYnthkTWecBpjN+LGdQSQABb3WbmAWgsTJuk9B7TOYM82wy7
l8qGZtyQ7PcsYhUGJZJQtOEhP1tnvoSu6l9RG4gTZb65oVbt0+baOPgfnoExnzsyuMKUo9OP2qay
/iqDkqrFffD/VqpPrdKDJEe3TBZC1xJhqrXlkRkuKIi81xpmGyEvpG84ht3+UxpqHCvrL8IGoUuF
/gIgpLgGWCs6phxG6GFJRe+G7vtweo+RC5qJcaQaDVroqG7r9S+WGapczxToPApbYToO0HyBEGhU
fUt8AG3t0vSWfYOzNohB0MMtToqEkSkS8jmxEsphaMBGjfy6Av2ncqh/iXNcaD28VQp/8pdtddK0
531qBn+4KHagvxNjK6mK1b4Rx+41W/dDoGu7Xu2jeesHycno/CpjjMY3T7VCN+Dik9tdIHVTC9hB
/NlSUkkpdA9ZApQP3AZHDOIlbPfktqNV72wKa5puR/T10+QSLE8FOcsNQYuIORO5SG/DQs9KnFUT
pW2x72c5YRsz2cqElTftX36/HSko/D9dj74z6ISGXXROtnmEKPCzQEz3i85P5vRUfINN2dA9xQkH
Nzi+BvbhUheJl0A5HIf5c5fp5A5xLOgbFn3imHJMf1JhEQX0TdRwEC12cbdNGCFxXYFg8lMwMSpL
wIloWX1zeOzYXOt1yWvcrYtEOPbMFcUKwbcJt378V5PuhvtCwY1cU55q5m4FepCMPjls9meJ1pgD
NlYeCIVEXn3T84PBHHrk0UBaNQAiz1Mx3+FaBTsXIAFeoWe9D26VeJCxDzNViyK8zzlNVeSle/Qf
QDlgSMH7V5tr0Gr6xzpJ3ZDWHvqpBPBUkssPuEMm8xZwjZeDRxZRJGHncOTqZPBzdViQIhRrOvtF
ccq7tlaVlSNCqqmqzAYMIW3q8tZ3kYWLWidAxVg6ggssFcD01XEqJJixMxCdZRQsTI87zw4V4T0q
lLTbYl4MT2AJ50tQH6OsfkxYAZjZtiKqfDDnWMFprIkeXCpVwzFL9cD0YByojE1mbwxxgLxCrR2i
JUoFgJPMqxbTTpRzLDVGjTs9m/jIJZ4nvilEk0CTHazc4mzyXEGVDE6Wr8gJYClaJPkyTLJcbPbl
ZWxRRVIzLYUqpvkGLRECBTkSnvuy4z/ude1qcifYFCeclCV10Xl+MnhyAowDLO3zjE9WerRbliMP
ezxuNFAbxwNPjUlm8FVKtQ6fr3zqegXK1XnmkuIoMWFMjPlOZLDs0HamegA4CRO69gwy0wx8gEXZ
7wMd3WJQdz8+FWda9CYpNl1NbALP5kG3fF5Fsh1HqSoG9z6+BY5eG3y9l/ELpEPs5fqNaxcmrzyn
1JbFIr8LPwuAs/pJkp0jPOAJ0z+JMb2hJUbdkq5NeoQhxktxhAsCSJBhgLwBUJ6tyRslMcTFRI9V
CKwz1KCZJ1DJ5LHr4F56Zg6Lc/8VNoDH4B9SlTzWBOokpcGF4gXF1wc6eakut+hWHrJoTtyPaXPS
JWbyutU3dsO4gLB9MHnSwi0W29Ptaxh3Qmfs71bOBb/116ao9jvaeJOuPbIq5QTlSqns4KqK9dsI
/XCbRkcMozEuIdgzJiSDg23Fc6x5IfLwqyarvv05OlSqP1dPB5NG4WLCapptjDX2CbVTDkGe81qt
CsCnSsfkE8KR3GBM8ohdLn3wodnPxBuHR6LxrxWgQgcDzt4T7aqYJ/VKoir4Vl37nOPZwAB+igGa
C4CVo7LVq2i6qu0sGolA0/EVa/1mZtcjnVOjs2CFGJcA3W6UN5gTYMTS+ocDDEpOYUWkac3jPGpZ
coXSAnZ8xdg1//yEqWOyRec6mcAbuMGEMUumMh1phm9p/56E+XlhbBROwqqEyCpPy8/4GdO/j5tf
dDIYnQckWWpZ3Mxf+F/EYmRUJQ8+/4JqfLvqEWideFpleq2Uit07N2lH38hI76UwZoJnpkJSBVS4
ZTuHVj6IAJ6jyd76kd4Rz9jkGqCO9nchpS2e0IEJWOHIADqADLJxk9QOp940pOsi4f9fysa5J7dn
2HHmSS8WpXdOUh6vB9GSZk/RpoQhcyWPj/R588ftRY8CIlXI4pgux3y94NYuqMFl7X8KnEkCuU5V
QyzT/hq/ViMx9Lw+tt+hTnPD5od1sJ0k9/P0SifHS4QuUd0ZF9cDUlhTXXopHv9ak5rwZrKkfv4c
VHdw2owqfdfSEX8ttx+ZiqK/r6LQlADnNzTjSrlcYshwnE0kKJK+SvU+TMcJ0ZYcKNG5/MxbK8AD
PfiPj+gHXuUC9pxVj/gVJC/GPYN0/usudurtXR5KJgjMQmlfk1qOyLihessP2tQ2oX09WupywqjV
sP6A17KYB2mKjN5h3wa1DvsyiM6WCu2iT6TU8q1vCbABc3ZbP4wGdmB6IULh8i0Yilf10gN+buIw
+dHWsshkPxVtmxnPEvRyv6ze99+dhdbfPOtdKxolSe1necqsylomwbgIDFSJnjJC8T56hkLGu/Ox
7ksdIpAvDRroIRC8Gd61McaPwpD9hKCcvcT1D0lKBBTCs3oeVY+nJNO1ZL1D2opfA+zWT9kn7i3P
UVVP2/ODcK0uW5aIt1ykltlN8wiu4fse38Jd3RsaFEFNlAxb5bXBHFQbTk7ddvrPRSZuvpd0EDWg
KeFybL19Lo7IXcpU1pgKzJVixiz0ZzYcNo2gHz+Uh5ROq/AH5u9TK6GcPYtz6KRBpSB0GqFcmQOA
7IdZu7HgV7KbYbvTLFT5yuNTYv4ElRX+sD9cXkeEPSULvA78c8KNVwGOiqLVtfJMOduNiyTOCBb7
+q/Z92TPQqdFfQSIRH+fyKAEkXhdmekmOd+oZhnFTIiUVXRKBH9WHobS0RfX3OM1/rnJwpqNHAcO
4SWvE9FeWLGooUPbUUr76wquH1qQ7saGa5sWVC6imuihdk8JF98afaM6J01+e7XH0dos6hPIChJQ
CNG5ittXhCpJVESXath3f6OljVPyUw5ZdswpQ9alnxoM1s+KO6F5Uk5kg3REI2aQKRTR/CzxUs3I
+bC/skiec7To2oy0CP06dZgYQ5wlQI0oP1+3tpkTNK0Rufx150b0fooc6sI0aYkJdE1M+6OXUero
inCZPIMRuHXWl+F/LcDUOIoeYOs4K0x5sjbL4IZ5wee5Tuf0DjTGk7KJbZ86xMwm5EAjsRhKZzkg
LYldp+LQeiC2JZi+Rb1FTGMR+fclQqohx653py7gZbT4V1yBt2Gms/adZeyvpIJk/Bll0sIUy1/X
dc5xQRlt6bS15sOT29f1tZ+jXM/Pvqbt82bV0lddSeJTF2rDXuFWsg30VlHQTcd0ZRqFh9LDUb8R
XpIfgKf2y1Qk22Zj5rSW7TJ2wU78i+uepaBdMNgbOa064iOTv2XUx++mepjsUQIV1zZtyS/RMk5B
feS1zEYhpInl49aBMNtcFKKGksl5vgbNq2qVpOZJk/cFHtweL+ZBWMJK1h7b68XqBM6bt53MU1yL
7TclD9dGHOfmj7Tdc+SKLbzEeodNLG/sMgDoltBeAzhL7JCehY3lQLx5oKIEl8QJJNPgd1298VpY
hGYxspbhbnFUiqcP80a+UL6LBSOrRUm7LPb5ERbuUDiZrhZhTIyTw9cxET3+MwxNt/Cbhl0k21w+
uqpeEwYV/YKK/EL3H+ntPkHyBiN6kmG88q0dsve0chJS/sVXM3E3WOzJcyRbVqPZiiAvSqcClO81
DTUH+b1HAHOSL72/91McR6trSnfkchNiiRKVNrKZ8GmbFUBj6YZne40XGhJSF03PlYScURUxmoIa
08VPbY4CrSa1hVTDB0++UXT+P8K1LI7lcRUwmNDUdsIRB6GF8vyLVvRGYrzHK/dfHaVG+bEl77po
qd03OaYNQ8T2uFJ5vcxeXZv7ICIPsrkQPi0eaJhlii89/b983iyV4f4Ygm3Bjq8qGW+/4ATguFEb
eci2r0aSV4YSxYeRDoOpNFpi6hDvy5Remz5Rvylcy5rnP0tGz5u9gozaic4DKFEGhzc5Kq4/VcWV
vbN0SiPi1XAtKEU3KnpSYgiohqbIhNMXFPmklRAOm2aIGe8bmCMZbH79GvK7p4w5yVcXBgOQWtVx
MhGeBtONOuvgXpaHzeyLcVhnLooH5XMlnWTFZyBXZ5H5YYW8rIGh1F3TebA8xx5/DMuw649oZ8/k
AbK6LV1/vJwpi6bPPCwCRP5sT+knXWQyDxWi+ZDigm8nGS0bSI/PQOD48r1b6O9Fj3r9X2fzGTD4
sdaNmSNuCT1b2eDh0EJG1lkC5ydyUmXmVR1+FotKHJDsn4W3tlw944Pluu6CAalJtQQ6qkfIBg4T
28SjCNhD/TJQS+r0W08ziFJZsTv5JNF6+1arPzrKwj/wPnTdmh1UGYIPfUuG345z+UP3jMItENfZ
H0MisOpcHiy2d1hPJ6+V8BfbU9eeyqncfgDm1FvsFZ6dGcHfLzNd66xyiuRFcUwbnGlMXtvjGRrA
rkL0hSFaFiy3bIgOGwrMlp+7l6EtTmpPaZ9tvHSYIbzYlclcyzk95VfEj4F4C7ZwtunCH8GaBO89
sUHho+qsbP9cDBxF8iEyebd6UziOtOtTtDmfZUmNVSD1TwlzbDrKYVPz0yPzLjNuI/t7od9DqtX0
soZxFtaYzrdMr0J0ApGd2cJ9JB+5tBMlfBJAKAk5H1aSWDOBohYI/IXLPMIgrerkGxFnyEv+9vJ7
MCM7xsNLBY2d7OnyflNqxXy4I1K2pRxLTmyRa3GtidlBKntfXRyjaXdUxphEWmEtiX85Xi/TP2cx
I07xRPy4J9GWqvzVLROmS2tHvP+ZytHvLGU2JhlFiOrn4rBi62lSGqU9doVEH/yoMLYXXpWlkXTD
IjxxI5YMpJcg7pk/7zahIHllxgBeLTv/gMuuJ+/E/Qarc54pZz9t/aTDxMwK9j7szH7kybOskhta
rsNQ2OlGgapL984TlO0fb9uPj8csFr0SPu+5v0RYNXK3jadnazo2O8o72CV1xUM1xqS6g0lap0OQ
pIDEy+gYZkfdC52PatRSgviX4P0wzIaN7KE8wL0exmASmVI1S2YqBwZBp/bVaPa8tk9lceolVD+9
i4OzgEh/v+wfNO8V2iGwRp8s+N/5zC5T7XdNv29qhoHAgdh0kx1Px5K6hIUCxY/lNUTqo+MKxGMn
2swoFS3xXq7AkL7Peu3SbZB7YuDN8JlipwxaAsTzDUzSVAoIRFIS+NeOeuaRl70WZkXMRbzk4S+u
cfpqX1f6LKEdFayCPFbUZC/QnruOrQxFOJWdWpqwnKiLf5BT46clQ2xTjxhBSroctM6qt66nJnHM
p3UUy/3iREsoaYlUC4Zd1P0Xq53925CH0g0m2qGRZ/yjJU3VQAamv4FDAxer8+4whucnZk56bvyR
b9VedicG1r4CEpfYCGdaVpr5zOalAUw3gXMQpirjStGvpLkOfDls4IgAGq6HlDAf2kxfPRNpjwwT
qULTmNfvtfVeIjleJnD+moMI8uipNbQ8LCGo95yJa/gWraRdyeglHP4G0kDRgYlgkH98NUqqFGx1
oBwP8fTtGKeOjEHCsOX0OVleXhfBdOGvb7FYrha7gg4Jh3SZ03YwdsnfML9ejcRssyMrvpRtvMki
aLYq/apenJGFjLaAR6yf0dkc8CIbbrVFZUFCy3+yyaekxLNsNiD0yQWQ9HaCaSyreSA0VLEdt7b5
bX7ym7KQsLpSf6zPgpNr/ZhOOppdrsISaQj01+/fbfZYhYfFnvj3TMK+1+TFkKEa9kjGL5mURONE
RGKIrAV7Ehh9RgyUE7XZi/Tw2R51lOm6c34q6VAsVq+jGfl6o25BFNaP9128sl26Sk5L22YmDRS8
22qI2gAEHGXEZHv7YV+9hY/ck8q3VB5gYMmQrEDOEd7zyNwqWPxewtl77sePiZIXeelcPE43cW8e
EQDAFpH7wQrmSXHKl+uTe6VEjuYzUNf+P2ndkQhuP/67oAtt3VpRkmNg8ZAqIxa/xpIK1hozztwx
Cbsng6U6rtAo+M6HcrhwZcgAHQOAXC/KAUEKK5jHPkuW6VcuuQLBXDsA1b4rBefF5hyo4yMVYJex
YrmhTedOdpka/usDHJ3NHWBKLie6MJ0klpXZVMBaS0ok3pbA9Fpk7LGR5sFaXumNLuE/gfKo4o4i
Lg8ZX0DduZNw3aQc7I1LFPE3awsHITs5P7RMv4l6+7BExVk8kDXKVd8WQMAC4+16VO8LF0AKk4Tg
T79WCw8mwlbXLxaXGukwk6tuRRGv2rc9IPlG/7ciFmrO3dMqytYwiTUvlj8qToAxkf/YyErnGrnF
MJd4YXyHF0maGIO2qV9rBeKn/nJGlAA3LLErirUjuxzH8jnmZWfU6YemnVRA2zXK1GwrOmNJy+ot
MDZqlK5DJFUrL/HN9gWEgF5iEXM+rUNCmh+MF1uOHY+9ZzUWqn07i9gbHX1VJ8e3AIM+ojH7UoN1
XNf1CfyHMhh9Khf3GXHVHMPXVYmJEew6P7tNrnR4FVb3B7LRpdC5H3Jr9xHj7zwZf4EEbkte7UaO
En9q410236/vcjTWiIf2AyjBCWLM0OYMfeM3qVPUAGeGX54bt1Yhf4M4YrWsk5ygKLrZFxHnOQ9N
aVF3XGSsku8+bEEDr4XPbObBzOosVe9S+V4kA8mU+bKfD2vAUaSz7A0Nu/ZO2c8jHyKfgkcfSDFS
J53DX3dg813By+SGBSRSt1ix8XbpIw8MRNOUe9SOHtTJMws8GXRzgcnca6sm0xtJ61Mn2sFS/Z3m
Xq5edB6bDJM6EtERw7NjC2l2BKYYgBsyNDUKW+npPPree+RFURdQZm7AsmrPl2C8xOLXnv6eUYMC
HeyjKJXLKvFzeSK6+jMcFQc7h/JRNXHOXa9A6pX7TtOdyBdtj+hxhAqZOq4wZtp6hBsTMLix5WEY
Je2hQBsZ0suNpK2WxVrgY4mOeaO/94jXdNnOVBpr1z2r/lmwY1DOrBgSL+MNTKCNQNxa4DQQDAFI
k/IevS06YRxPI7gvBuqNRvr2bLoHYoJdjLyixc6AaquzB97k0Mu8lNa/uQbesH5tEgfF1ME1Zf+D
JV44dbzP86vJ0ELgqX7kQTDDhRDMpQmt9Tl9tJiE7yF2EceeQuDyKrUMzS96nxDwU0UuHEBlL41o
xnTfdiOcXv8Y5tvwzfQGsONLTGzA0wIqpy1lYWwKAo+H328Qp1lNXnt1Ho532bA7+PpePXcXNZUy
Nsw42tSxQjTkTwYD9sFyoEjzhOKAeRTzmxb4FnR19z/igbPWkAukyCa73AfKBVIsLoF3ctU6YdVX
rTLWRMaWUpymFS13ORg8BND4C+om2GaIGtw98L9UCqNZGnCbYGZAnoIHrjJyY5KdtXGi80R4vdZo
2rGZY0ksp1GbqNaBfnExhRJN4sq791H2CF5SdhfSqtVU2/rY8+4ZIed2Jx9qLm0gUMhvZYRtLxOY
u6QCKmG4WnxdG3a2BjOfeKwDw8rHeMqVB3s/bz7KqpIuXkVDMRI8Pm2vO5YDpoG5sCwJ/yoITQQG
zp1chHOw44P8ZyHY0aPgFn9K2qn0i7SBbycuzRgTOKGQMq/+4+e7emH/T2Xr5rdSWtLD5AcC+zdi
L4EpU0QpVUr1lDtS80aKpiTUg9pX8XcsvDJk4fsFaOfknRSt/c9LGE952PPujHUCwVAiK4BFPYBd
TZiJaGRYHV/I2RD3c2HPwMfZlN+hxWJdoqlbjcI51Z1L5ImenAc8A25lRyUJroFlutBgVt2zQpIe
yz+i85gztOsrnYF7B7bGtpcNhOjGqvXbZuK6a4peSVjwm35UnJmNoYjT1M6CGkt+MR46Y8klodsh
n5boAEc/YTZIFVQcTrSrApPKfKNjlZCVQukomWbLBBGm8UupHnkZGBLlXPAeCD09pFL6NCZ5s13L
MnKO4FritsfF+4ssMUCg4Bn1dQ17sErYPFb5hgRfGsblfFclk19Pr38IsyPY2BFg8YdAFqnDoFLY
KS3cocbgibt7478nErqVcddTWrpNUGQfW6NYSSlwO2XX/e5LnwowIdmFOUWj60O2rpkE69ThpZRp
5maFstHsCK8VcvS39/Med4N4JfgqamyoWOsZp0Tqycnwrc8R4Eo7R/euZBFNLGPQExTrdhkVhaCc
TJsUmeupfySJ4RwzWueJwsxK1luWKD1mtXcBka07+2GhkJjTg/dxyYbuGLU1Y6zYcQd03OgC0rsD
adF1GKXjD1moXGdO4kKdANPb7G4c68bN/BJ0jzDrEWTM5lfCJ6u1L2gvFPW8CtYBAO+nqml+UfOZ
sgLuO9R+AWMlC7T8SjVjPw+n/CuI0seii4V96IcwNZ3wCimmc8GVmMchreGL1RX6gIh6P9YlLXZe
n+go+MS6Ke3YTWuBrebDl2GDyzDvHjOD1Tv35HwV748EDa6+rUcC2HqpsqZ6ljEtTdiupqD5RZRJ
+FTkc5PkobXdhyVHNEXzIfb9sWmVW5OwtKmh0M8LxEETyf+OMk76PeRW38dmCjJ5gahhlCpHkxz2
Al2h++e/tMNBDO9Gp3qMeantHhqA8hzzXdIRgbUR64rwUOL6L18ig8ZYePB8KMtwdvHTolzJ3Kzk
x+qa7ugmjKovM2vS7dxFyv/jwDhtLlIqf9B5+wIKH0WcujRXzZsZKgrYlK1NQs3q2GF3xvl6wBtR
M8tH86LOhK7qKw7yHx/A+HxkysiB2sXzYwIM48K9oYsfeCZcYCplIbxejVXPQxXEMTw/tIQf9qeg
4ZUNs5iY8VxKDytcIrdlxE2zRZFShxKFcomNjegbPrXfND/2jjTGkgv1B4c6O6BBSX0lidEZyh0f
0DX00r7Tb7UXPRVA1wwrS50kSe72vF7bgsvrzwaw800WiIZUvGgu61uISLVqgCydl2UwId2iCUv1
z9Z8vA/jzTYd19KXEQTThv7H8JPrw/QysKQRre0pBsqy9Cj3giuDy0pmY94PMirAdsYfKhF/2QiH
sVSRGdc83pW0IVgb1mCjPJhK4rT1KehSR7+uTSw31DbHb4WSsBMQsVJ5Gm5ZESEfgjnV9LYJF+eQ
ovtJAWXrqgqYnf4BpwHxZX7JmnZkwqAJWqqEgGZ384uZDH0xenYZdUWpPS/b7WGq7wZxubxYFr1B
Pnqs83IU5uXKGTcjfdRbN8yvg7VJZuSySd6u3BycI1MlQ7ujh9hp5UOCccIMpKhNbRPmtCP9Xywi
S9J+AetGcukax86XgD5NvVWf3OEr+O5xdew9WHt5cBg3tYXXS9V6EMr5QApawrN1Jhuad5Je2QTQ
8iFn78f0lQ29pXYQfg9PYztHBzqVEcVLQ8l876XuD4EbiQOW3s4CchF74w4YCiiReu/HNYchAhMP
Tp6FFcmleE3kfpyf6XrbERy/2Fx53gwB9Xr471Paxt44gFqxo8Hi9O/AaFMu+14RvbLN3JpckA3w
YyxmujaR/fSTgQ7CpPRBVSAqhKejjdCUypVau/zw7MOuYasyEvBR1zPoL1UkRB2Y9S7ncQSFQA6m
24bAS8P8nYOy41KZgfyXvtyE+G3rTHvxauTt0YorAHL3YtRvDGjOCJWuWjwYsFU21guoWrzC6WOI
xHp0NQo4cnBbu5lxF6JaB0MbDKaPjW+EAU2VsExBmF02JQ4c8KpkxpOuR0kENSeJri9R0ZxR9Y3q
JAAbQHcaLmMwaMQLAJ9Yek24c3Eo7JWL3uj0dWMfFqssBedkYlOES+KjTNBSUNqk1bz+iLPlxaPG
LaZ6HF2N6DtAvbnyCaOW1KXLcMyQqArl11GJt0FwQmXC0HY8hHIPDVVVtJcLnOtzPTFyxiY2KJoZ
p3PNKz7O87bVHn6s20bJdWVexsBfrp9bYIyzcRfkctYjFRm/tEmXgU/S/vFBXV41y18HLMXlVlfR
eC8kW7AMytAzoIZKZwxmjFUwnFROXQss2skSf/Q8r5118iST5CcjY5nb98OWf8myxwGV6GVtkse5
5mi8ytqvnd5KMxmHbi6IU9kg1Yvx/ubC2aYei0I7M51I3GEqE/KQobxK72/DYpXSISP9uHkCnYm3
eg0yO1vL7M8qKb7l66Gf46DU5JKCy6Gx0lOuonIfGIyCBa3cMTrLhTSCNexEO2jSX+9VCXQg8OqR
iOoxi/I7ew/JohXgDXb8hX1KN70NR3zcsTH/+xF5fL8mzMQ9iDrxjPZ+C8RJOSz7sMeGBlLAv3Uv
IGXR43J/D56At5nZ7frSb5NwfZYrF46DlHPvjC+gJH4nyVGGtQGsV+jehKHvYgWP8GIiSOZm44ZO
9jSc08qeOVx7zcgr1ulUcuMf41XMtaavYKduuZCa93h+2YMBS7Pl5BhybvSX888fy0tUE5I0zhwQ
y5+CHm8vLWaTS+Mzq375/WrwBBhi3PZdzxJlwkqKdLbEP6eSKbmPUfznXgpuvfXydAOWPqfO/cOM
1xNzfxmAPjh5Fto1VUjCazAAPpDHdvEWBdVUR8itD6a6WOgcGCR9mu79RJEl61QamwVO+18t+Mxv
Pgnk0apckeC+r52mB/KNJ3c+giaWV0HnZYe3zNzZ7HwU/U+7ryqO5ZHyRjjzDvgP0dPlrB4DK6u0
eneOm9tx3eWJc5FWDJSfr+EzddcVqg64UrIS6/QAg7Wbm2MpQWN1MLrARtwvLoAcKiI4RIjSsJ0V
w8Ya49vRuYp/v70U2mZZB3ApHPMdesWvFcDT6Q9UVElPutGPwhC0YEOEp9fnaTMYU1U206LM2jNy
na8iuhS1WXDmfWU8CTWzxaeW9/8NUXRCgSaoOYK7C3NfRFtegbUW5rvR2P0AcFQ0FVFZrEjGhFTa
PST8x0xViQ3OJKQ7tCwwMz74A5GwMhny535hW0F7ISN7vSRPcW6JtD+B7246S9koHPTHXieT+tKQ
Q81KLM+W52glvFII+t95CVbUHWBwuJpf1qzfwkkqkjhwibgWlG1SYcwjdvTT6eMwwVauuD0f8Ecn
OXf6j3I33YD1cY22axSfgFyWkBc3n10wjMzUjdqjRpN69mK49lNl9GkQSP7/ggFyfNJrgANY50hg
ER79a7xNbfNJnPsNBciu+BbDmjmsal9mUJhM5fg5ffpkwc5MHv39p+mdqxtw333ME7YpzBqZqCkL
/MgNQVZ5YL/cgzhsE9EsviGq4xDr94bzXYFghSQnBCoXhVgfPfAJxso6Uj7QEgMP7wpMlO+XV582
Y4LBm9WSpQyU5m2als17RJP9Owl0WE044XgfftYxZKoJAzQ7fX06do4mFlEMwm8cMMdO+1y4oToI
jwmeXePffv6ddvvjmqEBn9TRNd2csjLd99cLgjvp7G2nBdn5XhoACrRqNRtfISrXaHt2qbNXHjtp
rjbb0chFcC2dP58uvoyRQlZHZkU4Jw25ddXOoW9zWu5iP+2uwiND2t20/Uztw5cfF2X1hizDfiC5
0/JqAO4c21b/mcXwgfD6KQA5BzbnbTYDPxT2mr52ugzHHpREoihnpw7a7cg6oiw5FaN0N4hxQQa8
5YcADEuJT9focejVFQsyO0bQffhVumO6oNjtRLOfAbFmMgXr6fmsS2SbcVYRW8SXbCpmcSlHSCW4
bPEpgJuebTum2ijEuzf3cWU+FVyW1avnBPL1Tr3ahsxFWgHTHApFivfFq6PhDNvdzU/W8ln0p8tZ
P0AZfqwRZCD3C7xI5Klvt17stE02mvKWN2M/g2fL12up3nKD6+yF+p7EZ4cxaYTHFPLS6hxDakiV
hAgB/rLE7wSUxuMmvX/4YEisVeSQokhRE43xPl5TBxtfWZAKZlyYzsuLJ14KNqox0K6rkVgeruU0
yKEZLzVw2Pur8Wu9yYvqY1Wy6Le9H0K1GAOAJSrpEXksYjVQdLRJkWqIJQAKpqqQHzn5H9jbpuWY
9rLdkTkiw1EAtfQyUPibQQ+WmSBihBWYZeRttfC2ga3VbW7erqFba04EScJppQ3AOx/gE9pF9BQI
AMXd43D5FXJtFHEoLtrSQQS9fE/KMMQvo2DNODDHHFkBqWZOJJlsTHfN/iSk/Snm1zP2pcSDEuu3
4F+FCMvnz1HgkW7HIlksTgNwRBEs5qBZl9y8eXkjCFo3RaFlnKqXNN0JQA7+mKPAW5A3IgxWwKeM
1OMJxGO56ZJO5phSNcAQ5Mko/X+OTNdiy1C8Sc9o+6QNmeGvwq2aIU6r11JyXcmicA4Wi55F3N8A
bkN4brYYa0eQW/uMwPSemZc0nMswb5MUdrtWCnV13ScxAi3bxJUYmkmgCYkO7AJpDBnLWTSlv01X
hUQSGEKPunq2mB/rgzpH8CiqI78fuHFMHZk7PCL+/mY5Mrc3FfQ+/+3ATYKBQbz7WTfqoOehvXrF
56MlKIctTwuZLcsvjneeaitrXzvAXy6TvzZJE5prsCuLO9hHrdaUwPx390b2nPGujCEWgwLXsG5Z
ggkfR3Y4RezgZnU4DmyCOJhAcguV5OW+/RtfiH12eRJ58SZUzH5zPSeuDRYjh7DKsBg6RjFY3CsI
TZEQMkyp4QseE7lGU5d+TYnGO613gyjgJlqvdq7rWOq/iFI+q0GaMWmIjbuntNiupq8PzUzUbheR
ztk+WBCRPf8cRMlOJ8s0Sy41IbVF2Z5NuPojbOR+3QWuKiZ0eh6DxtbtUf+/l/+VLYRm/PF2ldvm
4phRd1cV7yvAocMm7Yf5HIUbVkFgMFoj6GQavudmEj8vZEip9PR9SYMDbUNhwaKaSwiJEGjDnmLV
i++MUqun3k83+dJfTfmkmHBJ/SW2G4BWZ6uaUxhbEu8UaOi3to0IresP5da+eMwFBOW0glPrmhwS
HMMLcnllvzF8knB9G7o5iN2abnuyAseL2ZEBse9WXLYqFV9SpDR3tyrLduaCr2yhUzNQ1x84myAz
p2gXqTyJ7VVkLgV4/Ot6smzoUnvn+IiYWm1+QM7COWCmfCVAffq5L70qSH9MnqkGqvnJ9JNsfEbp
tCDPFbR9p4imjzncNFH36BqgUdWA0rG0aMaZAJLTawwSQEPNHCIeiIFlBqYV3IxsijcpQsDGF2KO
pQUFrbGpbhsOIvGVtzEosUWrfhJz7iOsUhN1rrlenc5wHIgB+aEbMIdGF4ijVxpnBJdMls5xJHKK
6xo56wvAHoHxlXQRN4UGImOE7SLEp0w2dUe0lSOUQQhMgVjGaav1xV7fk0MAhxCkboW2p/U3foDt
FMWsNukt3DHs67NOYwx3P9FDP5N2gigzkIBzs6+zkX77UfkrSrgHBfaKUcZGm1t6X0bShEtnPLd2
7ytAVi/kZ1U3ykRaCP8Ga2kdKwXgsXCHqGofhwPi50654btm6d0sdkXS1wIVAfloBy+UMl+FOP99
VEpxGtTABskJ5VCbJheV14eAO3kLCM7puC/TXulGQBs8uJDct2BjexYab1ZP5uK/V/FCHPWFazsV
XhBOKa0h2hP1Y79uAxigrfzo5rNgqaqsyBAFy0EdG31RzF4SATF/B49F7Yw4jcOzxDvbg/kuoTP8
bS2HdleAqzeAFIpQBkfwxBslNufo/TBewIWa5PCOkqS3kqxU/iMobhaATdwfyWiojtJ6CEMJI3qs
GMgI5b/LdLh2XBMEb+O0uVTq+xA63Q5s8F8VkyMSKPriOaqb3pttsjc0KbD65QbkQKqJ221FIoca
ADZz0BL6keH/WwWgdu6yzaBrb6WkU05wni3zqhzrCtgoxC+thvfi
`protect end_protected
