`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpyGJnakVe4eFwHNRrtXIa+RCuZaQ0qVqBUYSuXeBLDMviHSfY1mCzj/qJyuFPr2ICIcOEezrjcn
MbxPF9P92A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jh3yASIkwwgzr/apUc9g+Ktqdivh6HjK+JJCNFA2kSkiPvq8guq3/lsaC7GbKg/5NEvb213QTPY0
NpnAUClY6RR2ov3dH9dPPxvGfehp/hqLFIhJOYWxw1bD77ybU6+oK/D52y4OgeSVwoBtJtFGk9LD
dfixFhvGx8OVLViTKeg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e975i3NxLBk1BMUUzRrkJfAcGoFyeKj+kFcMDH4mZzj0scrvT67hwn0PGdz8+dRVgR8fryKRATqg
aifkssK2giAkTb3yC1DuvJXSC3AMsnhiNS6Sy8VGya+H8Bljws4X+pe1HtzRRzuo+0rDBp22TIQi
L0/bFyYfTyP7D6ejN889ssZ2/ukbljoPx1swOnsUnlxwsA8pqFSO6w97kxPckife2KPcjnAYZKSU
s4W6RSxmY3lLSujk7q8mVCUbCP1kVFLkUivj8loLW6v/CVnYKpSBxfQEmL6B4Jzhk+hYUH4xvVcV
+Q8Id5Gmb0eK0HvEUZnAJBDVNYTP+x+PuG7rxA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GxU0Y2bsjWBVg8rJOCuktP7NuoOJzJE6OTkZud4AWKxcgnLEEMnRhCG8SWAdDCPdb1vihKYfJYeJ
3qphKALSH1b6XZb8LOuupIWTPWQHc2F7ulrntFyBl8mtoue6PiuP9Bt19FcvG1Mij7xJoPizusC3
Ih2ZyJBgc56RetQuSlE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G9RdG+dSoKCowy96fI0Y1/YdHwx3EZI9yTRj0mubLcYX1iSS9rpZZAWKkieTVuUf0caFzaiVIGD1
y8NAE+jmLKN/4V9+YYN5OLIwF9g5htPiyQ4UHRayQbf30FZFpgrKnFu5Dr48ff4Q0hOmRiimlY9V
5+vQ2b4zLIcjVk4c2jSrH/7hBeIz3lPFOa5NrWkqtd3sIsClvKV4ensnHUtfe8Bi5gjqGZyfYL7F
tb5zR/KJ1O8GPUts5kfYLnfbWvNb0tPf89r9SQRwbOy7Kr3172Ie4WNFmAN+V45aq6LKHt8mJRzb
sGb0DHhBkeZfnxSgW6BV6WX8CrYlM1Fweo7XMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10960)
`protect data_block
APWsJmm5d7bbtAZ09mYLoBomXjHha3JzaHs56x82zASpDO/fKS4DY9EzJ1FK/wamGneswwROEMe9
YAWwLOdGJ0zJlqQSY2tscOPyQiVRltdS5sudkTxfcMOhSxvrrzhX7ty4mJ8huI3g3O0AC542XGnt
qSHbuf/djPg24gBLeSasg5/aaVMiDsCXip/9ZSwsr1ueda6UvMgFL9OkITmYtfhjsN8c0jQRnkQA
6J8aeT+4Qx8HyZmRSllbSJZiM1s58wVnppEOSBK3oU53+IMEIjh13yRIXxQOXRbjU94t9GwRKQ9f
323qDnY2Da8u8m4fQi5CgokGLZQ0BA7ZxjO4tWhqmD7yhfUXs9haDq+c52Mx/xlzSLNvliqgf28r
Q8n8fMoePQ8zPWLSED2SgkypB04VuZNc2rTTf87YjogzIUczNLjKypaLkQhMtPYSfl6bCP6GfoH5
aSC0YXP6vExUzdMcBW7KKikkmH6+qXx0fo8lbr3xsN5VWvu20Kzx9ls/FIUtMJfhw6PHJyaUXruY
Eehpg57BBZu2WUkVsWw18by+I106P+z7fQQN1jWNxi5I4AeZK6wqwkp2m8KtGRv+ioOHkH1NBQg6
fyGZYhhO5xtcSProEcs213irV+hZdqpnfN567VwTZ5huFlgGQz+RpP6cBFNrSDn6eqpt73aZGA3b
ybYysE1tl1ertx1gmd42CVsfMeJdcCtUMQLxHMV5Hqt0dfxB68L5adJQP+5gzmH1Vp2/lyrAJQhp
QioLDrBdtNWHXRsUzBfvq/ueUx3JRB6TMUsb9/XnrAR0Ka8dn0r1hddz9m6Eui4IPCSxMjtv3CpT
EVuPUFa361oDsmdC2UEJ15KtewMPVekHtTWQnjNuqSwc+sXBNqjT2AwbGf97kW4YueKXz6vIi3OT
c0JXW0MV4rReGC2Njv73mrfq6kthuIWjS8ChfRrtqGXh6k4tBElzf98+ZTybGNMsFd9s3JaJiPXy
KKzgrN8v7Yw+smXbp1wOeyg/g5/DY/vyhnsxwkmnrrnU4QlTiXYTymonYN/OYWcRLXTMUtNv856W
nwVcx4iR7kPUSBE7gR4CfLfRvpxRJbvm2VYXHlqXNXOTMTMtA9LkNIDu6FQLTDp7BTvxpU1P4+GJ
aOQUkMtC7+vjQrTHAJvCUQ/rr23uayWgwXT+YXlW2QrR2JLYlWNsFxXrYif+A+GGsnqxaqlPHGqs
Giz9odPeHKOdBbXmGA/EIbUBJ9YAyHqvAx5LlyUPfcDgQQsHV2RImKUBaQ063GfkbDe49U0FHict
qhseZGXbeOmVfvHaL3nFXank1+oyF0k+aLRSnAAwxSBWy3kl19LXKn4Lk0ZJefeqIk1x6LSr2lD3
GFfZdGf1paGZf4lV+lEYsOBaLuPvuV9x0okXj+UYuqjyws0RpPpzOYJQXqrDypfNFoshzL2QG9ec
7l2gzwKW/de3VpE/KNPw4xgRaPaT7lvnm36LjfflS4akc/OyIACfQU5jEezo9W3B3migWzJyQkJr
CCbSKdjr3yPUmMKdG1ERrNiUK68hhfCHsqyHfXheXg3mJWsydwI6xRolGTAZ2fAImWAN6lQNHv9u
teXv9923744a87RLMLJ8m/o8A/ddZKA+00QWoGfULDFdq+rumXuYVEOCVq2cUWYKTc8Mim68R3fI
vtp4DdE3TIApjXHzzMDrOCIL8GjjpxW5P1/OrBSpXZzv5hYjoqGZ6zYyRa6EfGEIg6/aVN0P54Ad
S3rEtsXuYcSvgobTcOX4KLhk00MRednjslnhZum5Nl/JDO/NGpJ8uQQ38IVlFkHc7WYAzhZO7IEi
q01tyv+T7pcy2JPE0UHwB/w44/bZmUcczfCAph3Rbu0dolj84TIIqqgmFo+mheRXgPE9owZIpmhi
ZSYjRtVV5D9XHu557yhw6aazTVXZT5j0a+0qQ4WQwAOPEByShQKRbEhpwFzot/XC6iVmQSlhdcHh
2ciFb5cjzvyhJtuajxwbESy5COJAjsq9eUq2WmnYHrzwDf017ZaDIHXszHQPbjJopXUuCTlLHwLt
px1P6+61xWx/XqSDvGAXwASHWt5r2/BLoOERBbPEQLq8ZvYdgPtXSWHV0jyIcxhwNd7+NoXNniVL
o8F1xbTfEAXH3buyghhKys+hEMNfsMO5/4nfvudiKOnl5WLtR5+WKhkmIVgEWCPIOd+7sAoHIPr7
D/KCpvi/hRKQ1HkZ0eFSZDdob4CHsL/5QRyMAMxVKFT9YHZfW/UkNJjmrbZ1oUw7o3XM2yFAmX5Y
N1y7Q2gw1IiOXXdsqeBgXlFpBhue00T3jbdcP0DuYpdNZZyjGvshJdbOCDPfopOeDgYprWavRaY7
Eg+gOcxtsJSs0+N32ehdIifK8zqey74jK1DOymN/esrYaSLAvTtJ1GKuRRVPzYI2Sy/dviG0y3Pr
qJTC8H7lQYbBfg+kDmH3JC5QoziX/cJTobDYB/WDQNyK8i1qS9VX1a0hDhuX7pF6Kg211icHG5EF
x9zw9kpAQ8TrO2zBKNUSvFhShFDKw19wz4meBRrOO8zw7x1Um46i4x1muuQLfv0zaLzOjF+8/aZC
EjKCSfTS+7OJ6EwaqN7BkLbXqAznMbNePkvsi3l+XWtKSNPMF/0I/vOlnYznmxR1N7MsEEj91M8z
974HTSsvhZilBhUYvok2lvPz9loEziAaSkExpexsloj73GNZdGou8RVcU14mnwNC9fOkSE7O/2DN
7mm20NdrFRiHdQNMTrofdF0RkXbFxM81orUA0vHLDCPH4AP9sN9I4N/LWb/+wVx6q5nUrRQmwig9
5Y+t1lJDhKFhBn0OO/HU9yBgQOpyYvJBp0xhFUlSOsUkiRJnSBZ2n0arXdazcP1nBMP2m3vMMCLo
uk+eHBTyq2+c1CXHeJqh+qUM5USUYduiifzRmcq3p3Jxgfcjny3Hwm89AxrZVbs6RnKcR7pcotYX
sGKAvnxVi2pmWmqWC5qBCwtuNmpprteALHW0iTKVUFkTQLlAE1WNLJQH+yDo7sfg5k2Achlzt0Hc
XmknmHmwrFlD3GDcX8RcxKXGVGXSC2POHAr4oUhcr6TfFRzFN2L9fD57xlf4AH8ICmvB0y40rdFI
/I+dHSn0Emb8/6PD+5OFzpz2f38b3sD2WKMSqGdaUEBlCrtUmbeDPSLvXQtCwLpEkb9VRJQzKaf3
HdfEkB/CqCbJVvkw33SVP5lU5vCFiRlreoeEnn5gEsiKrQxqbvcljVnPqCQnHTLkcgnWWdYFsDY4
58SuZ/99AVwlAoGLWxDoROsacKoqYq5S9HcM0CFcqz6qnMLF/Zgao8U9PVTgpiUz3ZziUj4GwFWe
BBV6UMq+XL9THO+zajzDKtLV9HlLxC351P3VF66eBV33xqaJsefyS9sTUrm29/3vIjE27j6VfTUI
E5AHqsp0yJ2FwsTgvKdVbGNLJ88j+eTqlTh6VDeAMpAhRFkbZz2sk+AcWclny4PNUU0MDHcAa7Fv
HBuTBZPH8i4T0VIU/KA9spAcec3Qn0pr9iI5GKe45RtoZmHjC8HsRRYvisq54uLOpxd3GqFqBxLM
gifjTl1Q2pfGfP+PfunC+wEuKwmrw7pOlLu5TX0PprYsUYQxSP12rds5S8o5eCd+x/Dr9qiYB/Gy
0gcHd9as/1xbg7O566QXj6m1wY5Qj/8TGGIpCyApW80O2m1pKGjPFSFbI5FflcjKauQ9rH48EZEc
QMqh1Wiv4nMjLH+MA2DiyeXKzXWG+7K86C4Y3qCPUPEEBtjUPksp5ANnJwLfeMBqlCFYTHXWanRQ
ChxRo0lQbBa7Y1CyILxm8tGmBVVB1C/q902jpIvX4JxxAIcZskDqrkmf0vFP/VYx+o/gajbKIh8/
TyIr38iGAVUTZD/cWMBN23WKKgC/ztD8RYYBTG0tLqiURu9X9eLujPVNGTTwiMgreMlBWICbTWw7
JYafl1swcUoDPzMEhujDBl2VSsKNs/9wmwR9j7haUCLWidvFyyxUJ7GXJdGpw/wWPifh7+jPOJGR
U+rqxLxMFkoCa3Mfetwwe5+SnqTi1rluDzzt3Holm1sFrigeUsHm6sPsrjjpyOUWpZp11fU/cmL/
LhSJuEgGPITM05/lhrfp28UYnjMR3yZOHFUP4Ed++ksNO92eyvoe/Le7FbZ6dApzn78oFrpJtov3
2bKY7n2UYYDXJz9WxXOnNJ+o0r6/ddaQ2L7cZYePPeme2CV6IsobVoC1r1aBnYgdCFsvP5GI3EeQ
t0QRGwwyIVZDZ631pin7pWvc2CjTj6XSMjDnZUu4CIyiVKxZC0JGhYw3ksohV5QVka0dD0DmDgXF
8qvXTVmRKXAWi40pkVGUeOZSGwbvgr2igYdtk0kWmGv+NruS3A+KkIi9blzpMt8j7sK+U/F2dgwy
ndumq0BsprDwwmY6r/7ViMQA9W8Dzc8D3GIxesWLRLXDZJcE1f3drvvk5dtxB6SnnipwyDa4fNG9
FSmd6e2AvQtKZX8Dxdo4zzf86nZx5csfBnvzANrBUy9ji8kTYc8DFjjxiLBkrArXhvSFVlUtR/r5
yM2y9ay9W46ctUb/P3zexNNIcEN64lGIza9voCs+y6MNw3qUUrvUxYK05QHLSY/mRybYIESoiBpo
DOBk3CvZQsqrZsFp09BfAmDVKNnnPaikTQMS7vN4CIiQoFbbYx9mBgdfEN+tKYN5OGQOruY9/2ED
M6vlovLJHHqs8k6x/pzI7EcYqG6+M3vMmrf2roleFAg5hQ+from/QfshkCrupT2qcv5YNpkkYpqN
j6/nUmXWmVPpckp8Pmu2j9yWVxebIEWDf6aO5Esi7kykMBrRsLhCBK2zAQzvCAA38C3RLf1mObQh
As5Jfvhx0Yy1SuQ0/clpwZnH2ZB3OKExa3lh7kd3aPIy9o0W/SIN+gRZVcz3AZJrxck1GITU1Hxz
4+Prpk9gZAHP/3pHVplGneiNZYN6vsZkE7+StJiBGar7kGpcpRtFLOXzR9TuMQlcT55pnnIgCllv
nWzanVR25aMFqWO4EXftNSvi3PneT9SH/yLWjUFxa5fD0Zlu6eKCwUFB06Q2NafJAq/ZDmf4qclZ
cXlsR3fRblU+wcwo8nG+8cPCB3cMDl7EbYdhW14QdVxIB4xaQHf3zy9pd96uP3OPGmm1e+1uLE6n
CDPtfEpqZPCmBP4VSrfLW7o2xuA4fMi2QfArf/vvQtUgpefV7VAg8uLYxRF5UWr6/58aF1zImHKZ
g9O4CN4q+Y/hf/TMVs1490Fjuu+uOWvsak1IcW+OunyuhaAiJPde4/lyNdIc6IIruXRSHuHoMSfU
uuxqdVeZc+1iQ3EfGutsXFHV66cxBm/Kkyupj0PII9L/rowpsyw8r7eoJAX3VVJW60PZEVG1HgfO
pR2tmboZebIXfGxgDJl4Y3AN+fkDnM2Xn6GkVwIxmcU/6u5B+YF6g8RzC4M7dL5p1i8bYwwd057s
MNLxrEhjvggMT39k3RdqiZ3k4tXIAY5yWJns86Ik6Kw1QNtFZBwumw4bVhrO+vLwujn8MFxy+nQ0
NBRFKKtjV5Cy4HjhfsjNVyRLcbhILtccZGO0CX6qGxp8hc3H0RuE0JW2zn3/hy7pzwLb/EsCe5bL
jfRBTjwMYt90+fneVKGMWTTKCZxemQU9EvQb86rAw3jBDWLidzRtSbkc973gPjUk3dNb3ZEREo+X
VRSnfQj11UJx7GXnfKijSr0Lr4VwkyMP9rDC7d6n3Zfsm4YqSbnqG+eHNmDyFAsIPy9Vp6JuSpk9
AuP0JAv21asr+hAcGER4F+ciCq7Ut4Zdq8Xb6St4FzPFNzbYr2HUHd/Y8I/7z/xwJhKviJ7SUnVf
jq1TL68APF5ZSqO9dFysXP3TWMVnHO6rR/ToNLuP8A2YB6M/E6C7UlxpNlS4sWzFHgY9rK1qZ9iH
Tucs+CQjKka5BZsbb39IGFa61I2YTvJcvL9I3Sr0L1a4ZXN1AOwwhYKOEg26/p7CaPS0RVqC2QJY
Lf0DDopMweNqDbQhCp+pZ6brKl69BkXJsgwNi5FASBlPcR4IrweK6RxNm5SWyswBJQyv5wzUjy7J
0RYR5UEU645qhi5W/5kTC76F59WhBJ16p4AuzqsAfPSCo4G6bEkvaw34khp14W8oYDRVYqC/FL+u
fC/c31kGbr6j/1luCYWc48tVLEGFGgQNZaApAcn/mabEkta20DXZDo9l3+r2nvJP3KtjaPtTJdPh
2PXn6ZMFE2rCnljPaI86Jn6weFL9UmGtv8IWOyo7IVd7yFfVcBt5LJLowWTeWUh6w32fRs/cSqgM
l6H9+QhdktqHjfXONzVNei+COdyFoD+8Jg2Ij6LRnGbgre+LQj3/M7q13jtACZug1Omxl3AHzGhD
nArfd8jOPD+ZhQe5sl9Jy2U41Ge0/SDwrNyrNkUSOYODRkIwdeXB/5A9AeX++htT1LDLDCXblrU1
/9SHkSdRjx1hXi28GSsjWPsVO4zLhDi48PVaGAw7qdRJOYIcqCQWVwOzPZ4CnlC31XWeKT2GRZwK
E9nTTVRfO2o2aQdpS/3ahyWj0oFx0xy4Ll+1IWQrAmYE4Cl2cAST0ZoUzmcmwCyjHhf8EvjoOcqf
2kCt+OqiF3lzKcwKNOTrId/2yGo/bp1nNMBCfmVgpMcdnR167CBEJMv9uib5kwq21RiNF0QJdgzV
AaMOg+2K6yS3MLIDuYGuUW6tjdSZcXtDzG9UBKeaMIaCc1KceBgBLaKjJTPPwXUsrM5cR7KzkNRb
vdqMy5LEudQqC1br2A3CX8Kjd2IBrEo9ef2yqz1f9wLgxNNw9+I5MT+HJXrBJddvlJBdQBKIoqRM
00RHvhTLBS0ceDTjCeLcI16MSEmcxKuE4TXDr0pxC7Z9cgprHnOdZ0WOwNhqPCKy3L51omEiPnhy
gu5g09P1eCAGrcCxNWSF24sHyuoPJ9zerMWeqqfwbfEKNo1WZWvUBp0Ih4IeJQwvOIzjlhzhRsem
mO5HnWVh9sd1wnLUnJR06io7rLtOxmbdWdM/VI82ksOeXFuYEYwvwbIcC63eWvH5zB+CG3mgYaaq
ut0N42U0/9qyx6qjm//JP8LYwSCKAZ7B2E6LwDaAkIvyYmbfUoRDkSMsGxQYQVEbCHifzjxK3mYj
YyZSbYMIZUHKR3tdDH+4b8Y9T3JRMh3esytwxY3SnByQ33MqBeOV/Umc1K8fObCc+MEGYKPsGqSp
GNo27v9342bP0joswP1KRqxnXr7RXP3U5OZtYSfa2XIo4qtBYyIbyaXo2mgnintvZTShNxPsSw0F
4b+jBwwO2L8WqnJ7mnsU1YgPpm2xn/qehZHSadPK0OaB4odsOXoke24np13f2le6jU5O3k7oNL5u
xyYi8xuftfrHa2Iqab2gYMpA2DS9o1OyPyZjLW7pojiw2HG/gqtZGvk4BXfBId+xC6Vj9cir6qhm
bOY13Hi2TAgZi7/JJRMSx0+u9YA8w2C9ghz590iQs6f4j4SEAl5phT5BPu1OFijVQG0G3/HANkVO
JPNfmUIeRLT6swoOvtaXLFbMFvlF2fMRjNQmCx0M5yWjjSe8S8oFb6K0OI9tcUiJWJB+wJl1QxLc
sWffBLUXTVVQvEKQ66HHdadZwpLTTl8ylqlthnjNb28Ov9JYlcTrfvtcVEJJOtXY+4R9gHF2zIup
x4QGQ0oYRqQxD2TRkWuZigBh3TC9ErTQE1cruHvxNeOQs9/4UGc513MhWnQ9MN2wfZ6bK3B1133T
oqE7wJG2h/2tBH8iWAPGZeGiX14wzM10/F91f7P4icS8tykWMFjhHH77A9RpTndplV8K1UEa7jPT
lhg9hWT34kk+WIMxno/9RqSV8ods+UCdZuyilbUs+3oFO593Q4ZtxY42VVCekgYEtgu+IIOaxGUz
+ViU00edMvkP2ySWzY7xSN+ol+oD3sCxNi6cWw7W3DJNxKX+mxm2ZzDiqD58WQo5yNnj+7T11Nip
R4En4Dg7hJqrBQIH79orlP92+b8CwGH5RTKvbZmHDydEqqDRdEsS1qg0aXnb9pzZ2yBA9pjIXlWy
p+ullDf1rm6AeztkZ0hGNWAoX+3bDin1iYD1MUj+UKOeF78gPhIgAXcmipDv4HTneOpUfntEZWmh
k19xiA5uzVWKUif0qUfrZcoXAx9gcdmt2kWjyYZezUDOM/ie3SjaRz6PZCnqiDwA/N7Xi7xYNFep
Ce2lCnBOUbhPsSirYXWI0me57bBck3NNDIx39fJ3qL6igVpC01lPZJVZc1KGWEMqMGRfFBn6EJZj
Cejr4A6N6/mw2ni7WUR6hVTSXLL+k1eK9t+VZWXoqXJdEO88c7UUa5hpjbkISBv51NAiCVHpZVLe
NqZGNgN65GhdQ0sVl6Ih0lh0GTnEP5hdb8t9oz8IfDJGhm/dWCWkhrQIFUmjkMVoLc6W15kcHM59
hGGKaIqWfGLFK+vxJvx4VQTesPwxXc88uHPWie4AmqYt6SMtHo7npFtJ0p0woYAoapXN1Eg1L0Oa
kMOQP/bq13El/+8oPiXTfWuFbt+0xpDdgOkq/YkjqtVDzNTsEIiONg3CAPoEBWjEXBBYKh2NqQN0
nADTU8bO5uDNvj04BAmZlh8jENPTS2orTaUizL1sRPHUUgyb2rj/Kw1r8b6LRtdFPkw0GEsolTKs
XTMRe3CJX2txhLhsvhNIfEgeS/Gm7vtw/beNEnmBsCya6h9c2RvZy2FBf2d2iOWwju4tpzqQpPgP
62sOhzvmcfeDzVvviO6pv8xS/+Io10pAD0RMSqM/JwPMtDtNc997pKhMJh5/MQFWbxa3/XpHiOjr
Qla7LKYNz6KKUGdGUmTT/0kZoExrQV1WxRSlwdUJ2lZrRc+LNBLAf3tFuDcql6l/gEKSXRv5xive
53M4yHCCj4pa6uUEZJWAYwlC4QwxYFfF4yidAm4wwTYtzxd9v7bZUHZtNDy36LxLs1y1IJHgWPtB
OoEYX9WxpAkTqAA+5pBA+03OX3/vrGEfALfVoMagfmPL04z7jq/AAilIbsmTOi+u8Yyh912Op1uW
IACaJOZqP0F0bt+G6FSrRnzDXmjHnjA9x5BQ3z+Xah1O5Y5dceHD75Xbj6Y1o+XV0twSS5jT31L3
7GJL3cF+1AHrX/Dx/uandkuqY2p/QPNCLQZFJfYBscH3BOvnQtXXmPq0oKEDYTZyRzVR3IGSdE+G
gUrjbRPu75SaQVn2ZEYM3mOoSsioI6RMiyeS11Anerd4BVjsXMjBKpFFyV9JWrMO62cq2iq5rFMq
z9WXXitqa/D/oVoNE87IU+YMnGYLl7KTvCnDmOoz2S9NzVMdPXWiHq+CINLEyua3ye8B7UpWOytD
QXZDcIzT8x+NiY1AwZ0hHZIE2/piUa0eaeXEV4FD4KkWpxxLuYtzhxXkztx2zqnOTbhTKXt6gLx3
XoTY6UrgsCCzCzQ7CxyS6lo/XQdArWUsfJY7RYvHmhzYw8Av7tY84IHt7lkBEABdM5T+1DpRtZYZ
UgRljH6qEvHdDGCfzKPbo3P1IxdNePZDkwkkAS8m6lQ/V4b4qslks2npOic4FcOeG44cQL5S2ndx
LJSJYj5/A4iqeEqDCVteawkIUty8BJwjZpHg3DAG0xdt8sh10cWAzz7e9DPZHNV14OoS6SL09vTX
Ui1Ra1xDmyDaNwWwXMAw0/hc8AYCmpCnCCny95Jpp4CO2O7jQ58XXGlbqxGSKwRvbEBkRzHPzfyq
dMyTB1AjjaemjjDPshuFDBe0Tvyuv6hXro6YtWDz12MfZ3pkXJdr3ZWlZd+MS3aJ/q9t2DgclKOQ
Erxq7pvDOEaU1L4jZOORivCqqkKfutDKL67k3DWRLw+ySvAntdujm5QQVfp5k7n/k2FF8F6p7hdC
+fV0sIP+ylkPr+dHyjGMzRN13ygTPs4VCdfgMUejguKgb8tlrWy6pMKSYINBSlaoFCLG2Y2snG/N
XQzS0CCGrODHchEZzZH/TG2bSQMOWflKlrRgcZ8qzg42N90AvVSDzhuXwKIZiGst46YmGo8IdP60
daaje31zVCkBHivUV3aJfxi1/iU3qH7gEGR5mCQiEQqODJAYBejk+/YGO/EI7ADhGJEmhoW6sWlh
fvD/Q99SGI2Qq3hBFGRTbB84Io4gW/Vtvoqd02NfpEvM/eI8235fuzsNtuzzhrquQmujB3uwkQq2
/d9mPyMZWXhtTW2Wqj5rooOMOq4Bs9OOWHZpKMITY9QOb9K1TjC6ydMhcvazdpWW1oZ9UdAb4+oB
Go0SAdL2bDH0cPvh0E0PhUIM75Bvnj5fj83MZjKvbCDAHxVBSvV29cHUznp62Cni2ND1Ggp+OSDd
HDWBJcAu+mDqd7OqZfOtF5SW7Own3VLJh1nbc/BxLKZRpvQkca7JMDOMh0WTCGPfIigNqAx4LgrY
DISyPsRFKJasMhqdGmgu53R+m96LbBllpJj86UOohtFuL+NoH1ExQ3TH65nzKkuzJlJNEbnm2V82
Fn2W/JcaA2kpghGR57NAtWS87R1XRKyeFpwTcdQOUwsnQj6GKePxzUSpkPqlCOVObEhymYgllRMD
BevzZSufMQL3k70Fvr6cEjVmaPxVsIQ21GD5rdOCnM6U+DH00E2zXGVyLhHwxoAnB3jSEraF5FUQ
gq5NKBlWAu0yHRZaaP/lD/IOaUVoyER8MHhwfCdgSasbzunZjpH8GaXYzK2F2OZAZlpZOI5e+5gP
sFLbhyRaP4iCP5yUEyPHS7iueWT5t/tH+NZDwBWAmd2iv/gjstfarst6Ad1hvm48lFJnxiMhJ8GE
3wcEmbQI8iBaqNcJec3OWnupCgDMfr3G9sh4kqK2nQ6LuTNrq9XdFQL/gEYiwW4mlQUoUfHjhtbj
AZxWT6gircFujvKRy+IponoN0WhKsdqTkOLiV74jRBmRrzJ0JawRVoy2RjrQjPuobv/Vf3em7XTi
OGxiuNSMySG9uMegCLB0j7n5zHoP+F1q1G7o37HTgsCCCNoJLCz0svS+6d0CSjbdV85DGsIoITua
oi1h6damAaHR1WZ2Pr2V7yII4l6GHRddPB5Ha42hIH4AwKGg84GgfZO1YZ8uVXztuBX6xhp4zgt+
UMU4MMJ20lV2WRxxbJ7iQ2ZkGgBp5zDseBtDtb6Zm8RypZ/VxP6F15A4itn7mAgNlIlpkzTAO0Ct
e6+KWSm40fVjGIfYDYwCkzuO2kSUSzpQ70xALx1NawXRZIdTArK/S1ZihffWDc9bzyleNo/hLtFn
ij6phSb5fJr233alc2JzQA2IxvU3eArIuVdd//V+A/OtWLVT3Hem83voXfqS896aO4Oz0eOzBmmp
kCkMn8mRE0Y/iMVjis1i6hMzr1BMs+asD8Lq0IB+OpZWWZHaIlezUdTpwIpSwK28yFc+SVRzdE5G
Auo6VwMtZurLmdy0NlhGgd5gq5mmgJMV+pcNOr61mThl+/QlUgVwXkmKq/djmSLjSrBgv9g/0ooD
1V6dqCWNzF38ECc4Why6en9fl125byUHSq9aor4y3yIcf93t9EUyZkjgKe/7DJnPTpNmNYDpCfdl
ZE3dK1UESqFF+jPkOwvAy3NN09e5MH0nHPYwhujiT6d5iH8jCV3zla7FmcVLVuT4pAM16Obtv/FV
d21uWYYLmALYVZRIykKMOcA+3Cd88DQS44o9r9d6F0pp7nnDRRA2LMUdfA1xLBAC9sbv9f/WnvIC
xup0g98l8Q+cZNSM/PYY8CDTQ3Fibak7Lv0ax+XtqQMtW63FKC5GKlA+iDCxjhsJYCCHo2rOQ/3c
s/hJgMugARU3U8ZIx0SnAXP7CyvL8sVIKcDuIN+3IG9AvtfGqbxmP/Ie2Ect/LX9rF93K34SD1X5
OtY0BbUFPgimVGWSMpSvBYgKw7yU4VCi16hSfB1lF+AdGpVyWAi6DHaaZaLm4sabd4goKRFeAQIA
Fy/5uOWPVQLAh2K1lY7u6rbsTXXK/oApi5arO7RAPzj50Ft7vrrNMQsmlVUg7JpzK72THK3GLYID
Hfq9dFG1Lm3yi0xzWcNE2YNAg44uW0+6QuK0YYadrmgaivF6IYgil0fTOADsKDUiwVSvQXlNbl/k
PBTcxjy7+9X/vM0UAO0iDVKY15HFcmW27mjcSp5rc2x7cjSpYLSc3ibr1OwKfI93ZIiLofeer16d
NjYT/cPRILQZ8gwylL/EpNGWF7HrKObTlnBcJn4yxOvuQCB6+VJZ7SeUkFubobs6Zy+n952ULgVh
5BWq6OO7GVzhCHf5rscW0U/09+JSGRm/FJ32GS6x6QGjSM6RPDALggQrE/c3icXZukzOvWd2puo4
bslPayTfzOePd7qU3d/m890rd02kIKgVNWvKPuEgjjhrcVE+aLF5/vab7TAnsIxxo30rF/1h0rFW
39iULDjBB/HC8JHfm3vOnilwd7iWGnswhSz/csM9MB14rd4GtzScMaEX9roAHThUoNmyk4NpJmpJ
JdRG4s4lyo4EwYodVofVVRTiFm+gubbnuzjDRieKz1mqWa+4aPuz8NoeRXPrh9p+0EcYc7dAt2NM
aaNV+pL/9UHBB66+kxZn6IdgfgdTOIfXwTw/7+PLbv96krqd6z88pul84GUt11ekWy8oLqMK0uDO
I5TUUJ6EYRzlKwvYgSlc3BNIilxAwPsrOTADL1tkvC11W0Yk5mKAaRJXjDDamwS1pNPT0PLBglok
tzFEdDe0+FQpB5rTXnVG61pxaLfXcQQ3qbDfkkrFQTeegqdNrxjYr1ytLgBfo6vyBwDXzREoLN43
58K4+MxWKKN1ACVWco6wa+dlKzMtm8szXb1L61kIziqfRrsD6Sx/OIESYa6JeCbwtz7hY3tRcvzG
m4kfHaEnETYI7vmak7fUyd8TH+ExhncZUypzCjnXf18hFTAopJKBpw3yeHPmRAa4xY5SvPBQM116
Ce9BIZixKWVECAgvAH2KN3zOtquc/kyAYbWX/hK2YXY0vuBoTsUK/Z1JcrsmugxLxxyH2nDctizP
Ggbf0fC4/rISOwoBsjuHLAL2FQVluiC4rjUh03VwUMF9qOvUW3Z99Cz709f1SXmYDb6vNPr5cWBn
Iilz1QGq721+vJpPKjeQ6DAWRx64vpvwM1hcNl7e82BRl5Fk9gNmPWX9+7Oz1iq/t16BcfYFP2qH
Zv4X3uSsQb+RY0JDQclVgOrH8kzuAKQeazc3NrCXL7dZiHH6BtzSD4Fqnbxvy5ZLpHBKGd0feBPw
rd07eFedKyuevDDnYpv1hNk13YqHuwc3LlgnOh8lr9hyDOBtikD73efo+wai8K+j07+nStxoVyVQ
gxxBegaWyEFxQJFnitBz2u92NA4f96GMgQd5aFrECe/bEipjb/mxineMtb3oglD+sTRgAeZCE1wq
PLl9M7qNeRDk+m1YZWpuHL5uy8L9OCVKVv8+OOx+tl9y7/O601JShH/CDStyw2SX/4dOlXzyxuAe
nZgzdmRUiiIbvikQCHWmUXOsnUImSOPSgb9kns2ykzncPaJWqirYR/qPAPQppLuP0HrX8COldCS9
O5yxkmDw9hResVw/5jJvG3RQjX/+Q0HmUxMXOLO3Sen4ypC1CW6MjLQwS7WaC4Wbh7/bpRwrFWjL
srOmGJHBrk2ihzIEOi6mTMIrzjg9hNTZnQomWaHTN2UUQhktFs34zfsmb1IUxGd3WpQtcYiq2tqm
9uiDQ4G4ptAU9u67tAy2ECb1VySJy9HVWNJzLgVznfdmPM/4eowwj/8VsgJUE2/KprEoIddXfh0p
XUHnrtuUcJxCfzvYQUtobHSQwLuT2VAdcG0potMYmM7uBHPpdV3AeqKXb87evDrmiJb7TkwjHfDk
bnZvjZlDVDuq5/EqUOWKfaGR1yJEirKFlSyJmD+uNzpZiMLNmqqc5oL1A6qCvdRhPunDg8pvxzJi
mbw3slpaGqFxvfbHg9v66iM23zS/e4NaWZLlAFECaBXA/uddvJOiIXKn9RxWRuumWeWgw5lrDMLr
qfofrKxE3aF3YEDPEyN/hgh2JR2ig+vatWRBXUn5PNwR1Ct6O/jPhSfxPs2eIpcNV8iZ5PBAM+vu
qLy9hMPsGYadGkz+xriawiBUd64Q5+9J4RiKEp583PkR5kQA/I+YlXNhm0ae/9yiwcmA+W9+lLG7
QDyNuWGUDSvE59LyYwNPRuIepI0h7eNiAcTAT6jGtF6/YW5zZ/y0xTVokiu54eSBPLvjZ9zWV+yH
WUK4ZxWNtdHWkWN87gVuWenf8tU+0orsaGS2eCmbZoyJYW/tftXG+4Eh7QdmrzM+Ix4y+S6WOGTP
QHpz4lMNDNho2g/fY9jonkUv3wye6oQKMCIBI7pGSluHdTBcSeCdI7vcuIfRDckma1U36js1Y/i8
cwfMVjwC+4yEdgOQz+AYlFeaM4R4/kA1KJ6XcLUlO+0iRDMbmGsETkm+ujuQBaTtXwJ5RTPQd0Z1
K9FPDp9pHI6IxknTDWKIU3paNDdNgZp1peHB2kO3mUD0I/khXm3/BH5syUO1WbzuykiTf8pMmAVA
AzpqTX1JNO8ORpcQYnah2tQzJxPUyrDpo41T89Om4SWMA+OfV13jkwxagRBvKiUgK02hu91HGFxX
283XXugFpvFZl4EtslJvwA==
`protect end_protected
