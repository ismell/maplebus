`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i0Fk3zlG2MLpFA6wmhrHKvpEh+UGFi0qpKrewi0I6VnM8fliwhvc+jFFiPDtgDZrX1WYIC//KOOh
LGuAyzGOnA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gR1SN7ZmUiYRGxhxiCD4ajjfhcHvE01tgwv0wEO4nMeu4hL848O5WRWVQAMdMozlrQHaIddX9F1v
byOa1vNDGlXfWPiwr/s0QM49gIwEIIpHZlVqlXJDYFDAQFVGsIMV1O6D4TJ3h2c8kRjA9UfSJ8M3
AuDf4P4RkUXcUnh6c+E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eutnMwyDKvwIwEaRRIw4vS04xAz2EMQVqtQleIIGWWWAUENynKx1yxg4i+fwH/mReKAuubaIaIU5
y7tDr0T+u3qexJvw7pywADxxJ1oS4yr8kF5RH/e2hg7cp8JyxbYh+vcBLlRTyRFn9RO81PhEZgoA
J9NCmcHiUUrs4Md5wvcTBmJDHCubp7zX9V+XII3Mi9XOB+K6xJMPzjK3SugzjIxI4OaOmslN5CtV
/g+TB56Om8I11LzPOhQF5XK0Lys0fcvX3/L0/xaZLqVzUjEa6FnLVr1QQuCAxrcaDLrpixfXTMBH
2h37BNpm69Mq1TER04faARkg5BCdQv50mEh9+w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
esMv6rifp9c2aOjbm9f+WqIZgGfuFCl3XipiqPu+KbPiE2PmSJihqGwtZyHLy0ToXQM1nQCI1sDJ
vxhLEooWpUnVzDu6MR3/l1nGeCSwfTiCvgTJulzAqJa+b4pwPhF6rJEcT0GscvLnFgud7x3kuiQL
NNUve1c1FOfvX66HWXM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WzZfrW6AWNlUypD4nDmkdSlW0vKsnJHRe72r5ehivRzTism4wWlP8CeubzlQwm3BYT7y1tv6NmQ2
/2zQv/IcIDAot9KTzuum6+ri156+MxY++e33YYwgSy1H9wZIgd9BG88qcABSYDxfX4Qaz7GrHqJX
RyqgCRcKVL9qn32cv1JUkMLax2AlO5I5es1hE0yzF0ciE/Lh93D09JYfpMKffpezurExgNkevmCV
R5BSOJhH+DXAS0d8V3XoT5LTsCbkgaQ+vTCnbJ/4x8Yy0r8IZArZzwey3Oj+1d7a009O7u5J1jrx
hdK/aC1MR1MCxmC3VWTkp7YLpNrE//pH65P/kA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7056)
`protect data_block
BtJf7s4rhC7I3ERsD+YKEViX8yR58uJPGiNj0Y2ykx56ikrwIFwx9HIjoCGbz6hXFjXZkG0hB/3L
tdvZApJfKnmww4hozQiNuSSf37Qjj+TJmEstp3DMJ5fm4pveJnfOugKFK3+vAlPC9R23MYYYEzCS
6u2DwM/tS4ASonRd+20eiq49v0T4surxs47UCiLitv1B1rn5fvem2N5WXsUuaNphLINLAsum09fe
7ZOuMHGywosYi9OnTqmjWYxmNuth1dajNRCRm962S2/sr7CXz4M2cJ+HQxqdhSXod+/SzVT8cyO3
gj4JeI6fHlAd6fXrw8SzS1njtRLYKQYNtl9aqUkaP6aHBoP4ltPiyfufRzYsSCb2UjcNuaArO2ig
7rwPj3ePPW4C/Rsc7UjI3im7m1OecGWTNDyd7sPcssVSHcLipgzRSz2ZCk4MK+xzvdRJdtKpZ6t1
qDOvwCzmGV3JyeZpsLePVVeVyCLlXLlUOWA+3iQ7KN28YXGg8SQwqrw/ojPCF4k6WO/BWMXfwo/s
xB+TKDJEBe7XQzeCTum8X3fRpNalei8hiaA274JQxTiK9HfRtBwq7344ODs+v21bBoRmWUD2IIIy
0EuKUxMEkEAwkT0uhDEr1Ol8RpvLZ5Wbek1gN85UGHEvxxrFYlUF9KRFYmUxEHWjFM8PiGTZWamM
vpqdVZ96vRz+rzuU4UuQ0/PGG8FEV/KvlCrSrybZNMEcPNnKIjuUS/gCVRiSpVCL8ukdPs21BgHN
nkArACJorCpL3O4PrvIM5U/JeBFaHN6K6aFG5L5NG2hXn06A1Kzbg8RnpiIdSbP8bfBKz5DwhUUe
F0BG501vMYieTh6LHT8tE0r8Y5diHzWJSw05ILPKuYpPvkSSLMMFa1zvIhXapShhXKm6nthZ6MGD
m3M8aFLkxIBgdPPkaVZxxSMcrWMGG4gyYQxCNFzwbi12fINYp22n6FdqJEQKFSPk706RpfYHwZz3
vFzjYNLDU0Ry2yf16uVR++LkpP2kvFRvZVoClRh8HJx2h03eRK3muPzFIoAG72KlnCgRuBjJNLrb
bh20xebp8qg6CUOAtmq291OD5ahSZlcVzx9Pf4ZBBOsxguE3Ksiwu7FzfxzyI5Kbjrzrbr9AHlSv
Cpufz4Lun2nW6n3Ryz3Pjz2/Gq30ULDLQE2MopW0r7dqa2Wjs7ISmc/AcMJNZtBBhPSqvw0b0Q5l
QauJ5T5bP35YHVO2NBfkO5IjB2+TubR8RNB/lUsqrLs2e09/qZ639yCLmB+Az1A63IUM86VMx8CN
Jn/bc1343ZldoIf9A2oKbmboeEHMs48HBEfADE4Wp8Jj0YE+GfE58ZYRY0wyNIPf52q8Y9dOlqYD
BoOV6aTh7DTbA0mJvT+G/HwoGDT9UWViZU7bERoMhbB6uX/r99dE4PUR6bOMqhGUIRplQHMqFPBs
BKsuWXt2doDaXQGRxsSeyrLzShIWCIgORz32K+JPkdnFwl3d5IKGflj4b3R9MG6ptpULWEygRbZo
aR0dqcxJoHPEaRxCArF/RypbeXaKi0SAG9PPJs0Mg0dj9BxDLDitbqe3ZK9iYDS6IIYFbjm1Q0+v
+UfaVc4h+VPEyZf5uLHgOKUYHhoUDox8eombSLs2+NhWQZcdOjYp5Vy5vLwrrLQCz0Z3vNrGiRks
W9+sgkUVcUo1kl62w97C9ob25bhz4mstf1lms4ubq8cr3N/6vjhomp35OhLeaJaCZnDXxz8CyQVU
bvHfpF3rFbU7oGTrO3E1hbbslDRZmbN1S3wgmyMj9Do4eBuj7YVySC88uIvtw84Dj11N1GoElBAy
C9JW5muDVNvszhYY0w4c7txpn+PciwDDfAo1LYW8Bm6mAsuZMvvTtGpE73QueGaR67DJ5gKvjozW
DB6RRGIV4lDtsbVanlP19Gpwl3MvIH1veC32hebqWCFHYzHBdVQwkz21SKgDwmPEYMCJL8OA56Pm
JVvbrtZUhkiPAj9dPqDPM7tCa75HNtUk7/lZrQ6PTKs4URp02RIr6+AxTPbmxiwX6xoQcgzqTm2p
HkMNNiBlqbqSCu0/tYdfTC4192YsRUFkAyxeufrnNVX1T82Na3QarD/U+wiZjHN23djcqUAGb2w4
tj/ezF6Xevhr+Si+8QN9zpr697GKpzR9O8MNgUkVlZoYwBcLAGNPPU/QKYH5brCThcA+vOVMpTCm
bMkQ9i3wiKyj1onOSQEVCDnY+JaDRzjxTHVeDx56xT8IAY1L2JcT/0KpOIbR1MbXBlhZVpMM7MNA
Yl9KIzkVu4KpG/w4Z98AuPeyE47SsRlPF+nuO4UeIz86L5Kdovjc0iVTxnyr4liEg/Goxi9yPXep
5ywMXgcu9yk64ssE8IQKm4WxNCdH1rvlZMOANU/9VRZyVWDshJJmkRPi6PQ1jDYUvPdcNlwwgzyy
P4iZcqy1oAvXRGp8rRgWwpDZIs/wfFem+Y2ho5lZVGQ/6NcO/S5aEI4Wu0+SYVKOuOSHMKUb1SNr
BvN+F3aeCNf2XxF4uZz+Soc5U7uVcQxModxj4swuE7mfP4dByIHtcaxXvIz95cWYoUgpiwowASd0
ZEIkJMDKUwmXUjCDcLFroIhmxs5ky22nQOxJd/6g4wRMLtoQfYKCpvaOP6gTkRu5B/QLON9MIuRj
byjeUk+Nt1t9Uk4sTdN00T6kSTdLxHcGoXkG+QheE+/3554dp1gegXBLLK7vK9Q8ftLdtpTK5+i+
mMlml6LSDyTmue4PmBN4DCRYTvxy4P+RoEigym+8F8KSBXjxkTNtxM1eRFjUoQ8H88NsKQmpdQNM
81j/ccmT5jK+ZImndx7jnpBVFLS16qrLbzVb/BPcUgxJpD9b65wHubJBrqR1Ozgj+oE4x2tbChOC
G9zL48OiIAmfpOxMoUMVzu/z/7x1RVG2HFqgrd9trAI4CqH5BK+NIbKcgOp/Zq/VAsNv5cuwwCQu
oFH5/4QpHwSFLM8V1psYn5+IiDunia2OHn4tJFSE5UlJgmJjkcj/l2yaVL9vlpPs4Zpt+6RdlAP9
0NLIoXuEkGwyZbMlvWOYdMMKEmD4WXh/PLiu1jtxVr269R+8VJyKoWHKmvGxTtAPqCcxmg6CkYS+
07DMkQNXe42/HbARdVMPJlzWPI2gMJJrWbZ24sF5UG1Cx7Z9cxjk9pWatdFfLiHv6sR7dt2Q83sP
wjuFuGWSWZEmFujk0IaB+4KGRUxnFzmGddJBgYxOFBhRfFO2fZ0CjwmUfZjQkfPtFS59NEQHre9Q
fjhbZJFTx2DaKuVeJ/A5eN2PlWhlLZqbUzjiAsqRdYqiU5cIKuA03YfQdc4SPh6bsCByjP1/8wxO
ggoczDoH/L2Xruq5zKW8yGX7Lp7epcSFYiCARAtskdPUyUzFLZYxXNvfJYnnNNrQ5/c3ucU2d4MP
98Azyx8XyB5WQ40EZ+VhlqA3m9Zxr9JG7wZWJtCkmxgq8ajA+rxwsKlNshIdKmrjdrIh8BidYwX0
eETQEEK0WqT+FgegzZ14nBFwGgY/d4F3XPhjnN9smU9ESa+Izk4NfX9rJC7jVLPe6GUZjZDeJZZ0
YP3bpjLEaWzzwnyJfV8ECwE09VXpxiEBKVJxezr9m3ohVitBdqw9SaA/mG53i9Oa4TklgGCx0Jhs
Kk+fUZC0kIZ3P+mMiDMxi/3fWw+WtzDp2QfaHlQzjmmL/teyqtAqg6BC93skhw2QJnOHrMkW9iTr
qodjJDApYo/MSjumLMnqWiO+7bQlHSH5in9tbtMMgbkEUWM6gpUHa6ywqAMU7tgzVf12d7IdOHGq
TkVN0Hf1klqRkoeQfY6QDjM/9YKiyzGP/4K8PH1DFCTRXGZVlfnX99wDxv3C0ys5RRbj56isgD1s
ju7WQO9DvzGjcJFmoPDZxommZmok+83Z3A+UXJy6N+OEjRFbWKls9DsNl74LzK+X43VKTtFw380x
jzVBhriozKz6dhkhu495TNI5yALKaP72QcjN5WdEhjzvtzk/iiGpXRPSzU/mwHXfCRoS8skvcprB
IGWRSB/jEDm4MEMI3ziPOrG5Lxb4IRO+3iSP+Sc6Tq43ug9muUy41TkhxIqRReIa3O0GaIizVri6
7dKXzUjjlAfZDVytAt+r9KFUoGVKUzoBXoltGukfALkrI+rjpELllhDjMv3tvLfG9QMM+D71bo9Z
wK0uuOmEE1k3AUMfHHsxXXF16iZeUW7GhuGQULcHDIlW08fFkmVrjHElnPFsef3LbxL13u8zUidv
xI10p+x14i9fGKWf2AggSxDM+t+3hrCNLr4h9gvD/ovJyBZzsWb2MSk14igQu8Y9UMHu+2X00KIK
3hLM0oAn6XQwE8iqITfSkqONT3OHHYUmOoGonGJHz0DCBCqDlHQpOZoZ0P+APKeb/T3tSnLKANkO
hXl9NGogj8gzgzdBK41rCt33izTj3/XIM+fk7F/HyxnZK19hb4l2wvL9AP1y3p+5cPh6G9cB94Lt
Jl9Z9KtNudTQc1A2L7HRCwwg1NNlmAQaDJ4wZuw8NdITHu12Wy4FgYC8FZTjDcEixtzCSr0/4xNP
r/nTtQPsqK91PxSBLYnKOzsIv8SIxyw4iKOiNAdzGpE14MrQaV/lqziTHBMP/InX3CGtskvH8Ifa
97jKFRHE13yn9uqKKeks+6UW9EkepN2tmpsLdIlvnfM1S9IkhcieVmN18vo1i87qOmHL5udU9ATr
Mv9buZ9xNHsjjFrf09js+4H32E4dmpR+eWdzDpvYRftIfCfJoU6wwM7YjYZZFNuxJt8aChF/TQqq
1/LvIfBS1cZikDTCKlBQ+kANjui4Qn5pC8lCLmMn3jZ0ZbI+o7gtmebBPU8wEVJWpEYAxwIl5OBB
tFAMt/mPxhKqTga1qLL4ipcaihyvNSnmHF3AA6W9ahZbvJSnlv1hu/ma3mJa5KL8oWswFJcC8afQ
DO51A//yb2dGnEVIutrYxDincz92ANfHEetAjZtdy7Av2IBfYlPR5BvbG3OsdcvzBYS9CwsnEtyT
vWF8FIRPYvcphTtWuNcVPnjee31X9cplhzc+mY2jXHxhgmdx615yKG0lHdGly7wO0zTQ/GGKwd+s
xI4RXTu+chK3M69CPXA9ZtScL+P6ANPbeZN/C4rXAr0Oh8LDT0lUCiFk8HDIkUSIPKUbFKjcEFPH
oeKZVdQasFCYoZrlgLXNKhhRl9Bty2/Pc3aXsYZwa1w3O0qnQOxbBZrrmuCOW4J7SOTWrM2OPm4z
FzF729bkJcrhWAvfV4zcxlTB2X/V8XHbx0zzqtASnCPLFpVJ50DvcItBZBFcaiKHOxwX9dJbJ8Kj
TXfl3ZdwFsRfx/gokIq1uvAz9HKqXlvSFdhXb84wYnspviCHZ8K66Ax1jYNkZwUeBJzZ+gO9dKD8
a03uUeT3vduFhCrIkVWt0/jE+wp56jEVbqmSEtLSL5lPPkmgPedDDa5xmIP9yLNwO26zi9Nvg4Xk
EIKbc7tWF2Gg7/+CgaHxY/ONugH2dzxgbkwhoIkh4biCOtyD9UQKAwRivPfxdgdciGSzhVheQ4ZR
nahUZhRLwz47yh5giREdALZOt7DZSyCtFlOZuRhfXO9a12KW7UVAIbooeCxlEmIZjaWofiWLG/mo
QH/1A4Eww/6TlEfwHOIeTjqDnr2ASQ/tB3VlVhDoNr7dIGPeB+pC8jgVA1Rur+TiUvtqb+jNcdi+
5PooBBzSmMkY3k+3fGvPPAnGqYv5LOr2RMb1Cx/q+zDPDybHgnziNXOMApkfNxGH371rdDZ3IuKP
qE7+VY/+ECiFGoS2Q7htbZNKOK3i+kdjwHc/+StuKlXZJmoQaFnYTzkM7MtikegGfzieYVz018Uc
BAkzLCHpLOH4cQIQqWE/ncd7PtcRyMyi0M/8n4XblO6464hAJF7jEfR4yENNM9eOAuk6gvBweL3V
5FLyrQ6XJcbFg1qX7dOj6AJDfoWrBM89cZ5zWamaJwIpGN7vvqXYYZf+RTSNNjSN3u/rjTtakk4x
Sm8kwjpAajVnWxas4Aa/DUI3aPVKZrgfetCwX9cGDljIA6t1aLeMz/x2IJ63tONEKqignkKU+NYh
hJuu62eOJCcQxeH3Lu/JXNH9uFIrrK4AgP1YYnU7PgIIGTF8Yn5mgiscMTRKxWBX7zZdw7q7+xq0
cgl8PI4qXJT6PWrmp1g60RywzKPm75vyuvRULoDb2gS8mrODLWU2+jaSxNHVRUZ25vXWUlZJBnSa
1wifRaCtj/XYHAvDHX0M9BzumgMV0lwtO0akSZwtpMALZKRyvdmKp7SxCnvr74OscgAPn25tdu9C
z2MRrDyslZKEcee5tLqcYJDYvYchfHLWMjrMnsQBGAJIwKsapQi4SENEf59+rXALOo2Bx2oZmeP0
+jS2WGxy7JTA+a3GTiO5trv0l2gB4o7Hhc/uYlXMXtT2YIrnmnSYCWs2CQam5QAGL1jfqtDFo0hf
uDmbJLxUIZ3Jx0cKc3CeWyX51nBRfANM2x/CepoCWKL34iUdcmDZVzrM5q6RFMocDbjE0Vs7hTNW
vYp/H8jrYaxEEqCaSIkl7IOaMiOupXnDR2r3HAISYiBvD5CooTwgPEAS/cD95ojHbNQJQu0jud0+
SoGWDa9zpsGI8A18FgKj5l4d9M8A3Wv2DMwFtMoSBBvxeAokLxrea/vspnJldN79tCtYyFwic7ay
zdbzBOjH+rPfa+Jp4Ske4kqb3ubMUW5BNrWsSMq+qypIasoGngyXiZFkgEMRm11YOjflS219+mJf
b6swlO6qw3sCBeO8VCYetKCgqwqUx4xTmMlfqmcFsGuhu696sDnzK+o84koDNpehlNuoMPTtofeN
RV45jS8zRLN99GwtiPANeQzyvxOhE5uPh/gh0Vd35McqpvQvBhV19Shrn6ZGMWPlfPgfgPudEe64
PFINngj70vj8dlzSJ2sCTagKs3tZJyJA+qkyY9qDpx30rKhaLTJCD5D1Ua/7CRyHv1Xa6OG9GxPy
Jisv/VOyxvTHuiA9xuzW6MxXltxP/lD1kbcI13dTqH4bNusV0uuJILGZqASSH3i7eR0bjfDnE4+K
zjaLSMLnwy2epDwV2+7cU067RN4U0x2MocAuusgKgkO30SszI9ljI06C+PtTx4aa7vB1n0lzNnJL
fwZr0Irsb6InFskooYzOeWAukhFu2piOD3Gc7JZoCHL6KhgRUDf100w+kyjZoTKE8LaLs7DH0AIj
fjk2qDWrWZGcVkIKFksR4r6gua3LWSDBzzzA+QuBUIMqoWoc+nTYMdAM8vSm1rq75gGFRCNXjRYX
nDzYmZFJ0d0sGHpfx8b28ZI1MsnJ6nGBeKz2S8sqATGN7EGdOOIQihBk/rEw2XGUJtHKc+1cQEVT
FrCBomamMdnlxC8tnsYn6x7ATrXMeQ8grjiCnDN8Z5FDUdaxHxGEoIXyWhcZF+pjyG1r2e8FRj57
EDZDa4x/MyVvta+aqUKfUwKYtoXjmUscRGf99YIi34K2gxFlP6Gg/JYmVlK1+46ry1iXoMADyhqZ
UK/Z3wNmiZtA9FcWKSrF8h36JkBYaffje0qm4E38gfTPfUKn0mDYGU5b41Wdzeo8fh2wbZ5nZY52
mVxif16i7NOa8vXj/6zi8ZCdBCEj+/YPMQC8dIqTPOLTTp/YGE4SgA0gQHlMmw+nRZKra1UyroDQ
f3hY4Wdbpcn9AGSNIKKJ/crUY67X6lon+Fi6Rg+tl33pJlcBLUg5RICY2Hgj+VjO3TYY4KsN9259
HrfocNI9sBF3o77B6ETlBsXvZz5jhZLpmAer4gMqEYbtgw2fIv5wVct/QDdM0X1holUe9NL4BAnI
duPo75hmu7Okp0HYuvYw4za/SDtrAamS3nGV676gHdGJZ49sDVGonjPbC7EwKPem6uMjNiRNaAWg
1Vi/sYy35hqhLYamF3SQIqB5aTXfiM+X/dtiLCKs9jprwhhQEsUACH7mZXB4GKXSNVxXHbfZFP7A
axoBfGV04C4T5oDkehkLE7N1eKRUg9fszkStja026bg3Tijr1eqIEQ1zsAyZieF5fyk4YiWwpqNr
HrgQW1tXGlmQ1g3mpQ4szb9un8s0CH2mZ6ojB43i3IxFP7G7ePAQvbWEHwbPIHI4zBnPMyawFQ7Q
fOOSGXWwbpvAFUYOrNXo0+fEXqx35VZqv80CIxSkHO5dJ2FGk6ohCyk5gsQjm6aMfHsfOLl7LjjJ
pxFqc2zEVlPz9oAAx+rCl4oeKHkhQMNcIGt5JU238+7A+56G6ZHApJUU3uwWioteN9dRL5sP/A1B
ZgaFDT6poWMT/6Mk9inPro6I70R3TqwoA85LazLs8ITsNCcSD/4jkd87W4LI4A0Ii7oncytqYocV
h7PoTcN38Ae771hkQfNJAy575/ZrYsPdoW4OnHkuQeTkIa7v1/xULGrtKEZpzW+6CtA0oxBJ9sfd
8tP4QmPu1jzmKJo8DI/KwzNcKXGGpOZC+C2lTFuOoV3fN/+RtD2H0DpdpkFgO/IMHk9p9F/GIUvM
SMiQPd+zYCpnQtQUkyGXOIMskajkMa/2WC5lY1sdZZ2B82KCBL8Ttz7FkBaYL1+3tOykO5YJHO3A
nK9/2nug1wHj7bG9rMlHfdLXEWzUjT3qrYN1d1SxXo0kwOQ2ftHZS9Sc2sM17CQn+ETg40XBXglq
Wu1OwNOXERYe3BphsaM4t6eKByvE4+iCR2Bo7Ao6fIkyPNZWgBfBINl9hsvdc6BKA+EtvIZ19+M0
kHpurnFDwjAUzG0Dh/RFwl/PfZiaX8z/rlwaJPchGY4we5Ue+t8zdgxe64LWavekb3j3F1K/RrMV
AyK1jwDpL8SwSzU/OiiwYGMYBGovP61iQWXLSlHE/wQXyWYFV/gS6oHhz9noAG0bJspwd3XbEUpO
/FGUB7wWd9REko5AiGem0tr55lBH2w3+FAMuK5Y4c5WhzzbQ0MjZH8VjO7BHWDx80XbiDsM7QCTY
czuhBpWwNJq7ocLWqzq7jLiN7Sa+UqXb2hB4SQ8e6BFlkcJcxLOPi1royKv1dFcxoOhnRMISn1iB
tsyRpVU6XgTwVrt8ylohBVAmrsloErE8pKu2iUoA6KSz/vOTuBvm9nxsx/r1bxaW36jnbq29Z2Dy
pu+WU054h48or5YXL8u2KeyCqmQkR5xa7IsYLZD8GPoBLLHRlrs7VdNxTGcO5Yc827X0e9tMhJKe
g4QYnN6uaQKwoaotrRyVPRMSz27XRGbPlx9EbiSeDuev/QjPej9DSP8vridCLz1oswHwkZZJdY6y
nfYchqSoXqYlTdbDacux9ENlN2ueyTpBkLS2n/2iIbj9tWy23158RNiuSKBGOdV0xB3+jxRlrpqX
O0gUa2YOJQYLjE36pj3PsSoXmcu5BVXmgtGetiRdndbBW0b/f5RKr+lPFY2Y
`protect end_protected
