`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WjFxRci1wyJltN+N7KF5bUTxa3fUEk1KgggcUGhS/jvCTgYc3h+1Mur1VM5UHug5shjI/9Jstyn7
06WLOEG2ag==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EjtjKcJaN0zYrzSv29bqzb9YZV58+fu8IVCeZxvn8LH7vAAdZv4w3fmaSwVZtJSjY/xhvOjcnq83
bn94R6wsy+KVKeiZqH5HEp5FMqq1RCsSKc/6zpGuu0MzG40ZLOXfpNWXQPKUVEqnJYpSsl2+AXKM
ssJcnXF1WJvc84SEnjo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JD8vFM3HJP5VGcXm+p27FhOtTXbpjhKwYM5Sgie1kW6nnGKMenZlHZcCICzDXfParSRPxijhzhPV
rvDwRFWrRRUPyrwf0cvaveae8AK3uxQHbuwtO9Dr2Kzt7s+E82qkoEvUzGLQydiu2EJnhQsELgkD
4V2ceO3F2vZWq+yI1BXyp1PsDKDdU1DDPrBkPBGE/lDKebzuYqJf3viOvN0LmWNJu3C+PJX6ckE1
DOqiAw/ry+1mp6E0woM2YNc0wEWVcXTpdKRgBthQNCV/ZMC2fqCcm0WT7QZI5GgpzUE/LHihHo+r
heEJXdK00dbsrGeV6BH/6jf+C03bEJQjg1WGow==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GDpWUJqvxrIUtJfwOZuSj/RExwivhLCWlU0BePY1+GiMdEFhNy+YYNJHH2u5JpYuMdw0OA/ALnWs
VgMqiYbUucksPlCSKfZioklE63SpKyh/w6yMbBQsfUj0wt/AtT1ZXO1ZTUx3ZshixYXHClinkegF
7ZtggMbQLEh1kJh7TLc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bwzUeNxrSpyp1eAMa7QGW/KdVyK7zkJRsJ53OyODN3XAlPTApsm4pI+e+n1ZSJzR++oHih4kXMlf
/5fKNZaPBn3jt6MpSx+CDm5KhFZHsfnjBEU6PRJCCfCHz7s9xEZ/9I0wxa1Dm97GieeUh5V3MLcA
a/FEAsCvD7RNXoy0Xc3rNhFHpwOAw50pRksqLSwze+9HL7dcPiVx+3G7u1pD9nrB+JbNm/Npx7Qs
PkwLjZjQAdQXTzAIRdxdIq3DqLiEdCK4QdAdEcbJG51ogZCSF2JuA/qy0c0TURfn3eYrpqL3me1c
HWCT3wy4empHUWAxXJ7eVxbka21guszGt83yhA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11232)
`protect data_block
CIk3fufIKXSTK2PtPfXvI5A2rC+KMhtfCnjguV6Iuljo7x1JqILK6IgJCwHE+qrw4VFLXAa6nLod
tgIVugPaX15Tz+KksVsKwTQk/e2S3knYs6efDPIFDkB3AqRLUcyDKl1NGfvrCLkeYeuPD/YA/tTN
K2o7lYJCrr8HrdxuQUIWbUjHGJe+QC8yEvLkNRklpMj/lcCpbJwo0kADimKcBdql0cdrohaGsf2k
FvDIYH4EFAr/s2Y7/J5DkCb51o14rhdYG9MJY/5oAACw6Vt0cmwp2H7SV9GZkmtPv0+2DSH5r5Vu
pdo1aohv67VGBSl4rgeBZaZQ0EGd3K29tcd7D9/ZbZjr1wlGjRSDI6BE5Ml6GopRJIg+fJR08Saa
Np/3GRZOTOsex89eoR6POFmaaAB0kntFM6ioXxffyuvn7l5lZzlChKHJq91SZO+O04w9W2U8z5TX
USf+yje5IVlmNvYAi02qw6LLcgJ0wQLs3qDmmt2JIL7sGGNh8AYE9gVdvDhPKmmqwhhh6CdvLhlw
yUfXTX1PHz9DAVuK6IsCHe6/jRu5/5kdlmpFe/wNN1Qb5KDXTbpJ7CeeS1GPkxxxFL2Ct/msP86C
Q6BmqhYOfz/QTTqSplH/HY783S8eVJw3OzqPc+Pms/7+lLwJ7lQEj/IpZE/vQ1kiOVC0iNhHZGKW
GS/rlwivYFEQuCiuxJj83kdXyeCdBzDLuZiE+hln4ETZ9OgWpXJVIBVTy4ecKA+rX643FPgZEQ4H
0UbXEkbXOTjxdrZgHiTqByLBzXUC99M4BmypOD65PyImPex7J8CNeE+Ciil4LWpWjlPwTJKdkyaQ
okm9irrttmabdcrKcPjSKd+eLvGkj+ZGzSig3MbACW5yw0sG4yc6mfXeFfYQhx79Mh7bTIawq1Pl
66fyXNLfw3RKZBsDjQ8k9sF74xcVjqYCUOQOsX7VqKM4PJoIVLDROxuGLOhwu2gs/v40mhRSpEW9
qmmD4tHHFSmJSCWulm5gJoREH3XuGaZMUkOmtP91Y5rgj+1GWd6d7VDXicPypvQ5PGuBktTzbLQ6
aiyV3KCED0mDHf5K5nsIYoyAxRTlhrzOgYU74/pKVg+etVQwBbnxJmiUZHu6lBJr/HCkVM+HjXVH
UPzFQSxIhNUR6JjljI79/6B/oKDz3+Z5s+T9WNWQ0j9V6rXeKBWNE3xHf6xdgtkzNDXk8j7vSF5m
KmmblCqiN8/F+dE6fkadewxGTM82syvNmfYDTa+9lTU3UNAKBzu9pBpZxwJGOArRF69Wx1rpsVkK
yBdc1LQ1X8ClELL4ymi8ZGSkjRjaeF13aEy7rUbN8Rfqs/KtZ8RRb1cn05bpen2UTOX00Gfpy4vG
RlD1HGFBiVAMHWnGxcBFemsxyndHbdFPI2SWJmX2GvdbwMKp/Z+8CUXrxpd/ZPTUfkcmooRJ6q2E
vqNaoCTqWQwDj7Hv0EhLFiIPMwJ3Dk06UU/CTfEgU2Zw6fK6KdPDEmCN0tqg6+A4Z9WcR2PPdLu/
biZ5133yCRsyL1pYa00FoVUP0PlHqkEN+BB1rGi/2zNmVAjgfIbxSym7asGoOiiEunirdqaRx2WC
i3DmL+ABf3yNyXy6jbXFi1RZ8ZVeR0PYjTDgbCzsLnWyfbLHY2SDxWiG60fezLp8BtrFDkuZ7/aS
d75AdowNtglzNzlQ3zyeKeISd0ogHCuBv0o4QvmGEmx19RaGYgUa1SlcPd/RqQ6B2ci4Trg+QgEx
XiGxDPtl2v+4u6gPJutQ9KjyK+9lCJ1i17n5aENy/1vGv4Awam2uDtzaSPnttOdbP0BsBedlaySJ
zj/lSDZPIbycuizPJbSHuHczbOhN4vuTns8rHq2lkyCAzLX0yUSACDgVSiq1OnrQM5e3ifYKQXCb
9Mw64ea+R5j3opjlB7MYp4V5eExfC/OqxuvbdhUwLqOoH3lPhT7r6+yeM32IjW7PJrUAn6RO5eLW
H4Yyhi8si7wgOLWCNBclQ5KFOGkMlgnWzrOTp0vYm8l8A5yOSKSLJsc1ShnK/XwuP/DHixqNdAP/
VvNqllpRgfyY1IrsiCuAp3R+o+6QuBP7HbFv4Y0BAFRfYer7XkgbxUBkL6WxD5sCu9SGY/FfcOPf
+ueF39qohBnRhuxExwt/gB+bott6WwOY+IxHCSqiVzroYgCk+9iUUnazhPwQQrdiGEVRdUUxQ3DM
WKX14BPsTSI1ZKoPccIh65WO6/+MFIyQ2L+zoDT9RoY7qSR9O9ysxzwOoUzPerh79usq49VXeqHl
XDLEOAanvuJg/tNj2kujR6H1m07XYaeBsXvOHrrS185EGmVHSJQJgXm4NUCkTLN/1CGdOfpaBLNy
FxgPcxG4VMWhgwf7AKt6X6isSatVWAjp4w0qK2L+GllRr9H1jqPUqXkEIQ5ryoVKffJSnl4tYbNr
J2G9I36fbYd5ASPL1X9JbrYG4xIqX/4TfFYa8qtzfRFZL8Lv/uhxkiOrw9zg4AHkH3j8/YrmfRQ0
kM8MWtkhpN8k54AiSkefomgArPcEUKE1RM+KeJ7EqLXRgnIhpcwXu8ajO0l0XMcWgFCkXeu783h0
8Sr/wBjSVWb7EZVhr/VWMiw6rOj0B7QdHkM/wJTZtLU4DcFjZjPF4NoY0X3QFtLUK1txA9aRHCua
4+1jHuyppKHE8c6JXt4/a/2dvxwn9gp8EIy1O4TQeqxoB9YZ7nQDcjHQtl/9Ssz48Rx4ajZoq7Ea
e4JvlEHQaX3au8p4cdRe4o2nXghdi0lZLwLWsZ13IUoWBdsvZEwW6CpGxl0oQIlW4kGOISQh59g5
udjEr6gSbkc1ig4Tfr9N7suEqvhg4UKo0+DBHjmstR2Qsbcv3lmkCS3QmmOlmFD4wE6aRv5T+Cbt
rqzbihlr7G6E9CskJeUiR/DfFA43/Cl7fPrpLHWXe3q+bPI0cUrbwGv+3k4zu3h5QgclhwvijPME
zU5ShFCH9hyBAKtTJScJaFkYS5qtXNtsd6cVEAfYvFV8Z5XQU4p1PaMV9g0P2USBVrkECxrFvtc3
AAcFTrzF1KYJZjDi1oQ0VWzpwlEl0TKTU8R6xIEe5RJDxATOkAt1omFXxD5eFfd5vcU/DG2ERSax
swCqVTvB5Eeg6MSTxt3/vBzZdWp+HpfWpOf9HYXKzgRNR2e18w3Qlrx6q6Tqsp8LhjK78fbGC0Np
6seyT5kCBadhwwZcpbAncFqW3n7P2slwTvVT32A4HJoA5mhRr6Jjgw3YT7jpbMy04fInysVXQoeb
pzWVs6p0JVn5h30GFiBhukAL+yei5KWOmqfPoLA5FpBJfM8yJoSS33ap18BCC7yL/4yX+zxtQvVz
2ZmM2q2XqZQeWHbxdwA/sq/6pinNidyU2sAvhfe65KvyiY3PAcpWaju7T28XfslEMWZ3hi01fo9m
nBnvGagPKEXk8IBvtaW8bcyhLzyFaEE3oSwawMOPL5pyYx37KkpKXLTzUUVtHTFBHj9K6ALVzQDy
6AALYSGJPG4Z6qjBnW2sTBy5J7oQliRBo08ZXYlLrdO3ERc/NQANAMCiHRusp4fuEGnOEbf7Ixbh
ZBttrn0rv2R1tAhdvWxNiQeFxYxTZ9Yib8tzZDjzHcUhus8KeiM968ECY6+WHjP8QrSO5yA4CrEf
0AsOmf/XzF12Qb/XR7r2PVMbtPrN/Ph8x5ZMkgNFrVTxhc2RsFmpRSSIWsJqh5EjgZV9puJZNTcD
o44LDdAzUOOc1VNX5MiGFIL5hcPKQmgejjyENYq/R92A21kDaPtM2i9FyiAhL7doZX1R94qT40Ni
SAbGizEJGtLOYoQ4GYFp3Vz9rwet424ppYJUzhac+2BU33WkHFwPWdW7Vkq5LOm+0OJVMBG/dMAQ
dnnV/jdyUVo7zFSF8o0w1adxC6ff5vuBCUpBZRSDlxOcTch/L/KwayWZfqyqEtreCrru011u8v/2
uxnRVRHryhjs766GtjRVzcZXTqAjBhXkK6U6QcjChkznhBly9jn1F1T9o9WeUTuHCrDdDKaMyTfE
HcPRtKqaOQpukPQdWUfVsLYDkm5oYkMRsSoV+RzHpSYJIAjo/stC5eBo23K2G6jLmvnwniTsVNxc
A0ebg4oaJASqMHJdcPSGAS9CLajJc1PZR+zo1qoliKpKLcGutIly5Fre3qWDMaxWU6ev+3u5OIN+
mj6r+PDa+13r2kwGxeZcrvsXHuCze4/O0jrjQq+oai2tB3dNVhAFKluL8Jf2Wz1z/pX11nzjFFaf
MCuKKA/0GWqbSj4vT56fVfIApM2WTHOYy/9XQxjemf8tfa+8D5qTm4nmNlzyzVZyLBfV+9RBNSuK
UmeGyEdsdFheC0PHYCcEbGMWLtVS+fB4N7VHv10baDSY/WsJMlJLnFCQkiI8XbFnWVzl0B4XNBtb
Gp0qPx268GtXMQCKGeszc9C0QGhaU5Majy7eKDzhoJ9lQ11FiTplyjbghRlMVt8pUkJZPt2U4feE
rZlh9e5wy82UrzMwF0QDvhmeFgxaykVIsyszQApNz3cgafgY05ARbhVZ34Ww3sB2ypZ05vdKtRrP
khHR+H0SxuFf7OUbORdA+9mgdN9oEGC+tYRE/T2iFsrexnxwmWlH8YRZFS0EvmSYJUMiOY+/R0Nw
DPvKJgYBTgIQ0we4c137KZAvQVCTi6Vh1ut3hgP94KUW2bLJ7VesOJx03JL4CI7zowJKh1jdvQth
RtRflqyecEDzZlPKGPTDOQjl9q9GxBT+nf9CD3Wa1jFQ0YShFxd0sHBrRDX1wLURD/G715xS0XSw
XGwU/J1WmMxtLUaxJp91jyv3ljxmVWu+sJKf6DyQXqgp748ffz/lRdZzzMxhdeDmpsbBgzXzMlS9
J37wBUXornI4KWrCNgm8awveVWZFHSxIq/gtNOkASvLJ7oiSsZ/UQfRN274IZoDAztf0XMmmyPX/
VhuZc6Lr3JYG3kJ5a7mu+wFyV00rFjZJFtcGGy4bb5q5B1ibRudgzOjIxkWGfDSLnQQLvGSzmaPf
iGzLFS2+VwatKw7/Pa/B2MDyIKZ7nakzgVZpYhJBjsIogIhHajArh30g8JyIDPglnHRGSS99cq3c
uBcWtFsgqsG52ZSK5mPhkk9xZSl2rusD8hrJULjFhk2NeWYAjnzJQQ1waHCo1cquPfz9Mzxv2udd
N5+Ome8x6nd/4e4hvzdPfwl6lBDlXsLz/OR2GJS/RIJv6dAkywj7MslvJYOfy4GYvWMZGTmCgPyo
60oNomIWrqL5Vl1+Gv0Ubr4I2/l9UAF6RmxV0rUwG3NapMA/VMlKvPE55taKokio3kzxzt551q58
RS5pcGzOCqG5aCXLf3q8viQLOcQuG2bh9IeZmFwPSAMCQzEk/7+BFAJilMVNaxMhjZVLZwzIeBYs
qNHlg8miaxA0PKqvDJXxk4SbIq6QDo6o+6ErE4I0lsij+qIeXb/KxpWfX6Dce5y/dZ+pPvasfVkI
EPfocjUMlcd0iSp2QrGRGYAAN0N2ieFwNscDzysGanTIdHIahPMdeaRgKFzZzGhTVFdlN/eyINna
R/YQMD3khSlH+Bfwa/7Uw2aoapgyV1GzpYE/mlm+amP5Pq2IDbgli+HDBxZrOHnlqGxgQb7xXwfJ
8TpxkWx0Mqp3fgQ//8ojEsmQ74zwgor/5foSYu5yPyVkwSnmYnQYMKDhCbGUtB6ilY8Hr3oxcQtt
Wd4lFbcDXrwR4GISuUfw0ccEYwjCU5yuhzHpXRhga2pAAIIDzWlluAtc+vhj1ldspUuJp87PqV3Q
GdmUybAT447WHCGnIEF5DIeTnPElGCfDm3t5bwN80nChk/XJEajunPq7sYxdKRA5N2mXAvuHVyh9
p450Inorig7VUOVMO3/NAh+2y+jG7Y5J7oXWkYCHi8tESGOK3bovUV1LwvgHzJO98Rp5SJBO8RdU
9TOr7riCUnKVPg5017rMkPkB0QTgyHZWpa7cmo0f2GU2PTXTn2ZHrDDgRA2RnWBFG0Bc88zn4IlK
V5RLlEsRUOr1Be8zfr3+rIIvbs8HQzHhDM/4ix+AjxcTiqA/B7HgUW7Um/KvGhJc0KeZkr/pyHZ3
uAX8okca9Z/te1UJZTtPPVn5Eh8zMuFz+AET4gTEex2Ckkf3C5U5zthDsgL8xdGVQkscdqqI0rb2
PQ+PT6WWoYAbVyVeY3FRunT2GJTzrtLWNKoukJSPX6l5Zo/WDmKSVfyIDkKBPTWJH7p7nNnTvFDk
C14zRnuMsKryBxAwJG4lvjhhx04CDVoJyYTYcxEim+8GKO+lt+YmSoSaPmGo4JKBqoaBuqP0v1ei
Fk7iRCs3zYMa128UPZCfp9WKrCHm5lloG5x0Py+Xa69CmgGJ9fKxeDgyX2tYyD/PAvCy9nlSvOBn
3I0UCSeEtTg8VDLIRb3QACNzCfm0KR3rHb5FWpD1+R/x2QA66tsuszNn2Z75I47jnKqxCkpQvYi7
ZOI43S9PnRnTgoLSBw5JjvRz+HPAvzkFhwf0K0D+kR01vV+CJzgFt0hU82AOEzQSzjMDQ5PPNeFP
mx/2jYDv7FCL7bktHW4ck6XQB7C2WKmsbdBLHc0vEOIc38kAqoUpZy+uhPIoPrdSTeu9yb2OIKyu
eF0yGa4swN5DevxUMsLjuv56HVh6vWpr/3wTPa4hyvaF+IZLjRTWPK7knfF89Zgf02m7q0Ss58eP
+wH8b9Dhm1d9EyF8exwi5Rk2ocrmekXBTFfnlp5oqUdPMkzF3yMdx/SXVWSx75kRtSYS1bxKVzXT
5+gNIYu0QLn8qy8yHWAAUDkSIYSTPqs7d7G5f3w68F54qTghjs/aj2WoEyE314Xz2d9Ulj+MMMZB
mQEGoNonWyttJ8PZ20sY0bUfPjCJtcJy+1Anf87aunLZ1GrPaX7IUH2dUsoS1To9xqfP/0rosKzp
Jexxd3HJoD2PUBPttbRBxP2TycairaYWzPK/GTq2rlRp5xjnI0muBpXpp2JDSwI7ud2I3FridVXL
EPwxBW6aPJmG2vaa0OiWVAoSRn/UEN6eOeTUydUzxXDTtiePzNSM0KvHoDWPyiqsEPQVQvsqR96M
SrnBqrXjWjOHfqITQkflH7uqHGZ4jlYeV6aqxpXf8Xqj0L5H+QW08bMlMHfDNX4YpNO6XyaL9FL9
3XBljczsJP3XeRFb90MDdtu3+e5B4EpHhaBGt5yL0cYdXG6a/cE3Wmd60Ym491cuEoqcFc2IXsH3
4QsaouFRJVLRkAW3si9V5AnjZddhJUrTqfpJdWTe40m6qv5SP9SvargamD5GJqwJOI/SZKPq1SrT
sRlUUXKxf7EZ/SO397zaGD7jnCzpkpaslQqqGbRKpKU9Xly09SvWh6aLwc6RSBiKkcaK+kS5/o4z
lVbBzRKJFYFOdG27bnmbBonf7DS76eJB//Z1evA/L9LLD0iq95ajskJ9HyV2WacRyUrRU5Oacgne
nK5fHeNQWOj/gTCsV/VKUhRqXOtjgHDo8NvnErIs3n903bnepVPd09/OI1uQf3W/BmFccOHJfzJT
xg4wH/11VEzO5hzge/fCrjk8jUeqc/AIKPQ8SuEhzOqH/3Kh/E9gEDSc6WnrqeZAnZj5MBdA2HWV
qX+uJsOdEqZ9x4GW6v3oc/sATMfeyijBSqMKFev014EEZeGnIooMoQYGpRWkIJfsVRicp/o+4LIQ
ooIY8SyQkja3Dv8OGNhbYq+UKo+kIIZHqAF9qdeJnhlAv70xUo0VQv+0EBxRt5PaZ+ZZGsEDaIyj
LgaQoXV6lc/H5sz2fzbX6d7vpLtsF/jslJrBY+/kCTQuVNe4Rl5enVr1jG4MCm3q5DoSxeqFEBw0
y1XY8ziVUc1PoAPAeukzOV25KZGsRhH8r3M+aEGgYe2CYEITKzq8PH8tWmxceLG5UUPuiT20vc4p
21TS/05b92opiPM8oWyjNGorJFdXf1nj7DD2FU2xwdsKY6s5sc3bGK9KWhs+dRbPDbvOG8FkLP1b
re64XWVtaCDXcI93o8uq1K8P86jNV27EcCYrvHdSmu/L58xzRzxpM3XIdDDT4vF4UeYYrztkSFet
MszENO8GddS5Ao6LoXYX67SAbLxaBOQ4sFib95+KRRSUMR/A+xsqdN+G/R29zgIhCd1iYPmkXuMa
/U+BdNgsF11dv8NjRzxDyFnrow6vBfrFUijtXDBsW+qsp+P7THfNa9J34OKB78OOQ1O6O3yYXPCF
KGQdj0ZvdXiirgpqOx6208uZrNwsl1MHkyWxCdRD+NnvzmVl7GAfWPMMauEmxuNDj5I66dQqyrpt
zKshoBDb/aTzVaIAWsyi6lnhAyM1OA8Jm1lA91mvk45Wf1IUH1dQ3N/L83NceerZXp9v1f2V+kt8
vF72bJ5PlDUbn2h1EVJUHygNiNeGSgF5iyoFpyOlqfRkP+8LedItQYmMyogsGCKPUgwKMywIh1E8
z9hLnSFHa1tHE+Qr3c5pZhnsddsEnztVJT+z2WaBT/gBPyoFbdQvAybVpt+fDsuCd21R5EYcSnjm
Amx1CAwxXVDzUmX2Y3+ZSSYr7cuw4NLUip16H+1iRxyIwfhCOcQ1RErOz+PfoCtr6ZonPB+B6BFW
LMYlwHEKCJ7SumCGNvK/asvyfvAUbx34yTYScek0EAZ8qkaEGdgN+zEIxgeEv9ArzBtTrGfBZAMl
H5Wpsd9cnXIpio1laXm6HKne9lYcrJkim5SA4uVVp/4yuDdwgxcgiGby2w09AxEjUl+V32iOExPM
XPgjktWBy3Bt9S2HDWi71UjieDtCaU1ohfooZ0r3OP+Rw5lfrnV5pWjZHzisymS+JrcAzYjorRjX
17s87aRKJU6Wt8lgYiJBLpJ+CVQbxrgHgzKPx4n0zeyj9J4cl7r1mMBsQ+vJJto1dxLuPkSmIZio
ch58H6kABa9TSGMfXK43shif1GKeUsHKx06WYdOjai0iaH73AYy24Pc/icwnyxV2isnG+2uCzm7e
W7chiFGln332l2pz9qFJucrdI8MEXD36OxUQJGJ33iCi4O7290H9Q6xroM70mQkBFmgp0G3Xisjq
khFE2J0ZXmKxy+4yiogJHO1uHngE0KqtypfLhu0INJeAl89q7geqYZI8dtLU8TtG8rWAXjRRKhVO
blKrZGOPYH4t0Fp0ACSWFkjyh/+X5VSxsaeNYFt2l73d7DikuRT0B+6V1Ud/ohZvW3gHetVneRKi
1jFXI/7TGcythV45I7DHwnQ0x9ndQn6GARTQeCALuzjy/7Cvo3a5vZ2u6vSACzXQtU5fgbnvrGU6
wXkLG20fyqzZ7KYysnxcWuO3ZXOlZyWye6bMu2nPSSK4EJsSwQl0gISN4NCcHRGfVVtbcw9LDgKP
gaf96r3zBxxjZrXmnwXnDyVKhxHyopG/yvXwvJNAFuJElWVUUV3W5mSb4wCVZS0lZ4EYTdJb5rHC
djKk72yy9jVT0YhHvsg0GLpf/wi32joV4X79nnJ5VeASxIRdlCEgIdFVN2onT7C2Ln/vTqUJWc/S
6m1dtZjWlH9jW32QajLnEW4TmgfSvHoawuPBPNO6Rc1B2C/XO58t+T+6Yv7ML6YlHDcf0n1fifLY
rlR8w2creGAxFhooXkFUKK8wPK5jQCtXu1fYpS4fUf/jiwgrNBscFftvc7C1I52hOXrvKaufuHpm
Y0xPTFEV37/e5bKX7vYPihD5GP4Nn2BqL+NURKORPOWyx62UCEYfCmE/CRwcoQGeQoz/SsxouZmh
WZsDRorpSIzHpTymSj+bXo4v7COWz2ALotGTVnt0IuQEtOy7Az7PGXaKuOXGFUYyXRasWkEpqFVw
WU5Yl4QTiyEtfyh0e2ewrXYiSh6/00Z91h1gwZw1Xc4d9LoiCI2g2OTHoC5RX+yu8f4SgZsAaif8
+wDJ8DhCn+08+ywHXw7lR46UtRpJpaok4GGCQfrcwJkWcz6pmZdSFEaEMrlIpYXJbAZY3Yo/y2aw
QMHd49YR3y7Yk9t5tjZGNUYLancZ35wEZ9PFJyCpnkd3kvKpKZMQFH18QFPOW0HTutIQ3L2bSnz9
CuvYf1J8DB+DZmrn73+ZazEMG6PlOZTFQHl8it6n8gPBdCpRuEO0QYyAExPEMOLgkZ9TftxFmUbt
1iPbDmEEZZNI00YHaRJo0+9Idzu9Z3UiuVFMuYEKQs02F3/4jXRgN1I4xGteJWLM79KczhcZsLMT
pVUKWCHT95GIiMQV+1pGc7pab1YRO0RffRFHVGtjU6L5KQcl301wJjUPP6nUg1GGZoK3TsAVX8N9
i+C+V3uO8Ap19TqE/3T8Cpogxig944lMt7PdEjEfefgpPEEfyWhg1iT8c45f9uiWlNgF8SQefFCc
2GHeGHZMJ354/BEqYduhHt8srRrj6c8uPyqanSwAZK1HsUuM9WH4JdQ7MgkdL0/O6sBqj0aFOVAe
ugJXSQEmcdGWMScPiS2kXUpBkVykAijas87Vd8QoZdgkoOVEw87WVJf8GlA1q9pXcABJkUFg6FO0
pokXc4mnlUtt2uNfVetWh2n214PzIWpzpIeiVLt7UzMVAsEgWytSkBHvZyCht3kUgQ96eCp2CvAf
zWZR4LCZNP1Fq4Ln1L2meNVcHhti7qpfYPKBFxr8qalU0iBORrrYTEPoRv+9QzoLBDDxaA1M23Q7
O7B8FrqpGUa2v1BPv0C2mTgjg/DYTRN/W6+9Xln5G3qt7tmfQwaUjySBl3O34vK0R31fk0z0WKD4
91364Js/PEN9T05iJJR7k4IxkNp/YUlLvK7yp5k5HTjgOgNjeckEJ29CvMCrbLHZNIycfoLTRzzE
GWqh9/qoYKnD+6F8imjXl9YuIsL91QLIbTfmXTutWXPlqylSr0MUf3OVaFwnZHAhBZ73J+Em4375
fMRqNbKToQs7eO9gv0qyJutvQKj/TrupIYj06/T46Wof+n1SuHkwCw1GTjxMp2ECTgdu8nFVcmh4
olLlgQrIuRxHpYNyO3Kd3P4y6F40D3A20yvZ/seChl//NoPbfbvmTMqdN/NI+vdZxmEuII8v4hMp
KP2lzGrWOe9WRCm85xfi6/m6rJEsDEgNse/4D7DTywfixqixYC/vvUmzxaiobIUNczz//DXfEi/Z
mUyrdyHddFLbNrJZJ42uOoiCWradw0BBcPF1P0YdhDoZPFvG01CpCGDxKCjOjNPpeJFP5pcCHJaO
QGjtqYJrRF7n5Y8t/x0NND1jqOSCPP6m0HjpqNaRIPc73kzZqlGQBXVMqGV29l5OHOiddATE5cxu
oIzsxlBgQ0IufDOaMfJth70Lr8uqzFGHfTsrRKaUpxNmmbBp3NmqsBJKIXXnVzpG+o0of9gNbGeh
Dzo2WDJQs+bGunDNkaBxnkkXUjVCVZg9joStCsJm527pkD+FoSrObLNH+mQNLfLg2aP4A8zu33zm
LvZqFP73/D8F0D24Bzj3ybmGeYcLWJWdNA88eLiS6qq7Y3xgLJr3JApMQVOZBJRu6Svatdvv/ykv
L/dE3kRwv44F/Agx9/28WZJiHV0k0t/eWyuiY/dN7M856sk8cYsskiwE43o9XydqSGmPLBPvMeLS
37SnA/szlTWsgvzAShU/+w0xuTF5NtNha7xFb5h+to7g7dcYJQI2VRKfknbXrwkDFb5FpYe2QFUS
U5vQNfzxOEKfXTGCoGfO/dafwZoQEUUNWq0lWBIMuYh9ThruzzyMlfwvuxEKgRjbIqqKGx0QQYLv
+jcRT8DfWkeM4sdFtvaGR/303jFJcm1Cn3uK92dFB5kS9VrQIluP2J0GiyDvrsNZlroYoZeiMVij
cPAEzl2f95EfbnhkWgFjusM8Dnf+6o4bd0MkANJAHuxTUCCStQGXTsLQomrDmmrejJ/Y1imIUKw8
1STpENb+m5u3P5BzMAsIgXKNtRW1KJmoKi6IbI6m9I/gvZOFZt6HY6k8wNX7ZF+6zcrP5uBH9IZt
PNmfBu/LfNAlwKwfGSyPZJOjUYxRgzPGip9yEU0TCEnSR5lzX1P4Bai+kLWfNV+aaH8fbsL+doWU
LAMxoDz0aHNQSuRiDrQhyTXLj3w+UNOmMO7Fg3ovcmruUuiONVYF4aG2Hf4BAmQ/ea5Z/tydokCT
EDqVTpeWeogR49b41JQjLIl4ngCpwoJ/2/4lAuh5WILc1EPTSi/OuE/J54GXnNEj/syqIgKpraBV
CsIgaIaANyZlYtcJOJ+bhe4qngDaAnhLBhN7MdegYpCbFTWTfo1DixiExxolFIDxrSJ5QocKmnR2
YvXTJzSoD+VVRI6xTVYpGGO7mtlpuSxLZpdQFlotQ/vxQF+lN2vNYJ7JwuOHCPDHoNmP/rfsoXPZ
k99e1Txm28lmyeYAimNYz+r6WBWxOMrD1pT+sRADbAoIs5Nv98esx18vq+imuFH3HApcP72y42DP
ppBmr0NQ73I2b9f98tLHRdl60bczcpH3fWL01AaGc6vXuejn8pNWFo6JDwyJtfNKFkTCEaZvf5JY
Zi/uy+pk6LOSJ6S8+g+puqJGHaPQPPzVRj7+rMljCnuJGjK0pKBMKDfIBBgqLscAtglcNIGSevcA
KQI1ruJDDlQ5eiZxmYfT6wnUi9u1yx15/wXtQcKCsLwmADAkxD70V3+LjEhtbWSCVtYgSIzjYrAh
kLIjwZAJIzeuPwd6Tq/7wr/b7lj7jCYrVnLcQu/68IQYJcqajNJgZv9vC6EbHbYGaKb8DqDtBNp9
RQwuv0RQzkkx0wCDaFMNKI8MiKqpx1A6UeuBhUXYNcOFbfDTwM54RBTQGKlLh+TbFLi1uZ6d+yvZ
ZhkKlfNYAljrm5mK9Cwt+cdW9Fh1rEs5yl/RQxHtwX2/6loSYK/ZdgUi0LYPle8caZ8CBJ0ks5A5
Oks5+HFu1GCsDmVCiPrSG2OhIzW27AFwaICMdIprGHGfrVwEoVwFiFwBgt7+0/5VIDA8lyw+n7+a
oZjpCYuUvOVrWWSwgZpNbBU9oFENfhl/Y3W9LR0YyLFdW2iwdWw4Pzr6XkgV58gSF3n+NUIgv29x
coNHCGAxlsnRNWNSauC5Yp/ChZXWSb0fvllVxTG3FDLaV3Ce/k6Jyw3NbvWfu2gE1bCO0j/nAK46
oi1nRPGCMS2WNOoUMVmPX6cCswNR9kFR1/MefIJJ2aVlHTlB6UI+RzPNIje1pJ54jd8nXK+SPT95
CNjtj1iGh4NrLZVObg/+0EEIFW4fxYPLccEBScHzPZac8FBhyOgbDNBhXUo7qHG2Fci7nHkfko6U
M3nBLE4c9WFSiMItR4Y/ifS2ysBWnddGvYQewM4sEy3h+U2RH/ks4Ht0j8Ftge+to6rdqDsbHSHC
SdLpbUw+iaA9l3By6JzgV7IBKEnJHlo+Om65xn64bPwZaf4++47J9r0ipyy7yWH65zAg9PrW8uht
IxWdyexZK4UkgXoPANLt6quAlFCC7KoCXsqfCn7+MwuicHCHtfxAqPKBpUzHSgoCviT7uL3B5FrE
JIu6LCd//qvRcuefCqXkInp7ynuXxudaeOUSna8TEHdpl9xi8rlPzt8WXa2pA9VteSauCEbtfBjj
4mMGP96OF9XhxCZD4iNPy7TV57ygm7VQ0a9QaoaiVj1rD7d74Aqze+Bf+Ri5F2PVKy0z48VvsKPE
Dqrx0x50X8hc/zgAewxHhA0EqfcWcWjn1FvyH7yYbx5csRmBmVw39aJ0Wqcc49H6hv0pc/m+HODb
K57/6Z3ZBvIzvUzhMoUZafKBlshqPRbMnoHDpB+z4zoDJoRBMkZxnqYzI7eMHqFNCd/fsci/lq3d
WDE/HbSg1bG+oOPNAutw3tCHp4JcAWrkMDnSBueJwlhfnAtGuZ1yrzr8irIIoUM5mMXG0qwHRQUD
CihWKYR6H5bsGjHZ21yCkrNAl3tngxetOwqwr5vjRgOFGBKspp/7oRruDcsga67Zu3us2i25FokN
+BElW6dXzygdsu3zeG/qy0anHUU9iiY75/JuijhQzW10801+EUD2dEx91Lr8OrBomjXJVHul/Tk3
s/1BN6A+jX3NxkfR9TTbAkf/GZ0Hmk4X/y0ZHhD06ZuPiGTE8wzr6QDYuPULI8szPHEon95iKYSY
2B7IBQCRUYLfLxviT7KM5OF1HR4qx9DRW08WQKn7rK6UfyQcV8IhDgN+B6pXQnVlEKZSCnb14z/R
Fxud0VKdN+/5ahQtTvQM/kDb0YcmwE2o/5i1Hrb5j+qx9b3D6FmKS+hoTCieac2w0r7JacOl4u+z
Utn/Cs9NBnY54p1MAZHwdC8ZDzatwuKMXeO4PnHkz+PloRw9/vOgUX7CAOgfAIUE428x4rc8FEGn
k1rVw3b0/YXZHVF1vwwDg1U0BzAAfX6Njdo6FOJfrvr0f8ftjkZa9SffdXDSYiA1lv8gtKkkLpvU
lgL8uImhGigAxTNkS+dF2g8D69MX9/UwKfomJizNgwxrp7qK1lOzgPioO7QANkKR9Xuykv7iaMDv
TLZhKbrKvcn387oGdinwl/ELkFAaJ0Xrmx3xzoL6aReumwUoA1GCwGtZIYpNMHg4BLP+7JpUSnDU
6ugKholS2wJlt6yOqzxSfR+ct/L+GI7khU5/77XmesaIWGYi7CDzJ9pFtLPYzqMg6N5hRilKbxe1
C3M/6WQeUvW15WGvZ4VNGJEJtyvjajqbuLeI+QTFW0kIc2hx0uqGUMyzETvOzlxpG56flC2q5LQK
6c7D7MxaHpklWsbQaM7H9NkcihXWwUbyTbxSO4C7e1DNHZB4u8EvcHpJ1Vr/XlCa7e2J1UbsTode
HeO8orcxrJDYdCMzzbUv5NYfD/AUkVX2DkRvv5JZno/Lbm3gZv4szkOu0Mv9rhmgCSg40evA8Unk
lrrHP2j0mSEYHVRFk1olmhL8bNQO7B4kDC097GP5l3+DAtkiSeWDzjWrrk5kwnTq4LQO9pwAvfNv
vPEnYLUlyR4bXWN9vVuYGPh0JNDnzTqKK6boqFIGLoaeBIBpPCqQDkfy0zw3iZ99+KKC4raBiD0T
etrB
`protect end_protected
