`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JxfuObrTyqbe2hEA4QwOiYQWOPxLUXGFSYHQFiIaolfGxhZj1zvQa30JxIBd8weczinC6gIhKHYQ
OiZIjcnzUg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jn06LYncZ38HeZKnzdwXlEyWtMsLkGuKphL9SfI9vQ/nin3CMF2DWW0aaKDA3K4kLYA6+0BVaYBn
UL2RuFCmWsSlnT1u8CPdPkxnmiI/ymwfOFbHwDpi8C5zDfwlSxkcEmk1JF8rhnHEG0TJVtjtx0Xb
DOIfecnbTgrj66wbvmM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FvWDVCvPueXxVjxE73Hg+66ukrxdvjInPIExuSYH3rtAJ+Q67KaWRMFv+yD+oLMiZWrB+9ZN3z2g
HTzYMXv5EWy34j4bEpdxgtMV0THc6JUE8dSrC4UqQRGHZgY4aSlZo4H+4lAhkBWdMGAxJG1vLI8n
EM2J+2s58BnuV8K9ZF+LFzoDbDZRwhW2dReFRqmiqQ2sG7WyQeyRz02eFt/5AY/hAL+T1Xn7Abfb
VzoZUWM6XUQmBytIopfxBZ5q+H8MS0vngPTj9pIOgry5rmepVcRgoTrSqxAAf5bNJE2Ua0AlzVz9
2+aobB/Eth+AL66PQgnrK4wipZP8U2G2MXCZEQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ibFWWG1XdY/PW/BH7XKrn7+4Aw5Sq++k6GO9sQ+2cEkTOqBF5ivD4ad9Sy7RSJKysoQsrBE4Dl9N
fdl/3MPeQybS5AvDlaewDNsg/sr0db0PfG5H49Lgcc82rMjIrbEVeWjyAMxxEf6KvuqlW0Zwv9F2
4cWwSS7GfssRkUKfjos=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TBfxv+m64ke5f6OYO9lUIbDoPu+8GznSlDm1X4Lt/JkIOWNwtkGYOZhN5WPiVhEYzEeKGX1N6cgc
t425QQWopPfUn08uWQh8kMi5S78FcvcEI90+JHFJVB6NqTsw0oNCs9mo5BjDlYFNSawez/THWthD
3XXvU6FRu6JCeS6ev7Vt1NHW9XY02khpakJLLTdM6FIfjjYf+zNL9SW8h24wLw9c02alUQjuQPee
K1cdLsr6VwTokl9niddPPQ8yf7wJbI++74bTlp8ITT7V/CitgT6dAbG/KE1mPbV+a/dbgvK3T7/A
FV7uFV4jv/voXs6JQohvi+J78c7V81f6dbEs7g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
hzTcvoZR7/RRXogvGvuPhkCeaamo4Oy+4gprRvyc7K91a2NzHJ8Wd02xnkQNHGU6hnz2pPmEDNPi
Q1zFjb+yQpmouZ46NJ6foJLjuVywgEz1bNdyTmTMSJ30+ud6QksdSCg3KI4FsHCAOA1G1/VAYInR
hU+Hr+OQ2K4VrD6AmVWuaTWg7taKTZH5GSM7Uk+8gh7Z2zifD0hpG+hoPOC/rznu4fE76bYzj+wM
xKOr7rWnkuQ/BjemuvShDD8U33xmGPNjdeWRmz3KmVFXCWzBwB14hQTGSoWGQLK3VAxkvAElmwZX
Meb4RSEqPlSFa+8//VFvcNVvR6pq470+MuLh8ZJK3J5Xu60xc+kVZJkiTNYfWN80pnQHOR3vj7pM
baeLQse3ic3uTzEUobQMv2gi8PPZ8XoioL5kNv8Z+g5WTNFb/uPjBfh9gn+jf8djzxBywAKqrroY
w8aTB6f1WjanUmvPH6ON3xz0eiXZiYgHBakAH97E1LXUf1VW1ILMVsVN+ksvFQQRQ4wTGL7uGNbS
xOkSjuRhX0k0clKAOJhyvfHgGyz+d1slFvSvqoqfcn58Na1dkB1bO2+icvZ6vP20n4MVJfhsgq04
c2Ws+2Oy2/HZbYXwBv+AjVptbBTFCPs/IzeDfSMAmz2zpMwlbX5F5MaCnb6iooniEe+tCbWcNEYg
lLjDXHRlGPXnm+I4kiNeNN24kqIbU8gkOt8AHRJcngYG85HVi1QqDB/LBMh0Nsmq/pIz9Aj8QB4Y
yh03ib9GuPnWNXcUmiCbhYEAJ5tVfhdcCyE6nGTS/B9elqP9d4C4Wpcfgty/OSyiozTBHLUUM60W
/pXqV2grHeg3efxRVKee0hIML0IwxVTCuMHI90aH9n54nvCJCfbruWd2GqXLqiZhU/AX17Z7iKUo
SKl01i/L2RTtyX/NEWeI7DA821kcQP4DirAeCCv1Feqj6snnaqpUhRYlCOI26O5MixCcPlp+amED
P3MaYrl+ONe1NosVt+swARP42sQhbVmI6qxNko4XU4rlyKJcYPQV0lgq6G7MEKbty2afFNasxOxm
SHZd6TrtVelCF1i4S3OFGmkt2JmzbrgJdstRwGTVPulFxhdG3VX3GgKKwRFFsaOT66uU529HK7wy
kEK+RsK6vz/dNJnhf1F1vnObNWUBrwqy6ExIzckR7NrYPPxdaR0GgVewU2O/5FXxTJZTYKWiYeoL
VelN76eutw42leF4Dlee3ZKPRzdQz0esLdj+5Fri9RFoOkPBdi6d/fZLb40YUbr/QiX/iTfEjQec
1YOMmTTkMj/ETPk2BqT7H2EHEEvf/eP4tgC3ShLHO+32smBQ3r63u85lv2UD7JVo0nBaXIjIsiYm
z/wXcTxZcCJLQW8kcva58HLUvsRqa1BVhtcp8v8zRcPX3RtA1MGjJ1pnu6TjU60+14Rr3OrMjRbJ
R3B+/9iztcmFZukN/es7keRExMm90GpUs6TGIH+L3DYajaSEMjcjt7YHI0RJvnQeOoufugq4poMW
tgyrLic3gFDC5dQwqEog7hrNaR9x+ma1IAezI+irGE4cqvtKUcIwMTeSA++JZeEk3iH3eMfM5CH3
5IhJGirvBB4uEZAQvyZZJhWhEJjU8+9tVQnadmiyf32LraWPc9MgRBftjnERP7hoCKKamHEY2Uxg
9hGuNQVgEto+M7boZfsTCFqmbmYGT9yR/g9VPak4iYqB/iBHWxNQmSn8f23QrWZxK562z1NV/1d8
0T35z+8iIGO33uGjRvN+2gOP8FPulhm9AIHdm8gjZ0N6DH7mlXCG38YXoIBitQgUXhi8kgFcGk4q
ETDWT1mQdIZz8vYG261ELL7RptVob2F6txg1ncXhrd2jh/g19fyFJTtWtG1estA78mUpVP4WFAl4
gQKMa7TIpNlDFWnVfOQtLQVNC95J4Hw7K7Lr99v8wDLitDrP9rxqsjfGrq1fxZFgv/gSTeNGCWI1
UQDlIs0+Z0CF28JHn45VHqgS5MHk0ZRrPxImyupdGQjtNHXRqDto4rzKIJab40ZCj27I93MF91KG
nP3GZVwTUSrtDxzjFdrGIPbnW5F+ozQAIDRof7lSjbJSETFb3QKK0Exw0X8VH82pPRhH7Cmzw/rJ
2wdRXX82ETNeJmG4Aqt/cVokXlNkcBUsr2VY7NWklLE16U1dq8glESaIR4BvIqsdCJ10skJVH6LV
XxLvkjkV90KPBPDFmFWhni5rnub7kxtSMaT2/XjbyMyh9RdkDcW+HkGYK5Gr602iGvivkRg476rE
PpQ5+bpuJR+KU72LHK3ksG9Gpmrsf4Ykz81XZ68Xb3P45sK6CwH5UB2IPkG+zqRfoXUdVSIN5we2
ypX99vJGKOrKO/aoxgvzNIFA0tDndjeogtPAcqbHD5+qK4ayGf5KN6DCKV2VSq9ZUhdj9EeW/tsC
u86Kz8FatsjTvCCYRsnfRzahGWqGp4I6NkwTfJXni3zKRQl7++gbuD/Zhhs3ZZbwwhkcmF4K7+wu
EWuDzQ00flqezPmIYdzskiZVF6n9Ig2E4uiESeXL6WZiDpA4+jzRNhdbKKD+ZW8f7KlvtdPkV7Vq
TwQrxFOjhaeWIie3ZEW68rsrhcvcLMJrS4hiLqqQmTJSMS+t2HTzLvi/fNzMsODiQ4nwM+1A8qwN
LSa2Ota/EgRRJrWtZnI15fp3thgesi0dHBpE1/5LQaQFcoRZ1KUPBx5oZbB8qpAB+mVZjsX/GK5g
5sgcrq679CBpKlqgQ+1sXpEplafArGNpNm5CXlcA7dCjAWX17rgXyOn5pvb3aBVuHl7KDkxCXL5O
f2Q8WoOBeEFF9k8L3j4Dyw333PFqKtt5j92MCsED4TspFdXxx88VARojiwp3o97lXm3aFeWsER7L
sOGrK7YbNy2uwomR+V9PXiWEeh35xbEryz8QLGKxZZwLpI3jdf/ixNr9iyBFLud9RQXrg/cXhxye
OmF9EKGTRaBkmY+NML3wDTILRujMAnV1GNJ4Vz5fbni+AXl/7YMQuATuziD5n3Kk0UHPI4c24kP3
bmWejdvPrBYQNC1zj2aZ76dGNOUlwXXd3GUZUjGTeNdE46yUqUBPy/+JJfXkAgJiCB8MgennxNei
OjYvWWVJYG7xqXgTM1pHWJU6zypULdNgUj0HSjif9KXTSTYSJZkFcUaEe9vg7xhquKWI0+twvsv3
2LPy2zybOMCbjni200AhFHJGR45Jvf3rgsu8/uUy4So3KH/t2E8i2KdpCjOyv/gyTNnl+wWvftk9
blDBwDUCZ+FE3zEfXVSz1I9/+auAJhawXJ25GF5yjLZtUF328VifinukkT0JnzA+l5iJ2rREriQG
081N2mhGAZcTvrxRIWxJQAES7SiAcn5RHtvZqDjf+c/Kq9VeZj0ocqpiEXEbePtATybm1FBCA9Vp
uP9uagGFb5F4WrMKqNZg38C4yFW/u3Bcklao34ZBVF39OQvhfmyZUQpdWFmflXytca2A7ot41IH1
ZWdmP1ViX45h+a74lnlSA4konctqaaXldSDE2UIPKq/PPsq2FPuEh9aJfaWFWsPRa+tW5cVF2uJA
GN1QVOvrXBQgo36fOwKEYCT7nEMomDYKrl7OB9eJM83ERkcDeYp9GtXdiBQ2lORdvlg7uOY2DkeX
jaXtTqG0EiFfZ1fDJ47tGcD4j1839XBhhQDg7vzs4W3cjsUupAdsuHXWVpTmCeVecboeCZsf658Q
62JuJ3dIAOWX10EZ3/3hZeIC3hSm6N5fa8fOooPNuqC6xVOK36nhyOn1han1rpF1so64AIilRS0q
a9M7G9Fg69c1gmoQ8ugAoEhSxAez/enT+2qa3GjdtBSQeXOKmpP+ihtvTwJGBrBg7s2VPFGZonHR
p9aObMYr7qdBf1IpN2cHWt2JoB0caJ2YiQE+QSyQ05i8zSzfEOts2Qkw8r/9p1KeFqzgQYFH0R+B
nyo4OVL0/lzU9m74vqR0tcRYVw5Wof4RcRyyJXVxcPbsoHQ0T6E+orQk5NXQA3zB63vTZUM4WX2b
f+a1rO276zP16tS1d5U4J532TFIwk+PU/IzW09OlOLeCMCCep6Z20U27F8k5gMl5zNKru4XSiiGk
RNmHSqsQSChiNycXOTzc/O4jqnubXD6QXWD1VivQitDsTBJ8j8CXvrxBEsGsXeWOZE20q6eRAvS/
rLuaXkef4CBofedI1aJaRZu50OHCMZjGzPnVDcm1Ox1Jx+FXwq+0cRGwrUEQ1k8kFxM7eVkGotyE
X38OCJCGnyphZa+2vKkhe20VGIU/xwuD2+Gh4/aOTs452WzIGlQ/YhvcKPqVAEX17TDxthKQKKMI
m1eXggiW2YMO+enK7HfYskZP7ddGHVkOhNxFyr3kslfR3NTG1n8st54k0a0j2+Kfaw6Pnc5PKQD3
HAM9/C8/mN29t2PuSgwwWahuPZUjsWFlHJQq3CHLvZHSIgdYt0l1CIkFlxMuTxPe1kPIB2KaLknj
l5rhHlNxNLaON4eKCvlWH3OxDHGbl0zPmcWbil4/MqgK3OQmtom5u3UBihrFfYsXG3nN4eCF/N7S
W2KptFkM1OEvbP22RiYlGQbMsbG09GwvP51qfORzt1CAib9MAVYLpyRmg+M/OxW02Jd4pzuT6Z2y
Y9gxXwfIRG+ScLFetTVUSnLF8khfM0kCEr8o4Ab7R4jqS/AIAOKh+5AxESwyaxHpqejr4lj30WS7
3EegPNmWHRztSApskdoskkkx17gZKuCEhvSVPF1n4Chi69HSbFHXiDs0gUxTLR4KtstL8A75ioNW
A6kIGxpU+0h95JZyzbhRJyQp5fRyaGJkdIkpw3n8KTJ+qfB4hdaXY3RFRIBweI7ywyxrn7zgxZyu
KFaEX3KYHc+ODHzL4A5jjJ47RbSJF81aQH7/UJIYXXsnlRypMyz5keUQkSy/I0/nUq/cTIKSTUs0
sw3dKaxqNUrcHwt8C7aGiHY7vreJUyeyYH40LvajunEN9ZP7NqanX2bXhszkVa2rBaJx7PeofqX7
vhFYQZP6ZJ4Lf9hp7xxbQCCym5hzawuftM1fJzUtAjqdudHHT6+1p31z0g4ZScZYsAkmCFrmZ4IG
5PyWdfnDKRwPJGpvPFN5A/VlOyIbpP65rDIlLlJZWU7Vgw6ORzpfnxnBGSwgEyHZR7YPVECvfTUa
sw/wS7tjD8j6eouA37uRwKrTtZaHJ28+/143Cyj9VGDYEkg3AwcoJQK5Xsq9LJgVi7VWFuQxcY9y
LXnQ426jwaYgZWuw9zY2quPrDzjXB867/jAZjA/ZFFuWmFM3jKlAHozc5ppukUtZLZjCeqr8dlLq
jPioPP3qp4Iy+SXJ+XwnyJYvSw/dkFl4om1Mp163cVaKHOUHP+6LfMWIfzqwZmHPblkIX4j09NtK
VIXU1GT35pYuol5okmJDP6u2LYUvSyklcE0YvWFJafI9WoMbHlU48EMln2gH0Vf1iSwo9YdcoNoj
d8zAr03wxngCV1WYYS8r5tBotrWQq4d5z5XNYhVhtHn/FKW/AJ3YDikb5CnHZAV2n28UB1HktJj8
qQO5FAy0DGOo61sr3zDOkAkm2FsHkq+tyBZI7xe2zeOEaZRNT1coDfqrsDvivzwkjDCpVf8f/5Bn
WoNRGuaczf9g9nhbh6/mSXhhLxYeOVYB9VkDB9Q2X4lmIIUIcYM1yESjSHrzAtRtC8sT6Njc1N41
f9gH08Pu8aZvvIpGPeqxTLXr46Gwf/Dus4R7JJ7ztu2vxYGXidFEBmnhsMxMpV2Z4BpBNiPC+TXG
DCuAjwU0nW/DmnQonU088kUD4MgPUQpsz6zjC8HYquv6JtN7DB/kissUMMbM4kpfo52XiqCgovqL
HEmqrXWbWCgHKi5y4JbusAUQEB+OjqVH3d0taaYSJUfUv0wGlo+zh13GlK3in2UOIXe9g0N9vDxZ
c1WC+YYYF99kLcOJ2HSlJJHE79EHTYaitajh1PPdvDmS8u8TUecH1hfHSmRI+WlIxZGsoBTWtdhv
k/DqPg5qzB8KV0hc2ikZqUVXfXAyRkSC04/szA/IsRAPhYVilzbq/+u1wKq6o5c2HjGWqyE2qPbX
kf/mLyQwHJOPASBbg2KpC8LHNgOkR7jGgoL0T14DsBizYOrn2eaqY/HwRl4p2kUSmDmXAML9rcj/
uzfNrRShRCJALVnemuOukjmfTT6NOHBi6Yy3GN3iMr7Xsn1PwJUbNfNEUHRGcLxlp5OTRv3PFgn5
+LmAW+BPn8UPsagDRlA8Zk9rHYLIIwltYZftAR0WUBrvZiAxEG5llaCs+aZ1kwhhOeSl5LAJtKc7
k+4HNW3OQyqg76kLdFoTGqu+futgHwu0tE08Prxl7ofmzuj37MAVAs9hrelVV3dwRZqxModmYoQV
O3kgBaZDJQ3mCsF2xvneycTjF8S2ttvsM2UG3LRccdcyEeH433z9QRvvfjmAqseTRwpukD91D35x
uXEWTzF1gGGEHXlnIQXuh8xRGWkIHmEzULYqAcSpmOP2yGzMzD2eQBAcBOm7TZmRdvHSivjjzXDw
TO4Utsw0fWKCquC982axAQ6U7zZxeTLIV6g6YmhA4hQD1wZmg2ZMGTNLYGccrbHI7t/Lbf4YEqwH
VHUlsAMeUCT0FVzrBT4vSKu174om5Ma3jwnPI/9AFiObZUYHh5APfQW1eFvBJpV40BpqRAb3S5kl
mCfHDOfwcQouZvkNVqs3hfBfxHDPoUoQKzWGQ++E60ncmv0BsWcC9yLrtYAA1axVg+bMWhBJzMo2
7wkuxeaBSdezNmuC36k5koLcymiqTwWLF/eFYAqa6lzslzZoA4ewNxQp4dg9k4CqF7XgEJHYQL2z
WLO2sXG5sIYfLJZUX8LkeDcDXGzNrjDMpkHAWk+kTFhWlUbYOHNhN/3PXcFn6+2bBNnn7pau/8PN
FQRdNuQvl9iIL+94AOsNMXs/ysmr6yIHY93+TWioXJM55eVHeVy6G6/C7VmFGhAymIvABun3xJq/
x4THPSraJ/6UY6QHAJ2KCvAbZd2aO0n21vTiNdEtWb0cJNo97mS9fna4jX7Tw1+KW7QuIy6aNigM
4VTcQwnNvs33GHFW1ctqprRVTD8yCNcaZ8y91Zhe4R5P0yksqz+93Vfs1AQVr7Wblw5A7xG3qOjJ
D6r45fwEe+zQR+BGkefbSPNaVX3z2yrqkkaZX3ytSLWtJVqoWqXg4aUXsZSkaMf9Gpi14E48CXAb
nVfj8Ogn+osud5LoBN+fR/5grqtr7/chJCmjIqVjEiDq3E0PGgQJFr4y6FCbVkTOf2zV0W7YiDPL
6d7B8CwfshNoePv/cIblBZrhZckUcI420P+IijZ3UfXn6C6R2sckhedBcRLIIj6Ub0VekI2+5Y/e
7+cxIea39OdPNAK7Z7XKbtrSkI5ci9wK4Ea/eWIxEHnxqGjSnn7YIbQ/ypF8ePgBQ0s0/HN5tN/r
uYzhmK3illcrSNmwXYSi577t0Bv/i4cIzI0NtwxSxXtgZCPqmQNuRe6+sP9NtLHtiwfwaDM8B+Hw
7S/Vnn2HV8rVWKtkgqD+/oH6fUmzet0ehVQkl5KSeFG6pxUs+fjpKE9gCvFTTDtaSkPim8v7GWBB
OYtHDfAwfjNnD4jwvYrIKRAsunrK4Ohj4x4xCWBdgXsbmKJRjCXEublcZNHiOD8ywDOvvLYo1PDq
PaVgunbTxsZyY2PczyqgBGOW212/QeJyVhOQuSfhv8QdYpOyAO/WLrZn2+Y6Lx1x+2nt1I/bUAo+
kJucTb+08uMyTtnT1Swqt+QZZGXyM5E038J7eEbsqJ6H5BzcGz4zycefWOFrMq7UongZlrgrGbwL
4haiB6ia5dWRe1rxJPRQwG5uJYBv9XpLJzIJMcLvAOzZVMt9mOMMsLKTac6UNZtxmTACLVTx+GLj
pDPmEgQPfbPcby+0boqgtL9lC16zhTeCqMl4r3XGvh3U1PixLukPftAAS0f7ey+YrrAS4wPUbwbr
Ine65TldAmPty3F9+acD3EpkTIo21NdX5+QRJfKcmy08zYvvaJQ3UANJQkvhMY1JtT7rWmAyABkt
TO/jHWFH/ZetKFJsVJBHhwTxMZ+SP05DxXF3XpN1smpLjK/p3RyJWpzr5lS7sKGsbDX4q49Tkyky
+VJxFHyueuozHIBI8xXjbG0uB0Aey1cKljoq9abfmz+sopXdmnSZlVwb8Sp2GTJOIu0SQAd/urm5
EfiPSpPH4A3NTAxaH7BPjn/Y57R1NRV/ZbjXVxY17A6eOOdSn5JKgbey2QTevwMmSnpZ0ukzpSht
XWxQW9DORbNMyuAZZozhC/Ez1Ke9EBbINqjtyasD8COgWQ9EKsgxTPXxzp1kMG+ZRZdOgV7sRYVW
vYgaeUgeWwqK4bZKQY6Uro1i/Ses3G3LYnzWVjfRHh+q+PYHsIrUtzTPqKK179YXkJkRPI0R1YGu
TKeoEUSWNFhg86wYi7AOcP1dS51VgE5/CpKUZdFnKwBErsPJvHhUv60FbkiMlfG99a54SYooq5xV
Nc25xV9aMwGVYOx7J30WlPk0vrG4204yc/djrOyhqzAPcwJpdyQssNGBB9LqUyWJNtJ7yFWlDyFT
bwJLhe2655dsZ/NJXLu2s5ZOJqqmRcJmXP6fNquSJjj5yHq/SjvoVErAWWuL9v8+IXFL4UaXlwLC
msnKfJeqI58m9DeKA52iXV4hEdHiuhZbS0ZseDOhrDkNiuzYy47ikhmBaoa96g9lIql8J5XbMA6Z
pdHWtjYzLj81sAYmE7NXAU55i3wVPz5lDiVW4qkGD+Lz3zjmgCRK3AOSzf9BPqcjU0qjtqwyZGyf
ZrvYTYrhD+kbmGHz3qYEzSIOkK/aFUcL97Gp/qysGfsukTaMciChlBGtMZgPSTq0tBCoaokg2zyg
7EIv0Dsm0BPFE0+EvqrJwOU+2Qfuq/znt1i2WOTcQa9KZlZdef3mJ6Iv0auow+Y5R7HSo8ANmle+
XDC9wWKPxMslBtl3tLQEQTy8aaEHly9YFaznuIiUpirFnIKjXK/39cgev3f3dzGytLAAaO+YPFsj
ACQcncCgovP6CCbLyr1uprp956yWJFbbAynFKyWYiNX/EsCZ2Sw77RXI3NHBUR9vejtp4UvFwie7
NN7tdygnGz+AknHBeAyEBoDTMa8Jpv6EV/9Df49bhhZOtcOcwnZOqJAWLKmNEFPLm0TZG4SIzG2G
0GZoXaK7x1CrMDTyVb/r7a5QmFZTbAn3W5u75iv5SK4qfiUw1LhiOM87xWLGLGuBf+WjMNEo86K4
LD0XiFSwrAeR+/p/jUPRXWv9eM/KJTNGsyb0Xi32xmy6F2klACMFt4wF6Wl4RRHxoX7nb6WwUPMl
ZftJYfmYYGr1SBz0GvZDauXYjcLmWD8w+nV2RonnuAObPyRz3nj1mhM2LdIUzO53A3LdDCABbxWL
IXgYBPcXMPQRgqKOp7g6PdV43Axe4FCnzQI6944S4Pty/7X+K+8bikFWhvH3jUMG9MNX2/YceD2i
0fPlkpJE4Zil86qG76YKSBp/+x5VtF5sB8CnJdZ/wjTUcM8UFa0RJKBVdGoRuK77xyPJUSZIPBEa
IM1Hm+/Hc+iq+SQYDyi2OY9Lm5b67L9Zu3IUqy6A+CN/epytRGbhjKvghXknW/3phmsrPsMUUzs6
CS1yUbOoAFkqg2F2IKAXcmB7bPcF4wwO4TAYp3nCWKf3IGGg+rJJQ39nVFniBnjXlme2z6tJttNv
YR5xkUxX3EB9yhhQxFr+/kDsm9QS4EhO3UzNXDnTBllOg4VGj76bRw6/D2UgAXiuaYKd0/2PPOQv
6dLnsJzYN9Favvstiw7XAxENncl8PpoWwQnvmHFMjJtFnpEAJa9foaJJIalZtyFWwey4urpGcZFD
tKjXk3Vf+bVxfu5Fe+Jvaw/ra37cYEZgwWduJ7zbrWvmAdAF30I4dYI8nqfauMr8xnGhhXFJB2Ru
+YhyJiMXm+odqs+ryqUonl0vmtM6rEnuMbfi2A5jArPWsV15rjVS7WZ9leJMt3pjVMNmrwZYc5aB
mCKqcPZ/AkwXhX8rkQsW4C2nWq3gTXUtGEi6a2DkTOOysRJgNkdIcyTxS8VpDX9IAizGpZveTP98
LUPDmm5laGx2HfGxJ006bWY+hnC2AmCR6FuTZOHukKx4iE73PmFn6oMQ3YdxXaQPMxFSWUuIkIfK
fNdfAU0kU9muVCcmF4XTN6noBkiOCCTRe3AcB79mZlDi8W9eSVTwezjDF88RjYoPa/1DbD48bqY6
Vw8ViddXO+2gEg6f3Lg87ipmXSf1JTl+tg19NYEM0oC1xkDQ8X89AbpRj+o8wIDi1BBChjDouHbC
NRSiIyySZKjW3Lex/IszqlcX3NaoFSaxh2CDJLp+g2O1gNcdiU/ttQFMm8UWV04bva5L0eniHymo
Z+jWhpUCqD1Gd/6f9J/GkE3BMypE+Igi06cGaEbyFfofi8sbx1z228iGU6nouYi8ezgCVtVI/MQW
zBlumY4wV1ErHsTpZ3eDa984UlG5hGiSlmbuu6fGHqVB+g7f1Qk6UEKLettHXnpqB6tVjpJYKLBa
Ir9sPeQGAabWLffx1Y7CoEw11xaK0tXOA0GtQs7KzjoiM/BLIa6s/t5jHPO1/C/7iA4ZLJIDN3TG
vJ/bY2XjpIBfsaZ9PnWdWlxTtuTQzrvBAKN2br378l4MZxEbRZmF2Gr1a1Hp5VYYJYuynBv5Tsdv
YL2hKTzOE5Ntqy2JnVzuhpM9NZAZoGaj/I8Q0bexwwGf2VQF50y+zOJPyj5qGJWm0v20FC6YbHvP
H3yMV+zjrT8NXzarBm7R7LA8jT73KV75+KyvQX6LFNBrzHZ9jIlzsOKoOgwRkx+B1Q8kKBeUyO9X
LXIBm8nfB3K3XQBjQEGLgknzFSOITHYIDXcae5J6ExIVvPutjbG4oq+4ZbIze+9jnIWbaWrRzxvw
EEW7gkkbgVkWMSvuPuQzQUjWx7kPN4CUda/v5wvyI7UeHzxN1hKojlddYPQQc/XVx4r9Kj/xKD4W
RI1NTvWdwZDLPXIhI6oXbPdO2ES05+Btbu+QGcog04CITJ/PKKo1vdbPZh4KQUngt8S7FVv9JDtH
8Gc+TmvvDpMxBZuenNnKgXlwqz5197N+HunaWlIfwI122n3scwgndLYUiGzeXZtsHpsY1EP7nXHS
1ckGK/7xOUoRMVOoiH5z+95/7e6hLTs7Ubar2yxKjK6D5sWb3GvBtFnc6mDRt9VqFulo1B1Gdd54
OvPy5aMAs7znwu953Y1ZRao7kv+3EXNmjyS33IhYWYHf3yoBeOWzv/chtT1RrNfnVFgxhyyuvNF7
4H8eHYze38chKlkpUW+7TXWVquyY+OR3/AlDw4gUojVg8/f0whaqFYpGGRj09w7AYdrPX/3pkGQk
h+VZ17/Vy7g3WocTyG+Qt6jIWKQ8vGSs1/2aHa/C9vxk3UoWZn6Fz+t+Ap28A4gVLZQNc7/dHjpa
k1EmDlMA78haDxXMDq7zG0XfXUGkr6PL5vmQU/nG6CATbrujR5mf5h0y2gVwQqTK1zAnzIcXSkFG
EH3mAUMGYHz9x5MsTH3srlCJlbUyq3FGosDqaTWCBdWMBuMHd1BiBn6sgpaWQVjAn5cs0RhxOVts
3d1by7nJsXzLuMaFHGf/zuwzAJxP38uFjGrL6XhC46rYH+Bigy9cm9MM4LwvjfXcjgiT2S8xWWB3
f5ewAejK5hyRFVOAzdSV2wU4EKKnZL22wSyndbz59jVTAISLoeYr1+HPirOyDoVVCXhmfxzTz6YB
c3BH7r119Y6tHnQLiERS2LoeVyv61NUtSwM2BhkQ7MbVLgP6Bq4H0lLJEZI41/+PfPGZoI2Bq9dQ
O3QDaAzyzNVEmfyPHn1293U2PS5hvM321GifxYuXYrssRT0Xf85Hzgt4vhMi6BSdacSrb9Tfh8FN
vdspG+xR82suxaqK+0wVHjaHuCdfJ7QNHAqu7sq/L6dUbI4l1lHQ8Uz16ypT+uAmZ2Fgr3OpjSWk
zHZRDG+Z/XsrL7oVSKBVX9FCBdbhYGKDBrVQ1G+9+U1jI1xw7Xsfju2AmVYZv1V8W57zImoAKjR2
GBfo105OvBkLhA/mZRDR0ZHqHKFQrdyJqyqBhMKFh/APSTNopXoWEL7mTe/Mu/JHO9l7LCtt2bmX
4CDP/fbvbTYBwo0cDyrrB2e3kmpTCl6OeAIDNX2cNFxPrmKX0gQn35l/cCs+ag1Z9FUxQvipFsAL
uxutHCggstIo5lQ/SInEroY1BTyBH3dSt3tAPLbFVk54gsrLX8zYd0pee+xZ+jPIPDHDSgqCCSav
02WZGj3TO7K3i3GEOd/+Q9ZZVi+FipnA5MvPf8hhnQzr2lws+gNe8VqsLU8NjkzcrswkDT9qxLul
nZo8cFl8szHxqxde7S1BXOYvCtsmwBEuWhm4tHgGt1hM57aCq0OTg1ZoyYgOabcaHPWERbxKKVh/
1fxeVhD80avDzMEckXxMFwpmps6Sqe//EpuHhZiPdlInQfT6e4b+rdJyFoQVV9VuBs9eU43Hc6ey
kroKEavOqapTjiFNTLi2lpe+nYLFviafmfGMMoj8xbZOhxA/E0qoOoi3tLWMGBE8U8/Ee+fG0d6g
sEyllMAZDUIVdhX3MOuBjWt98Nb80HpL4+CTDJFUFNUEHA32BVC7/URPdsNYBk4c3+WYBn4tzubV
gQBy0qp3b3yjaMMUvf2fldDXjH6usNV2PcCUsnaQmW22R07w8Aaw3QpO5RasmSw7Tm0SPjGmkqaj
q7REsQF64tgpRNS2WoB3xWzEra/QVOSbweWQkYU+45ZXvFZRTGb4Ex1pSsMvzatHOJtBaj4eur2p
SomfQoIZ+uun2i5PD6qH8d9Ux1pl70X6DbfLaF1XyunIBe5uW/4o6x03h2lzwIgNNQZAx+Od/ao5
WVd/5jcVNtPGvj+g7rx9lh7M8AciUH6zSpnsEeDzwWWzPY6Zhb4C0IXntVcsg9xELL+FQ0GWEKYO
ICBzyCdDTnGWkgFFpbdHrVWetx0sTPIqG7dIwC4H9dJc+sVxZJYlzmDF/KkflheznRIz6SEfC/E1
fFt/I2zGF6qlkK/WyKG9hEofguAbOVIuXZRY+gf65SrvwJwxkyRJ348LCjhJDa7J8NaOLJLtBWlc
w8n4p+cbXx3zHj0XpwQPZpB9rsKaX7CfrCDmr9ymKl9ZnRMcK6vvsFJINMjEfR29S0CCB0modI+j
fzwdzVKBSMeInfhC//s+PmjuwcJafrj2bOlOJJAqG9GvC98+ugt878ST3uOOTSZwjNYFLhG962Hx
4lCu6Qcnj0kvqSLLp3qnMh6J/Zee+/eCWiFjKZAD6D0yqfMvExCBXigT8NT9ONagmu1lYCWM/fcd
5jZR93Q+TORYlC10y+N90ByZT49R7ieni8WgZ4HgQrybDN7kONUkm1SNx5ncC0hds9XZnLUJ9Mjr
pDdk+u93ZnjlDEu5E0DwB+TNDE4lb1GLWTDWGlsvgGNAbE7Q4Rd4ouuPXHGgmAdXHUvUNqkOgKqz
adGOXncHwSGd8EtwnZYHxvEVU5XTaERpQ+NEhG5sjGwa66H5mTKOyR+0NzQCdJerAoWQqfwpxHmW
Yg/l1XLAOJBb3YR40UhiTq2EmSmYgYMv+LKVbYEKmi4S5IdZMXRXmGhNXqt4Kdj34iSKtRixZKGX
PWpGrIsFUMdf5Ba8giRhzVYO67DFzhxFTIOZblubOccItt0udDorcfAqqDpQ96K/19WuLvbCIWwD
SyiyULgNoPIji4tHr+jMuQTRLZRvUedFIqtGl73H+TrnoTUZigCKwK54tni5wSCNdVDwkSOs+H5n
999qgbGF6IboKqRi+O4J1zdOTW14PFATfUAF+MtuxijrVOA61zQ+8OK2xLUwC26l0+hsznhwk+8x
SOpkEp1CxTxzKUA6PPDGAVj107htiG9xq7V6HooB5rqy36nmi+UWqQ0xoFP7lSMd3t+YiIXVkg8L
YvgQDP8DyaIW12IphqV17dU+TCbrCNsJBKQ8sdf1iL/Zxr09z8yv+S95WLH2TLLmqjPParuMjDWU
rB/dfHLpbxvbbiGSnFPK5OEhEUxKSS+dbtZphgnBhIIVd7URdpDjGllspVBxHmn1p/QU+saQabeH
smkwMeGZhIVQU8YvqioTIb2rbaTzi41Bl/7w6eI8z18CPzD26Ix2UarfW3/Utw0ndFfnt9m8bAr7
HeiJsq4/B7p//aCeYrSXiiyhfT5lAoUT2l742b8alrlnioLfTaUDAkk5o9I4SeCWskvu9N7jNnSp
b8/YGyXvp4xpbld+D7FZUgaoIDrQPdVqxN9eM/yq/hTonOp30oLcRsl4gDCcTRiujU7rBkN2EmmM
CV9yRD543GG613wRODI3qXyjctXIh7J2b20rb2Jh+Uk42oq3wt23ljvBSGWks+5nFpMVVGGbrZgE
KjJzU6MLsxZY6s+zS0eo1Yu9C4U1d0lkqxnimgrM7xOl9ZCCCP8xQJKqRUKqLHInSyNycFazGTM1
vyEnKvbdfAvoB+3x++boui9aX1t63xcmx+8U4SuoG3y1M6SdtS7ooYe9Y/vEH0qU8Lm60PclDKTi
CLJ1HbvrCQCZiceWWQ8SrprmwjRvVK3m0jeSO95y19iSxyeb9TqcndCGgmM//AxWzFUZBIa5zc0I
S9bw9bYU0qYR27hCGvwCdDZOwGQcO6fmv28RJaANKM+/La+8CtSDUYroK41tUiV+OjiaQbgBwE9T
w0jb0ZkW9+mMdeWa5I5XskRLZ/wTV6FR3rUbODQ6mhgSmacZZbiEfjHRA/PhhLxZmRcPMYkjjDw0
a6+TJ1kwF14WM1NILbDvUcmT48XlLEsD0m97JsfUwPdz7xuPz0m+Gx0Ew+b8A/9szh/Rrc4VVnAK
mb0H36E26Q9oBtgdpnLvyqhkVLGlLE648NxC4X1pn5sFX2rf7YTn0U3LeE93ywtCbw9CxHRgNRQV
IJ2Fnq6aYlb0ewPN4fcwzmpaeRZhjv9ecpe0qX5wuj8jmX2MW+Nsn6uWnnMejs6iGOCMRGR6gy6P
b9mbdxCzriHDXi4vIlb+Ioto8kIbg6RnpxmleQswJvlO6nhiArCsTycsG2wOWR0liRn9DNM5BzK0
IxxM4XM/UBVugz0ck/BOWdklJAa7E20ZS/tfUn+n7teDJDFOwHVssbEJPf2Q9GPtfCsINbyVCMLA
V3RwvKP3cyWMd94xvPboLDFqMSwTJ2qEBbRF7sNz2SxF7h1FlRMrmlcub7j6PNZAGDODrkQT758d
xGBHlJEiAbHcKx+Ks6RwaRsb3dQPckZQ4n8acpLMocKK26DpKH9esgAUlSw+3r97BIEqaNTfqOCz
x5lMhisJZu7EQYiidmAvnKac09XNJo1M86ZuXi7y6tPEbQKPGdaWzmMfQ3KFAJA3vCLOjjjdXzGd
DURn2H4hoqj29t6C0K2LWTlb3zLSPk2mwyGG+M9POFlil9IjM3CZkmCwanThDq1unsk2Rwkc6ouk
lxOlfsQIOBMKFkiWPtO5tEb6r8JfS1RBz8by7v8xeU/JjuAk4QyKqdoD5i+hG9YW8Na/8Qkhrmvw
quy7cCw95HdPI1HobPdnW/vUp6biC3/19jGyaa1trA8iK66ikJhsF5eGDlgGXURJQBkVriXzTDI/
ljKLmzbKo3WcsG21p5+ofDQJlncyd6/Iz4gcQ1WlwHHmdEY1K+2qe/B7dXrMvQEX2FqNIefavrg5
VMp8CUl3nwBnae40+uIbuDqt+0kZ0Hl1BIF6mown7WNCVcgr6YG/RVEeYx2q+R+4KipOYNuPUFDr
8iGlmcNn4hPndXb+/dC7Q890Va8zoEUjf/axB8XDyrmjBhCODASOxLj4gJl6InvJXOL3bj9dHGmI
jiE8Hz9gQYjwKTXlvIApXzKg+eXzMe9lX75FJMRfQqmOdXPIhryVkQUVNz1FEIgbGEFaHbiqWsYE
couRMqlXrEe45kMZHsrnl5DBbM0SaixYOQvx35W1pMOYTdvOm3lSIZ5bujg0c9CPNX3eNFEGUBsH
iBQ1XyHVkYUA0OsHlnC5eFgrObCmy4znGqzaY+aawrNM8F9o27q8v3rNyAqUNWsw6Jz1Fb3gjW/J
LnUICAPCHWxoXHQ+uvj/c53jHktI2iLlBhMeb3ArzR5CtIE7cs0Ei097QH/RdPeKWYMazera25wN
dc+1Riju/o71MLZwQ0FuB+XHTL5L8rlvqycHIFV9orB43yYb2rntqPF8DLn+6NnRE4VFEWRFWwHJ
IttlnLH1EzT6DUObxeViCxpwdeSiZWwfYswCTG72knqJgbxWtD6Z+HK5WHThmyhGjYjhsxDxzwHD
nU2klz3e4fFSuCVlmwt7x2Ff+zl2IgoHAJaodq0StWxSCUzdhaN6HfXqbWU1TIPgtiGv3c059S5W
LFeeXPZmz/2kYSUSQRQTYo3rzvofMoBhBiWz9NP4fILMPoNzr1+faI/KtRHIRGld81rKyDqqNl71
4Yd10WjfX0vJQ2CRe6g1e7yVcfTEye6hI7cbh7LpArfVWNLV/9tT6nL9OGqO5ad2aapSsSwrE0nR
Sw898TH14P6UBG3v3iqHlauQQqG9IyLYbpcvU07sPbK9xEUK1oysaNW9c4Z80OJ93sUmm6O5NM+w
hGdKOAJ4Tz2Izsp6HD5yUkzbo2KeUVIuvKuAqZkabAB5jCObCQTGkjOH4DzAf0qB1QIO9M8xZwX7
E9mHadAJ96X7PcuegkYGBgecDV0cmr1Oghwa2ft6VETJPnyImCdMwYbe6WnmCfZkMMUEGtXwcNoy
lk5SwwkSpQs1p2ciOERu4iZuhWnDIhW5WEZ9XMscFIbh4gD72c6ZS2gY2pb/q+pqe6pETSyQC6Hu
a2IEBK+r8WvPrFe0m8AF6hPOZn1VKJzQE7aBaCD8YigpjVkuP8CUnGHk6wYBAHPkdN40wvbhR4lh
frTKv5v90sTAyPeqgJhtHP9R3LlIwhVd/C+e6Lp4r6w1ANyukX5i30uihMTP5j4BlCeAwNpm4FD1
7K5jUFd/gB1q76VlJLBw2f8lXSW6zNm/ytsquI5E4SVXeaX1deD4nYUJOVbogGSAeOTTsDH0+GtY
IWYVXavAUIQlcK/CxqNDnlj6T/9yuVf3lsvKXZC4GzAcq+sYGjj3WFtjwKRVPsK8yD7YuFTtNYJ8
f5vpgiOrJDsm2qjhFD7Ekr9RlwMwuUR2hx/Xb4I07fgeLsTpm3gNQxKGukZBTkg9qndkzTCobiEw
MdFFpwU4bnNGH744Gxlf3D7ipgYHroy8yELgw/KczbTyCAGrsKrdpNTO7Xb8AP8aBMwECIljPo0+
2nslUgXfqSbLkvRgLv+lZnIO2U48bQ7zvHcsbuZRutTjYg8qs1epVu4YHao0r0ckOFnpDwS8BKOC
5kh3LoPJt09WQsu/SAVJF8dELMjkqgm/E/nVNF0bHOf1BgaCLulnqZNDkdZqIVs0px+TAk6a/U68
MhKeuagMXFagWX2jGBC+cbkmTcak2uvdasYOQn8wejxNNRn/e2Rl79n17+HSqmIKDxezyx566z58
OsuyWVtdJXS33pR0Oj7O8x2TxCEnULA9F0h5gufEH2Ua5D+CndIe5bn2GtifLCORxsKVHF4FwiOW
AtjUBfPENotd/ESnSZ2On7AyD8kAY3GFwZuT93E6XWHxANAIft0E5sGeXoScyb48Watfl6FoxIx3
yTQ+qK2F7n92hFugT5s7umiwYSK02DZo7Evof9mVr2Ya1UFi65aD7JezdzdYoo0cv/rDG7LV+8+c
mzydQkJd0Q+c0qQE/enGk7qO67n/UnrIceWD/tKapo0lDAKApgSTz4OIDpAooA9DGTVcKN1jj9b5
5NJCGmxrwJ6MKqb2Bdx/Uu6zz6M561FYnEE6buP+LP2uSHdjuxibeBO7I9e3u9sWtZKprP+AoMty
hPiDs+LQIg0px8QGU76PxImD2+qNGzOhvxXFeznSehEwW09iiKl7ymRkRd013nub4+ZLMWO2zhA9
FQ4p/S1EUVIKoQp6ozRq3fYRuT6P6jY8cYzivCUx2fZ3kk88hDipnZ3NHHpEww1SHO8dBFEuAmUV
z1I5bKDO5NqLiAAbN5u0ZabhXvbrOUqazk9kxJ23XgSOUrALMWiuKxEg5ljJIIgFiMowd7xnnBE/
xng8SQJcPGeOoFP6Y7FDqy0ASuwAwC2Votec+XXQxrD4ZxpzKQWk3h74atXnBkPSNCf2XAG1mph0
91yW7SEL+KaodHDBLIG+H5KhMoMJoAs+SMsUpzXhgYkRAxQq169CyO9Dgdd0lLuhdnXfwIAspKSM
SQG5j5ww2LB93hTbJNFa9WEsEooJHLy6FC4wBeUCRkJzdVcn/Q+OBeit2tVP+6nFlpEbNCl7/P/m
AGHMGY85woK2cJHaNJqGxKqywI2KpikkgfeCoBz/GQ8yntgszTWt8Ms4PihjytfYPpSNnp8HDzPt
XFE/2KZYnu955CYo3S0lJhyW85OzPe7RXSQwrYHz+ToyoHt0ygi1FvX6PlvshIY5r7CWswQP6Bk7
XU4KKdoi5RE9olJDt6LpkgalskHwuUdfa0tEOmvozOMCcyOx0pJqGkxLoLw3dD9i+72ova7xNWl5
zFHGcucjMbzuGBtEf81P5hSkOt82Y01/66m2hB/yEk5etQebinixyvoRCRmspnc1Xn+8881EnUyJ
Zxk52Zxhy1hqycQY2sdaF+e7DrgEN9tyyeEWTKvLKBGwJkNy6KfQBCvEGO1qvB65PhW931DEB077
6wxNyx+hQGLLJVW7ieRRZqSXnQiGfZ4t6hLLjdoesIufVnT2MdIwJ3zTEzy8bixGL0YO1rFYYuvL
vgiC+TnCRgPK2eLCAjIyYHEjE4raB/IUZBX0gMT+UdTzFUP5gzopFo1IDLECcDrX1iQAuRgfelcN
VAU9cQ++iX1/azhwIpYO3XaVG45UsIJ0pjYo5wuLeMMFLgd+Dce7B4f5QdXWcWR7m4xBkA7bkhYQ
ntjzufrlDfKcDfq3M94ivxwQtmkRBuEWcqYUxfFftE9blrN8GcgCrOyC6uyf8OO90gXzK+Kh+UaX
OPOo7DqKYLOLqmhnfzvrH0yLhPBTA3sQTuJ8EXB24RGHObIm3YZo2K8JxO72QRC+xi109hFRGDU3
vNkuXAn2OP4/spLXlbOq1qDBRLV++gK5qk4fI6L1UAdpjhndXVQfi6q4D5vZOMmpgolATM1NYf6a
fTUM0RS2oCxp2CmM7Xr/leFZ4/SRPAwU3NyUQz4gg7eTmuYtbhl2evgORnKMCVlJEGe1nwACKPn4
qgUh+vh3IIrtoam9mCu/qHhI7zx+CSHHS4Pu9eZff+xsTrkxFqzBkycb90TyeEVQjkqhYAySyFw5
LwWxdeepNP4mQhaxv9kUHBOUHT+0BTpELL5aPjBx2kAqrk4b11p6Z3/yiIyS/IljS01hGGIA7mDB
ecmlx7E0VWE0+RwVhiNw421HFrSOeHcy5vWit54fptqjiGYxi9NHzpawtTAzU29co3vfcTiVMpkS
vaDNc+dTjy1XFEr+INGetLzPMU3G051/uXyitw/zbjOl9Er6s//IsemQ1kOqi1fdqwnogEa0xCEI
mHGcfzIYCcpp2+iLUZw/JCz9SYBJvmkm2F17+Rm7gHrUozPHIBW4+g4U5ImEIVO3rAOGaFtbZ1ms
7EzPxvQMoY5AD4jMWaeTOUugShijhBcCwsuaKyx+fCTaNrtEtW/o0vxACSa2/OQozvanuPszmtRM
8d5cBqELo9oaQCW5DOwjjI+zSDpJogtJ9G71qQzcIIkAMmNwZDUeHmD/+DkOm4u8LvPnvRaN5as8
eOAzKIo3dSJ96eVEiYIpSVezkRgE8jUxqiR50T2jGaKM8HVY4elCv0uyYcm1W6lXhAG3G2nxI8MC
S35XmnMiFwcKuPDEJxpEaxlN+iRo/gi8QJ8cVjLqDNdoF/IjUYphG8j7674Z4a9kpaGj/RYBl6TY
QPGa2wI1uar1vPrsjHe/isSOZmMTRFUTyxRrAIIG8p/g10EAJq1E8KKR7bNupWjsWmX5z5/eDOPi
HFZb+CdLx3Qoakl8WW2qiG0kmWERiwa0ILT0r0UjK90rAy1yQMmMDdpDyomlrv3uzecEUcLNE+Jf
bWoa6t9O0P6QnyHguaSe6akQAf+JcsRskopEYtt7DvLT/n/DilKOfDr43wLw2CfamLwEzBy5H1DC
LIP/C5zlrl4ZTgVSssYpJMWFXTfShiEiSYh/O9arT+oFDECgTuBzjZuOabT1hUAx1rZwadaRoAFd
BqWdIOuvCfgr8FHszLXQznl1/dGiQj45TlEfWbL8ECCZkHrj9pRiNH6CUqsiRyehEaYluRNuXUpd
SU1U9KuxANuOLOC6BvoqEdWakwvX1ixNrqH600IxaLrWKweoUv6K6Nvlk2dfvmmRnkgSdGBs8Knm
1agpTe1unLR21VVq/kV8FIRizq9ZkN+WacEmqIdw4EcAJY/BOUR8Y26KCSSHgfoJbbY+/pubwHa0
hpcUTUQ9Zm8zNwdJnKvXFT5XlvIhBPQ0gOnp1vtyb8BQBUwrX/ELlnm8pemv+xXRaFIjRh+j8Myd
YRW9RIEI++O3tfYlj+xdpkyIcJXyl46EaSd9PFykFPj3quVZUY05V+EReBWHIiuxMFBs+qJtmHrx
RY+JZsRfwTcimMNjd9J+viWILbEfxcJfRjtkhW90d48+dhFlc4cYvbwVoONG4M7ymR41pPYPOO0g
Bp/jXocQ2s2H/k961kQ3aKFsgfLf5G4BnyRJk3GaluWTcoCRSh6ebVlReJIGlxFZ2xsBBu8SXqtj
XwtMLuHskJJwAmZ3DnZ+1QdXfBy9cTlETntPkcewREBKsELhN/G25pof7AFmiVNhAGf+pRPMzilU
F7zf23zFOkky9QS3zMn7xGAxLt8WsIKuLUk1T+ES/f46z2yZhePHoGEIZt38UtwH+xgIRDuE4g2j
sOAg8AltBy8S6be0Mgo7Ym8tFoN3X6+6eLwK/V+bJ9/XI+sYLVIneRVnLyk/vneIZcM/bdL64ziv
IwIhriqcbYUO8zs4uPKpxalqcuH8hq2BPyc2gpiCYhfg6Mewen2sLfMpHQQGZLD3i+/t6u0hzNE1
qk5ugpt3ugfzDZtyLeWxn5IFSs1XUjhMRWYCdirS7tLVIXazID2Qs7pgeNoAeNJN2qkex3z/noVs
csqKGvXlczCY0Tcv14gKHcb6Tx2em26gqKAU6ajmyc94OI+tTvMCXXYUrGWpIiS3e9dgjw2XuVm2
NDzd/cZ0L4EPDHnky1fVVP4YVGPA2uVYjLA5KDui290LXgAWWGYFG2qum/n7wQ6I4UrdvsdMkcu6
bCb5NmMgt7WUOY2fS+YaOGjk37EVu9o99TwtPA4Z1tkcYHy1Vamke3sFg2zHUGT9dBOVX6uHeutA
OXGSb6JjNowX6S5/U3pPA10LIbZk9+i0yCh6diJwsm4mtOrOIHy+r3YaxnBHvMcOk2jXBmUUYa90
Ruqgv9L/xzkVynK1AK58FpavtHd9vkpkSvKUbiS7botrfIbaq4gRmpW/tlc5rGG8LTRdVt5/8wGU
AssuVPoMiE6JtGYLFJ2iYxfAcKI3WwZYW0KlqQ8SEU1bfev3TTJ3CCw4XMxOTPVVjlmTbNjMUS/8
0NvewYe96sYJOoCidbC1fDoItEt50tQtWtFnLFbGnXX4F6gU+hllqhBgfFWC9UWbqsazavTtBgfp
FSskdxkpHrZQ3R3NtYcM8FqYNHuQgTquV0k9T/tBucvCVABUr3y5pvGeL1acBw1oDedgAP9U6gnN
GmkHM9PsfVcnAODwLEiYxM8zRhk/JvN8tcwq7Nmvb56G4xrNDVKex40lPD54CqbpYeXxLylEmAUA
KZKuhnNT7K2OlDolWXtBLdug/rwtpsyUk7tSBj3YXR0q2fYw7mUeyImL+vN8AUFuOwd7d60HcSbr
RSpa7+EXoUaNMjODIB/GdRTiFvBc6zcYg2yao4hMipTnyZFdTJnBV5YtH7yG+38cpDnfjuVLkfWJ
GyJZ6mlWeHlaNNjjBHbsnVXf1LBl4j1TRgW8vOw1ra+Woq2kYnO4DVS9HdVr/zhJY7v6C6B6zJXU
NyJA6FXSp4OpLZNeaR1q8xDo2pryiVUFONRHdV+NxkACj96uULOnS7rgcaPLOeQgHz3TOcjxcUa5
OLbJS2iqwhJDp2P03DpDsnqSRxnbtOlqp37/lQ==
`protect end_protected
