`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SOYVpLO4bquFSzdYRRoFUJR6R1VGHI2ZHnJXFJeeBsuoDRBfdXEWHORahW4A0rWgjN8aMxqnK26G
ZRLY3P3SMg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dNa+su0lFKlpb3yzn/MeCLuMa1m2nviQqs6wDH2vpYr8aseY5omDbRfqTey4y4neerZiDBU/I+oi
EJWIIj5x0QAmR21pyVBdoG5HGcdYghrQk1ER3FOkyb5E1kSGx8taYfs++jHGNZx+BMIlOXX33k8I
esAqtU7bjUww9e//E1c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hOtq1t0vzh6ioERKB13p5svtBYs1T9WkbLbHtv60aM1RhdzL9DaXckQtYSPyG2bpGqMgwQ4guxt+
yzSekaMVPVGG2xSbzXkjOx0L1PK4tgy72Sc3uO7Adnx7Syb8yPtrQZU018ba/GqYHKbgmA3RxMaK
LYxQ3MfWvwzu72QliyVY9x21lmsaCLK7qRIX1lC8LQKpwBL3jZbcEl/VkNGdt2RC9wBfHOz5v/WJ
WP+X8UkkVqRN+j0L+bDtPermjSsP7k/KToPqOMioeL8QeH2H5DbtlR7Aw6hCK81tdcOXtKwyYcnF
7uBOxJjkFwZZ1VUTGtstTiUu6Mhjo94EEgfc4A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mLq/sLLAWOJLJ6eqKJGMMoZypYneRQpmi8SD0LfVC7FuoVWq0qj+ord9MslpzRQaKBHqHXXtK0ZL
8LHVkuowCb7LckiOTeZ1z4hHYAkSC98b+sIH35GlLpY6GK/LEz4kjmLQTgYuLs6ce8aZpbaQl6Zw
ocUb/yBYwP6SS9z4Oeg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eZBT+C/pu9ER2iL3EzIRmJYdWLYV1InlOdV548JBQv5AE0qovtprWT0gQ4dME3Jnh3sPAZNgKSk6
EJTUEGlaILX9ud03JCFJTvCeylo0P/3rZ/xjqsepu1/+6laGC64ZLwZ30/u7dS49q7G6ZQ4SWs3Y
v7IvZnT5u2KxPJcOyV2EJtfAqNmZu2Y8CFs8ZJXw2jFwTM5x8E+U33QnaJ2RSIFL5Xk3bGlX0vDk
WHuN6xMEvnUaMFqpNjesChxUqWXc7UlGg8Pqkw6QjSa+WCsAxa3qpNrSW6t8HLLgZrTYruAjO7Fu
TaToDEJrCrpUesNciqaJXiWD7TaWQyU9B6jA9g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
f2EOJO+2G8kQ/UxBY7TFfEQE9sfbdpTGAqtjOReNFOPxGANIBBKOVp/g+0kGq2oYqofJFR2bmOM5
zgpygDH6Stqb2CV7spMnwHSaQVIUHOFh3AVs3pKgpsKBX/FfAz5A/C7e3pFJrHfb5CLOy/wOCC9E
TomOZ4Y2TJvssfXLD+DTgUrBJ1UoV9BoiPBrck304S3kFolhUTfrpoui7EX19Qd9g/VLWuNNat1Q
xDhFGiRDj8bQymh5+QziSSyyVZdAXu0Q+7ccD4/+Tp8YmXoz/qve7udGiYWrjFf+ZJWn+fbVmR1e
mPXIoGb4npaCV+QdTbZf1ia4GXVaJuVO6BDHk5UvR6TV/yDg7gSGWRGKSE5G0K01T9eFosmHS7Ga
7N6fo9KRFyuSewy60P0qfIzaOVT01b5Hy5eCzFg6aqiHafnKqsjN8uAZICqkwYDx5bIGbvtYtUo5
ZdiO+CQ/E/KdlkWElSDbGusesR+/DN7xqdby+qRsPoOGgnvH5aMXr5vNdQFWGa1W8TOAcO5zbonI
CaUZBiYIBvR3leddWT5OYZgZknbWnUe1PQ6WPasNYBOjgRgLkRSp7bAYzAC8oTi3cSqSf4uKL/WP
msORC9hO52Q7vdKPwtXzKt0RQN0OG94uSBSBK6OGtD5RxlWBPw4lqXVrFsF6vXi3BtmpWVNLoFv7
lm51+1+YNxgmOHbyOhNZodxNLQfvch8PnOFsDB6wTdi7ML22UzLsiEzL8+4X4dA1iURrDlAnBXPV
mn1aLz9hXAsWGygPiGJKJW7SkAe5szVqONVQuRywymsEbNzaXP4EBZ52oWqpskYSZroQ9P6s429n
8a1cWFz3RJOFJwPp5penBjpatN6RWRP1rBkjRs7xfmnD6lkHrkflDjZmHCxmPh/l0Mq8WKGXgDLD
+c1dNS1jWJTRNH67uc1xHWB96kEYYr3HEdWUAYSfWwgvOg1I0yvaHbOSBRxpFWl+KGyp5PaZ6nMl
yiMHaTcz7TXsS2L+aQXSRNWFJRg6KIMxJaEwmK7jtk4Nd13nwHFyCXdj/SOqsrwJVxQan26JZcTa
3W8Lmj4bh4yVDF/qANzuwqEgLK8G1HjjDScwECBLtbg/Z4cyR+1vsVrdsSTZfgfC189hnGMZNc1Y
BgsIK0BhnGHSmdY8OP93VL/by/GuqntHem03gL5nUs6GSX0L9nttJTjea78WKSofPjEEqoa8McLh
gCesouDAsr7DKIuWGNP7ZG0+f871IKWn8/2SDHh349pUBLT/1TN4gQkNVMavXGbGV/kO4d5fuKnZ
ybzUyoJFKAgWyFldEzVVE/PNyQFv08LlOFKOGb8u+jeQ8GrBzBzHSq72LMNLVRy3Zi6FcCs9l9Fd
zBa5t3AUUGeoud5KEX/CjMAo1LlHDGVKtpmX+cP6we02ALC9A7fiItBUCVtAQJ59dDE5SaZLWBFJ
UpZlq1Rk9ZPby6clGTIb+Ukcnxr66Amn4Hx+8NsiU2EYN9AleBkD3Drksvxm0ILd8yZd/MQd/Zef
QkVZr0lq9tUkQlrfv9AL/eT9pVnyxXLq7oYbQ0P7TsrSN9GbsrE6XFLpnEgTmat8/ex3pLDa//0R
OE3nlBwTrZmXzMVMMAaElClRUwGq7SrHrlM6ynl9sbOFuBuvUktPiU2pHDq9JEgke8JJJ+qBmexD
rc0JJsv39ZARR7GtPxi4uryE+ar+lagrg7Cp9EH+55opeubmZC0aTQ1lRlcmL0uk3mEcqg4i3A7e
6+GT8MoVJ3hkDv/0AM7q1JvE35F/Pm50aw20Xmhap8/Wf71Y4+k3pcv7PTF619lhmF+d/9NOjyiA
4cXp3ZsjNwmKII87Wj26esWzatXsHOES3J5Gb/tasqFR1CBmLRLQRpI0vhnQ7U62eP3taNv8fhNC
Ph1wZrEaa4PYMtkmICWfhiKRXh5sDWBB7K2wUl5IVorUuxeFzU/ZzbyG25I9In8XLMqeGYq7RtVB
50cPVX9l2+RWl4A9FfpviKm8uXRzTidqsqD6NL1upjP4lPOWl2V1KdkMZ5KzkIKVBfTl4iUNqPl4
yJQdA3L8zk96OskOfVqT8vVlmlllwoAzq2XTNVrVbbrSHzPI7n1HdrTI/9rWM2112qtvd2sQs9/0
evIso6cYwrY2rag0OSAc46iayr8lZGl8EI+LzvLk008uo+Yq60nEi/jDXmEeQr9W7r1BnAzqP0H2
AMItYT8udCR4uX0o2dBt/dHbC/lgWnsNRB1vY72udrS860UEj1LkX2MeDQJ8YBjSPlBp8M5t2Li4
pMGNAsFGEYiG8lsIKWUFG2+oES3dh4VJSWw6KIuKQZpxmcLfRZcBVfWSDMhO9ihvK/Zc3B4jQ7GO
1yicdZusY+3V8LH8/l9IHsNxOt4SLgYu+G/00Tbc0UIEQwYI73sWTVo0yqDqrvPgl5wyMYu6899P
+61rLb+W/srNww2Zk3AW+owwa0iGw/WFvFY5LeR3isnoQSTuxfgmd0Jn95xZzQW+crdQqqooVLCe
Fj874sILLHavLcz2W+4UNgiVi6AbQa2WjG8tI8HTo9CsJ2+0RS03X05GThOPHgLDJS2WCtB7/noO
LAM+i/KEuEKr+8wnB5i1M7CSHFMwtCi+t1HFfUnnpnZ25SD8SEi031mY55Vhf9fs84GKNTEObRhh
M+q/K1NNnhbJiY/Ndl/eW4ddcTumGQgHjG+wBRduOQnOp+j7XYk9u/ARaA/uJ5kuZAJNKh2uTM++
jcJ7wm78RjYqBGPoA8LTBvMD1YP/SAWkUBPU5MZ6H6226+8jpUVxP/+lra3djswXVY+b61jjHkAF
/SVVw2WfQhOlA0sXMGVRXO6ruV3bHeyLYdf1s4KaS68lbDi8nhDbaB4MAAP9y52eTe+w+u2qS5jG
lDFra+hjQvO25vMQx7rxsRf//eGv9Cpf3BX9QtbACzdc0cY6ixUsPGzgUS9sjc2DLXi1Zye61k9+
LuFECJFUrL1stiXnnt/nSCs3pf1JZzurb8bTH6Z/59aVmSnVChUGjgICAeIiu6UqZ+8yH2Hu5Ydb
kPBPXScGiHgk3zhPc2v9pJ7LAWyKZqRcI1IcjF+KF6IKNbE7KSVelbrHCsq8s/p8jWeFbJ8yRVtk
Gzw++bFWaoLsRuzz5zr3n0upbfLs0iAgGTGA1YqpO5vmaCpkeV8QRDYpeYfjFaQARZSNactFZRxQ
Brrfdr63SU4z+i3L2QqxrqY4zhoK9uOiWomqXB5jW0eSg2JAPQEg2T9PSos/yYWLo6uwFYZTFFSB
dMtswUNGPLe2VGViZLv/V4vjfksm+Nt3N8oezq2YR53Hj7bdo1R/Qe9xZYPiNvr/GCskFUFsm46O
uayVk5qQjSNPv3X1VZG9lwChD+b+w+ROWyKm7ruE6bor5FyuP/H3IPGvQMbveB1hd3QiZ5UFpF5V
W9TncgJ2vbwVuoRWgBmyBkV7GSxhwlk8CUJluGbkYwq7wabnlpXoKLy+blQwQh0xIIUfd/poHWeg
KGW7Osc/l3OeEsrv4kcsvtNV4uEqr03/BGh0vEnwpROuDxHqqgftdDZ7nHx1CisvbIKHVYZhEQeW
4NGvTatEt6YfvRktjSOD6/PvS+2yjhfkdTwMEd2Lrin+0rD5zvCktugqzqUtrBRmaHSwI0qn0X+p
ynf/hC5W85snlwfYH8QVtwdQYtNbVyhD3uSVLoDx5rBnEWrYxqbERdDpRck7RMhg0uCi3nQnK3SJ
z+6oumKRZZnET0Truw26VtkbVnRryQVC1NJqOehO6plRxN+WxIdD4p09c3fFimfF+3QVn8/NBlo6
vYuJABDZ0wSPbWbWMRy6irYs8113zNIKZp5e9SAGIi/4Tg6SMBLG0qprCJPsuKFZsNWR1Tg2hdfx
PhwSDwhzd/1w3zGwPi1kc6ikLM5jNIRMBa7ddWPSWKVvJRnw7EABQIhqIHoGg3Vv95XYcFgPHjQs
2AwmxS19fW1y1X7SHfcRnB7Ue7ReXPWQnYvGN1yKZcXgSoI8G44/aQgHeQXWc+5kKXleboVCbVJL
sUM7FgA5mf4ciaXfzHByC6WXLU6vGmZKoNUvVIS3JltyuUdyNanrIUhIfDrCGmhL5EU0DLwS+vKG
S0VdxMjn7rHyz2YYh4rB5OvYZRPQeeg74knsBZ31Ie5BzbS/BOuPok9aiZRNpvsxItR693WY20kW
er2Wdl3twHNp3lgmNkfgF6XOU53AIiVZ59+8nMvOZ/u27BzJf/G7rjrsRx1mZxdsJwV/JUBGpS54
LR70VE+HGNug5DKfnCWCs++jqIagowXk4NVd6gWlOvt6e/CytYLJk7ug8NlZ8VFGh9p//bovvdlN
rvQgoCJjH17UVkP8hV3C/U2ur3ygZA5QpUivW6u5mZAcVvwN37zTL4SSRKyqcmtUX9bUysnS0pnc
Dz/KMKex1bdd3NAut+W1HJYj71MVjqdubh3oI7kQf3q65TmKhBfkIYr++/P+hKxXwIzbJ+joE3+g
OeSLhV3USebcQMxULIJx3WZviJGsEKDkPPfRV+ftysC5qtqoe3QiCp3AUnhNRoVbdptGxg3PWHsO
3ahHAoNbtpJsw1ikeyeAZRu1sNP4Sm6Jp3atJYGuM3ticPOgew2dZvhyFjPGEi9wMMIapWcs4ICN
ZzLaSh4DhS2QONeWWI1ECQmDBMXy8qmtO+0ls3wdjTGhwGYdyCBNZgniDuJR72Pky4Rreoa5P5PN
zPg3mMGN4s8xiqSCfrXuvXSEWJz6kg7enY7ykMoQwO5FFNl/XnTJcth/yFPikeY8kbv0M/fMqFlc
/icQAWna8gBbq5osO3X6AbhYhSjYQh9pWO87ianL50cu8uB6MxseM+0M7y7Abqxo8Ruzvm5IWnxg
Zm1+QUetMW7EbJb/svouhQmC9Y7bFhstSEsXcB18GKi19of8vxaYNIZ0g/6CX2ekyfPAKMJWk6P6
mjI1ibiYPailOTFzHj8vq+1q74H3GY1dln+xb1LIXHHYlM52Nnq+P7JVGHKGzPyl66f39IYjqV5j
/wYcBzCYiP8iGmzZEqj4hVSPKmSKK9dKecC0V+OKkvBKOd9LYhySOsEGxTZ14h6LHc76PQJW9E4F
4+Q/GsI6yc7YumH5JFWL5lH27zqx2Vu+k7HdtvBB16lBEX42UN6QFAFyLvKHyNfXAqZ2/faYimVh
d904jBAjiznnXaXIYoWEHa9I3vHk0Xv85leVB+3tDAI2SURv61SEetSZUfWFooqYU7vzl9g6yKNQ
8h5F/uAwVrHs0IL6khptORK4js09lLPMgVM2tqCRsYDDtRm+7xbMwXfJ6EKTq0dKVTXdrOmIvWYq
8T/E52i2+Cfez5WYA9P6EYC2kCBYLwRq/0ypsMQzPwQPJBjaeVkEGLC0VzCQ0Uwmkdcp1TTO0Odd
+TVua8v4og9rxe5N/V0/CP207Ba6JkqlXAGKSoq129dE1zOCf3HezfBDgjOUOlQw2SZV0DA+Irn/
rdMvpYnRQujtwCNunBGBtZ15Iqfbf1Sk6Kf5aO+phTXav4k794u33W7OoRlSxf/FtHtnr2D3TdqN
nU/JzqiGaKjpH4WL/P49bNtRDyS7skpGqaJboyEO6NF+ZevMfOqjQhekiTITbU3zmPi99/T/EgRf
CszTqn43HMi20z/qmjWCde5AQg5nIVAW/HVnhLYpbOPDX9252jidlzGBYM/SU+bVd3cZMlXqFSkF
zlElPzc+OpyJckZCsJdT9U6mOK8HC2XVJiHgqNnhYZAGw8Z2Bsfwd/4wsHtFwKlTpqWHRKtYvN4T
OGB2Z7p76uDxKtjzVs/mYAdg7vA3LjgowA5Zx76gA5m1LmSJEzr0a/f0OCwApJMtHw19RP/D0Ehe
azLUKqDSofX69ZI4OEJ8GpQjpFUL1YqXekoIWBWZX5ogSKR0GiNwKJmLDfcCznUIGVqrJpQhljHG
RpbLdc/Md1b1NGyFqahdbCQpPDoYdxE+pntPGtD0KR2iNn79RRkVg0kvkC8BGXOvsSek7S69HQP+
ZlKOwO4Pj5DfcA3FvtXc3W420TAicx7a2wbUq/mHwk99HWcaePNZ3d2p8JY7koOfelMVi7eYB46k
BzNv97Ik1bgoRcEbY7s43JqPafKbruKq4huDUaMvKkFZV+tcmZz1lTTVxj7xyvj6lR2XCcVFJpuI
gU8tfuLY1BAGhfl4xJvwTeF/HWI38fpZ2YnRx3g/1ibevXjvkxHvVA3Yk5OiooWFdwmsZIxp0CWM
ZX5orpJ9/EbKd9bjkzT3gqyrN+1jF4GDjj2m4T7ye9P07bRD1CoMssQ/asXkuOviXzlQwpKpOzUW
cLTOk2V0ad6tyLVdjAgmmD8BR/11Oq43AXx6LZAkKJ7SnMfg2tUxOojrNtWCLAayzvVU/BMMg4Qw
hMnI5CvjADM8r4Z7DFx5Y8HUW5O6KJOwlR5zq2+vRNWp2iu1fYcNF1UQAhwhJx1jnr5IYGOyDe74
wE9N2VgDx8rTjov+qVko95OWhryzic/NmBaG13taKbi9fwTznrSI+jWO0iuONPMiSNDPnFyzxRf9
u53Vdvtiv2Fpd40fhDnh2O+hovJKTE2FCeUvCfGsHuyjaWsPSBZhamVruk5koKF2vZvRerh0vQyu
gAuDf+9oq+FkvmGhQiX1leYEr30ZHC3KqaaVHnizlNputI4OTrkEQ+8KI4++HIdo/FnNXELHhrpZ
xnhPpJ3UJM0xJwd2FneBwM0pqk3Le7U2Fx10jUa+UDRyvJToKURyEqXQBeH4UdMX64aUDadFOb+U
Y84AhVjOfa2lbUN+x85bmULac819DjCwKE+sgBX9GHWTHRrCpq2AawPIyALehk/eWjwJmr00PKAE
83zxvuuYthre7DCS1oCqNTBVRfgPwQBeXn4N496bJ6bjFhrwWjfA9+0KXubKCn5L6IPIDfnRM22u
IXSR8Dvhz7eRCYkWtWY731ScHyvrWB7yUQOnP7qZY7b9u+rdFrudLgQo/stpe9lhPzUCqRtLxe5H
EFH5yrnXaZs9S8maM61iAOWg95T77nkouGph9PfEtOqkfQ4fPAM8zp2BVvviurkUk9v70lmFgk1X
Zk3/OxCb7q62kuEWGNjbX8q0mk8I829LRUwU
`protect end_protected
