`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fOPvHkkMeoG2YSxpdCiiaIsa6OukwnK1nUpGs+ws1Kzx3puslJ7iKn9T5myI9VkVUgRFFN1Xfit5
dX6F014IGg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HgNCPi3QHpb8dW9RkjxoUGM5YOGOMgLiuLQefgSbCuez4Gs1lAiQxdxBQhTyXNRS4H89tPbEkHbH
4Kggyvl0Af9heeHWsTafUvqQuQWNgivzOk2qQ1liLSXiEJl1Fyiq4YsawJBYE511/GABOu1E9kTU
pmHAixKjBq9m5/peLok=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ACyuBPaQ3cHp5s6xGUvo899vJ+G/MHO3F7Xaj7MR44qEHb8iz7UONlim1fw/l+q+pLsNBpoVE2XP
zJRxKhGGODnlablcYtB85txWJY2O5wNxUYSePEkcSvh0aNjf+cMEMsQNe2HL2rZ4QpuBDEvwlv9s
WW2rOSkOtnkb96LcOQBvhFfaOnMJ1hyH3fZjN7kEzqhyOzx1lZ7F40vGA4At8E6hirc5xMjqdEgS
nhipIIHTzkenqLhApVGgUbafRQbG8ESyjA01uFRtZ25J8+Pr4cs+tPGobm0XSO8t3XwLVZapRDY7
SXW1qYkISFEa6NBGxO81MTbzFuTQYdh3r/X0qg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JF/XJkMGoJfUihOS9R76tudD+YiVNpy3w5hfoZ0y9FCS+pWh3V2jVVw5cst7125I/hGyQ4cnB2Cm
MpdAa/YBtj6yK0ds1YeuSU2Cxzm0w9QZ3nLSon/2jE9kx1d54bisjxRhEcKKKTSHuw6W+FSHffj0
JOZyc8RfIJ5IeOr+rqo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T1BVKuyJOlWV6bcI3uYrVButOZWbfA/40bEMumgKuFASXUB5EUZZP2K7kyzSOvm86sj9UL9ICrc7
AvTcJqoQYQhmFnASRJLODgvNhDHbAg2lnzfWs6NJAS/1X+/rmymQ74dE/PCMYJ57I9d++M5vjskf
w0OpYjhlBVYSir/Tk9MztjSWYD+sQILHVjHe47WzcVPfaW+EotqO6HFgKqlaDo7HehG2c2e3vqSf
vOR+wJbW5Wf5aDiFmC5wYka9JsKtHRwx6zm2OF25VJgE3xTsK+bAIDPdQfmE1j88uDe5XhfBnRre
CJ9sWYXEWxeZpiUuR8hxlglo6dezNGJESHO9ow==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
XOWtDNZRv4FbcK5HgglDAnuoXeeEtQzM+5dwtbTltQeOcgiGL0ldThovapKXwlYS6j3SjEpt1ctW
l0HJEu5CZQbd72e/yXjziCbCs84D4Hl2Vork8+ulXUTominLbvkE4YkL+H3FyGOZakEzvv3vHoQi
bGRSzkjeHwbXiPYH59tq7tQeJMQxgUe+oj3vs74AkG1R9+2YXPdoq+c0ike49CI+BgwG1ugOKpIs
VgL02xZMnagJKOXiUgf6pQ6HJDu7a4cb6y+rbPzvCZD3U39xEI3Y25hhH1UhPljfkI5NOn8Vu/l1
pd47R931h0LHGQ9zMdTwFILbWSSgIXW+Ww2X6UYKBg6+XDIGfN9yLUc0j67yNx93C6w7mxcdUnEf
d5XBmYrPp9/EcMoTf0aob/1TYF6e3buFL344aO7XizDEZRYc7KG+GUeDaZr1RZaf39ICNvcxuUup
fPl6qYVf8bE9LBoHxQs5BKNxGe0s69ylsGwN9ne9Mu/voJBkPMqFF2/pXAkTAXy5CiAyNLz2D4Qj
Kj4V0wZXh6DUewkdBgOgMdnG4/SHl1hzGU1DdVr1bgJrunH3p4DNx7ETzJJKPsKmU685dPc30nwz
G1ysAPjxF4rsT7ysCwcKpFB5BSTTWnol85/tmFsSpvgHZbfkKPGr9PEQFg0S+Nth2MZL9N1sC+eV
I65XtorUCbUU6VD3zsuk5T9ykchUyiijID+xcwuAAaH6QhEosv3sG3+v4M9FbpyXXU2dv+3hmD+Q
3qI1UDa8udQd8CyVOIu/DMs7GWf+DfuY5Neb07hYJcNC12Web7v6KPXVxOxGkE1kdqsK564hww9I
7if5qaA3BuMtfL3+lBhZn5GKYywMy60g2SdSoxO5GNEuBLToM97ulyb91wYTxuvvcJ1nyjBVlC90
mSw7nXfXJjhsbDlqix6aaMoQ5mq6WniCyO3s28BGiKiKbeuQhEmN97BgNY4qvZ3ZxA+oM8ipbDzv
OypQL+vvEilICjXzp7hJBlgb4Cd1aCebECNJrqe/AMHC4+pHwAd7aC9eMinjkl0PDhteljDSS4SH
SI0sNHQr6d0Jhzp4UrvhRDvfJ9nxbh/F6dtS/msNc+vgGt8T0wmN48DxMu93EAv6wTDclbebzZFe
iYRCgpUN+wPNk1rZQ6OWwU4Q2uE51AjSfHdzUotLRFgcfVYCKBHfqqt1xlPe15VS1bRsW2tteYvo
a8vf1a62LKECyibR5UbX0qp5OwFpQDxVEu7qWqv9DpXrjTpTPEnCw/er6wej0h9FGgxxiUC48PKt
t5PRY2pjB6y6ZEO/wrO3MUfjlx0pLCSBOOfRrNwzJ2g20gkUckYsJhph8I8mBaprd6qd03rmM+H6
sZ1QapOO1+AgxxoWxm/JtLO4v87aI/k7apNcMnb3rtdyX+nQlkDh/zy/F27S7SK+sxIXnYkiVjHU
0c1Tz3ay5xtmN9oMRWyPcehQ+AtIS/aGm5mQxSTRqgGTlNmmXdUm7uwmk0LMAJMx9IEVKD/T4G/e
VkFj1wXaHBAjrtCIsk4mpe4/9OLRtRTG8931GbjC7aEGAFl49pXz+gEjSXfgR7jKMASaaHekT0Lf
VmubPldiz1uvAREwZStCTrNJ14kjJew2u6c/gzrPyRT7hLC8HmeJ22Cndh+eMAluZ3QjydEftzRl
6/swDB4j2FO6r9VquZv92LAKPVJyjPzR6/grSYjVkPbydBSE2qSkJW15/+UtzZWdDqgFKIUDi3MF
WV80epAX0xaeQfJSwpx6bP0Ag8srHZhkfU+taAeA2JjCKfeyErzjt4fwajeMkrb+v6rTZqxZzovX
flE/bvBh7zd5Hskf/4gONrf2kiudfSC8AqaVFxEXDwg1zvtUTwiOunUBT78AehfyhdJuv/e5xY4k
L6VuYh3esIUF3ovizq2tAX/P3X0pgcgynUvLg1ctVuJKtgPHFs8vbCssvzK672RmPwALLBmR5uxy
fNuRI7fWrXHd70jRFTnsQk/HEyuNyTQSDly2+AfxaQBNohUiWtZnKDqfAAy4feRld2qMQyPediJb
a3r38TDceZ6AZNVhrpp/JrwZHbLR1zzBbkGL8BvLerH3VpGSRsZDmTOmw2+QRYQ9IlnPbNUAWBHi
IxQXruHEObmJWgW7PRh+5qxIocXp9CZqjojH/49FnYhpbKVNQqVb0gnRtdyDz/nCusx/6WsjhECw
pteSfnlYktSikI9/pRx0jEc/APbMNAwm1xHQzemGr0L/EC1m3m90wvcT7RBsEZlK6juw8QmMraoW
l9ywXqdDXM7Pg8z8eSMiavXwmG7BPjFM5bcsr6ys/8raseJyod+8DRNSbRVLBMC+x1YrqEZBwnGr
BuQ5FCnaCcl+NV/i8bIE4GCeSX0TO0z8GE+2vEfD6a3vN50uDN/0pOuyft4JxTshOCiTaDOT9cTK
rMfsE9EGPuPUUfmss7tV45kYpD6MoYo6z/+7Ry5lcWcAwffYgxPD4K9BXBurqWafRoWP2l/+FSEQ
V/hR3oiEHA7U3nvfM+NZCXR9pkKoH9ELa4D41lo435K9b4GK69JWNX8VDg87AOmjGLHh7SRlddfr
En/wyvAS9aWef7b7diP9yLE5TQS2kVI7SlMBnvwJaXkSYLwMn9wnfpo5JhosST1yRkqHbgTB0gP4
mE0prXfcH/Myaf1KJFwdxXeIHCOp+eEyuXUgyemHz5wpwY6xrEJrd194Ew8tdENtoTXi9cfpQURr
O5m7wA6I7ZQdifuT4d1NftZYNxu4fTB6P8j39JJpO0aaf4ByNs0KpySlCG9n/Mah8hzV+zq78tTt
fdhAnZpTDEqolldjTIGsvJ0AudF35IGFvmA9myx76yXqXo7DZzaX2MghZ0eBnxzdNeojGuvL658w
WyEi1jjwZqUnzjhY6j1EhaoDRXID0IL6kjlImg5/YdUvU+KkaqhrwA4mvrbUVsXFuWUBiYymIT8u
ZR72/bSZ2qHIj8CCBvJ86gUNhkW32fwivTDIhUbEqVMtsy0sbpE6fHF+AZqieahom+MEXUbCBFYB
8rJfKF78d9GDHzrihX6cerqy5UKsuMDSle++UYgB/1HS+6hm07PjEATky/704K6x1LxyPII2d4Nh
HTO0znYLeAJITj6X1zXFBLRxz/7JK7PAgPuH5N6hrfA7ZgH+q8VHdKgdS/c40obQLdFKTuI3AAud
2NltlIMYtdAkPBXf8U6iQkucHZ7orFA6XnpsBUn9oY42x6a1mFZJgxB9igPiKvmqsveCtojdMefY
2SibinbNAXb84FGbpehLb2PHZgD4pUe+Zhtvk2qWyHnsMRbDzaiDhnwPmHdXJ1zinBCvhJn95gre
EE1L5i7hlB1a7Z3Lndas2Dff2v1Ylq1f3779VnPSdWh4gm3eRwasiwpx+wQpWIMHefNZ3ZFi3j9S
yAJk+gdQT5iBsYHod3H9fc/o7oaXPdU9T9bqAhPpIUwWg9k9Nqwx03nWngl85fwsez5rvKsAMtcY
94oas6UDFJ3qfcEdxSu9ZY5e4XS8K5puZm35BnSWjLL7DNR60HoLRn7Rl3otax7kXiZGyojKx3xX
AZ2F/XpnBxK0FBVxDOxXN0JuvSmccBTp0SE4qniOq1hobl7+J/xN6bvWvI8KJLUFXrWgayB8quDp
wD5RAYL+hh8wKN6cWMn2Pp2Nyu/qBHFO/yTdNQ3ZieLTyFMdHinetRZGalL2tiXtn7vljDM1HSq2
TD3BZSJs4IdW71hbVUzsO7WwtaXHu1KnPlyV8WuQBQ6W/b3zRy8tJoJg54+SNYGo0nQvzH58D465
ZNHUMpvGUgBhmVr8u2wn6x4vTBOqeao+PGh2zcyNYYuNlQFnrrdjUkFNd2SsManO0dLjZkjFTJ4J
65PTBo9JmOnJj5Z6m6YRVsnnHN0YX9ZkUrHLEtSlRkc+VBKPPPQl9qh4Xw2ETE0QRNwMsmcAY6m3
Q6lPZEOxwJU29Izx8JpmnfMYBgF40jgLHevQNzkBquYTF5jUjwwxPD0nYmett0Sd0Z4TlKyCa2pr
7HCbXu+31aP8EzOufHPPn9n2NVHzCgK0mMDae2a7bjzHjpTjOM7EK1SdZp8U8mflFR1LVczaABvR
m6LlwFuGPaqtAgV3qwJpGsditX+6iy1qdsDdTbO6Ncv3Nz39ozjMhuN+45Sz9LIi9SFhS5U4VY7B
KB3jG1IFu0VmqTHZA39pxGSwlMMPi3sljSL2gGIc1/A3UWcuVPB7v4PqetKn6j56wA5V/7URLTBW
surtCev4U5MKJGKG5Nu9zBf1+afWTuOUzeptlfYO00jidK5FexQ84gt0crgbR6IUWhEawmroqPhM
vRNI5CMzDVmS8Jm57mgSXK0H/itUFURaTZrbEXoTMjblseGaZOt+frsgHrbbyZN7kziPaFdm2hZh
/VH1a27IrOuSEiQnj8fGgRgIOZXxymHqEGWQtRR0/vg8pBaLKg8VbC+FAato9y5wi/V0ugT6IHQo
pb6K5lA+T1nfglPc34nWxTroDt5/3S+b7fi5c8A91AYX15Jd8OI3UVXuvCDZv2yoMWisyhbnqrq6
ArxW4Un7mWWwqCT6z9EK/B3+B2mbIY+IjxVwk3BHTc2kL3DV9oOc3Z/INEzhAUXCTBHssWl+01ZZ
oCkU7BQKf4ikm3RfoEr5VTO9WhwrLGhsH3nkr/chCRd9xdQHWTIqLKq6AgxHLA3Ljm6BcxZCSLyr
tJFd8UqA71VO1VMpCQ9co7imT14HxQ9UvcDORi9WKuFeAjCAMW2ZTzoSuz4LDfwdcD9LSnRL2YiX
VLV72Vx4eY/I1/CyQYu9lIF++jrljWkPyAYwWoJc9cheOagsxtpd2Vbyy9Re9RHw93ovsKMV5+W8
DtOy/MbMkBSvC3BeyZWdwFTM2s/fi6Dr8yfOeaJPlIslxU/WuMGyl85DAD3SW2bcLF+STvPbhAPN
ZWAnU1jFPqCIYPcRlTYeTpa7OFz3VjcZ2K5s6qBzMDZhaqaYr/Tz3TL4m4vQDbCg8EQoCCASgjSL
DP6OZrdtV/hUUtWk0fMhxXKfJdPavEFpNZunrOh61zReRo8pq/f8Yh3J06c6UhSKr6WR2gTgmczo
V5MVXlDvDyQwl8XjZWQNZH6McAPu4x+gAG9JhdljE9kZDmDdeWDKu8K13OCT2hgMUsbIb5OFV5lq
SUUpRsu7OX6QzVe5ljg6bCWaE6PCEt2nuC39ilO+DYbe/Pb/YE+/3xqUcNTNSqeWqY/2FU6KHNOI
nV4Aa7LL2pEAb9Eg7vzHIO+83JG3CdIg3L8uS0u4C1iYAfj2nUFi9liiuHGNth741sk4N+u3BVLp
cN74fqTs0d6Z522ewbQeUR5nRf6IUpusjxJ4BR/8FLYp+oRG7S4LAXqqhX/hdn3gYuVSfy4AUSHr
AyVYX+HmvwTR0GjLtJO1I4dAxGxapz4maqia8GQbci7XniTgZvNiS+Kv6lRfopS3nfvl0dAZI+Yq
Pb2Eu/4YImPUzzJPqC9bByJwLjoGJSqI5EaKjC7gEkqQlQHqQDeki6pIMF9k4B5XQQl5oLaE9lWl
iH1eTpe8xbAC4SIxqceGwVuGF1RVVfwIkO56XhuY4lsClB4WDJRL5FZeWAogtAeatzJOexW1+VNp
ESAknDB0K5AwIwCzWO8KaDyfcwvWkBUNrb8PDEhpj7HsVKgDgDwhB1etg4ZVVjM68EOSS/RMrWhW
WyZD4pPwSDGDRmz3+lZYYp3NdlYfameAgA3HH6zXhdoxSuOzotOfNUYo5S37Hvo4Y++1J+2nSOxs
2gtu9EozusMtsVLu7jZYMBKmqwjIim0nuGe59PVkW4TcoHl/6iSWbE+yvTTqtRBu/xFlQN1Iju4n
JaegefML4jqwM+Ecov6VU/EYqExp/swWPC8qThzaVt/5q1g7skIc6O/061HP1uU9mL7gl9fN0QMN
pnwz6YDYJnP36w7D/5f13DAiQ7C2mcjTdiVOhtfgNtTDA5MAKBodIGz5zXZgwYaBwBJJRQ1cvqVi
MjwErKt/3/U5/kQ8rzjQQeq7J3ssX1Nky+P6JWEQ/HlNtZDxKFD5KTns7n+ovEUKqyseJO24qbfZ
sdJl/oXftTHG3I7Qqw4nlMLszeq2J4KGux9k1jzKDOar+qmEpR77NjgSTx2Ud5QjP6OjAjdS0dK2
Kt4HzKajY2r62FQqwLFnWz5M5dXAYfm2HZVsmV10JL39RsFKFofHH5dFPvbPhMhYAvyBaytYQ/59
2n1+oCG4Xgw74L2Yv+Yy/NFavTYZDsVlxGhnVIPCE+kGLD8m+zL0TaXtK5XOWfeEYiAZw77F3Zb8
d9HYYRKEGxHmNHuko/FYrnmGpwfl7qX7bEpkAJOrQDa5lTjyKDg6W58d6BUfMI7lBOqGblUy2B69
44th80thR5xfYL+qj/qtIjEQRb6oI4A1b4De5BvZSyxOsgCWfmcD+hEbGaQ8c100NkALjzxY3VE4
xX2sCOIZNpes747/xq/FSgNas6YhmaYpCCNvxFOFuZyQAWRRqn/W32hrg+50CE4kHz2N1QZpQDt7
AIdwAnt7nhf9EFUwvzQQbcaGA5i9+OZMWX1fSbM+TfmggFKMLZleugCack5qSQhsvAj9ItOc3joE
/CGHE4l/pfTWtLvT27+pwLJaLk7VnxNPGysYS8k2443bvIj44/uJJETgkRcGAZfXBarJux0qJNum
PNL/jMyzgmHV4ZrhiTjGDvHuVQoZDFhT+dbl4UOFs2u3OZMMCjzIp8IbNU1FN1RZepfnyz9b/Xo8
65X4wvFBbOIm38EVOeROS8DhqdnSkOQFyHuzLJE6e1Q7i+807FdxaM/QBeUCSZ3+QqO/oO8lp1BI
l372/vfrlFyGW6h6EKF9LJaAIpGjU8uJpDl0zqsAJVeJsGiEbmqPoSfDCnDV/ubNdyAW5Y0nPlY6
Ixc9a/x0AfGS+NoyPwEIs3zPArevfTTFxBx/G/dXGpTZ/JoWAZhXrwlF6MaWjkfJXTi3sMR1b6A0
24TgYSofawStrJWTe6PqG7Je1X09BeN0RwltNOeOCjEdiko9cMqxRvdssPNtPHACvE8fsfJhzU5t
RzojhSHQsatlFZQ0XpBUPwLxbg6nFgz0nJIjA3Aiv6yjfRFBAbJED3e49FaZoCi/E3xel6nYYWsw
AbCkd1j0u4OaG+PxaEQlxOUXWHvnvjxiV9LiCmnFEWfHnQvUEoi1AIVWC8NIyMXXCapzBBb1KIwq
vYIDqwU1ljZgGZ0KvG9pr1HdB7BBm8zvcjfi0cKHvdBdL4EIktAQPZyel5fZe9jO67tNmsQMCi6x
ZPO61n8dHbRFSbtmFkbNcm+GHjvzhAnYnoqpYCQIIH03389hcOz51bFb2sWSScMm+abt+pKOwgTj
NLPWeNPuQQbAbdY66UnMbm01h7oGMv0rqw+VZ3aUf1KkJtH7ec0SCKnGE0HWjLwiKDDV1l1q3RW5
KtaLFIrLIDQUEBr/z84R4cZb/CridLnlq1y4IHRLn+uOLo8kMOFKah0wypCBznwce0PBILrImQl+
i/70t2XsTWsAZYKUtRPfj+qJ/Jz05ly7FOgqGDbmb1zF04QQEKKGLj16RIjZJS7EuUknReM4U1R3
cBYdV4U7V9+jK3JKMOGchnzgU0skNaxY5G0XrdR1x/luHLxJhmDxjazpBbaXFjfVwUtFavdgviJh
CMWndo6lU/i6/mTExKCdP5hZ2cYXHJ1/39hY1LpWawYEkpvBlOiCauFMea85wv/Xrfq2dkQyNjac
VrvQHyMm1ZFyqp2UZLu6J6aDEkeLNN0tMY2+A9AndDetKMQNzxXJ7QiCsgMXpz4MIiGQB69bYtC9
muiyCPLe4qW0T+hptBlxmCwN6RMvDFyHszppMEDGcTTpDBz486h1mZEwBqRWgeRAT/jdwrA2FDMc
bPlEW/oyHg4UVueX0IEKRCMq2ikeX6DaC86bbYICX/Jbq6PMyH5MONkAfiRFkvJJJmGbKu/tzT9V
fPF+F33bOZUvdmUZoTFcPxDnJIHybNsSyaJXAtsS6ipzuqmxilssdKe7FvRBUC8m+KPJPFffWBjc
WcMcRvyOMPl8nfREfUk4ppg/U4P+4bkvA0DebS54pAA5oebK44vIx7f0rFz/nmc7L+4J3990Toe9
iYTfxihECpab8G0tftQFR5bRkcipoX0nYwhCK+ShV6QiFlTasRTJsiuLYDX00Opw+oJNmIOq31SM
clVuJ9WT6zgzLNSnjhg7r1pUO/ROE9M8zec9+GhcTEMbiKTEl1MrvwcHAb2GM5Oof7CMa7bZaTgi
Mla/r+wgO4az9k7tisE2nYB9AXKPamKoB3gOS5MX7HhXlFl5q5WLllQYGkRCEUBisBFikG87Akqn
oXh2vKamrv1nnxWkLEbtPkeU82KPU5lpYHwkjwSzXa/aaqjAOsaG7m8OFp0DjT1nfMw2xS8oeRqT
KuTrEZ9KKMcv92HYRpO+AY2Myhhg3xTXngkvusqQkbXHms2+ZnrqNQZhHCnjiFXp8TaJt05TqXQz
m8azVa+EAY0iDdf6qpRX/5dm3Ft7HzCj814+pqlA0MMXET5SD6YGYUIxRJabkbbsopPULhwV597x
ouxRY0f74WUHRXhezjDkqMQTEj5qqGT1wmWcSvTkzGe4eaHAf9GLA/m+60WUiixLqRyaJQVJ9PxB
eX6iTHsvavp7Ur8LrWv/EOk14PdYh3Lh/62TzqaSjnF8jC8wYUgM5vlM5hl2DBLlzps6AJT327yX
0DutuynuZYYot2DRFzK1ZzAkOS7qFEt6eRCjIZqSed9cbXbGve4LKu2t5bbTKn+HAVwek45FFnug
HupFPoZuspncnlsvBtnhEuHWpviUKZNdxjYxCFWGC9ehytQ56O58AE4lGhit7WRFaPtNFKRvY9sW
GTMnF7j4zyzgjH7k800ORzaorICJfQqNgUKzcF9zjFDjJ4DybBDOiE0LPJ8fLuL/d0BdD+UPdycJ
RwV7HDDC7fFMYUGfC6RiF1sWczVmUEDWm2aQhfJ3RmjDMkCNZWlYKLJsemYeSw2f40WPPuT9Y1dI
adsHQOBkM/W/9ZJBFFp0Vw2xFGczHguu6aAE2yX5k78V7nsMW71xOZFZ4Cb8R6nahNRqjrKK/vNL
MXmQw64iHNcdowrUjSwpjyEQP2LpInn6NESlj0Ryxb22/pfdM6cdZ0b+bKd1uvYvprHC0u/mIg1B
QY468d+PzwWHsSLKpe+t2nMFHo08V2UprhL0XItMtI+XIRnrlZcCOGRfxJcv+MT5pjMe5QTsZEkg
tZnb2VdD1h2gNyBpPvKWSzy/nKtGRcNVY/UDwLz+p6S4SVPvsM+pi5RaVkmaWK5iUK8GrnCyu4HZ
pXyhVetR1cTLUuyAu4a/GoijB2iF0aDHj0Hs4+4q8ihTeRi7i5pfBecCj76pmHULeKF4DSPGYoqB
n5cEXFBoEiPULoAxet8UMalRUyc35As1pFR6m31V3K8IvjuvSqjk3vI6E+sf7OZ26ePWqr/2DH37
28qFQaIAOJg7L2W8GSnScxigbiO4FC0AgwLVZ0dYVRXcPIXiEEscewkwRTwgd2ny+jvyWfbeJ8un
AiszR0g4ualmQN3M+GJ6U5IGlIbVzcQ3MoXwtA79Tgkz2GIAYVkSsPVurNgS27fnw7bVIDDtEmeH
tz2ijpacJf6eIc7DuIwyRetPZUIjLrXOo2FRTm0IueiXIMB6/qwT7X5kfeDK/eNLe8aCeDu2+RVP
610dQKmznv4WzrmX9Bsx7faur+gUAYtuKtz1GahhWIdR2KBSbk6wv5kYifFUyPzsaHV9/OMUrBu7
XT+8Uj4cDXBfgrXzxAcf7d+Ew5gVbSnXA9UFwOtRm2Zb0TEWaNR0bClPIqvXzBWEWsqdYKQI2o2g
sghie6oYQ1X8k+/QdElVgmAxb8/3eAtSvu4b0XltOGz40et8ofuvQJrMKlNPjmwBSziwLmgcby8M
9c2gBK2N3AcsV4C8A1pMSur/m6IS0GFd5QHXiuT61lr5q3BNCa21I6w9GwkZrpX27nkUXdlbghoC
pvgKXMbDHQDFeYLORaTRpfrt4+nb8AA03V9HYiXuHJI7BAADWYUUF6ZDDzCls8uddz6upQGA/iR1
DHE+vHnb3amGx/SEngZez/60NokhxCL40RFOWBbOlBai4sUoZO1R9Z14e/3h5m7IdrfxQArF6oYu
NwnbEkbOp4BS8B2s4LC45xqxdqklxwTsHJHlEuGkMEP09E1RBSo2dRm36takiq69045JQO2jlD/D
ZL4IczKtrXydoMvO/p12KIR34FbGrFWMsU2PKRmQ1xhdYwQO45Ih2SF3YS2Pv6eqpUK/eKtr4o05
Cs6KkCuxqvlsPsxquXsM0uRhOB+aqxZV9InJNAkXnoc49YDtOooVJx2kjq5T47MKA3LfGTPFuVVl
HJ0TnhE2xY075qP4sVoT9X18w5Y22BSq0Md4w+z7jXUG2w371uvuNK31tNMa69M2kSg+89acKdlz
C2E/OAQ2pa3x26n/yK2zKJxTW9MToHCWsDv386tkn72QUmZ+E3Hu2LpFAzHGsBWCwkNCfU8rxXpR
piXukjtkIVzhLHBlGbc4MlRexvFwP1chN7s34Czob+wmYZeCsdlyRZEkN9kNcQoAP4i+yhuyT/yc
V/lC4tulnqfnoA7ZjTuotzO2kGUjIL37reUgA+NIXdusy6xNcV0RbZAR3yXmBpxrWshf2JMi0259
+nYjIIbYQEOTnXnZ4J0SMy0+/XWw69NRbTT04wa0U+qZ3pfVO8bx9KMHvgqug7wWEqyHIxeilslJ
bmFK7NyDhjX2m/py1dnrzuDCSh9f71flOdcgtemyJXDsPVCTHgRAEPQ7v8VCqIpik5FL7Sm18I8k
2ydYUEbFTwLnHY8sIIXmd4FcQ9R3B+i283c08bEqggHpvpj2aULyzgkgSbxLi99oKLkH8lb1+waA
XEiV63Th/rqHB7/nIDpu/lSYwgu861PoTFlexiE5ut++6ZdfN7C6o5AoR3bxNrio1nrQDsE/XoRA
E+bvxUcoOonUlL6QfyMdetYFN8zjsEg3IciBGN84QfS6P92wGuQCB+rT07n3dbW5D5VgXgle2K8Q
ELZ4RSg8kZCtySXh7GMShwOQOJN8jLjvRE+v/oZz9GVLL6teFijtDtyS/v7jac8dGMg87qDwyieE
Os/6Iz92z9ktym3nz5sPR9N8ZsHF9AAJUC7iq0Y2qMUsYm1H5g4TWK/t9+D5q3Xj2GESKfziI84d
fGJLSSW/ISzuIOPtyEDb4i2erVhtKO1SRIusRTQJzikuyJGiiLjlhwz3tvcWj9hWi5t//FMT5j9P
gey4tkbJohzRWnYXNcc5Uk/ONivVrcsE022M5gZqPMxGgca8W0LXMLY06xk/EylY2lEFahBT9m4S
3B8YQa1wNIQHlSS5qDULnqNHiexOxKCI+kHCl0xvp0uW8eTdo4Iyk1LMO8npQzW9RzD74bYhi4mU
1xSwJ9a5m6gCaUJe4ngNElHBsw6IxJ2jXpXMBizLQEE9YIo0BdhTagO83asIdDh9/fcbh9G91iZV
x77q0oBu9BYhrqs9EqvR/zWE2DPAjlLR0HbO+n6RRLOLmB8LB2fvsMOYMJU0l4vCO4uh3cF6uGYp
5oGgkoLro9AH57DiF4+6jjadIUMivBDp+Co7lLNulhmU4nmeCjBti0R0HwMvSzyF4L3wqj3rAGf0
dncmW3iN0OltcyRFMQo+XxORKO+bSDOZAVzAK8ZqVsh+UfgcjAboJ6hUC77/oNP8howK5F/i7G36
Sxgm5dwrok18WxFg1VH8ji0GrXzLpwMA7CCdCr0m7ZyHXwyVZ+kXXz4Ts0U8mQ4nAAu79BiMxVTl
cFFAYTEv5tj0rCGck93XP7A2U6xEMJsdAvjtoAXN6jXjOgPF3StOAcXTsDNLI+QDRSwj/NqxbMih
ZIVnuCmoOIktmVsfT9qdUHKGNX+E649k/TO/IqsG12kFzCelfNeBk6vq3Aqm6ZSNV6bR786/OxSC
p5XkcpFsT5Jorf/UoJi+j3SEpypQFUhUfpFsWkWEQWWmaa1XC6D6+jzn5BmSI+D+lx0WNp7+oLkK
bpOA58hLqbR9vpJ3gDqFqut2S99yS94rmfgwbYF92qnOHOQep4h1TEjgSSvnh0ApZLQjXp7uzxYu
GjoW9ndJi/ppKmsxLfUItG4ctUWbYKVTej8/mpN/1rnvciFlwVjcWFP6J+l9UqoqzcwIL4iwAukj
m5lchbhgF0FBAjq1zTidZ2U2GaLiEQEVmquz3P0XqGgXpiNf4dA8Nk/L7TZrOuJ2nM6mqzx7cEvP
KRHLWOJkCZu2xKPSDwHDgaK91Sz9pzDB5ZviO8U+1m5Q/Xj4mKI7YA9Y0fH6eRiri5smiLEkCfD7
28u+uGtHZjAic26PQ0c53PN0IHdeDn7SsrUhWMbjP8u5sPxcBdUmTQvB+wb/Ya0KCoOgK1gKL2cY
+TBRFDt9ACl2noFeudVV6EBk2AUj4otaRIPnGbi3cCrVhRF75VV69bpyzKmCC74kyvUXflIX+m85
ouJxK8iayCLSe5eROn+0kDJpmkTzMIl1vrJ6jnyIxcg1iQzul380xSWcC1z8zEOFc5K9vN6/6GMU
rcKSIazZe9HmXX9S+YTdZ35AEaAX/RJ7RR3lOhtjIY8jyQhzPdUoghwmqOGyyWEgOMJMnaPt+J2C
g9D9i4zwdd/xoOBq08FoXbG+ilCxYpCuHhpTjUw8hFw8eetqZsxy7CIkO3cUnROzWX6jJeckJKNZ
IkekzPEUUeLMnNCwKsvY0TBg0g830zSTcFkD7J8zNBNQNgFi2oTH0iq4ZvSFpW/xTVJMQGu3ggZ1
hlGYNUTZiwf8q7m+OtikTnL/RuEn1OsBCoKf74TxHyDFcaWYyNNN9FWhL+QIphWi5gKt7/XtmXQE
nOdyTqzNnFvjhnqlu6Xi6GOc4MqqRY6Hl9XBXpn5LkEvOf+cFikgnFvVPlU7sLjG2wbY+IlF41MQ
sucGJODsmiRJNf7BX1wo8gJCeTmKbMuj9BFhw4IzcYtYZtUWZChBVW5PF4s6z0IK4qeWZUk6yjRD
YcDxcvc2COnsalAVk6wYlVEudxuVusigUYIOTNGybC3o+7HRXY9vEtMD0ZH3wQlA6MoxoNwHDynl
RJaiK5cVjj/8ruw8LXPOpqm4rZJ0Jk31zCKr3Ib9VRPGKkW0h0Ms17xFlF3tITEcAE44D2E31urU
axXMqEWxT/HH9/Ba+FI1lOQDO8WlTXG/TOkPwKM7AIP6y2T0ZrN+43ckHp60NsfUIGHMOccBjUeO
hWXcHl18KB00D313tCTaXwa8zZ//gwFqoN/0EPZWDa/k70q0KUzcsX7lbQPlzC2M9MAbLcL2o6ZV
DYS1pV0geiTdicnQFohArY0zC702G839afiK3wlV3D3ydl367Yx+ssGDptp8RP/T+VopwRAs1O/Q
LvVF9+T6JIA3zS6e0XPjBri4TlyXarDtr9q6NuiGyK5uXCMb+fHXRwaZ8Fvi7ALKET/XvhCvtiB+
tCEbf/Bogxl83Cih0Lv5nXuBCd9yu/BdsmkI0rvXp4CHUbDbCz0mtL65Vkeo3C2u3CGaORsO2+IS
xmPPiTTyyArgns9C2OXPrUQF08EHYflVF2C7L0h5QBQ7zlWABlIE3FNge+0iJvurwcwCyUuurRvt
xxaSdrK+rTsT0aWkGrhV9DPwYMv0GfhtE/cWTTtJHkYCz7ntzKqThRPvnHAT8HNxqrrJhdgwgiAc
GmPuBoBybVi5TjooZNN1GgqU6gD4yuiUnwsjYkwNcyX0EpZFSS91ttvJ40Q9wHcoCkh5g+W72YuU
WdIV1vRoJmzhcJmmD3/0abZbJg0m/GI+U9Ld0MuXQmsxkuZvVZcGm9YvilIkw/tVbBxHQzLFuuHe
y83fCBHUrhX+5aVp0oQ/xKzv7SAgYjUUvVK54xCM9+f0I62rLzR0noXTXm8LhXK8g/AdIjo8dVxF
LNNUsSzsv7e6C2r+u7LiO5mg8366ZeIQqfY30TZ9Porubd8h+fZBm+SrKf+k3OF5bLvzw2C9Xh1b
DN1XgHAZobO5ESsWhdZfGwwFSKwNCb1SEpy1Xu61+4mDMtw9Nor3xMjVRQcFJDKfOfv3HEFrb8GG
JtnOxre0swLsZ9a77m62ySn1w2Fc0NHL9BK1nL/g9UUBBfDj34PeEVLBor3RoPiOQtnciAVLAOjz
aOC1Ke7Ef/8EC8Nxxje1WeXDIo1J8voygjyTpPm6HRH3sGm9Ua/w1B6ssTwrR2t6c+XIhbZx9D59
ZhX0MpGvxVDdpZGhn/D6qX2rgURptZQ6yPq9smFwarzpc26kG3ZJ1dA5rwzHlYex1Aq+I3/TOCqQ
oSbwSffhhTGfWVL4d6alrt6lWnkgSz6SmYf0GoFLf1ArpaYsT1meT3Wlj8xN/qdsChbAoVNH5czw
ipj4BVzziC04ELaLJCdbTGfaJ5g05+t+Obod01qF/hJ2Vh4xosD74zEBsom8RK+0rnYI79rqQljm
8jMrB/KiCGOHa6m/XvNEjSMDvYeRSLnKUNMvy4TJ1Heamzs174XWlP1uOyJr6U2srfB5zDaF01hT
VU0gQXIRwtamaUPzlcwL50oK9DbaNq65g4vkvwTc0UA08GUGCqNXyqNvLHmg9KE+4dw5USswRN1x
EBzJgKhdyoJuiWi39pZFtLIeWiB1vbbG9oA2TQQr99lJL/DwHrTV+aT9/ZzBSVA6yan0o8oVZnPI
bDIxzxOp2Al1aKZDj2EBFk0e7qj4S4cb/gNOWSuUJD9p9eRe2P1LsYbuj5OowBsoo3//BV9mvd3p
4BgOuNhgDhkzuv7oFD/UmtZhnwsYPL6OLbG8gAqNR87UbEydaYjd0t1Sp0sX0aB/h5SlX9Ar/Cxc
MJUQwJInMJ0rCFkFDRmzIKLtOIWYzEuGcdhIq9e/HNKBM5LpRal53roPGYgOLxMDYDkc+kQzI5FQ
D9tLQBAPNFRBrphY5Sj6ChWnhc8aeDMR61NTbrONci65Noc6a2f5mZKkOd99g/IjMeSfeJCCytpG
7+2pPqYlXuej/U4GyeLDZtlFiEXXEMAjynY3lPmLXPmDERoh6Srs140pCLIaCPFdLkgK08CLjXU9
kWpOrKtO15UtWJ3RegGp9xNnitXspY9AqJJU6EGf7L41yVl8u5eIWe2qdUMU4RyMWqM3HIV/8GW/
+ZHrbUyTxmuaZEMYNgJNLfT66CtYXJRsY80BwvJINvyTU1K6cmudreU7xbE6+ywGT3Zq2uYq6KqK
ZWAFwT3JRdYihXyb+9EMRy2DIBsWdHwvyaFb25OdB+QGj0XW75/3rNr+7pllg6ujkbTHt57/9SqZ
SRJLvJ1QPtGT1F/RGoXfwpgd9rgsxqGOv9oEbM0gMiJA3QvI6IimF6X93Usgz9cqyQKQ4JfGue8L
RUkM+HE5iewMYx1RPhkj5LRdP/oXccgatI4POJsnfvTY052IQm6ebgEK76HvyTO0YqFInlHYd/cj
7Wd4XMLkAjjWbfTravvDhJAQe35wvrF/Ltv4/ECS/vkDjCiRfCNRoW8sdU9Kcsk9j8Urgncb6oSn
IA5Rei8sL6lCK9J5RlcswwhMs2LP+VcJQgnzimudafrauXRTn7h/4odY5A0Izo7ruO+PEMh/kjzk
aDd6P5kINr1WOb0ZxGf8M5o/vmJEmrDPHff1qEWjudqaAsX8xBbLsnj7/Vce0oFM27w8T6W5wda5
Uj8kOOf5+6cMqnsMsOE2FNvmmmMQqV+UbWi0mTfoY47VmssCIWRA2GTOBdXnn08ivBrkMhwrK/bw
j/mwxPFwrYZdfahfSeyHSYL0IkVFoL42Gew+lI8hajz20O+JykDtaXGuYEzDBO07HBWJVj4qywty
WNKt6OFKBrk+QIeO/iY/iELeOPXvALgvrzK46fEhhFBrRgedPMMo7cX3RUweYvTYYWt8QErVaz1b
YHd4SzH96qA+/vcAShkWAGdObyCMT5bdYGeDKIKqbdlZanUCWtJ9m7DuaGMhl/m49yOiyKQCeNnq
DRS0UEH3mhpmKJUs5mYw5Ti8/RpPCf8NRGYD4ArFqdNafsJ4st5KW9SrpQDXzVtGi/ukdHATOLyk
bGdzPU+aPCwXmELjUxOeiSAIZWRhsoI3Bhht670gtQTiFk+mxuBxfo1+VD/69WxKUpi7NQYzdbpj
+SW87PdzXhL278diGJnbPivjaiG72mcKf/8cFgK4Z2ER7WTe/HyGnND/3vMTeP6r0SJ4KhusbArx
4HsQtxS4KKEHMTNr5AqRU57BxbLZyohF97aUfyfSOMcoMh1oo+uMf47DyBZpoZCz3Vyo1sH+AYH+
CqmEXlMT5JjHdyJ1jrkUgmgraZ6tRxY2Cjy1SoDGVwNK3BaSkTsDAzixOrqZ3qjY6F5z/FSCPhRu
eRJ1cJ4rSxbXNDE6/9UXbIi8w4ayXbSZ9mSWT+Zkny9g3SbZuG1hhcqsbpHJyMc1g9HRdkbfMtYj
Ce0nO4V2R98e60KBiP79DXREuxmCMYrC2Z+NLzWaAFoIvbtpsMa0wgjpgU91z9Ea9u5bUlGzGoom
INTHJDMQVbjyYYgl70aWiOIy92yWFdkNVDwcI590eTUxllEtqpGb/kjJ4kRoZu6nHzBDhNeIz3AX
5c1liG0VWl7+vtXStNnAGnhK0w83J5P/iz+7zyF6PXYlvCGMEpMrTkVHFcsZgEiI7RUvL95zyzYb
kMfQB4HRDfU1Ki98LfdDX4aHxu3ytB3xkoj4Tfe6EZomsY/vAnMMoEJyIQTYXLxykN753uKeUtMA
6icJzSnsRmSqmSOkY8z3L2YZcSDhOI1UeCd481Dh5Cux/qNcWWW1nRiR7Z7OcAkQBnD5DneWa+2C
5y7RVjWTuF5ICG/iPRgSpVuu2lIyVEGJpOKe+HJmmFoOBV1wxKRItNIUDbcnE3sQL/vrjfYWfZ3a
0o5qffEIhvunKnQ95NGXO40wFuXj1mnNCC2DMi8gV2R/xSn3vSXGxDPYVfM69vDTYbrkIrf8M7fF
XqhqOZQRmZ+nFqcR9kIz0Yw1rWPliYfMyvnmxn2r7F7yzKjmaXma1SoYxw4E3WWEJAdByh69Jnph
/4xfq+NBO1LUXgGDMo3n4htdcpTaH5Xt+Zsp3+hoHu9LPQAI+eLZgRmmPehuEuuCrpeg2tWDr3B3
Y1mk74Lvq9gIr7HSkIDZwr+UHwTiba8Db6HLV8KBsOR+afRvo4eCjZpC4CSG218nCQ8o8GztAP5l
fZyqFSUCgyIyETZWGGQFhZQRZCo3puBXPrUkkxqBCnsAAVi9KD8LEHXuREb6AUX2T+zKacAAavL0
wpvBhyLcM3lsqWZ2g8DyDjbrMiqpO3FkVvJ+X9K7pFF2d4WDlUefP8Dyc5CZv6yz2s2WIyHMkL8w
vRr62JX53ynYVYd2z2eiX9T6TxwIkPCyu2iLepF/QIKOpDAmUamh0YOLFKcLLlOYmSNXqGinlsWa
1Bm6nuu3jSHt/Sxmb32WM4YyvCmE30N/wuBZ/OswvWS5a3lCdoNMbC+d3Oky/snkZFms0MWdbTeF
RddKs7/tbLYcgbtRyQJFZi4EZj5MmhZ2iVjvThwxdxRIrq7jUp7lFD6tS6krt6DqazvxELiXadZT
NC5kOJJ9ErjZTcV6hoyANZb0WBx6LHbR2ZgxxOkcedH7DTzA8f2dCVwZVWlnrAXuKS5BjTe8RBrL
G1jPAw/GtIILyY57KdFw24cpK6OG35xI8KfqtNGqFSqmSswxzSQmf84cOCrgIXlm3D9ZoCFKA69S
eO998PM/dXqp1sk/ECqsaSN0IgaShVRII2/t/R9aqG/E2eayHrFvESZqWYmCBCu2PNLaZHy0WlGY
/LWK7vusAphHgwxLh93S4psgDWyv7A1dhxii0HAbIvSo28RT1yCHxJHvH4jDuuMjEF3NL3Cvc7tq
D8Me0fX+99xu1gN/djT4j8vMBIXX0UtmBZuLW7Q8rZYjxWDHEepie8dT2YN2EsUAF7cSFW18lVP+
ubtC04w+9IKN7njywZeEwhACtrZkxtnl8/LyHLdgu9HDv/jq1KFQrkvqbNt19UZOzVP0RYXwi3k3
HkPSxZ7m+6WwUK44sezKtdTuHMPQrfRy8VBA9kdc2z+dI2c3FDc0/B82Mnd5ZV/WOZ9rz6mfECFZ
ZMTjWoVCODKQh0QEosKKF+LCyQ0bxpq107lHHO7Pq+F+dTfHdFOu4XGLe5inV21AqyPgYbqmlQFx
adXbCnXfOBEokbmafWu7fF6tFCvndt+/kqkHqE9V5xspRjvrZ8pf5nrRoIkPP1b0
`protect end_protected
