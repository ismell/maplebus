`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mOT0ChHz6cehSpiLELxj0+iBo2W0wxQ3KDdDuko0XAAnU6xBdrTgVJ+u0CfDTb4Zl7P4zVo+9SdV
/b807CQOpQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TIcQNAMAySojflD08WJVTUU9TIju9tl3W2g8zvY8gbc1G19U84LFJDx/BCiaF5xPqjVVg87yUgP2
09TqxlZFyKabmzuwew9KYeR0jCYUfbw9LnykzrRmL8VwGZ+R+KKM6qh3sVi8kjlVL2vvzDa5TEBl
Awc1nu8HIXY2tCzJxYs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gDZhaaT6CUUs7NnIWeXm40ShkQoiwW3ulV3VTiLNOl9JkB67JiQncNfcedINRJBI0vrbIbe0VuEm
nGWVSgedEkZjaIEOLxHTzpLMo1F60XQbe2/TPwLYooDvdzl8qLzAmFDYq30Ba/2aGCezm/7vOG06
Dm5bE75znWK740jCPGoffZQ5cHij7UEXM6PI52n8olxHh68YkWTVyaj5hiyi8PuyGG2UrlIptOTi
D1+RpdGtVcyQjrxNNsGYLGgN+kuJ8JKutFcIEuspR+pdN80i9UD8VUs6tay8+LYMP2VIK7inJucl
Icj+a+DVFAuXh2jQLFzSd8f4Bhd0uuKVL0bvAA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
phGe6+X991WkQD2biWWGMisWc9bNa9/igwlr0eXn8S/V772jk636DvkirbzU7VGsfiTnxrygxlvv
j57J3a8Nt5UpmtdXn8mUc4uUSTzia8/FbHQO3bHpHnmXbnQEC73toicF2G7GUsC0kjGzRm9Qo3vn
adTUcOWLpYL/4GBEZkk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aS4078q3A9khzx6QcF9V4RShLeZGpuFmd1jFVkWlgDkOt6ay4mSLBwH/sXI6cnzi9UEFhnxS//IA
wrLO8rlxPXye2TeWt7OMLZoxoieAP4pqHBw9Kucl6CezJBsgO6EPq4FNpLzmDFabGsjkNcdr4Dcr
ugK8/zndRGMHcZ0sbKLJ9waDZ01Oz4muR30mJ/UwRz5b+1m05nbjDMvgkP8glnV9YsHgfFGJo4sF
IZoWULFK/N/g2ML20rfFUkcYFYf7BzItQg8e8ht78Mc8dO5u2afq+FWtvh+3qghvbZprDmmsz1ZS
1pm8UMJMetL7M99dFr8DjqeBexFg7nc+9NqI4w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
4aRq6hkgCeRv2fEtQSIZk7TvWcf7GtHMUGTGO6SfzJ68Y7xUq9AG9O+zTBxFhaSqWcM+BZFueRqa
OJgRp18o9aOoX/sX6PjUvE9196XVlQOITY/A/9FeC8gHBvwEjRDYtiFd7xvlPjvoFdnTyf4UvfSO
pw/OHk/wLbPFuy/obYln6lFgwNMIOjO7D6caRQoysyuguD/97UylsnuOjdZx/bqNv4WEQyzLPFL1
UES6JA64KzrN5675GUnLCP7rK653tgrdcEP7LYla3yYkhTD91sFhzu8phqG6cxPg32We7qmv+RYI
usjtH3Rv0HCWXwQsfBtg3/cG6O29ZZIVSWzmYuaI9czgOZliUsBq7aFhhJTuVkyNO9/9oxISmynE
XqyD/HLPgTF+gYzq2jJ/bIdOwFur9dszv02KacMTKb+i1sJ5no6U3M9CZosvdQ96L6jLWz0TuN1P
S4ccOzozOhP4/nXgdqnNPIHciEHh0FEl6LeUHYlPl1xvBfD0wFxPwykFai2pwCuNAz4moaMVEaaW
X0L2E4/hZa2Dj6Fkc8p4FDgEZX6axG4LeGIduloryW1LqCoElQj4sv7mWWHnYIU2W6n47X+wa5us
XHvYQOOy7/5m8yeoRK6jEX1QcK+lAMu+hosH+jPtcoTFk60h8DZgjJJRsT6qNapl3tqEdJLD2KEI
QBevJiZgtI/7zKztWgTDEouUxIyU/d/7hK625qk3cgPGBC9Mi1MejCuXRSCiXeTZ05pFTR42G7pU
cbwK5yZoZr2rAb4oFn/vFOTrdtFxV2UMZqLcbmF5z6Dptz/JmFu9CL5yDoeDGjiap2O06O+ojuzS
O2Xe5Y0XZZO6ZsELH8bLAUfrd43M2l84E8dKvJzSdktxL3q5Yr5RGdMstxbexX42osOomsHAUnAd
kTCOtl/4nHn1u9h1oN2qVhowJRPrtz5q+0AgMmg8REr3AC3C8681cBgT7hy+2FkGU7Otb48yF+s5
xaa4lKdhNRPa+RHBdS2HvwHqDPeVwQ+9wxge+t8cCknWFDjSVAI1LrS53KKlxXzKZrXWQGoBvNsd
ohaef5OEUEE1+T6/eajorS+HU/0nYb/DALqZVqojqdpBGUS6YweTWo0z3ldp00Z3UVIlz1t22pA+
ge5q2LEtc7jMYPPR97t5IvowoC9haLvnNB7+jzZm1VF+0tUWJ4BWERQvERTSMVI2Qk9b1QDoTTOC
wt7L8lWGkh86SX1OLaKEkXNhDjsCPFcO8z2xaM6odb8R57hYs6Ekz49MwJWSPNFwzI0X8SLcgPGe
+OZ/m8PEdC2+4DhFNfOcBcLyv5uOXlLoucDAmiNxnmvpgJQ+ss2+c5hPPslVnqKmfeuUcqeLhc7j
JnFZ3XXk9iITENPrhvUnYj1cT0UXyNdSInNTvT7hnQF+ZqxUUkyxtggFS5UboBgxk9iSNo/t/saF
9mi6QEYIxRw2fPFK2XtML3vnDiNBqJecwo6Xus8ZrX1ewr2s3U77lii3Ep+hmOydGoFhhStQU96d
/FEOCrN2HRdHGxPxujeHXSBCDNYg3Mdw20bucmjLTpAGWFG0q4EVbQeU/pwMTNhZKi53ic0s7fgk
v4NamZLSCUp4DpvOL+xSe7Qzu3wClo1QTzq8Bi85lrg8lHGrU6owNEBi5RpejNRRXnk/UBr+20bB
spOHnaG/TGjjWir2VKflzMRwEeDhJlOsPGFWeVOMRdFjugk7GaJY2gEXL9d9PouccQUhGVuWvKlp
6VQ5RZC8MkYwTNXRER7neqbFthDmZC8V5SzFzUYhc9QlawzclGm9V0xZQfxTORNG0L9KTjfzMl+o
aFqvXYRZ4fV59DPTI7tOQgQJrHTSXQO7LKvizIG0/cj3NZXN2+WMPp+t+M0SwlDf0g/Qdfa6InGO
R8ImNgasi82XiHV34ApOq37TC43Yf3gCTH2OEQOIvD+SZYuyQaFDYgWBMTommyAbUawMOBh4eVl0
xxJbHi4LsFw49PxIQW1qaONI6U4OCA/XUnz1Z4LwP802aS1QUHL04iJqXsZSy1ciVNzKgx20gYYU
8RccSdToSqJ3JmgOzt2ZX1S/wetC/JnfXt/+dFw4n2nJXQy4GsHErIjXJ6xRfnxdvdaeiqD5mkBs
NQzpmrOgtc1wkxShncndO/hiPdrJhKoC51/GsAg9+PMQBw87GTbCzeHgbWQXvbHDuXnK6gRolC4V
I57wXpZqZ0oG5x688ccz0DIG6Ke1Wh2f4G/g2x8JFxEGBRHU1dE2p64B0S8ORa1qK+NEbd+3lE+S
AKkpEf3VfLqGLqkvERpFY5dGQBYZRc6XiOHOY0Fv3BJ2hLfAhd3Sje2ryr5bNN/FAN+0ZsHSamzf
KoAHvI5oN/BEl0xE10g9jGvO2k05fmIb3CyM5pgb4tbbP2z9n4v00z5SlgbXNPJr8+kCBhAmZ0uc
jZl79VDPZMn8FIN3AUKKB3Yk5H/wQpx4DlgB8FTrnFB3dznGJyxbTl5HcwmCtsfSL1Ryk5HnvauP
Euzg9Wa8FH5lJ+Vyu8NwhbnUtrnEF10CWHmXOf9eYgkP09EuRe8jPqsE0xUd2i+t18H4TZQFWjHk
J/jKJSdMB7h3JxxaReGZjjBEMAM+eI4TgikC/pJHHbFbDrhdsM0jHCI3gY78fO/u/njlMVgPUweV
CWV//AizDqF7C4H8OWD2AZ6nz+zD2OFLv8xNenmFTLIdXMj178PNbRMyUIKU2R4bByGbXj3TrSxQ
SbeojSAF5TjqdFkNudMCMASAsFeLS9XXv5bCNbWdmNOcn6iWunv3vRf2nRyD1sYYTHcIiPohrYzG
3AvaMeSOgBlI92+EESyaxfusUGdYx9LuZ+CvoI5Jpju3sxGTJ98KqS2mNR+btheKcdLdwyj8A3DZ
ByTYHLrHu+cFD1GwGZ6rajle2ReDRu1nAY92hgphQd2cwAuqhr4CN22QKElrS6I7QvV0//O68ksq
mLG8BHe2I4EKnplri+YOIjtHSyaEj8nybkYKYN3GY+mVvX7W7DpBt3bW42BmcAY12/h2gG6hpSAA
33VHJ9Rps+gzJYVbThxwSTD8g6x+RRNKJJl5CcYjYJjw+zU8srqw/9f0A/7bu+h6uS3/FWAxorNQ
4Y/i6pRsyDS7KSFxfwqod+mfHQ05aE1N/I/S+hX8entvwztOhV+zSuUnw/+kSwjuuq6Yj3FCuocY
tAEoac+vBz3ENgmr1dHSe2sfQN/rG1wUITfD7/ezJ6LjCwgV3oYXKxVNgmHIYLNVoEUIftikY7G3
OI+MVb50JJ68h7iUROMLhDltjmY/mnO5E1yYqVFSnUciRc1Thocay8BdiqSHx9luIkNSL++pvedc
EpG4LjCfZuWffiAQx0bxV2IIv2pRKT/67hmfiEEzbjxJym6pwb7ZpjjFEffuQjTwoJvZhASRJnv5
jXBvJGjouM3JUP1j39Hk7UGxC2ZK9R/CQj2kif+9dGhcHFQMUg6wWp3trA0RnYXx0Isna2hTFGRc
WDeV1HOWwlapM3ouEwlwadCuZK/ODtTRqMzUuiiJel/BBEGDAjSZooQ7UbHqO3p74pF6LG3VV5AI
cjF/Bv6Lwhb/TGdlvAZgBeP3L48Lene2ApbcdMJzNQY79YUbxJjPRsZkGil5UMwTflksYFRstnqs
as6hGpZVw9oQmqztdVs/4jVsgEbdnRMXvgM2MZImXxoYWUZoZT7+Qo+Pi5Eps0TLEx51C2LbP0ak
q3n35B1dCjSKM6J0CHUqAFL14Sir7t+fyF3YstQ0ZPJ4oHVZ/alrcTu5CBNrO+Fc7jonWx3ob8XQ
2u/MthoH6Kc5cCsQvkxGvKu7dFQSPngmYz2gcvaMSzIX72lAoMSV6n2+KLMl5oKyZvPKhCSqhLz3
hLpy672FJyefC8TJrHDL7e7XnaxYHGNZp1q+5KZ9H6tDJ69hJBgSMl4NStRyiRzXF9lMm0r0XJwp
bv99x1XFquEcl9kTEpFlLCfESO4muzLetbpAIY1xOvCHv6pzsNbBCPDhbdZb0L3dzgCippdGPFR4
/n5fW/c/JTFBsDOwe57eO/cR2A38qB4dXa6bn2lybNqTZ6PcVrTuS2sOg/+jjpYKNpbklie5E+Lp
Chnc4A0lHUrMv61CFemwia8S4UJ5FjVlC2S5BhFKzLCUmCp9K3lKOkwqsf9Jeu+/Zw1oxYSKbvFv
W0hLnFHWw2Z83Lz1tNGt19ppiXiV5yC+3sNZICkWD62gfxpxVS9m0UgPiZgjyCVREgIpNQHPAf+a
6izxksdohgfOpiZFgoI7te9+4xtuB8RT3WdOkQr0g1HMw9U5Ibdev0PsLAvkLS5IFUbkjy74+u1v
3SoROBm2EgRpR0wWSXn7D0uWZlkwLELaw4P/bn3hhXsm3zqGS4m4xg5/KgTucoQsIKwQUhhzjNml
OvvXcpLfWaX8bpoZAuq/Y/QA7fMu55RkFFPWfUCGx188BwPzl0ctRvLf/ewIVHnBNPaBjNttaEj3
r+lcT/L0SCIfknLspGcGyDxK/Pc704/GCR8mIuVuPwqYVvjjmEkr0Vb8N1JAujfWb//vD/NCx2dy
/oxAyKF0LwYbYhb0zXJiPYMwl+jKZTUztiV2PL5dBuGp/jbW3cbc9F+RXlqfruRkc48Xw0A7summ
KeavywjZH8Xg9GhQ0HH7ymRHXVdtBIKYqUKddfyLYLxzJ1tBMRKpof7jDV1+Ew02qNV0qnaEvun+
rWlvhnuZKXufRVWm7Z2kadu1eTdzZAs6/7R2sOCXVlYFUK4/YwmoYrccwRN4/Fl48wahsTftRk3f
Ib45KIyfrFifbWDcCSAVqQBHWmcGJA1NaMsekjIIhK7UrdkY2F769y8boxFN3nKPUK+8aeDoJnCD
tXBp9/sljP4E0ywP5di7cdvlZDI8hJQ4F3zXbZExWyLwNKKAXMQwy1mfjjXMN3KUjPujQBg5AwnA
QKqBNBWa+AehL3gjkSe8U/Xfz9APMn1clpCMWnbWfGLwECb10yMwpISOkQYjI+CRDqj46gRI79ig
jP7FhRHhF2usnwDe0sJ/a8iWyXLpTe5ZPmRFfIQQE6JypGtZjKT4DJFIpsDOdyYOXwMUwHNFDufS
2a4N/4OrENNkUylZpF5L+z+WItyXOdXci3xpEx5oj/GK8AqAcA5s/tjePT0ze1nefKHMynjcLOfb
l+qtXrtIWTmDevSiwPg9fZza1+ls5vSG4yhMGXEVgCrNfR8mDALsViQ6eUS9HH7K+FObPQGv0jyS
8O1KqfBP6rcoMX5kKD2v5j5EX3D53O9VY6k1otoScv1VGoThYfWoj3+RI7heEZgRp5ATM+pMRIcW
OODQHSXiF3JE+g8DJMKlHJYh10oIw9FGX4cMSDN1+7w7or8wL9ADvWwEwzD+5U8SK9KuYNiFzCIK
wyekDUY1Nbpq1ZLGzpLIKoGnINxyEC39OxvNMIMM+oYSgYbwqhm0tzm92erQxGermkbVAp1Ve061
gEdVOo8T4rp6l4rcSEx3MrlHBEE1ZLtFA01X7CATrUn0tBoz294FpPf+qbJa1YBT6imRT0zL/Dt9
C1u5xbZU0rDDBbbSTm78XtXg587tTVWXxGxflLT7uAYoXvPUfO2BhFJhSja60B1vJkYUEAO2fizw
Fn1K3RWQRtwv5BVRqsvctGHVRB1K91CSIIqQMhdWqmS5oefm75dWgHwVznFMz+OfphmG/bI+u28t
5L5KYiluqHbpbA+vwYG3uFOn/DXHf9l/OGvxm9knGAT3quDIMPq/eU7NerU5D7aUpOg1AbCjeCj1
2KFtXdxofXZJS2n7RFl7B8e9498fZ6fH/vkw+O4RWwOEpvkntDVjpHKhexHCsml5KnrvIVIWCo57
L2JT/pOwpfA9UMoZ9JKrJnqYOrgnNki4BhDkRvDsETeYFLoL5SBJ4zdj2Nmoo4sdhfzXqvEjJYlv
1PsaK0T+F3wQZwNyNgupl73NWrYUKf/kpFfltmezR4G0Ooz+9gsK6vTHB1+f7Dfa2RWuknsRLImU
TGkjq1bimFfs7XqW/k0TmsQeyj0m+MjOAdQPZskvUcxdhLHHrMD2fkueZSf+e9feqK0Pd+eLmsI3
8+vFT+nX0e3T+oNml3IglN8OVFz7CCRHoS5ONkUj3/Al60X7nCIITgj2HsKsh/L3vIPr6bRURYxu
eL7ST/1TpYNoXvYr1rrJcujx4wVdQ49pwlWTh2LlKg+tzDPcnYiqneh8edauUR5ftWsY4GWQ0P3E
65FtgVTWuq7MSP4flDBoU6+vpGiPSxrjgEmWzAc5xTss27aZWB5AMZYts7G2KysnORW/Upojqeoq
f3hQuWp+Yc5cnpDD24xPE/Tax2cWstjpYif7SWmvu/msW5ylYn+FAozz/BoNgeUz63GAQilXZf6g
mLqhbcD6UXhwdqNZedM/O8lnb/wXV9dBzHXLxgsoVzrUWHuaSVJAtYyEPXPcOLAt6Ym/PqMn1O6Z
a0pdSK3tbJQxqM5mCWcUkZoyoIhVzkvCxRoaebF1yLbOXKdAVmY2MniMz73C8lPueFykDtXh92K/
I6voBRFYrswZKfxpFGR4lPuwQayTecGYQsfAXZeO3Wnms67R66XmT75pp6ZQEUoDrXXqouPTokG0
EcGhhhkCH1S9fHy08LYFMoRbv5kvUF69iSM9hNmFPc3fbC0lcyBz77+W1FTJok3N3+ti6oJzFP3w
CARHexVePBXDpED3j1GRZfolaRmST8y7cUscKiu1IYSHOiBJFKQDAzI/sAE8HtLy3fBxHHmk8iAv
npsQOMKmenrDwiUEfCY16Ldbq5mVKMd/EoiNZ+Jxfsp5wXppeJzQ2O5vybbXkoazI/jRecQ5fxja
jVVSVYA/EX31yZjH+M+vAk5oC1Ow69BNVlxs4Mm0l3morvctK7Dqrs0pP/wGwyL8e8+lt9Gm+9fp
MRXV5AiOj4I4xEw0IaDANZ3MRsn7yxSvlrgi/0ZWPblpJ5hIxty6jips+RcGrKDJMI7GYGKD3YsI
sq7V3H6Rowe1WBxr7jr1cSwK3+V+/z3OiwBLlsbmZbP7AsykqKukwfQkp30IlstRtajuOlKnYzTG
yUyMirsrlM3xTued2JF4i+XglDoQnM/jMvONgfDdP7BDZqpbLISgurHVw3MyPUH7+Zzxz9nl6S+s
xNJbCskctkLADx5nqrn1JHY6XZF7pZScm13NdG5G5ZEg85LCyDLNE3WxUG8qbjQcqyguttngPOtg
3DfoxbPR9h2zzPqDRXdVPhndjiAvS4tBkkJP5UwU/2XUT9q0IysnMLoMVRylKFGR+HcS+3A3cVuN
BQHI2Im0/eDAdI+X4eSEBV3roWffEqLTL091GRJHb/O8TSgmVhHxHjUebJSuxPlp+WAI9CV3iOtF
HMPN70ES9gl5mi5VQsEV1Du17YgzFgTiJ2z5TtpzZAgOZQRVwPXIT1BFOdyhCJux7x9TSs5R/Xwq
EWPT3+KsN5lrwQzqwhg21VyR+yDSlcPW6z5wCQTnzK7oovFPLMVr8mKjC7n9NTtXWkZctbqN1W9q
UR0HOjpVkgIbZEETL8sXM0EI9KWyUwv+AyAsHNS5xw695DqszQCJV6ZDbxtmsYxf3GUNzi4eydTJ
06yvrW17l7Q6+Gy+oKxR9mxvi6LjGSrsx8cDJcdjg5B6B9XfKUiLq1raZmElheV71N7wQSeBdaKe
90GOArBLjTr3QIyRfzR7ZmYndcgvMUA6OuyOGE1UShgO1+H12w6jzBZB47QNjqMTy6846HGFbrXF
xWgnPzetu8eMMfzISvI7PiCT3J7gas3tA9dRVULdOFldzl0dXctd0mUL7WJtMBBqZ7ZbEjwgQoJB
zhH3RaUUVwPuWlAuFBl0yaU49ob63uDFM65VxO2f9lKHm76wY7UQd+6xS4qGzWuQGz/JIeAq5VAB
UoHmTh0QUx1TxXxCL/eayy91C9tlOSJfTtwqiba80yOMOcWWgkNLIS++eGpn4stytuetDnFnIZN+
59FnxfIAhvZ62BkZ06C7HB8Jz+IeHr8HsO9QljRlY0PfsDOBYLJ5jwkqh4JnD1kRKXD5M0fIcpRa
M9URmDF+Yf5lFl+AczYT3yJ3Lx4K3e8Syuu9Pi25f+v3pdXRPqiUXucCTrPsCPXIXBK3G3wyzn3W
xeT+ZsoQzvaFqvsPt7XBivK7yzJ4VpZodQFlgxUpjR+DH5V/OnRgRunwikBwqur1BRnz8imU4g7n
xdfBVX4uDYdzrmgoGVoI95X8YeFzdCK8Rqp7yZKDGDpnrAP+X4RrQdbdGHZ2bkVB5ugAF8/f+TPJ
vzTI+jL4wzWKjvg6bSox74yXCeLj7ETul5DtnzT50oMeG995cD3ee84VzeVosDAOw+ZzZCEgg8u2
jwbfUzq49GGPRAmjnpC9jqpkX7KHFa40xapxYKsXU0FWgSKFcWaij+Qyv5m/eZ3zkzE0ZqlIjzTo
jviFxo5SgAg2lHeU5N6lQeJ4muw2b3BNKuApRWb/AIp27IVv0PhWw6Rq3G1g9iirEqKcP4eDCxp7
NOtqyNKBOHVTtQQOcdmdH/RG4ZBBBEsopiRD8TbFqZKD+dzao+hYzD2qQnDr3zllJNZ0ObiSVwj3
6XzAIXMANPAmBBKW9e/xqtREyiCWJpJtehwSe7bHEvvvRw4hGjUZIts/gaSdu+32X53UjDJzEKA5
ats30LoxUgqWc8tGc8+xT2ANhoEtaT1XS4ds9m2Y8816vdG/oeGlVJZy4lvPb/3w0zjy+2bclsmG
1RST/a7zMIOhk/Tw1OeB4RWsrikFZgw9SBbFhvwKnid+JR+yuLBwRGn4Fb82eS5BM0cTMPy21lG6
vLgGUgw6P2hAqIi/zYqXQCL+C7EMJ4CA5Oi6oJqOgJejhZARJAU5i072yrmTSq/7+iRW4C07Dpe/
MkFx4J+p/BXwBTymXon83wlBkAUaPR+SNsZlUEGOxG7lNNCwLaqgxdwOQHr+RHZCiruAAo/NQ2EA
BBodqybIzt2YzNycTMjo2wKkkiMrLtVJtKTKoiClYq0P43SGqGUyBhkZ2i8AuO4MKjoEdsuOLnwI
0vCKBnotoUjZ6Uejjj3oQc/cpuqYr7nXnKi0Dt+lcNuUufP5iZ0BNtTo0pNZ36dY83XEwkUPUTP9
eTBWqTkKoNau9IiXC0tvTSPhZBwSrldgoLuqsGUnDf1GR+1tHItDSNe6o96/zyqBS0UsE0IUyfyw
akHzBCeu0mwBFNcEFdOp0/asmsJ+K6VgEDqhmjj31JA0kGC/IEK6P0HiGSw85GAB+rE4XLM8t5Hh
ludBjtgV67TNoiapt3w37boYPgApVAj+9lAcEto9FGRlgpHcuzE/UFo19UD38oTwtX6FaHlv1Rdf
oKwHO00po1jfmkDIopF21wOZOEnvSV4m6flAHAK9wN78huTEsTnTTA1Kwmg5ln88wOis4t9i1ZgQ
LaOdsNTrrHi6dKAk0sCms8TuIptC/I9nxAG2CGgyh6xX2QkEVAXmErxVjg89GiTUm6RuN9mvFYhg
qXXKZBuL9TyPqbjU6foVLdI6245SkeiY9WNGkPFhtx1ignYkqkB2PXQZmqhKHap6tHeNxmrVz9jk
AU2f/Z/90N8CNfpM5XiVPZ5E7usgvwHfHXba7LXaIIYZAfwoBbI2HBcFT8CuC+quWCyoaS/RR133
KkcHASp7Drm1D8JkcPXNw/RZ+kwjwTgfG98BIalsN3J6ssYQkkDjHr37ntJ6W/e4/RPA1f+QwJvX
PlPD2P/oEcZpknSSTJlDCsyJsV8sp0olTHPBNVNX/bny2LIe3hWZQPYAhyo1ERKPPSlkdebQ9Jmy
0Wa15y9l43KLWu3sq2G+H4meHkXFZpVTWUAEXYuubwMY6FrxFGEG53N9NFUWS+K/gGHMnsATQXLj
tVFDsrNRhf0ff1IM4A1Mg3/og/bXooIC9ZtcvziLSAH88hSa/OUxYs+s93V6ub/hlxkIm16rgNqB
JqGIxTUnGDdMozH98KLIgIDTCJdkNJhtQygXh3lUSxlveHZUmfAeSxrE4UfNyzKpnHa1L0TF5zbr
dN9LEdGUGJYLlpGhpkMs3x8HYYa/bESQ5AetMddttENZc6rCCRziv0ZGhonWa/bX44AV30LZZ8x9
stm3mZiYdws7A5UXt+mgjF2aJTSsOqtNQgzo2Q+PbsquLA4fwd8YrQw/g5lJ15AOWgc1c7NBHNdG
XQ7gL8DszZLu3YC3b0usChwNPxK+I5c1US0P5kpLN0aCsNz/UaC1hg15UmxIhrrhhWavzw28pwGH
aPUZ+QOuMnA3nGG4s70pBRFFzR33iiw3VObYHv0G/5zDDyCGoLajDEYVTjq6JXYwCTUvzN6eTMx6
wHKau0UBhvUrVzJUrHkeyncXasTddLRinsJakvE3Awjumch2hWRDVVf9c66DWHbq2kGNxPLBIVYk
gJyFQMjL6OYmZU/LrZQ7GuL/lEWjkdXwoHcTbvONbC8yJ+airPLlX0WSDy2JNMfSqaxjdMYGk3xJ
K6rFRQgUKT+DLalqHcnihPuQm3M5TJJvTBwlmJ62lrDviARa1CFQQ6oToIq0M/rzBVT17S2rxBW7
N/nJU5xZBgAwmgw8oe/AdwqrYl4RrhGGFfQ3d3DJ0dqyJFixkbM1U0zQz2qPxAY1bowlZSGwnGjx
IiM6wTqM+eXoMKVI09/ScZgBRt1VYrtCAhbmhQ6yWXattj5GF3AhkXUKiNAN6PK/zEEKu9Xt5S2w
HDg3NbpcsIddwncVcQ16sU6mEQiIa2Bur0YG0JjrmC+uOIvNHtK//QPeWQ/SkD9Srxb4iJmcRfZZ
k5FM9+AziJLPdaaPBHSc1K+2oZZFIbG8kiyntuleKL/Z6lcjWqq0t2U1ktzu5BkzWqeciRbksn/A
6psIvUMPX7z6jTCpen6Htxax5nZ8lXTSt9mh58TV95RuURZC4ZGef5WpXOXjxd7dNSTThaILph7D
OvHZJHjgsJPuL4W8TCO6/tMLr/UQHWUm4IqHYG57bTu5SznfLrTYP5Fu/m0832jWiEvVg4zOg99r
H9/Ne52MF5gCtJ1f6JURNgoW+1fGH2aiwXb4ybmHO7yn59MNiYizLJVXrbaa/vtB68NMUH63dzfA
XgzVCwHmpMaNAH6UCMzHsm2gnqq8ankvgOCuAcVwTPDjOsAIyOUmuKWuyCAAUTEoTnjA4PF9Ntyp
D22vWsGVYrmGqfV+FNE15723BIdxirB7nxpIu7ty+ekGEJ7a1JBXT+3wcKbIXVNaly0UiReK9RVb
WhKQjDNl5Kzl+fksdS4MbJijg3ZN6PidrYBQMgD4iTrriagwFAxM9jNtHlzrD/Cjou0MO1CQ3nbw
gNWoxuujlWl123gKNs7s0sbWrR1TA9wd9jpVjzjyiCq2PX1eZWgGiaoUj2RP37k72T5nyMlvpkIK
3ZigHtGoQ7F/HnePVjZAMEYpx4bdQCawQwBxpBb/FhKRgGYqd0a1Tk5JLgYVD24opYUyL20l2g1Z
X3DpnwUyrR9e+OqYZW/kMsY51aGoqcO6LoHFOwWSZmkw/zgkuraUSE4r+5AScwdXdVNqRR24D6xn
49l4nzAxQyG79qU4OOIR6uJGba40Lc5OpIqZ3HV+zH/PRiw+Apy+EZlDqIXEerlCH7T4U2LlXsDn
1lQNnRq0yGbCKIhC9QFCifQ1RTbH2e32wKV/bF73//KGor0lrS2fxA0lMtyIEkZObKy7gpxTa1bp
pMWQV6rGHHsLCZji3o+BaDskatZGLmaUkV0IOMn+ejO2bYB4Ui1fay53H63XGiQURHN7729VApzk
LLkV3QVwdlqtQJZsH5WyTWXtylgwkazXvLP5qiDTga87V/ea8BkRcPWX58sbJtZQdoBQ7JBldIOS
4DiYPagEt3YxNPN/LCitZ+cghMwgA1M9dwcpA8Oh2al0WsVopfJ550QCU+0toG7ZVXhGGN4LqxUc
a4bjXQfMws5Jjtj4HkTzdtwsQrfJpXlE9ROCIyOrSvhQTMBz1LsdCD7jPVh2BxF/2i9zh0VxpcOJ
DsUDXphMY0iCJhrVrcxVjgk+oYAHHD8CW33/aRd2rE9nf5+6G+r45MZZek4s+TG2cH7hgZ+O7HwP
3z1DjFUbtjis1FttindaRg32yDarFutnvMduKNmDuwyOfD5HKn50N110zx0yVopvLb0cKXMpZMxK
F0NGO8DkbPRMz8KwlDx8TAb5sN1+km/qDfpX6sY3CdDisLybvZySCCLozRei2V+6QHwAqxyEABXy
+ri+h/ghJ3LgsRITfF2fqfzPybnArwh39wKvVTOVsrReisAXe7MA2yWRjVaxYEN/qhBB76noKpwd
DXqJ0ezrdel4zAg61VbyQix4H0JX7lrjxxZA//0wCUike5FifMYIHSt7czRGqAIgO0fXXg9XEwpD
fFGCPw9hUJa/8LANd9Rq9ziwjGzvjI+kNsQIxst3/1nL7V0sT3s4SJrSlhW0JPROVUwPjHyV/xie
wPrYXTAj+M6oDJ0oyWuUOOnu1yISGyN3XIFtp4ZhyFNkNV+6VtgZjb1q79BpWuiyymDY8YS9KTKl
nSBPCs6CMec9G0cUYOiayvsNe5Fo/FvNG6fUjsP1pEV8uzT9ViiA/ehVxwwQc6QB1pqOlyD77FPp
PUMY/f7ya3wEYlxi85R/lkg9AJ+bEJYzMgFgjDcgtX1M9QdW4XALj5ZWqi5yPc/ZaVMf1sWtf0w1
5TnD1Dkde2oM5TO/tsbJX320S71sK3mEYoE07ydbzyhShiejN5G6yRwYJFqytbLcpqkvsquAJn3U
WwB46ApLxe0UXgw/HLO5HLTqDaEcG4bI15XSCmRK/85i0eB4RTuGhLMZ6gRuMqrvRPgAJr+IEc2a
vLuQkGs1a83Y+c6GfgL2py7nWyULC6ktUmtGhvhDzXl6ds2NQPtfIeSytWdo1nfazFMXuWYS6aZ1
B4nbdj8/p0qyv0gNlnuFsRdE/l+dM7Ypb1TTVf7Q5mWJz5guS/BMXvvcprOgGZ1X8ilaMgG3abhk
SsyN9bVHD2F2sWKNk5/qiOepmV3fKSQBaNALNpRIVrHz2hHP0eSFgT8lySYYrAEPfPVlHhdInGsI
WJXVzCyRC2UzXlr1UJPTlWHwF605KHoimF9P10R/b5L8Acchg0OnLLAUVlYJZJnAWNHoq8FEGv2p
VKxB7G61nzuCy01TvsguLpOfjsqX3i+NfhswW6iOXUMKo9L6/+JkBkgNAhm1WhppH4JBZg+rJ12+
/rs8f9jC+qNoPWDo398zyKi5/H2Ba0qrmtlCyMidrwnMbxFuXRDqnJv8+d32+DqQWhNAvzE4IFXQ
Bpgly0kcplZCd3gLNMfm3mUdi8CNoEZ+uhFZGoi1qj1rQkDFp9Yt52l7WhdWXums/+4zGmR5XV4L
SyVF/r3tJX8BBdEWNTvA14WjZb7M4OVUuvyNspeDkMmOwTDCFip51CPJKjWIj4DLmnkbEby6t/63
nzd+uDbPuM4OxKPzdWDAvsl3l5c5Bow7OXVrT71dYI+ylU/3xOyes30OBuWjxDV+LxDreja51OLB
57ECUpA7jAN8rWlu8lwjwJmpKY7wc5YdAM/dQGpvNa3KA2XupLN0MqtHPDuzaWFZGEnJ3+4Rs5E7
NFacPDU+GzmAQYEpQ0Oze4H4cwatBZ2B/pWB64rsPlsSoTgQGID1Dq3utuhbpWziw8ZlL5MWI8tC
nOBpuZIWg9pjM8SUN8NbexJWt60bUjw6cAb7kAW8lxG9Ih5WPdkHUi40pQZibsjaHVg79nHDsx7M
R/CsAXgvQk4roWGBPUC3qm1kzU8KjKEGjw5DEP6BRkSbvNvxbeYNuWxn0nBwjiaiW6heQX+mlXHn
vC+NVpi1t/J7pY8Di3iDozSz12wxwDm3pdAQPk09xHVigvUH2kbERnf/NtRsecYGZl6wj++IgEhy
lvc8J89lr7zjIelNzCCvb/pYI8iq9zan2Xd3R6CYT4hRkTeG6xJtAbcUd8S00IE3X9trbGpdzPNu
+nWBqBIuC4ZoYistPy/1FOgIHrbZ6fHjYvFwUuJbPK6oIAxBTU83EUmV6uRhjFupdweITOHorCOC
ldRrSt0xdL1ShnKgqBttMwq42BMNCTJxGwaFbU8RLwLHsCkJ9rVbk2Fwv8+2wGyZOOi58wSODJEm
b0ZvkJ42/bkm4GLYuQnLCD6vpDP3TwWXQ+rfiCC4JvtUa2G1Bp3RUw8wOA03oehtAEih+P8iiBEh
TB9WKTWl4VrRtN29SBXO7g48XxywS/pbjFUEkqeVwF8+j9XhBM2S/Ju1UBk+XgYNzhjeWI4HryBy
A6MEUQ7QdzfXWXGJUocxyy/GcQb92fVbu6yRA+c3ER35vpaLv4SbNJhwEjgAVxcam3ECX/2QoIDd
jrVqZei2RqPS6QJ4nbJ76mCE3iHZTBqz2B0Q8Kip7/d7wc/LmtxXyuZZ2DRwOduQ7oMRSa2FwhRY
oAxPYxgWYGEzFdfckjWMo1tSSxzNAYNazKyUsPNyILL1TTXJpK0wb/8fem6wx6DRhzljIZjNQxoS
NgP4erLOuLPOzaySuo8LiUxBE6MkB5SNhCx56VSRFAS5I9eeeBXScQwrHNofwHAcZfwFc8FIYWJ4
LhGOTzgGk7b65mGsZ7Z++AgRrPg+2ekL0pGpBU1dB6eZFdiXwr/iSXf559HJT+Cxt9CyOLfsSMmA
NgtyD7Bt/JWDsWB2otHS4WNvtc4ppWJhclPVW1+pHv7FIy09SMm4InWkr6vEcK3ghCclbmORoKYY
ScaAZPn5gZNdRnFs607zp7gmrkQt9IX6YCJOJMofl3fwFFXcJP7DcbDVvHbtUTt9Eadei31cxEtf
TDGD86SmTyZrzQp+wP1TFI1O3QbRGp1EFzbjY5PyhDxTntPq0touEWIPV8PKi9mqSpa+e22UASyP
pYrvhyhFjoomCPAOm83YduXBoUr1SJG+tS4CzErA60/Zj6dXO5sAUQk/e05nFn3GnxctKUXTexH1
7lEQa4l2J/2tKHVwqVIVSgw+O4dFIwGI2iiRqP9ObJ3xN7H+JnWbKy/QxbWauShmKFN6BnCafdgO
k0QrnO4R3FBSUD9RuDaiweRwLE3+pRfm6wzUag0zqXgXQs0LmD/b2T0uZTIzlCYcU3Mt4uj+q9X0
BsvvH+YD75DygIoEnpSE3sWczVbMOdYn91PfDOEGsJdqvC6WvPhnJ8EJNf8t4fzbK7FRi/PCeN6V
O30wLMhzBw+EYJ5E6T0I8fQnRdWMwm6/wV+3vveNsL+0T2PvYY8rFitAXqtYjAnsOxgrCoXWOoKl
cEAv5FMFdFSHpyFprzVd4fIQcvEsH/eWgDYvEgwszvwV2wNSUlMD00LhtOB9Ztl0PZNeezQppIJe
zHz0UaZ0s/JIirn2n19j9t/oDvZT7KICOcN1PNEw3BZN3BffpJKChv6LdZ6Sl+ECxHzwyZZ3TGwA
/00ltLi8THmUZCQ4+DHc6ZTlMDpi64bYKVxMOnXNFB0LMkEqnrHzToLEmFO6YWipY4kuUYmCVn91
9Ker2bf6FPiJ8lLZBenrkoQC/ldtxsCv3L38xduwrIg3mXhNGTDWbFrW+BeZmBcIJJQZ/fM+mepC
NH4XnJlI6ZZEVgbve8kzCdZNHY7O0vI9Up72MDIrNoZB7lVTKGtZP4HS9WkVl7j1CFCeONAg7XoN
ReYRp3yEe0aV6wA+GMS6n40JLQVuXk3FCjhSHDv/7b/mWK/WVqvmX+lAfEnmX/+UxbGRtjywlB3p
cjPmS7m3/QgGhezAI9LoYmkG75xQR5tyvBAims/qWFnmyJzMI/rLECDC+oLmQxiqOsd3j3HRRh4r
ajhvY5FAp4+o5qkE4uaZOAUoj0kT0pat+iTsn53Wy3tJknlw6aXJ9dflS1oNDoDyvxo7NWW0by8r
nLU+AIAXsWiAQIriAHAfoiirGvO3Rwhbbi05HEVBelCOMDCjWD5TdvUdc8hdbfZvWZdqfz5ap0IM
xhWBqk1I5B9gJ8wh5HjmV40gQSmP6steyGwslh+HHHAvhli15cc8dhTH47PyP1JwRNs9OH81gvLM
eY2gyzLENoO6A/NLPBmOM1ttbOqu7UnBuRh9URAhBmwFtEe942KiAp/GIE9iYWNOPxhEkbsfPmKZ
hYd+P182tYXJVKGgrGNMktRwCfrFNMaIBp778bwBdLVkZBh/k/wF0GQmGpn9OUR9Ze4oZF9kuFkl
KVn9eEbOtkERIsYUNuTI3zLfQC/SK9U2Oey2IQZSlYzvm9RCTTaRk9yEug1ZBGS5LlqTZXPoFXXo
6MuIrXSD7RcUSVoxkfVs53XTm0bz2fGw4yCEHHB0Rc677MS9fnRD7tVtGTaLXTIdN69cjiJc5R3F
P31wYwXgxjnE6Vk9y6JRh2LLgeASTVi61KfZ5MnekWI1y3hnUho7LiWJG06xExFHdLRL7Q2c1wxt
b/xtYYIc+6lqpXVu8prT3H4daFJlRxyHulEzynczowad3VGkMFk1KpHrChpWzB4PIszyT1fLRdx0
eu+zM49WFAobFQmtBoabkvmvcca6c0dOK/Q1AftPwrMrxJrocMWfoHID+cg85htb2E+ujeUBooTo
RGq2pCRRkegyX1Fqjq7iH1Xui93fsyKiRmT9nKH++2x31bpVl2hfIQLDoDqg+ax0cjIJTkFcih6m
rIxz5ImbCJYrO51WmhYywndh6Ruhe9ExeVs3BoDjY7LNjxDHZSJTEveXO8NbdiHJDn4ib9zq//sB
4IIklSW1OIZ3TOIUlReXx2cST+PgfZrRY5NAujqbtAqqQTYr+fcixOesFqyfJoovW0eAAe8aMkMV
5c5tjmoWVA5pCbpP31EVlSMVLpYomvTw5lJj4EiKD5b0I5wa/hNcczybPaQPsyPu+hAbacMhVIbN
T/01P0q6A5x6p6RuECRNSo/NpMaqr+uee0IpSPgF6fYeQzyweSBNFjxjDxqL8ZZXffJ4S598yBDP
GeBULUotTwa8tR0WP4fk/upCARXMuP+ztbJbMOLyKxbBrUCFbKrAhWYL7XPBD0j+7if/B4xH+ew2
1/IhvWVRpUfywXs+FBpx5ZWpkMGEQ7FbU6rqNNEWglnIn++Bh5jmBFPZgc0kYb3nXn5OurnhsBE2
/kURTfs31I+3hS7gZwGsvjreuOJsfKvJSt5TIjslWEr1/1ODGlqETixy+Vkry0223uz4WGwgqsjb
Zg1zir3Fi2sulJWnGML5Y5ope61HnrE8QuMrP0CHgO8jJgUkgvqU+L7rCZ/Y17iCETUqZQQ5JEWk
volTwJZjZuSLjx/RFz+7Gif2TFx6WhsSozw8HgGJg2DIflSbFRuEAyvAB9CFfZycDO1AklEwoIt2
fX6JY4uqGiQ6sz/G0jPl6PQYefHFLtHaXxsh3CjJJLqiP/NIxBXBo8IVp1bhqqfD97cqOfPD/7K6
V5aQudoL3DP4X+z0nOSG5mbyQlFMU+pWuS7DDFarwOkGm6XxJUEi8V2evn5u781E7k43FDhli/dZ
dYh8pTKanuyuzRAMKaR2c4AvzeNrgAqNZ28xqfEZMY2UZi3mmL/xhJtIUgb0FjZJpp+IFscyP4Dw
vDBMJG0KMutHyfDfgQq/G5AiaucxheXjAkYKnKymRsgNy4ACTFZ8hevPKQmzgy4JkyTbWu/4IZsg
EXBpEjkwYLQ5O4eBUU2mBRlGyMLasAMZcNo3soLYKP2L0NcsN5z6jo+BgBKJINQzuqldGGEIqao+
DpNikjyi+ihTqp6yAN5laYC4LoZnCCnf9w3QEPCv0MZaX+MY+nJyeofxPeKx40/cbX6NT0/bzM7I
laN7W5uPFIPZufqeuZioVH5VCYrCCWKdjIB944DjxbZLbzauR9sJ2F7hM4wHlHGqFpwusJGjAOeB
siKv6WWkL/pnQbJpbF9gsZgldU0TbhVY2Igqk3hqMM7LE8NO6i+aPq06CxXPtxJrhOq4yAgUZewA
SKFpXra4Ph0YbCf8wvgm0YbiR5nbtNvYOKwnxjm017ZTGTZNGVVw98rQU5C9CPsV6LErMXtqvQMp
jlAX/GCbMKT4NSpBt3srhav2sKPCrTZoDpmPYBEsPLVNIkNg90LhfPorD9w9oCS6OlrahaQzJaQs
loJJp9nzIFa9K/cdxxw3TVItmHYuXr58XJWjhwaT0yrT2ylqwn1x3ySyYpF2YZp7I1wFh9eZX6Pb
nnwu7oEuBi4nPgoe77+Wwg/eKeao06P7XsOXtlTXjseFzRTGcMPMywgmSLFinVFQc+R2e8KvMuZ+
yrxYKs2YBIO1Cl3DrtGF7mxhJC8yVDSSfcA/YY74yhjvHy/Ay2n3BEnMezn1ftH8ilKvZGOfA57m
feA9xu0OICdD7eXi5xxngA+38uRGgh4gyNiaMC/oJ+ICZKqetMIlNTBAaRdZO1GoRLt8DFtB0MK0
fUTbTt7/HkhPa9smT3SS8SRVNrA1gWWrVRYhCX04Y3hXIv08sdWZznDnKbkBDVganLk6ZdjIIWka
FIfNUZ8qV7A/fx8C5EVYFKz996QRAY/Gm4NlNO2tL+GgkV2TPyanmebE6IBo9Px9KdEtd4iP+oLj
AOf7yMYcR5Qsq15bvPoY8mrxJJHRvmV3Mfr08LkhvioDus38jBSPD/fRzmS7RrFJIA18kGKQmTkR
2DV5aWMzGoWESJdZPF2xAdzl2cnf/ULvIEO4KAMHRlTpg+bK91F07WQIw/Qxk6FSzytMRh8mnV0g
hM6+DJQimGr7LdvoHn7eXEbGIU7XCYPtzckYsS3mleV7s05bnecSJd3IbsCJz7q2V1bkGP0KnAcF
5MrhVnHhPgCHnm5m9pitOqc6oU9nR3HCZgQPE6Fh7h5MCjTMK0LV6THsQ/Um7Js4j3MSdyGjq+vk
RvirirI8c03GwOynyWWIGMoLvnZ6MhWJv74rwda2hav+kou5bNkgBBOdu2UcAbJ6IZzzaNhCcGaa
cl51ufhjivhD1eAY9ZdEwrw2Gbr9llWwAt/5iQp+tjAq5DYJ0gErclGbTG4k5dVX1LgLsktvmyxS
hhFYvaddSpslSM28IMFmxyfBokXQxGtxJNBgXdjAGXSAwEb5PAnzK7FG8hlPCeSY0H/kwb7+92hs
1fnIMrCFDLmBwsXoyyzHNr80YPP8ZBoSEAD/yUxvKAVht6wT0eU0I6Uzzov2Xq8JcsNUFjgoR194
pEGR3IEDCfpcKRjOII7KJ78jmw4i00Dyl6pVUWjvyo5km5NSYFnRyHsiNyLZiA9O6sF9WlQzWTY6
6TcQvZ5ErxOiU/OaM+Yo/6UrSNj9Gkt4pfCA5O7//URhBxWesHXmL1xZnExvjyujkMEXJmOKhtma
UIseMYPM7AAEYAoc0YtPVeY/TDsBDRCE2FgX4eS+8/742YHDTFovesACBUnT36dIrlKHEH+4TZ1g
fQ7sEgn+tGNficb310INzp/xJNvPOkPnJJmujOZBDDqQQd27K/W8vH0B/HrnNjj+7nhwTDnF0qGr
EMnSc/GIC5ukqKA2eqQ/dQxEPDIZRjHKS/XCeOa8N3hdRRCJ6E3pLLnr2BMpPQLkctyDnxA5NCyZ
qIvzgHiGNmP6dF69VUt1AEo3wnMtc/IqCcUdbHMS2CdbtJ324qJiEc/1PpjMJ97vFp0OGZYyW4IZ
JFfXX354LOwgSWBtxVrZIK5W+eNU01ywzijyS4VXD5fVeyIHp2d8c2P9iQLHSnKTsVJ6VeYfWKLj
9McX5kBPtLEcU+SSbe+E3dLWL6OOmtQZDXhXfGgnEvIte8EAZdeXOzV77CwzikHmNGONSgATNkMu
d69vI1trGZIgWD5ngFx1Gp/GWxsU29q8Q3IJrO1t/L1kAsxM+0UYFeXpvejAnoyx5j3gLWfwj/hz
yOYjvBSOaHmInjN+EcGlRhncvsvQDfhppPakHesTeVUg+Xoq71KoPe1tiE4x6s9pzqetdg6pW2Xe
4iEiRXml4ImDPNppbLgQU2UbVoOhtjeX4DzrSQe91HUv+d5HAcudxfi2ydD7K7FJ3OvEjC1SDrmL
61KAv1OYDziIBkgXZgeaE/Z6QKZLV34w7vzVi4DOj6fwnqAjDRLw9h7NadxkFpXxYHL+BFmtNO7p
zIYNpANNfcCO0KBaVwAX4W9RYrK7JELsUFhQjvw+hqEN5m92+1cLMSFemybdMNqTJiaYPjKYpm1i
SbrtRKcjHjvN/L8UnvXywHl/beGyOk+LTyC9FnFYSBysBN0PNOxkwSHxSXn+qvj3WcV/dqMkYsEL
JAxBU2qCK+B8tpnXMjDJrfUw/VjFM4WDNXbluFTcQozAXY74vfwPRhIy/1i4XZDk9AyNWIDGBgj7
3JxMZeflSaqzYfMdhUhsQM0GhYoX91NzmnUeRoQ4lnvipEN3DokwEpMuxPlR9COfyLykMxPNwUUr
QAQi8xGnMFtzMrNVtbMrlAjcx4ZH9lWFGsD6UseqhUQ5+BpHjsE7Sy2LzmQB3Os90j8ZNnHby9LG
niAWE5ANhv7J9n55TGj0VFAb20Roch22L/jmSxrbAy/B6Ja3Vjf2ixheeU/OIpOcNXOgFQw+Lh+B
Lr4ew3+EN6ZouYNuGbIB+BXQ13KFj5gbbanBPyoRJ4sRiNja4G3oqpmjrT6pXzVodGXzjh3ji8Sl
gu9/ZlFr+nefDBROaXTM2g9MsolEc5oxGQYf5G0Zy2nEO/XhA78zt3Pxqvh7LrM7e0i4/UG5SzHE
xl6a1odD+sEHGi4e9H0qsf3K6wYb+jkiwR5UPJ5P6E4Z2xWr7TDPJsTE7pOp4G9a2+nv4mSD81W6
er/tHXuOC6q0pNxbpnzt7pJZ5cHrsqGGF2shJBaOGKsKZe1pCO4LR0abzOVDoAw198Re69MqMEJI
H78RINGhdCw+8smF8ZlYyOcVQ3wzEfplJ2ZfMT393/4TeaMIDGB756xVOaDjqxwp+F4HljDMjfwt
V1YMIbqm+VTT0ncLscZ6YFvz8enx6Lmr9ny+bP/B06+Sxxn+6XYEqcfzOhC+yCYMw/LfeQdZwFRU
9hx4MsS4yb7EezfURg8dNmfqCYlvu0ZZn5T2VcKBW3fsMEWrWvDipEskyjp1iTozgaLIiZlBsvsM
V5Xc1h8jK09YqbOYRe2OimzFuEruZrtWPMe/sJekxMQEbRo274rF3Hxae0PdzGAiMQpWXCaPPPr9
ZB04UxyNjGYZiEQgkChD2Mt8QJDTPzqtH5cV98rfy0K2veUc1sTTUzPoftjcVftrNUak6kbEUlSj
BwGmZdusyRmoppoWKJ18up9YkWVjserJ8Cf5JTiUq57bafzKpGh5bjA84kLBzmOzZTl/k4IKbDsD
34+zsxj0tI0Q6aGb+ShFOGBTbstF3ndcDbfCcEoDSJfhM8hOOLKYYGIz0w0Py5VR7/Y0HDF7yd+D
kQIOAFiBR8P4CmgFJaFmaNfrhBLhTdw6R4SGJeoS9CnUG161/G7kSsWG8+psvcl+SMmZxLtDSlWY
n3wKKcfuVO0U2DgMg2wXMPwDRr5WVHVLl2KM8qGpjLNnZoVTBVg9QEbUc/QC0U3PVY0chX8Kck5a
cVvI1mZ+j6UgQpI/vIULH5Mg2uexi3f3ceOFJIULS5oMEVf4/lNbG8a5qWrH0pg9QCr4nv5D+2cM
LGhh/+Vsxj5uN5JG1c6B0aw6Qn7TbH1KIf4+dXksR2Y6iodUMUnQHanAMSKsjNmLrx7cEFx0Q+0x
6/2Ry2ZVAtcLad2ilZMe02GgigJbMYRyqHr7dup4qCHay1Ac5lplI5+mJyS1pJjd3zRi6jFFb8tk
V35kgnmSrxUw3UYh9gaDmSp4uG+qYLC1lulPvrgm+gbaQ1zxIPgZ0YAvEr1qAi4tvZdhAmEjpG7x
PIHOlYJgbW4rL8ZCRWSFLmHIoLovuu38KOSVOtyVqRB9vHSERLO1+7fmot2LDJYEUYcN7jOYLeyH
TUCLUqbnBj/qY7V1wpu1MbKoNVHhybb+XEhlRtzn8YNG68KvGp8Q/4V2RjcoQUKJmQyEHA2WKZMm
W+egHo5LM7rs6rCz0sPIaZ7+fSwIWkV9FqfVboNHouwGCEepmIF+vfr5sUhZWUwKmM/P0qki84MJ
4P7SJScXiO3omVG9fcXI0gx5W55UzhXfFHaFwViLvqAXtbWmk4dQYI/bvHMySwe+OnX+ujjC3tc1
z59SPZglFEVi44H1HIxcBwwZuAXUAD70CnibIIX5X+YjVkXBFRQYo9/T5oPBVyAQ6oqTxEpdAUAm
641nIkEgPI8WTLkxQEyYhTKRS8fuYgcsSktQL3OATLsK0CDw7e8RzqobwhmIVkWz53Lw8L8oOX08
gbMQ+hgp1V52+pdhoey/cFtvCoWSzUFBlcLWvIFlis6ZaLtCm539ea1QlD9I2DXce9/VyNgEyvIM
JZZzumcwm1i5AKBEMw3JLzstBM/UFctGrS2PjGF6ygrly5bRrkXZJlUzZ7gXCIGhM9z+pW5aAcFH
N4LujjYIm5NEpAAVC91F25PAaMuk4ecfO9Ik1huooIaY52xmqZSlRF/hT8ER7xfh0baesQlY+2IN
5p4QkWOBf8OAQ2cGXU+YnOCGRZXkrBugzdH7PWGC/rtw8DOiaLVzDJllyF8yCzX/hPx3t+YmCgng
JmryHMu08LVBgruBupEYNzkZchLmUUxXp+ap5qdL2qa5KRGe2oMNbwx0WranlKHu2K0ZDsfcp/gQ
uiiOxYA3TrMsJiZYrYHvVBfjuRyQqFXbm4EAgfauKUupn+uOQWLL83MDK9vP2ibK+AKnr5DD4OOt
cRMicBK4kC8M1oPMyU7EOD1MlwUt2LWWyIbQ682SKyXaRCLEiBtmMWI32JIpoTmSiy8QJffCCYzM
tOG7DIYVzfuzIXxrZi1FL050jBjrJuxv98Hyh53jvRQCqTvcPo+bSdSFfRRFHqhZ3e3Y750hAM4W
S++qnSLdSIlfe8eqnFMVYzNGGKUnQL6ztMfG0HEajMzmBHAoBJ7rqOZpdrK1NLoYaUmJXlBSSNfQ
NPENpecQ85vEtPN7aDcocKB9Hpk/hJuWfdxQjKKqIIk7hGzi3hxxs8mBraZe2fq/vbKJRAz3/HOV
d+rftRtA9L42Ffy6w5TJoKx6sNQ0pBdZA8H00Qrh1S03/aoEgUXgWNmEVZOu+7eDHLefk6lusoQz
m0GMQM8zoTD2tqlccN/DQ3JlWQc5VPGJnzUCFqKFJFeAXpe7itPl0K+vjG3LGIims66D6H7knGsU
Opck932eSlYTS6YF5x+1htBZijWpLmDJBqpp6SC6cRSc5r8/C4zWvv9VLP23cPAAGm9Z9ChtmOFM
6T1/JAubUREIt61zI5km5sXct/1y6K8UZi9YFUZQyAxNelHpXvp24Rk4QbF37hUA96Z233d52gt/
JO1j1M95ahWtvYJ2OYNxYJwKZVhO0ydOeTWH1Md76O8hL75TSbyF3iuigbUACKZJPhwHqe0FK4tp
ZTGnPI0Y5fGjShCho1HCkI0Ft79m/2jkMQPKAhhGZ8nskjK1dzyrwkkZ5t/m+qqTnu/UlbcNqFHB
0LVXW2S7/hRcvNq5Y/Y6BdVHfXvrJ1WDtv+y4Ij5fYcNdar6ioeCB27nj5QwB1O08FdFPjxAT/U6
BSDQ4dtDZ2grQ2TPWtzGBPubC2vzYp5jkYwgb+eDiXIl1oeFWUGD7yF2D/T1jNUdFlhvIT5a2/Xu
9OrLZiqtEvPcFfiVsoJMhv4U1R/x7WyKfA1Gde4zP/9Z6Mfj6bfHj2o4yX3CiPEplOsGDzPd34Ge
LbV6kGIW5lrJjng+k0nDpP8RBsDwLdh8GWyusxY3u9k5fHxHT5vO4MA8IahlzrvbATeWKh55CddR
TR3c+M408xdDK8AMF9Jsdur8dIY+i8o7rCGvSYEI90wRHxfXTv04YhFmSkfl1YnbaJsdk8vchMqm
pTFH5aQFUuC3MM1vvY51sVUyU48hGcA2yuVLcBXwQAWuTOT2o41EBbLzmMy1rHiOoj07G+M1tJsM
KomJvZomwmtk40dCJTPXisKgKTJaZ84OxUu845rjOc3UKYyg8s5Xlkk6nJvt96VX3hz3Xz2ap46W
xFZoo5z1NaBxfF/8H9I+q1kUOipZi1p4Mw8gq8VeAJ6+hF9DLoVZzz2SsGV7I5PkPXbN24j7Nmhl
GcLyc72PV3d5q7KbUIkcbuIKQhJNLLFpMn73M410etXxl4Fl+lnURgJOtcWuLs1rb0SWpLnC9fiA
omJqAA2D9GUJfUQInWnA/o8Qm37zvI0r6S6T4ma2+Y5hjABzdthC8R2BDeVp5x8sgkH9r5i/2/2R
j2LiI+fPaD8Uv2BIQnMeeBr0L2RymLoddlbnembQippPi3Wbptp02VwOdAya+WO9WPVd+GQeDzre
AoIKfGwPgTo074EBehWua1FJC0eao9FAIUmuqP9PLqTEJmc0oUul77EWq5oLp1r4yc/s9FGwo7Bw
I6ppZF08bAqVc+2d7m1oyRHAGVOll0FC3Sn+LNIkcb80n/PdGOcmcit636pd6UzJTMBoppj7GgfN
GU+ukvuYCKZQ9gy3g/7TKNdo/ss2+t4RQQKhKg6rudYBGmY2AwK1KrQGbXK1VauffHM3+b9RNAk4
jff/6DnRcjed3VLRwgkAMJHjQUxQkh4Pgd9BS6JDqCGS7zfSTcia1YyGQCQWSkLQUJvVFx1ZwRYu
tp2KD+3X0jXkff30eYDZakojnbFI7YHa6uAYFp/WBgZLMVUxNiE+PUL0Z7kCH1dZAgzRyDAJRLnL
MxmTtFsnF/kQ6WJ3tdj6/Y3MLDbSQjCQqw5GfA25KDpU9Rpxijmbrch7o8s9eNPjQsJPvTyFkWco
ZtnlGQ2+L5r8lVJPAp/fjeZnRMT9RAdgNZBoPg+9R2LdneXHIv5oQ2Bmr9CnAjJgJM+1fOKJ0/Nq
0zrI1ztYHkimujjstHr0QQsvwsl+h/tcAmfZLFNwFbn5QEdRNtXjjCfYc63kWvwa/rQXBFyJiWBp
G11lTOtXSF3kaZUwsw6kpahGZko896IGFxEAf+L95GNmefGpplweYvSsJYBQl6W5zSGdPnirQ/d7
/IC4Tq00P39YmKRNrzdmyAyno1EnZWR7pDpGNkjEMXCb768iBmb+LoUIrWjxKiB1Q2ciwxU001YE
tSJF15OwZKN1Q0xRu3O4eLYC/yhI1pGvB1gZhOcCjhBMyq0T4AmfpjHyOt8nhSW8ec/NdvSjq2+G
GnE4ism3WXQpE49Ms0wVVcScD5ws53fIVVnfe2EI14r7w8aNzCezga8dQ9f88xx3oW0sHr74NU3i
CcFJrTWBeSVyR6UVLgBapmvyknepnmGOHYkkC7OxYKC5aJINMiUshhlXod2hJxZrKw6TzJ3yiEXl
L656dbfFJHMdUfh1fDGEeHoM3k1I4YBQe23d8RM7Uc6hegPTb4J97v2F60C85CdnzqgYLldtg/Rl
UalFfoMVab+A7uU931fxw+2MfLbWd8k+1I9HESLj2N7MHsNYY6cZgXkcbIePT0OMte9ojyHqPu3S
+ZbC/eJ8LW6kuuGimn0f20UuVh4mQNC47S/Tr/32QOngOMOTUc9rhffV+NKDXC1kpo7UGtqXTmjM
yNUW82MEkCz7bVO4B3czArqKsyf2mBQ5zC/I9gTTkO/YzNcg8u0F/4nLsT61eb4vmng8cnCX/tI2
gwbJZgJG4a6ncqW6hgHKH4lJZ3O7SlDaALl/vkjUlW3riJkaQkxWnOSngkFPDiDhdul0011C+A1I
/Fnhr5Jl2txPGT1BOo7CjQh/S6MYIaFkQuKxvHcj+mrdbHIcVRnbg0c55wDa4ZOM60V+60tjjwXQ
A9O12JKcaNUyxkX+yxepgCsUkP58a4Nk3OyA0bSJlYyvUVbeHf9v5edLGtdh39t+tO7HWUmu1XVK
0xUEuGRUruG+QJENreBbzmMdEfSbNFKH63i7BjHowkab/99etowwYVdNPX+2renvTjbyRjkM+6/k
Oah9IzkraNCwWqUzsSlAG1jbaQz2XOwb5DEt7o+EOpMtE5rYZ7YNEpXoPiypk2RnDSK3QASrQS0y
E0bjOd6BmjB7S/MRluDe7PYYWVqdN74G2LrMhGgDevcFYhzcw9RJJcZW+xaQkDI1wq7WU/xR/Zsf
yHdJ6nFbOsqu0pUVmreBDAyqaUL7+Dg55FrEwS4W6JsUpC/8UohCCSRNV5j0wBXm1kKPe3TLpthk
5lk8r9uKR+qIbSrXeRoQTNZSc5HY4a1m0CD7wvWAP7KR0igQ1pQ8EEc0YEoCAgkRkEywG+CZ++XS
IwStRJOmZAdRVMJ8GzIvo9duftj5E3IXri+CSejgt8xRpWtXAx42DlL/CTA7KBFtSxeTAa12YB7y
U5DsNX6Kdg+MBoGM+9LskFTaw1zXN7bUYvlm1z2fnofWKyd3tvVltUXSgITb5gGNE1yTsIIj61Pt
utrNQ9Hauuq249kLA8OJis/uBFOHKfmZSB8mB3+rjsJ0ltM/oqBnzQxtZdUUyjugGhGsJcTRy9Gy
geHy7/Q6Tn3ZYnFPZHptz2H/zjJQji48+qH4KMh/TInqGWvsfoyrj/Nsyqwky2I3rzLpEeovnH6J
CTWUt1m6FtjEPDrI7VjIn0gcz4KiQ1eppS6RVttl6Af4kB4Jr1K+m/9hSvtKf6+RSS6YQn51dDwU
7e4aVEsuOLU2s8p18zj4Q9/QD9fmq2jYQ4x/wrsi/b5apHCgGJKhoa7ZPfVKkQESWZa5E575Ktub
3/5uAdKpH6/m1dtLbBw6sJ4D2f8DBUQ3t4M5MQ89AwVUn4xjMMLp9bilJObcv08meHg41C+hfv9J
9WhwiKxkazx3tI8wLY86usV2+ESB5vt4mThPBI6kxzl34QsaYINkxw9iwaRjcvA00TryJ9soqeqo
sQ3nQsA8bKxgHWC+vD+GLdnzMAHP89VcyxWO4VvLQaBCbufAp8gpL0O2ZwAgECVv3cxP5xKtESN8
LHnLEakdsSzLUikDm5KEr+ICwbxz8lg06FxwN9STvS+y7lzbm27cX8UM/N8yKqk4wfSY+fyf4CC6
HC9UNmWdt+nWmOe4D8j8WcH27Y0f6o2DOSHhIBaJaugb9pEUW9/QzbdkayEO3C4RgdpF+lT28KgU
nKZFxRfWSEHHiiayMmje+l8jh1/X0a3Rk94f5eaXHPCxeJQQErEIEZk8DXPtB62USgwkhnT0598e
pBo3ZpwqPUw1Z3H7fgtVQeEnGrmR2FQUuidwKc3kuo+wVT8TdXmwPIZpYKdEwEog+2YTR2qW1DXk
sxFbdWMkmZyCZWpgLvtL00goMjUcRGM0Xq6fko+eifXd54WJFw3YvPnzg/wkQk2ns/CUgeWZF1Vy
1Go+hwhqJ9MEXVcoOTWJmKLDRhr5Pg1v47rNX6dW5h1+qV9AyOncskqxIpaBkzkaabkaK3oW4LeD
oyWcljzDxogDkkWktgmdFAV42jRaEUm0vRItb8LLKqjY7u6UoGUb1N7jqydnpZI4TFauXttjrUs=
`protect end_protected
