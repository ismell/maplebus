`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ccre/mo4iYR6ZSgOg1gk/7yavHm/Tab3ZkZcYFm6mHsK2rs8opjY2zm8CLFAxyKzM+XWqIQXr/Fc
dQ62SDu8pQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WyYd7hG/1lw77JWK+H7uaCTBuAtJ0TBNBmyeEHZzKg+QBt3Cr/4H8z2MUPj6pZRjBIIMcBdDyWAg
kFxba6x1wM6D0583UJ6utRg76JBTYn3hze0vwLk8TflbT8BIsLMY/07o7U9RQLj+Czrd4nu/GcB9
pJ+rlEp3a0iAZrf+WXM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RfuO8rrKLN6nyJNR3MR3coxhKut1qVIAuEdjKuEt9/BtiGJZN+vho3sGPhnXGPXiGhQsomdebq5G
ubnDKN4NlrU/K/1OyNtvkXiCQ0yq0PS2JdWUylqpjwB9ynBw5A57ADeaCo/udDuX1y5wHWGkhROQ
fsJZ53VGKb1Op1Lb3r9BDB8N5YilEmUvvtSyFbdB+7psIBAUYyMVMn5URNhxA4cyzgpgQhfcULcK
sD4UNIk4VWttF0vTTR6gUts3jmAIHyHf3d6WxdEAShshX6o4OKR2UxT4uLzQata959gMnHWV1u8z
szCVxPR8xQQ0v799z81NPg3yNd9QbIa33NfW3w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vxmmKikWOvh/MtjVuTOdXUEizG5j31xAKxSiM9Xx8aixITyV/shFEvsvoImS9EU54TgPNBdxM8IR
npEUXOOcVxO9WfGzwhZNQ/ZK0jBxGyrb28doc6RBBBRFSLq6zp6eRXW4db+xriK9oYHqwZlnFh+p
+PrqAo/I9KP6sZv1oHU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kSh8dathlvrCSfMnDfy+H9hBRQczNUVPEe4uv9JEwCAa3/2S1CyBPGf5gqqXuNXvqHZolzJIX/7w
pSnd9F19rFWLAuVfzyaIPlTZrAsax9Nea4XwtEczdmi61CkouLWxlFuVwoM1bzkNI5RFMcI3c+mY
VVE9udu6in+oPKf4Zn+ElbHY3V+cc76JILBdVqpMZqtx0VT2JvmWZLAz3e78avyNNr3Xow0ywIGy
OdX3dLU09soUoUFPZH3IK98LoelBpKnR1+HxTI22lPYimCTRIAx2buuEryXwBu5wfWWSCn3EPtF5
HiIi9rQ4DoAlkBvN4LqTfIdUNmzaJr1QCruccg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 90000)
`protect data_block
lvJgp9F4NgHfQyd0s9WfMj2NKmMmK+cVw75XRIANBEFXjAglUPymuokPQnOMfyJFPf8qKWlwo3Qe
XrJHuaeX6LKfO/NZ4vjdMRky3qPb7KS1ZDXX1CP1z1s51WQ9aTQO6BiBoNW6ouNJWTZmvWcHc2Ln
YVf6M5x28gNptT5WNP+UIgu92VricFgiOBR1gPIL7FV+IOzcJznZbjyvYSvlGJdvulnhubW2D3JW
KH6ybsV2LnM8zlsz7L/FyejM4DfPUIqfzrVM08P0bR3I/cxLPH/mVg3BsSIMreRHxSyPg5oJgT7D
cAJ41+YIDsrJkB5vf/CYBXpOcT06iQorhXtVQLq4DPxY3lzIXuYlbAqYKxPLcRzPrr0e2IB0CoQJ
MDZdgW2WWv7T5W+8mJ8+hwnyhFhP9sv9oMmGA/gM9vaCyFFxsyh0ybR63XJXfPaR35uhG3lSunFE
oaxRIYv6LaEaduqlH3ZgH2OHX9IkqqTK3tweKgRuAfXLoGkE/6+tYPmB5LuBmSif1yu6bzDGIATx
rauJ16iPQRnnBIMEReZK8gv/30XfdrH9NmTDag9LOnv9SCeZv8slp6k1WjfEgPI4gQU6AiCI2TxT
AcwN8eSlKJ6i98Rw2jb8N16ORwBUpupPRejyRA21l6dL14kBHeZODL0LuAcIalmoMdd2bw2YRzMP
R+kO91ZduRRzsBM0mnr11LFV/OezvYwU3prAH0gWn95fyGniKpD68fYmccEtwa751Tce455rDm+l
kexsscg5DWc4PRhHqYCHk4j61IISlAqaYbn+WU5gaGNFp7O8UcY+n4AUAQbemP8fT7swYLfGxjQ3
z1+SUbUzhrq2vGFr9yRKAIbW2YblXIshzH5T5ezD8kQu8/qP5FKtwRQ9PkYTv1DKVC4amA8/9NB2
gq8180MPsmlVTYaIvCso+6Ohy39QEZhX5f3WXf9pqnMDxipiq0DVnoWHET1wDzF0Rucv9T2wnf8U
2/ubcR/Cv8DE6gw38amZ4XlnaUux5M3T2ljijEPBWN1TFf1ofwQkRafL797wlcpsKVB/6twM1021
Tvi9zxbYU0jnqqeIjZnYCZB2+MpPO+CSkSSW7IzbF0Mx7mXmO8ytmUe36dFEMa3c1ehkk/V0a0OA
BCp7bxRJoRiyzLi4z4cSvXPPjxp5aYGl/RG4Tf8XDj8R7BiwBl6TYf3uOHUrKUns2QTV+Tx2aRtn
okV0HBSuheoJNBt4aKG7PUfmJ799ESS/o48TBZ7rcxWGj1Ln2oII3pBl0AQ5+zD4lzbM0kktTg/f
c6Fhus0fkV0cdE2B+6awb8jenB2oo9At0esjmrCvn9ixhYQOItm2Mb9/t7MsDqThbhUx/E+9yXoz
Iy3BuZyzVCITVuN+4k3d8BzMqIbvAp72Hqbbxcq/Oe86UYGbaALGa9UH2pMawdeidGIeeK6csm3y
+KAMEhxzwHP2PBNr4aXiTId8+tIljBF/B2AOfDtV80SHz7lpSuj4kdbcSyfDdwZPsvXKoWnlRxLi
AkOJfGgUVLnV/bRY2BnJ4uQ0ssX/gd33ANwScw4x+hHdeQjh+OuxYpfzwvLPUpeY1jqCROIGODl+
IaS1GWG73dhWFKgF41chiVZAHh1e8jJx/u8SNs7DjMot/I+CBJPylr620/R61C0c9BNMJv8DEYOo
XM3gTNlCf/KXySjYIwqu5eax9GuRKHU4knBwJnqEgW+EA8gZQNRuryAyu8t7aze6YGgXv4fYn86U
+/PFVHMO9HEjHWeAKBwwXiezGABUXEaHuwoTbzuIW9n7u7sfobAgnjX8GFqz/aKaoV3MEVI7Zv8+
kLREvGPymwmhxP3VTUcjjbnFhnrZG/pBECqS5eFgWKMR7nEYRNZBnzOqZSyxk9ovt9MVi5w2DTGL
XyBTLyDfkljIPB20BerlXHMI6uuB71eWALT+IHAP/uPBZMvQFH1mktW5JQqQrqwNT+flWPDgedNN
Mhn/bIyEVZww7yGFdOj1+qBEUC/Hx4vE82P1fjzQb2q18Vqg5+fhn5HVQjoR5na5YSc3NG3rmK8e
ZYvGkBiuWXH9HlCUNtSSpru8h4idk7ZGLb73Ff1QzQ9WOqULWs1b326ghEp2pfrNAZbJmhzj5yxS
YCWLlQZDYqkGQ9DXZfQnU8sDWp5eIQLieRWHpKVASY0ckHpv2lbWp+X8UvoURRhec8UFL+lXpvfy
NV0Ht5J0ge93Y1Aq+h9+zMLaUIlwaGCex3HSyKfUpNOc7sgsBYY5bAGp5cp9hWQtz1IFdSIYPOFy
UCyN3tsgQ4LnjgKsVMJasDyCwk7NTlpVRAId8nAdlDEJ5deRVpwm2BKbyURzbAzPtt32gZ8fhaNi
7RHtR1scsrYFDFdg5m0UaJaowk9y8khkPN8tHbbF9ClnVXe3r7Xa7VoJ8qqrfGLfbAWaG8Lp++fR
wucf8SrgnSdZmbsCsCoVtN+Bf1z7I/I1NH25bIKlWfkulO0FkAgr24q0RMIgh/L95wrqKkYQ9mEk
9T3mnz59LUEoNBgxFai/PM7IK16By1hAUw1ufscArQjNEk5ndbzHqCQz2jzLOOsIGuIpqtDsJ8P9
S+eByrwbFio4v3GOvNtoG2T2aJpDUR5frWV9Wz48i32Y+dHb3Jl3DIfrGPFnPzKwi3vch7A+U9Dy
Jx8RxBl3kAz53wsTI6ZwLRZ7nPPIMObnvo47rCCnnEkMLuy3CXUiZe26c+C/hgYNBG4waSnk2SiF
3lQ3+imjn4bO1njhwI5o6v4wJrsKwTkyCZyjY3AjzjJqxD1BvYbuO4Cak85fXwsdhDSUypcId37D
kJYMgvtCMsMC801Uo2kET6q/zFFUjxHdR7XESXnNIp+KvfRA1kBF6CUXjDExyBTO+J5VLf8t/gWh
tihxBHNNDD4Cel/IqM707uhZguir5/6/HeGNcOULBKU64JaUO8C74AMbsfHiNat/DVS9CAhXqYUl
mxrphLZF480SScZ6o8qWXgAXl5k8Ogv2gDQxnn7/phON01yzwh9eedJSk9RWG+bxdNcO/01whxaL
1Hvp7+tzu+NHHjW1l3haurDqDVMmp/LLLPUE19eJUER8YdY4DqIJGgQvQjxPmqg/+tbbFbeFjTaD
Wk9AvRzP+J5a1AoDGhRLpcBHpwfj+51UJUiTM67VwRC/BSYqF5nJGtDGAXRJ8v+bfcXhNbifszi3
yvdW4B8eNFe4H/lfgO8h+qXSEAOob4zre4UBdodfqaUzq1S+qtqZdGmnHio9rN/z/RUMl2YDT+ul
nEIILSBI1xSVExKpHRkmLwGdyfNQtxwJJkRvnaoDa6yYejpEtRHJ4bfqL8caAbl7IEJgEtwUBTh8
MVjay/FT5USvbIGfU/KQX4ptft54iaF+5hIJ+eJE2ZT72SWFgy/tqGzKFT0sfSqcAl4uKiH/DSe7
9YoR7Wgga347T4L/swBR+5iguE8Cd257P90h4H7pG9S8wkuQJGzAPucvMaRLuKr7Jm7Cyms7rnxp
kxh6G1pA88HHmIcmt4/MWaSkKyMYr0aMS99lg7JcQ7RbqE7LtKh0pKVthiUTzciWiXExcbnNPv5M
7QfSUtQtJSJiTrIu3P4mmnhxgPgcrl9BQZp3iETjJOk7eDfJCInOhMEwETT2P8pvT8RPUUSyRbzP
WPssQ0OI1zqmP9jsOpHzyST9bN4xlF8OxmaLFFEddHelzKwXHLRgPqvH1+GDkTYzTZPIZYdELWW1
0d+CEtgda1eVep2JKkZpHjqmD2z5AZpQwKVkZ00T/1p73FoqvfHtbxBgIO7XKMAQWONuRktcTW5I
7lS4rkerJze9mrOnsIqX0mT9dRuY2ZBhALupbTvIg+4FfAXk303/KvnexK5GPJTVFo7ZuIC66LfX
i1CxAOmvs9sj7iJaJy4B2MuztvDHL+Rdm+ga44q0QVqkBheTT+wLAcavq4uS4aqk8dcAayabtYkZ
wRQf5uizuL2K90zpudVZMj9puR2DSOqW78ttFegLgOvQGhfHA/e2Vw/t/qlQrhRLGd6KuvIo6tVt
q6BYNMI+xNyfV3l3n2EC1qMpzlnTUcutOyPkywXhUE1vsYoegO3OR77Icz5CP03FIb9bbKfjouoE
bTCstTfet5CjURS5Jf4pBHH6bOvPKKjdeUyAJurr5ZHn0K+WgpQ0oPN+sMINyvTt2W45TxOcEWXh
krsYMNYe+epYAAbOMWhRCKGVFfudZpOOD2WcqNvDsVOmDBzLtgaM30ljpOTA5a7+3qsvdzxe3pVC
XvH+O5Hfr4le+Zy/+eu2PYwTysrmTKrnq7OcVNGMQPvPmuQdcY6+X8YVshGjkXnNtK5qzwMFeTZc
1j2JdpDoKsONbLJtiGaONZFLQunFo4aWXX1YO28V1TxyFgxGGgnGYzNuISiFE7av92Bmt+X8ex5s
r4gTpwBQnVXlp7tK/0Hmqu3wJR7cjsbEVFOqKe8IwYqzL57/KsKb1f6hLaJ+aT+KRgauATiSKbF3
G5Zpbj+LwukERrhoXKrGeMFjFlaTfD5NV7RDQhW3brZu+4drh0hQe8jUhxPysVPH2G2hSrnpTr8i
cwLKVay7ZX+IXFR38K+HHOTYAH4hMOrBLxu2Cpb3Yz+DIDxTDEkSyEiOkBt7X0aYSuxj3JD/J82K
bjktME5B+v7eSmOucz+9Vtsec/uPCgj+BcUPQ2IqkIryNpZ5wRPUuRjiVGDu4zHncX8D4J4L/oEc
LY94rzemfNaV/XMie8Nki/rls77rtdOXSgEsQrs+n5k6O6iEfLEc+SJl2OcvlRIbPjGGLmSv8Qbx
Qu/9llVSFow0S0Q8cqOtNrUrRhROPd9tfGIbKlqdpdG9Zb00oPXXHtC5KeCjokIUYjC0VrdEj0nK
pSRTdoi9EZ9JFVEcdnYvAo2AOZkSoXytlMFq89T5Qv5qLfybNZ8NDNGf6zb2YLAjuQ6QY7PKOCgQ
egzmwLkYZlU4KcODH6HT63tpLfz97OPXiRnX9lwAFso1VSUyUCpGy4xxjs+kVIivqg/Ho9SbHnx2
jRPYOPopVcXQr9QUxnHYiEVeZt4h74VpLGTEFICsOOsLIK9eujhu6kdZyClRpsJHcmv6Gg0ZnmGr
CLFBboFURI38IZAbpsc5p9T2fo+TXwcwGAqc8A0SkmPDoAziBBmEmmUg96em1zE9eGNzy/cJyb4S
6S80zn+i43Zr5qiE/ueCHjrusoJfCKGON0JBfQSCTAK75f+OXeauiTKyQX/PxvLnUU/Li5j3PqGN
z0zsRW+k3kaw5PCK/QUDXYOTcFGAH7/s+XsGubgaRos7bOP6RyQemjtlKjWhfvWOz3xjvfAdby6V
5/fFxAOMFwjNfUkDHt/wLwVeHs/M0LdiTtIutNLphfIWq/d/lC08FcM1afEgnTuhnjIRQoULorIl
tQUhekskQUVM3bHah8prXmR/N4qrhjlQJYcs7yPx3U15pG9U8IM3NDQiwKYjrNjxWiMIH5A2fmuT
RGkU5/92rRXzBcC3COQQv5sqjV5QMv4HG0JWei++MuW1hCykWABG3oaJgUkAx7LT8EURA+ycsKh7
4vD4JGo1vLBJx2w1XBX9Ddkg6cYPlAHFAaUfGmP4fppXo674p0VjN/C0Uqn+HiWvcKjNmE6s7mvB
MpB8clwkmImH+TpU9doOUKQxkvqjjZ+bE0kbhiYzXj+5N/bH6K1VPQFFvFgb6Izl3AbuM8OJgPAs
wNbdBXDHOXo9V3GMu7GxxBA4jn/Y43/6HRPLPOrrgao/2VFs2i6V1KWzfFSsLXbGEF444GshAxuv
8Lbqd7rM09SyMcrYIfli2SBsbETLRUTeg7MdLMfV4SKPipLSZX4paPphh46oiJJtTFfShrM8h8eB
0cqvd1pwpKOwPPqX/nxBAPtZzTnztEhI4oX93whVR9+S7Se4ebLFOYhjVBFANHEr34UaYU7aFj4m
/vrCLCp/E0CdMjwQ+kF1EDR5sMVQ4jEQgFzRn2DNFeE56OtoY3TobtA1LExfbvzBYBZwSiiMaZYe
mIk6G8PDBLBL/YbXW/5IMPA7xK/hN2zjqDJSPoS9qYQrud+8BzlxFmV2O+fKLJY/PKwxX/MoJ5e4
35qAR+1jODCBlpuzT2Be+mJWJFt2/u60t/yYehLUZy2GNC/BpQ8TAslP1wqgrD0AZ/VftWRWB9wW
h9yBQAzPdldRv+EgSTCXZxDXKKmbTHNseJRctPEN0GMWW3jL4FGXyR+MRBKq5kB8CYFPghT/FK4i
Vaxv6FSv1roGWhXbh8vGvqr/K0b2/3TtLdIyTx+a1L7JFTC5l4fGVp8nBd/uFy93WIXQGwmhB7Gp
zpEDN/hRi/9Loc6VDJc+HzncKQmgARUf3f9vvYjjzQY3u8KU7NYgWJ7cjCKM4DbVhmNvmEscfDOj
TfEZu5HhB9q62Q1+qAOcIRwUr3PrniVoXa1klAxS6StyGvNzEDFkIfZNgYJSCLw+QKC4V4jrw7Df
JG9DkAzqqYpyBWIoOugs7Bp9qgPY1XlV3ioRKMh/hYHO37W9ZiC4oxkGkAC8CqfCLr3dr1M1H2Ac
yYyOFCJHCkhsrizfak3lGyuCrX333tcftcCQKacOqn8msrQka1bN/iCbAB4seqMaQBnuB3206/rW
RCQKJMxoK3dqD4niSi7DirPcmkgHVkxoGpwD4a0leUc7VrDVSQ0Lmg+34XW5iCN+prjX75GpgVef
l0lPkD/D83mbtJcqFWpzcqiIPzWSFBPtvDFNsFhMQ2gV35HrwR0DKR5Dw32jN/UA3aJfbeAL20Yz
ijsLY8wRMUqHBZrKDZyEJkYoO6519tyzQu7aR9lvkWjs2vjusxsUBRmjMmGSZLYddGuvy2Im1mOS
PwNbAadcSqpKSHpb3gFSw+hXtr8KX6kikUv3GggEe9vj1B+rXH9CGpZwFP6TOs042GoTvOddGCNl
TGHM2ExiqnGsAaCAm4VF3KukzqbpFCaW1lCaV/s6UjO/Mfhk7SdmouttxUZArxC47lxewGB/+eDt
eWWJnWNAM9RTdtCe6+2LgA22pcTpi2uZF5LAgW40SeoCJZYBTqE5BpKde4Rrg8BKE5RIu0A6W+j3
YZoXh/8kJ3Ugu/RfovALpbR3HGBvwL3bwZREJKmyYGaTTl1XscwUGyz/tMGn8FCBJsLdAyVA2+lB
UxWJdUlSlt7lcLluSuyjLexiQsIxhCZ2vjYW1pEWVZomQggeOYu3W7tmdOXWXbpL3b3QOOsiv6Kr
aVfI0g1MkkWF31fr3lklvg4Q02fK/+BWmoaRUysR0YnM7jsUmKOyfFFKhd3eCQ+ohqA4EqMVKRpE
t+AIq9mCVv7tASWlEOExgBOkiR3UW9XMBq7M5MX7ddOH43niuKM+/zUxjvnRRpIDol5prLMZ9fBr
UqnAAZmczr7CR6XfyPdeQn5vRgXFPkMeY27H0mLB2xBHpRnG4W3Dcu/CfGbbVEMgG9kTNYp38HCO
4t0V8IILAS8yJ5scVmeAsj9I1laZ+nXv6sKmhmHnhqhVrp1bszFbPLv8BYSUalHeWhCClTnSer93
zNYOd8JA9wOiNxIXidgzs2uuwYKPQTqS08pbnVBiyZYrkBUsHebT9pW6+me3hebo80grm1INYaK9
tWzdaA59YbhbRcoYja/K+KCT+YaMlZvrK0JVHdVQxnsR9X8QkWh/CTeGuPRiM0D2divRb3LxDfpV
m5hf2Tji3hwH6plPKphfEn0WT57tBCES9uTEyJN1ET94gaCm6YY/w24aGxgffb9awF9+FFrRGLMe
d99JbQ19WCI6nJwBMFJlxD/1VKRXF4TDI77LCTcNb8i6+L8LPVEb1uOnu1I18cGDX0lzvrD2kdF+
HLOjeCQphucECQRzTFt+BzscLKFzZE6B1JtGx6EVT8jaoXyz9hLsnfFsAmUnssw+CwdGxe6jUTMI
NDcK8P+G+aSweCHlyN64K9oDlkdiIVzM9xLK+Ahfb45WGNkaTPdyskoKWThkAjc2ncupXz4y6/XS
s/U/LKA3226yDpTsPjL/3oZ5hu4NWMDVHNxKiu8sercAxdYQd86UM3+it0/q7hEmN6CB5/Qwnc9W
xIQfnaryCKvhFLu3Hf3+XvBTmtvImRxqfHj3brlsFacMUXPeUNZu2TCHxLWUp+nmLRm7t57pko8g
HWLKbIesFqMp9HEsvGsl/Eo18R3+QQ3ROO5Dzp+/aRXmk+jJka8n9CVCWSVJfToZotS9Uyln3ZbW
OAhEVpTVbXzUbo6rOgIMgohCBYOD9d3rzBHjHnI3tEzgnZzZnMh6Q2ZdEJMNr+lduN2SLwAENdBz
n2dPsFMPfv+qC3kab/MGtYuah4utJAQfiINioDtuS8aek6akpE2BkpUOqjwhq5GTEL9TvLoun2zq
Usw26kPN999H/3LvlKr3CPkN+Ztvs34IkREEONJEUqJCsnukHAMCmJXOCv+JkPhVHhIIXtMAieaN
kys9LMf/5LdVLtRMBNXrnjOmHA4iT5bm5l4ylcNj+eOAHPLmq1xO2oCBAa041KsPR0A/X/4f1ogS
fYPvxzDEHkeTmMzu6679hmRF0e8AFzs7kkmF1ooBVC1gCG9m+5+5OsRXTRKgEGrpfdYfrMGMhlWo
JleGrs2+1VQFNinj5BJA8zc1FJVh2uePXh8+2xiqRJQkxu8eXkt1xOc49t0nP2Hyiw+Ez4F4umsy
L8yYEWEsayXgMCvpufM0dtaKMgKgDLs9Njnmeh5KfaZSVsjcpTRYaCBMpKDTQJZ1N+vERWhs4dom
dkLsrSacPwfvchMRDK3YzCURHvf40VngRgKjRi6UgVJoWFP385PrjBEtLarbCIHkch3sW/W1e5KD
jp3FVXzcghgBYWPZYHSbcY1/SImnhw/bEmwFXTcAlmg9TbcWbLmxjKZDDQ1Mjih7pH1Sg8cOrY98
amGAw1yeRtQt4H+twmdbXuMwhfGCMtTK6Hylb4C1nB4V6MokBYhT9KAmAYdB0RihX7jY54g01v91
S47xpDPygGBt8lC8qODz8h3qMDjJHq6bqkqtQSIJ6HtBuF2aHRJcWD/AEGdtwc34Y1eQ4VuF2ir1
/4AYJZ1AI2ojRVel0AvgMyw7fN3ZXVoyGZ0Kzz2w0qINhPvpG1ibI4ulElnSngzK4S2irsiOGzK4
DscbatywJUfgsP7gj89FkOIEKp+stC742uXDJczZs6njfSCxLsq98evZIjfJadi1lfxf6PcmRz45
07MsvxnpkXNQztliaoaurcsyjhUeLeKmpCEyMCnOyh9mVwJ0Ym6XKOK6jQp7Gwv43GyAIqx+T3f3
x1vyFYtx0Ra29uWaltpeLLkigv4ol5ikuxIdzvcchM6eufLFy3IgdN9FOrCkUvC68rzFc597FzXb
ODUwroV5cAEQyuxtdmjqo1GJwqTJ9R0f6yjP/mUAI52GAcnOHFu9TiOyKtKuhNjByuEIwHKnlE2B
E/quFr5SSaxPURWtmHEW/3ePkow0cTGiRcpUBvGAqIlVRVdwqWn3HWGjDcL+1U7tb7Ly91WobxNN
8lcQfLBy3Sy2uMPzZ1X9s/bbVFA/ZAFlX9KjUSmxOgUHL5MPNnQ+jMFUecCUDtbcpiGHSuOcyxjq
GqKpSyoac7jFV5gx0G7y4YTyGfhxIbZUht/0ooDAxHX0dUP8ba2XrI7YdE7b9u+HPNjP3hV3kY3m
cYGkJCMEnqCwv+bzNKd1R1P3T3RTu41fYimwAtuGU/PR2TOkLJpgvXNOaohdDe4nuiprMk85s+8x
cnx20fiCdlJz7qp2mLHH2BbvslY+Z+GBtHoZrJI/3lI2kdIsGEnPFd6cziV1EoyIFy5R3Cj65yxu
Vb39GulT612eJKlb8Egx2Jcs9GaE46B3CujxeQNna3I10fSSzzF83jY8lVcYsXmfUnwMkwrA72al
ZAL8feURABA3E8SnLBmTV6JPhI1lxpwlRzAXJtAMkeDgalkSpQb/utfxJCSTFfP6ZL+J4ZE4Y+SA
eIdqlCpoN872rrWj1xpGA0TjR2FiteLRzoJ6iAoqJZU/9CVCqWOUrkXq1Y6oJkOSd/GjXLlb1Vee
cKjhOxPNIE1Rv/Tsu0t7VWUOtWFEz3tLWhk71Uw0MnYS2coYADNkFFo6oBFZN02YczAMeP37NkgK
EBujWtc25djZ2+6UheOX/dtl4y4/T8bIOYD1WQXTQ4SPBNKrYu00qizF6rkHlKK6TiiVGCUx+JpI
tvhHxMqUzr5dp42iP4Nu/plUTJmSqjjzCwrvNU2vkfkA3qSZvHjzh4eC9Ye7ZMdvZBx4Klqybut0
14gukAFh5vdtg2uN9gP0dmiu9oh4PVB5BVI1EyW3JQ2mZrn4y49e3No2R7CDlggeM+UbSQalFpqA
ZkcBDocyJvUi54qCUrXt3FrCW1sohJtxujAereE51MjGa2u/aXG5gEuKsZ0ZmqTl3y3yV6kGDNDJ
7yaz9mDiOrKG3er7hcMnGPFV4RPEljVZRJHZmpWvGan8Chx8l7vlFL26l8g91pA4d14B7Ts81fXT
fgUS+PkebqqR+IxmDNXWdqniSFNJC/WK4McpBMJeshohk7EB1YfmfSMmnhzqPvz3L8RDgRJzKC7U
Uatntfx5xXf83ba/dzZFZOVnvRzEVN42J9oCDVYR1xpUrGoR/PUJgz01Q5H4Cel9AEmT06VzTt4H
jNbU+yQ0YZo70n3bNk9WNC7u9FarbFKUV3/EuOHB/1JxeCM8x1FXp/AZK2yHvs8hlQZPuR346Ujd
dFX2y1FsH7FkIo1ursbnMeCgGWADXj0heaa1P++0OGSG0QypzR4+sByA23c3attfDeEKdzYWajPl
WW/vc5KJei4GTiMFd5wY72ALGBJV9bX8GDQ8BEV2cTyW+vEt817D80Ehbr+GDfWOHpqgBvZGRgj/
Eo7Dn/+gy65Yd0frADJStWi8ZRWTYFMtot6xzwV+QiYcj9e1/X1LeQ1vHBDQTTgbn1CSDIhV2SHi
1k0MXJZWaThdO1tLLJNPQcKgRaSWgHaWo6G8Z5GhtgsJu9NIlGTffzTEL6j9UG5qK6umMcH1m7ir
mG409fT/fiHlHDtf45gz1LjXu20SZZ7Jw69xIphzjo5L8bhi9X9HZkmZ4JoQELWayT4oJmgT0zdN
HHDDSLJR9o5AF1EdE1RbPKj+FDUOoSa3hs+ljTtqQHdjPD2M+AlzyCmIGy9shKQ+SMCy4ASjIxBN
BGvmnP3iWjy2kttgl52IgQs/9149HS8dzPgtyb4r+zXpGzVLOLYJTWzRrmt2F0loshZc/rTSLVpz
LWcp+60mAwjDF6rqB64j4Kpf0VQOfSVsvxK23dRFsC2SaBJ8bbr5l0uUhLadw7GAM6Rz1LXgmJtD
EVEiYeq2aqgN944SdaZ6kpG2VL8/REnGg7F8biP5BxhfCH47nmsnqPmMIPyrHmtpHNTrJ79J7op+
HFIqo50Igpjj8Oens6b8DSkmv+5zrAdMvbogA/eFXEyloQuMjh7B7pvH+boC6puEtGWtipfPAoeK
f4pMK53rmWbln15vxBJJFpH8UbOyTGMpD9DpCGjjKNJm6G4ix7kDfTCCcS2yp/1fi9X7QrmudEFb
R2sRAcyrLtGUrnP6nOlBtVGvut8biyZ+8AMZlEQI+TaEh2ZpyJ72Q+LrPuGG3c9SQzIaZT0ZIXSr
EHX10/0UpoiQixDoudtUyVxhj5AHYBRuO12vHq6OE0R83KrzkvyZ5TV97CEyhKXljh2fTZ9Bs9ZY
7I8kZu60r85fhzZcKoNZHOcPPw30uv2EurU6ilxEd1FY6cEA3qtQJgjFd9X34vgsXMvXVF6iXNb4
Qywm4NdcSalsWZ0owrIQh+0/gVu5/AhTEM0rk+/rmXop+N+5ZNRFda+XGODFlUx7j3tXl5RKS00M
yA3nio128kvLV3rhoVdSKcNs8+DjSuNvttTIwSbDlMkFBLLtgoNJzDWczw/yeD3pAnWR4bDOPhHT
BZDdR5BGmavuQm8FYR70OzX0LsTiNbPgVlOSH7ijvKAnRd2O5RRWYDnUw5H97EV+JIqQ70iZA55m
H/+k1dg939k7sN8t4ammWXFyo4cX+8DjjaCMC8BkUWttL5ExeDjpSzXAYMfIr32mfMtcrLB2UfJX
WFM+3CPKRZxHqfVGV0X+Jmfyydc/T/9GCJuDV56QzDI5hmGlDclLbnjrkeIuoIQGVq0WhNUgerfq
d5xFxNA2dJjhLkbA3SEFKo7R3ROg5QuZegpskTiAVYs6RA54unkQhrbJFZ+grsA0DI0eqpF18jL+
DOXQMnwUx8lHMl68T+fePgTMM9+voJjCXKv2BSRHu9lgiDSGa9AnwX7alVrxU62SB9ekpTQGrp1e
niK1IaE16fNp7Z1J90PhF/WUR6+ZcSNB8i0gLce+oCBvt1rvaK26a2ZpESJaoO0QZ60kzoLNRvzz
1bNN6kUOFDMnJX8XT0IaEOolXyivopvOE8TdiTMOSI7b6Y64+5dd8Cnl5ecYMgjReBIIWRqvfxjm
jGP7iwGYibm4iZ7YsPiKCvhBpusYbVwBrd9VW/mDUyUCwpPUTkM77ImYqRBEflKq1gYKBcgNpWvt
UutSP/WyJz9tWIyYkMdvk+8uP91JCg0S8B2DKzPi2KnBtiVOVhMH1ovcl/qQHm0OiL+9jw1K51qc
ikcxrRRQSlnAhQPckOZ1YsVPTXT5axylr3PcqDFjzydk1x3et5bNcveVT/eqhf1nVvnLKbjBfW82
LC9xBt/h1w0wkfrcERBUWUGR3CVR7FGZOZeB12jiRsbzsXsSmNcfdxGd3G4DrYiUYLm3y43Ycx1g
k9i0l0NwwCR1a+te/xVGqh9soBeK4w6/kDPQf31TqUT9LvJOAnVDOBQ/ESuS09qshelzC8oDSUXm
BnthkFpNcmEvAssr0H0kudLy1MgkvlhcloHacrPBXi7hXARlsodpP8LfphN0Kl7eUP00WYLcAyf7
RnNJv2h0EeFtnuUcafxsPyCGwbBzZmDd9CCtzIkRUckr6+i0vlIzNLO2sjxGDOhlQSCCQL0nsTA0
95UxC1M9Vhos8B/4/PJyIQNQDTDvTgOn7vigaSB7LLkjVMNiTFr1rGM6504hdHlMk0FrO5yNtkB4
fuKLQ1aeXnw0lEiCsRHkxKcxCJDFKSOQZtVbGrt3DRWqOr0AIgCpfDKn3PlJcR7UDmgCY8V4t3JM
9aajrLm9opy9qXM7pwXCDxAZnDxHX9NPhpojyU8iRbxUxXSjr5KEwadAUssNiwEt3/Acf7XH0eq3
qUgNVjwu6llQbLarHuUlVXRZrPZAQbL5jmJFPhDAUcvtonSf6frvm1Adeq/v9u3Jql78Qld16tX4
/vgfmPS/1qkdcKbCpWbc5PzrcdjN/L1aLKIynB7CsRvtIvUFbzRQ+wxMxTzjljwxrew5vBzkvXvF
v0Bt/jxrsAuz9XEj0KciDaDr70M4S9b2sC5f7HVd/82bQ1HGX15n3dMPdMk2z97Ryjd3EC0ZkI8X
6mqlV3PV1MGt/k17LW/l+sn4pWe1C8+Dj2um57XNjElp4fjCumHKTqDKE+uPsGWR38OiyjqTdLge
SzS1/JRQIlWq7S4dSdCDVMT7hTdwLQRSvim3z/y9Qt9Trn3Sh4DG3ZmgyPkZUoQkH4OJbySiTzBW
Su9aJveU184sVYPAhmmYofmbNWt2dvmRq/y7tbbtyEDbdVVzeagAfUZMUWszxXrMKED6lY+OFSyc
bxTvdOXYrO+EmhApTYd4CNy3UxPpbVcvqtZgnXJOccfjwVUi8H4MMDVUlv2x1SW8pFGohwusZENi
Ke4ALQg0m27AhXCLVlh79Ge8VBsMQLAK3u/2a1jOybW6cXMQ/6bv76pCOsFOTfZKB1RMTzhzfv0a
vgdxiLRK4MWIBjYqIFoX68ESxavhR8OZ0ETHoIDpPeOQmx9ww5I3or+KRQBVlRs2MSEyNHIEVX8z
mqJfcbn6q6Vc1AqYyaBmmLYuOnxaC4fcBuOwLlZ/1iDq7wl7+OtNh49qPani4c7juV11Ojqd4IbG
bfY47S8WmYlgtS4xwzXZ1oseIDHiFUahxGxoMDV3+0NMlM8O7WRy3w+wCwtkG+8O0lusXuOOnNII
d2cHx7PJeBcRKd8XBi6xNGBvnos4sEQ91zZDVH78vFlFHBmXP54zMgA6yPFvd/K5bywma0BQt3Rx
QkKMseQvUHnuI+FNcViAepoLtnDtnhOpcPAaM8X2y9OYZo/1M+FR4C7ohLpdQoHFJHkKKRFTmMeP
Tzkw30NHbdpLTz+8XHwB3xOnB2mkPO1aVT86anNGt6csJ+EDaAZZ+dGtVvZeQ2ChTi1qm6izjibb
9m42q0Bn4pAPP6HiBjzVeTkUIjhZpmMhWyBPTzn/XeUr+A7DnVOCJzZY9UhRsuk+i/JKvhFL5FyV
Bckrr5cXIPM8i6l+720T0v+ByogmSCkjkJIbVzICx7MCpwt/VsMypOqw+qv4TRUGjRH3D14BYI4f
b+XQx+F358cA+a57r28Re9USKSAh8YweBV9zpY6a1RuXAWP6M3+YpjNKoXVMWvu7K7mSqzJ4cV02
J7GqFrX3637GsVv5lfNQ5OUv7TPQJtGVgWP69Qiq4RBoTZh/jUfZIIIFwNFXMIqrMPFtLTpYfymE
/2Ok5qpw/NorvgS4bGm21sF1hqQ4wU1Nnw2qjeepgbGssRz9IQb92a53vyjvuRmV/jPvHSA4549+
gezYVVAbncKDOHsR2HoZBZepd9bUhZhIsNDFT/AFJH/GMc3ZlduG4KDXW4JEOk5wYvVB3Lku8WIS
Qh7UsGqLKvmTDhDynDQHjANRSXPL43E/NiBtRsPjkG4GvVorsqQq+Wg6UZjWr6EPkPTDiJ5LhyLY
2V1y5aj4WepUbYV3dKRm5lh//wCQNsh3mXSp3nX0unfmWnnoZxmVS2dCLwf90awds1DbeP45JXJc
/wF9mFe768H4kNkH1iVY/U6q8Z5y5F+r/C5xPp5+l5clhqI4b9ukfg+CKkuOdyBWNG00j8A5fl6K
eyX8VY0e+8dZhCA97p/7BCqxHh43VRu4emn32ifFhkt99gDO4EY2CGc/xMP+IHQEoYB7acCiaiP3
JhHxqDNX3RBqYporY/+FHn1yj7mp+tTf/ROdRAADsnTZUhd4ducQhUnoRQtDM6C5SVN/NxEEa82c
iAlgDZy3HhiqbsBTVaWxVFUVn3R0mdlkMYc+jQEJxI2QQUYKKPawYDEmUvrcpYNC7RMUjUVF0g6n
HNQmoOO+WVftnZfy8pHPYHLQAerQMOFMRJB9p2+BGWtmPyBgrRVotIAKfTgzty4VFtfR3DoVP9gs
3ACIlLwIA1ae3ntQpEKYjeMpR7uMMwsaT5mMEwQ4IXj9Bj79/8va/l8HjiuoWZoot52gEWY2sQWy
ZJEyaR1s1T1mb0zZqKh5PaXu39J5h3+ZZBXYpezjEMJoV07sFmOJgK2SSVVKcmrJal8jw60Bcpoj
SaOmHWHo3E7gptzP4zyAdebLx3p0SXlgfnw7gvwUjuMO3SxUHKRvynXcMp9aTfJYKVqZByf6ioX/
n89m6uWIDpiecTME5rZomNHIGeoChTPxnwUYQsgKuzU2rohucmnQMdurjTxtdC/I3iKNsKMVamWG
j7buNCvi7LlmxsWo+p/BkQADh1+AK2YpL9W0F8+6/EjS3rQSIi9ml2AkbacIx4HLR/VgRvSefm+0
DRrtcLNu6x1zz32Tyt73uj6XfyuV4zKQYo2SUhncAfqlGZCuj3wUMiySBNsK5BVIttY4FeigIg2y
jk04B+cmhg2GMwMePnxHhDsYGXmlroyFWvQs351Qa6QoErf5uMMc+JZ2fMGOWO/lukhw7oIE0sVB
TssXfkI7v3WohE0jft0WnxcsBtL/s7VhU0Oc6yE5772e1p2zEF93UHFI+zeoKfTMnIMw4haisPBI
tODuBC9cj6Aiaxv0bmp7T/Q39S9eoDnlqPGOHeKEJfCoy2yEpcZ6x0F+jjQYV5/vav9x6M51oXLB
Pzm5ppEUsWvVxasLTstqE0Zx7QNsz4vT+j3i+AQdyvEfiS5HOvHgGTmkJv4AsZL6jdrb8kooMFWT
1MOGEO6hAt3lCUHXo3SgreICtUtKdiAgfsuJ6ZisgenD2MC4gpJyTUWFauGIjFGVVoNjT/vPz6l+
ZovGiSMFZ4OMBSVjz7b2WWgR02ndKNPWCUEOWddZMr43o/yyv181qhBFb0K9q4vbi0XVJGNngAZ2
5kL4ais/DdBY4EY86SzeQvhVy70HiHgaUmRIbLEhjBmWrwxhBtrjmIcDYlKZMfngKMzQeymarmeI
8f6EgDbMiBR/1V86cmmXK3tambtMDcllp/ckJUr5lC9bRn9eDKnLpL1KPRZNGDFp/PtzTmvOWax5
lfj+sClOVv384EtFYtnSOEBwg2eGpFgZFOcYC47KqAFH8wsPgIPmX283NeooSHkwj8f+kSf9hXKF
jJcE4c0Zh8dAK2ixTf8cwmIyEpA66YcQgmcO5zbn8bxVsi0vn0r+wNS+DQ+nvEGLWWyeP38zyyHu
oTXZuYb01ViXtyMMAWV8uHKIApJHdPK5JdEROL9ogfnqv+IVcoywAOxPw79jIRX9rir806R7wocG
JHjyeG3OjDe3NagmWBWEAelmtXp+witAAlBTtYUa3kt58LbY2CdEwFTs9V/ZBXl+sr980WyI45Z4
4YIBlaJSVZaART1E6/J9CeUGOKPTMXfHaXvIOADORfJnmLFrKS35p6FrlfNWkPTE7NHu9S3sd696
Viw/f7y38qQp70vQmaYSfKFIqehSLLuJnZACcL9wtzB4BNj2vnEenum5sDtViE9mWTmN/B/c5utn
9EKbkwgnEhYANKBiG7LdvzHOLkcAdvCcEQy6WcZpma1R/T/0gkjHYjjUl0MdzVzOlNGYFH/16S+V
+l4cFPC4aznB5HmQAWHay5l5dISw5P6KqvGtvXdRwBuN/0f6f0AwwPBbIjWGF9jKh9nZau6ZrxBx
zmW3FEgl8sBAB2HrUWPGizxssba1ugHm3+UaH4rfO22s1gjAW11sPFhyluyIgF17BgHh+fSHmjtb
5JUyPa6N2nZhcAdHuYm3Mz2tDphOQPacuQj/TsLcCBwS1/jpblt+VJaXzPS0497rF7ErwYjJXe70
+Iqf0Z9I/tRg1Ep2/qq7C8nIjwN1lCm8mZI2cwHLbB+WdqILn19utqQHxgOLwj9HnYzf24fpWs+a
Ublja8W6z0u3UQ6PCtSexi5X40rSON1p2ukMJ3+6nptqjDmX7ip0SIv3a0vZHx49RFKdw6amlyQ1
WHKDRcPN+h6CJbDYrhRo344fTu4Btc++OzDZFrD8GzULtciQfAK7Phr2PpgILmsWU1JSr4tUsWJN
xZoz79J7zv+ommpZoIBfUi/GkRT9rJJ5Y6SslgGS8Zc8rAJUs0J38yNHwiOvHWeSXhf7jAqPz3Nw
+5XEKfFKXwgtRGWrgXBpzad2LoqJdhLDXKwqDQSXMF1uwcpkAEe0BRd0GI9XCoyoIBgxN/OoFZGv
IYuc2MHLs37CMJjDGsVEgy8HbaV3oT5IH+cZrbqHh9KLosurX2FuwGEjUyZD+5jWYDIrCi/uI8/O
SbTMYYWorfmrFnFAd5UUo5dobbvuZT5xRFW7TUnMcO8zKPlRdT0ZDGSut6nPBjpzRgz4prc/e1g7
Qk36acSHaTmnzF72huOAsqYcFLklD6Q5ebofz+1navGAsOpfSOyvDamx1uRWediZ132xs0sD4rnh
STzgdXpUZtL1tcNJ7vYwEGr385k2h8snG4RZOh3UrI8jAGxnLe0BrTVZFM6hXONaLGapeFST7aLk
lQ0jSJ0VjSW5zIe6HwVRw9wZ2o6ETaStq/gzKhxVFa6/DJFFwN/LmU3aleWqFb8y2kVzZkBaSTyX
4GmoesKOfPRbaMVZm42irJoeKnA/4p5G45Bxo88w2TswgEIGmaJ0J0YWujdzUrKzZd+1QPgjXeUr
KGdRMCl2AskNTiNEWNY81Zl8wZiL7Oyc9Q/B8PFI8m0wIxIXcFUzufQUo1ArWxgQTLvgGC2krtA+
8a6jBTH0jr7XDzQAejuDffhMMuLhCQNkrDN3TrseDpxcovyM7dtKLXtPqjMc1xlGNkSQ/SIRcNmD
hgAebhITxmfWfbdEk9JcxIR+BJx6RQHYUTTrNfVqv1FjquULS/+nTSvHwjf3MACVbAwfd+mV6dgF
sEDjOwwHlCepOsmeWsG7bcrZHtmPnOY9ddJkpz/ZlQKqNEPlZmrQg0gnpPk2LcB7GITKG4omtFPT
4FTuktjdfP4lCYLdkDcMAX1gdqyrqxbMLnKZRTN9RiWzIMsQiECKRp84wO4UyaFtDp66ItOi1fTq
TVypuDQhLMLTQo8iBAJcQJ6iYTFY4+IlVilKWPqlfUfRnU26SjbBohwuXMkzm7nC6MvCrddZ+Vhr
I8esKh6skT16vqUvh6L9DOmorHzIiZ3g8eoo151G8aA2X6B8vTu/cp2f54y7s+JDD8mnc+b5JT7G
gRQqwA1wHRrjiz8Re2bQLNsOyonMjvc5My8ZLImTrmun1l1i+wq21qJmJsYQstaLZDkBA97mfcm3
nLaeER29u74yzSy1MIlaCb6P00A+9ryFnS+MSuNwd1lHbyVGu70FjCeNbmJvUHfE+qFrauBriduy
uHPetJrSy5yyzSxE8yzF3B5NTsn5vvd1JozlcB2zD5tVcmzzZ0xu12jwJDMEKIp108HwuJmA3ZHg
IrZTpZOKVF6ON1JA1tLUWu2H+NqYiAKJfOzIvCFCZ8+CY0tVTAJrAtc9WQAg0uLt+C5RxgTTJZ8Y
KMwbmhKprOn71xsRvVS9lpB9e+6CZne/J6wfQqNquLKqS4R3NA4c66xT0yQD9Hf8qQVO2mepnmhC
UdYpfB+yB7VYikC61kAs7SlhWY27KQSqJEZPtbXrVIXzXAuJl69hnPsJ6bOhbKaF09ETurLhHbQN
hf0QsG8rrOOkrTBQZa+2HVSOJ2pfLYYrtjaob++xuM3rFtqK0QUZ8D5/8/2WhueDSbVtmV4c2ZZP
PrWNwoaKy8NiVectIHikGMEzeOY6J8gqO/lsIHqpsSRy1b8OkWaJhrWlDAtd6DiatPbqs0KTfwjw
ylGjuLQlM6f71AdV8wtFHcJr6Oh4zKBiCkPT+y9fJJfDWOxmEcel9pKkpTE+zRprkeSpuzVhUFyE
o0+XdiE/1+SnhwOaFLbU9RFeK6a4TLbTiXQjA6Bs8tydZyc5gEE90FxYm/39dmYZXFm6A2xgJdHv
rSg0x0Nu3Dra+YaokKeTnzVTrYJHdEEW0VZnbKaoKSKBBWgrzHGQCqpllpqVsjWwMduln/o7kt4r
l6eDAo/t59BgQGtkX2Er3l+tXawVdSFKPKs2C9D9/lQrHPa9qwRGV88LpvPg157YKLJWmAwKch9B
Ir/Vi5td/28mACftDIlERjPcXJWzkphBSjw1t9kU2gO8scHaUoJ1FmfnnWxdjXsilfvRzRt/pWaW
dAgue+/F7RVFRn115SOgBVF854qeBVqXJwUCx5rh5RvT6qY73AYsL5kDKmWH3idDem97mNT7wKXr
RU+bTmT+N0J5UzdqCaen7elFVuLuK0cYgfkjiDrjttG482gweDe9poRVFYhwhzbd/Z8KbigNUXny
E70CzG7gZAIjDmEUeHXFcr8tCyLh9FdIUf5mxpu3FbLrGuHPwr55U+tHeMBwBdjgtHLZVA6p5Lg2
wFYJ0n3lmjmVGTjV1lwRXjPO6WvpiESBRuFiKl1k5fIUM6KjsPoeNAL+RRaQNudl1uFDdt5ycgii
7/iafbU7c1gf3lU76gbKO9bribpP2NM8wqKYEne+0TRoTcvKIrGbNBf5dorx9S6BtJSpJklzQD/K
WdLZ8NawpTiKTQ4C5rzKKV9HN4XKontaHv8I+McTRBSUG+57dbakTkjgYgjjWEq+Z8ZtL3UIxwCd
SVYU7qcWKl1lIG9o/hHo6toWauxJUbUYKG5oCOIlqKVgktl+F89U8c1EMOILPnQte9aNe57GCck9
P9q3wrS6gT0oDZKzxpRxeHO2FrKHsX1RxzbQ1eSkKDZBQxoioEhWBcX9jCRi+B5/SFSC5h64PHs+
rtI4ICrXvuAFkV4rKbJ5Y5pKdCgiIOCEU6IejSKr3Y/R5azsUX7vApfgGBgER8qTKAuJMF6bmL/S
4RXEjmf2bvEq8FHb/4rMau45GCWz+K8mPOPX7wamynGV+GxJIt9JAkeP8b42Pm82IOTsnXXqstw8
iWCkcqtbWi/YRdfC7skPMLsYvvORfwrAuhmzxIA+fwr1menRedpzdI1jCa+mngfvGnHU0qwqLm7M
I1GfvwHPjsFoVNV7kSUhSLPwQFmIZ5bk2rNnQ4nxWx5Vaqu5zNyrSIdsLtfgcqfbEXiTiwfJbsmY
63/mqFRW/nzcyRoh8M0FB8wO1oV9uy5VgUz4eKRYdPa32e9puUQJkenPTYPAZLRAOnV4rvQ+c4E3
hAOdGSY3qhRALtvPBNGYp42cwEiA5S0DHRP5pvJ7P2iXnm98FkDtdAWmV725tUybn7GZ4kxslONR
he590ErT2jcVvmPrGWYRFAZwiCe/0dHwT5S0Zwd8a5J1KE9e22vKsYqeuM5+Y9BtWv4tZ4TnqMls
0joOV9NBMYzmL7lkZ3YX//g3e8Dv0NCwKwn9TEY1b3sOMj1CoGS2V5+jAJuQwtbAf3AoGK+EnC0Q
LaPc2zA2G4G4qCgpE7glH/pCjn47PM/dw/IO80D3siE6K9LQjauc0R5UOV754fwT0o4Sbl9gWwUJ
u3NsDkf7CF/nQWhPJNn84sA4Mfq2mmkZVJBRNHdm2rYha1WOUTUI6lnl1d4S/xBCyD64wLMe2Uvc
JspAxIItBcykgTVKSPB4uMJbNxixfNHaiU0Q7po3l0Poy5igBNMk7If4Egyi2C7Mr6lG8Zwhol7T
wedAJL/uWAJ8+ibN28uv0a4+juXUp9Kl7dX8K3jAn2qSARbZfBYaB/SKylEgjB7B/DpngoJ3JEKw
Gjpkw+qDGgluuiH4h5IwKUD3GB2W7lwd3KvQUX6Y0Ep+9b8wJ+17kBD4RFyMRoABCfGRL0EzOrZu
ZCpCmFweG4/HP8LaWQd4EXkeSwq/2lJty0T5OTy0JQJa3K0cZ8JthKUDdbmyJn2B345XGg23XoM/
vKjxIEQIDI0Wgs1Nhs2YH6AayHwH1MqsE/DkKkm5yZFoDE+HUQdF++u/4euC+nKa0W4JeiuaN8RO
R9rZkkIK430m2OGkHsT5LOm1iQQJTbL8hqogDXnsP+3l0ETAIPH+u/5BKVBQeNU7nX50ZOmKl3se
0vvjXl4iq2/UkZIvt+CPB6F4NupkhaA8XoUdkAB1PuK9gJHT+DYlo1F4QtR/eSjturwvF8W2fVam
7zPv5J3zN0E7+nkgfxF6lp7/syzJBsSYghrrYcab9t/cpdarygz8Z/4+m/nDCW68lsLhUxhLTRY3
QDWjOLbnqtylmWy4ZwdLK6aCrybGpbkF142Qa9YmG6LQeAxX080KiVdiDUoIzedveSfjuNyU3jwu
QVUZ+1RBGgjgBljj0zSweZE1sPlnfthscXihbcQkCiIgHQi73EruBdE9oGSNUFW6p+6qwYGgygv+
55s4HaL+d3vkXOJZGbYLNM/FJcid0qzY2jr6MtnlgXy1zZ11//AD5lR/3XMW9iRBKLKmwP91jiKu
ngfqUxks5+14clO6PORDspu1FKay4Op00n3Mba0gr8QUmpG1LXIuMgnPIiWRr3Wp/bnGgfYc1moH
7vYRNHYZfIKOM6UZThjoyVGct19H3JXBzKAoh5iVBFlXgPOsRpXPP+Zh53j+T5H7jKY2Xo6rGQYc
dai5svb3GV90EIGT03i0efGgTfHEMvxJFZZMlXeNiIEFhP8zGT8nnissjggaQVSFwf6Um/ehhRiI
yeXVLj3L7i2HlWpG3SOWNB4F32SQTfj1aoczJEQxah51FW92/aI0sU3A+6QadwIj4uFuaq///TnK
pDy3PLVNuviQvSex9rv3ZO0Xe62v9ce+VUnHgZyCraoIc9EJyT8vV52YrehcSp6Ae83UgeKDukOr
Z6WQR97GJ66zvehqigJSuaGQHvvMMiN4L3uM2N0k73wJwdWwBzJfL6AKFoyhqD56lErURMkNCxIw
rAh9TzKdzJ7+zlgDF5M0FFJuhhP1dXwDHubFUPchq8/AO4i6R14Lf14SERWwRVTsozAfj0AWNxiT
X/ByZbNs2RcIQpq3GIXD6LNowq9Ccllm+S1tR9E23EyUTZXfTwd6nUmsjsp3MHD3eE8I+WZpW868
pwU2WfPwWcAw2wrnBHQPkKN6gkfzZ7MlDJjb0iRJMqdd2aAhi58uSmVvbv0vMxtEcpceqfmofR/Z
5/Ugrs8w39LIILUndOCLB5zLd7qaqi0Teg9UZH1ZF7L2gXl1F8L/N9Llf3rNdwlPtjIcA4oAJ4Tw
RANUQU3snwcfjEmEaLpJkIi0Wy/48jvZmV6EgVT0aOTvv616ueR2RHjmSxnrdakzz0pLpKhYcEWr
VVWHlliGsA+v/6MAjLpLHtxsF3S+JBztWaGP/1dE1ZrKcvBzy31iIzZLc6aZ+dibygOfyd70VEKB
We0q/gXCn/+jegFkU5OGZiAczI9lv1fxGchw8UabHgPHuGlqeEvflq/I/xkth2vqGAPzyxsUfHrP
1txSBPalibisHYfiN/8dJ/uTysFp1UA5wQphxCfEIddDrz3gFM+cyvbGu2rzz9a+DcntZL9uY3Od
dH3HSUbbk3mfHxQK176tZs1iL/s7G7rrv3WvLSyX1muqmAT+aAwMgw4to+nnrgc0mJFQVF8nnjff
0Sa8FjZciTaqga6n5VBlzERbG+o4YaqtaIrwZGvd5S42ZPkPVb9QK27Nl4m3UHcDxU6Gh7tzCHI3
V0S/CSQ8ecBgIfyN8gu2JgNd1rjKq5yLiUFf1G1Sc+hDDQj2AyMuQHR8FB2rdnwMreo5576ckgSU
fXR+L8+fhqX7WIO2e2BF3BpthIlmSbLOI88ajhTX7dVgJL3upNU6vYk3wm+3qM+CC5A4CuQ55ylY
DN1FwK/AiyuwgArpujF57/3YprWws6vAgnAxe1VQu59Unq7nApIj9rqYauN7yVrY325SBDnlUki+
6E1jcHfy8kBylNI30h1o51Vpa+q3PdEfOPuH9Zn1LY049JXAVXsY/YZcBBh5/Ofi4lFGhDogcaWN
kNLHcpXo7puwbLXEnnuJZbJaLlP6znXq2vZ2nB+QUaUSHMRtmSSHboH7udIudkIVX1ZTa4S+zN5l
FIWDdwoHDmNXcWJHOljta8lLQIJOQ5lP9LV/+9+D6ET4bz6pHs7u0o7862bJ8CP5U3Te4uZXQfWg
S4i+d713rMvVeZ0sg4pLfI1CT6raGKfFlTkhhcoSq5Rc46vx8V0Es4xwokP0lPIWZAc4Nj3cqf0n
AArsGjP154WkijhHn/Eo2xGIRE6CrL1v0EYe0t0Laq4o1KvAlswIl0AIsdN2MTOmWHX/Gws/ibO8
NC5O2uewlvVCZmFTcJTiGi9BkLQYeQ+zfnqTxx/A17mfg2iDjQVlyWJcKF3RP3woxlM+v5ny0kxW
Usbu35vgr9tL/cpRJGtdn5qlWS4f800szS9EV6HZA7bZ2n+s6lfUqXyJ21D0m8ZWp9AQEuU702UM
zBcqcBh8wVOJwi6kFJW92G7Q9DKJAcv2lobApgLV7SISHr/NQJ8iMxHh0g0rm4tY56QbHgP5HBiy
DcvSXJS1M34RzIJ8CMLlFLJh/tEbbK5mvBMY2a37GZs90vbmvuq2mfIQTD2O3htj9phqsWLomKD8
D+ZH/QpQ4lmglturKbuU2iiJaVIgn8AdFXK91/PZwjoqV/05lJrgmtnGZZV6cpGVsek73EfeosTF
maR8BFzOz2JQ/V26oEOML/DMa+hUt0poA0Jjy2gtzmoX/WY7Tgpin1vO81nX9KXw+HAulRzWVInx
+C3hghW/4et05wJFlz0WIzSP45OnRLwsJ0Jg03kgLpte2s3dJkgrfzDfehNhCzBD/ehpOJTe6Iae
3af1/wu5EhZNdks9fEppzZBxbEFA41fSLCp6cAjeNtpspoOzflzJVDehM/QY0zS2dJPNX3ikiN8W
wTcryqVl7A2oxFIbmyJLngeyiQ3xEkRc8or8xykgYq4T0BntX68smm113P56FyouR/XQAhTfS5cm
2luDRcWOUO1Hcs0UEvTT6P3WG/mZ8sA6eoYYaAjs4SndJnX2yarjzKbXf46EAqxJL1PK3YJI4Rc+
7O503HppVgSQBHgZwhDMXJ+4R1l9Z2eWhpkuQCkd2xf0RMH9PP3uScCfenqFCeFKaZtgp+1zPIcb
4vDOFpOlMX2XhsO7Lyj6N7NotM6WQyB547i0pIlAYPHNAhtPsApLOcU7a2KWkLSdjk+SpyoOrUqD
/xDI4hOk8Hqd0YsQuA1beqXQk7Yt+WPeSOkuWJCjSM3z9Tv/Q3lVQKi2D/I6aWF7pghl1/o9dRFd
XVwtAU2s5Rf/gkwMfyKUN+deYyfsTPtfZWWhgkb8Qus4E5Lr0TPKqh8tSzNbqM2KQfnuYsQNdG7s
7xR/+YykXVVoynwBepRoiFqdjqPeWVjxRwh98mXXmsDycJKhZbMe/obxVcoVwFjKvVVAqDrIXXBi
uplJNdLDpYNbwfNg8ZOpa583Mfv86tElrVPVvni1egA+aW1rnXzf3lm9LMB4FtM0Mhp0BfEshndo
8miHUSKyr2qVgWMLPkEQQrOObI5kH1t1qac4YtndBrOgSZah6pqnHDLQhfdI29Q/AqS9q4BBZDhW
nPcDfUmnqdyP/rzgkA+HKPIxeGMzsLFuFUJQW3rRWKuXz3SZd4hZMsHgZoWPIV1ZwVZAcEQyjEOt
ZdBovJTTuqGnz2zyaW3BpgvDb9HpJ6Q1LqVf8OYCxex3OL+bwEX8RcuyNRA9mpObCez0kOOrYouW
38eDQjLk6cMj9ps4SKJezn29kXr4jK19E/YF5t+LtD/W4P1zyRQygyv/exd9pCGKsFH5fUIGZ35W
8BWWgyMVXOsoAyLPAq68mioDKk5fAMTtUxQjjAmWbbABYc6czQ3u5nbEsX/FRsPKXItQolfODWev
BfDxZ92xhFGKWJIhlesAqvy4Jycj0pBUWNgYuBjiw26U3NXbsl4mijbciyjM3GghJp9qUiOcUiXX
iZtH10gMECJ9cM1WCLmUCzaiJJfLfSqRFT5k05MGlL8B5dhqybTxpf7ZMh2ybDXu4ohS4Gh39WrT
kpjC8e10o3TClOhyKv9qqX5r2VO8634wvKfDjCyFKDNOxckqJG3Bzd3WxKESinhuI+l6kIQ2/ovq
vA3e2R5GIDeTu0pE/vNV6xoHuuw8A3zt1rFetxI74JEWFEeDqV4+0csjD/fKkHV7rskUH7UXLAFg
5UKQVZYtrsLpnZ2QSl7QdVCqZQLCieFKtfF/ZXHyDU4GhDJlzaXEHgNCTsYQ6+ZnzT/Fw91YarZC
sfpaie9hAgKugyoormbxuluE7IAN9MzFlhu+IqKPHMhE9B50MF5ozxVim6TCdVDKfxmBjVrE61qs
1vIhH15PgeMPi5OlU3ogFHItot1CJFiZEO3lUHx04tLLRoCPbQkC2tjXxWXmexojLe19DzNG16RT
rI++UlD2TjcAtiA8j1Fcg/d7nUXjo+N/epvkWPuwmSS3J2tJm6ZqWB8eRj7Hl1NexZGe4JsLXSrA
29zlDsV0NsDEPRDsmcN2PUde3uReKYUMEUUB8Otq+zkyh+p92so2OkSAX1FIWHk/UnuwL+yxzXcE
BpVqAEkmVYNG4jFzgEA6EVr0c5BICStrG7Fl/ME7iqE1RM6Qj4IvM5etyXQRBu2ZbAlixpR5EkNM
26keDSiIcgGaHttIhY6wB3SqjGZly+i0RzQyeTRRAPjFW2+JPCdneYH+WutsUKPpxn9PAxcPaIRz
mZNUcu8cJ7B5dH4KAdjkV6r5a43hmhoHaOxDpKSH99sdsBBSOwCMcZkGLRlcg5PDNKb5W4o+kHXP
jaZvc0w+leX4cfJEUkAIkob6STgVinFGYVDQrcGLlLOrWiacKrkl5qlFffEmNKdaTvrj4CWxC7nv
cr9k+4mPc0Vg2adfoVH1Byk0f0CPIjMKgzqVs6zkw0I4mVD7fz6Fgo/z+hd/88iXTmxWvw+u1NrQ
KWhu6KtSxMHEC9fdR+qo9e0yeeBW7pUhbbxhllWBL3aRbHOgTs6Ynji+ubCYqavHtti1YKqJGOA5
OiGEJ6+EuZ9btI1102d7hkpr1fXcEwiE57Mco7i3FaeXG3gc3vmSw8TFCNvewfuvqLMmEzMgDt5q
R9o+A4OCwYuU3loXziey6V/f7Jc6xwCcfiK4ujXlGjkPtOCxBuouFlm+sWpUfwEPuWhiSpFPXfZk
0yATseOs34kMkui4wJqBhroBpMYglPx/vBRr4sRik7VPCWNqZLMYeju9KGNO2h8hrJGxOjjar0hR
SglAJrw8CDCGwaL09n0hvjPkdOTR9qPR6t9F00CcepFzQGPNGULv9q0HE1cYCo9TS+HDo+r7DMW/
sJrgXFAwTayYxpRDsrz09dGGZbA7vgYj7wV1WfQdAO5ZJHcyxduI1EXBWiMYu5lY0ZCuJla8CIh6
d/1SZFfuArlP5dbWkMetQFPzsjBjSBdxC9do415t5R9OR8/kIzf3I/Xxl/MqWba6C8LRqlKpb/Aj
eo1pePKuksh9Q+VnASLroRa4Vp4CCuhNWHbtyyEet9HZpPksPjepc/JjIVvPeQQas1SHmts6ZeAK
EccZHVHxHy5FZ2C7AqOIc/oEQbWut8dGxpwH6kyTgFdYKKNakekDqYqFFrsKxlsCHWGSFw9HSIzl
MFeMdO9/bRI/f/CCH8IdXh6ZFrjyb7OCuH+S+f5uMxSTV6QOwsRf9iBWowmJUj4KJBuLXgMa2rgM
HNLkiTsLBvynRcwb1rLvJNWWA/JcvV/wKdEHwwiDORas0Ux8RxO+8+2y3k32XM58+vwJl7e8dB9Y
hrCNMI9O0cHeLrJl7zP2RLCZkXO1s3pShur6XRpxl39e7j6cYvikKFK/hXsDSGBf2qkZbW8FEf89
aJfoSPYWtbjGx8EKiPl6mCgp2F4m8Po9rPnsvswMloPNshQUGzlC7Jv0ou0cnpUzgcTp2Gaa8nRM
YiPOlMFtnZuLF3zoasodRi8FN+3RI6L1RlSaO11PTPMVxQhVVy4crkfYK7JxdwrfgflB4jzcOQKg
jQSNQyaZYaveuNcYwTajiYGAjVPEmXJ+iT+wLIwcAl0mICyM5opiQtYEMV7upjHmS6G0/9pHDo3p
OY4ypGZN607EAz5Pi83VveQjbJ+GvHTle6ju2yKs096tn57GyiPnu5BzzmO5ZjE3L9mW83RGBhSK
V7KUVChRM5nPyMAhc8jpNagfSpRtbQ/PdnuUTE0q7HxNrTv0MYAiJzt73ppU3dUWjK5SlZCInL8L
BskEjonN+s8KTCWbZgH96VGevfb0xDq/thxeBEHaBSfQIqh76x5BQPRblErWVn5kBEPvDuUSKGr7
Vd/oVRsrBl5zLm/yj5OwHD9r2DYKv/MzUQA2gMcRUV5Us5+nGlOVJs/5GtRIkvTr13ReiDDxy9du
jSQ5EKQ6pCi96khxc+LU5NpHzRBVwOnSVjX0uPuNjvP/aqM9jWZ3nufifDM/36uj6WNeEEmYFtZm
gfPhX2JA/zIpGqU1COSTfgikB/xGffZfBy6Qmyu0xi9ayC2kBsAOe6ZNQKUD1zoUtYGTyIvEdDiQ
aNPcgI0wNRPfWGKBOdj4YU7R1DT7uNTVesNYghn5Q32rPKWIaKq7eLRG6Aku9Qtl/Ped2xfzJbHY
uY8U5W4+xt7/3NrLFacWbH1+hecthjwvvTR5bRPMZGGPRCMtmLFD4KhF3yxRcpbJLo0ehum0H/Ar
Ipnd2YdCjeUFgR19qRCkIQ7DefntxWZb3KtNwum6HKYT8e66heaRqm3zk7TgMl7zBgrRaCXT4AFp
eWt/bt3MVlMYXRqLXPSCRzW/wvbRtB9IcW6GnNBKYiHrL/FyNzinULrLvtT6h//R6wShJznPLSLR
pVnAxJ002dWD2/Lilb+cIlzot29CQkj/5vHuBrGIzD6w7YM7WeFP73d6Bwbv5wNctPF4CUv4u+7f
Q/gLTI/LhBEUqtjL496Vczvm4nnS1awwkWPlI+xG5B+5Szw2zx8LbvZJUvv5AKb+JS3qjwY+kDNT
9kCL1EyXrI72jXQq7fvq1lPz5tnm7ITglpv2TJBjRx9l169f0/N5Ufc2Kccs96SJx251sM60eJ+x
l1lqSQc5oOODny9LfrHZgGnSMlVda7/Ww4wURzvV98CzImQOXUJMbPm5gnDsHfTxLHsg726Bz84Y
UlojlUMhblB7DBl55vryDG1jW8rN+kYr8Z6cd8MtVnKKKAYRV6VNaUOU61jKMDBQtN5NOA6iXWYC
85O3pGR+wwY8RJGZR9jpFOGzrnqp48S+Enbva06xEN+fgJM/V8tAsYzb/G+nocMhwD74Z13BNN+A
7uZdCUaMug6hKyo985jXpaygOPKlZAo4kFLkjAEC4FDmtq9jv5Nuo7yJQQIsd3+pfNaxsUyZTOQ/
QbNw7v94jqbnd/ObSJuVtIX5x4fdvD/gFWijSL8QA4SZu86bCgkX+p8zGPsVmnkJdwnU0BSn3/m/
AjsHy+8Gouu8ER7qfGZjOcIjt/8INwfKkmjWCKAMn01OoP6W/lau8v1yw3czjLBiFbYpFU/GhJAa
W2AJn05b+UljsO8lYuhwSFGr+/zg7WdLW2j1EO4PB535Wqel9jFS/nXuUH2sHPc9UNdRLpTPK69Y
yWSH9Tvv3XyQBWPo6NFmaRpNPqqVfhfQs0I/JJP2oD9g0BTmYa+4C+WWl2zo92PVD2ijqpE7gBMq
z+au1ZVVkcw3Dbg8hr5U7d3zvhSY8wWW3TE7+Qx56uKr03UP309IcrrCPphTGr9TN35Jq9WLszGn
HHD37hO0CRbiBSIAywbDKg80V7cuS6dvN+udrKt3L1LY0Ld1ANHi6sSqRvC6Np/yxMdZ9iKdvFRn
uPYvS4tmbKVdJCzr/9DhCPPy7xy4LFYpJuvrC+uj7ggHhQhWECadGSGT59s3kruLrEVOVa4DKbrI
b0pzKAazUViunPt5HwhDP5DRyPdILILLHXXWleHib0zRwHWOZTqnRfZwkL4b7IuiP6lBSEKIG3Xa
63B3WJfHdEaeU9+ynYr30vcZja5IggSqlB9oTcPdQPwr4V7wv4M/S5Z+JTvyaSUn7/0K6Ig02Dii
lEhXGszyJ+WrTcwgPMAXO8PIodNp1kOiSbY0cUADdbcmHl4u1Th20t4Um7jdKGVEv7mZYqPdfr+p
PYVKu0Up+cWTlXfFKOKONlvce9Rc/HfPJQwfhcGCaxKv9qe/J0AMfD2YalsT4eY6YRVbq7UQruwp
hRQ1VgJVsxXbZqVoeZHb+DL/BJ7hvMVHqKbNfFH217zTCNsJy3seE6C05WSjgKltWgihhTWqMp1/
PYdfesm4ZzTVDYmI/AoTua+ikrpXTwaM+Wi7VtcpS56lEsbJ5uexZuJgO8HFUSbdq3hPoVrMu+bM
AcaSoSDC1WCFI95ugHET5XQYd3llsnUmDwrvMaHVJ7tY0h8bYVO0QKv9D1e8YJz5WUiYoRHJJZq5
5Y8EdQIT+YpX7uEyylCbGfiWNwvxHz01Y8c8YUSuvMeq26XfH18qMHJMD9sSvSNNUrHDx0tbpEDI
brMaqxScIDL5RNc+uzvFnnrr6yelTiSPLt3N6V0XkZKDXrGulrjUPmMAIp/IACJlO1fqUZ7dOPSp
iEfKF3jRfBCFudXHYl8MJmJxmJa/lPi2+3KirS/GAHyIxm5yrUQidd0F7kjaM2qdbhcyFidf8GwJ
5LD1VsW8caZtyC/uAA/ReARWS6j9AMEMgNVw6GCpB095qDcigTdpxbLAu6Yy21Jpc7oTGgJmz6Bh
wlXrCrP1rU3aQxyzZZJvQJEkoIIa9MyosUIUHowyOl6C+LWLWv0ELxNSwLaE+lmlIgnijvLnyR5E
LRYW6a0ewSFjQ3IyZuQlMsNn5S9MfclS8d6eYom9995TSNCRnKe8QEA/LS62lduFb2+aWB3RC7xy
XUqXBTCa/swpZZ3LVwBL97xASdH81KGdhx4PeC6WjvvnDDIAFnt2ydQ9GpPFw03YWMkqIDrOIaF1
SF2bQXrxYHgoPVY62Xom6R+8AHgBCyXcGDA4ElEhL4irEJH1P+iIv/ZW4IQk9EbglgrqcqIwaemm
0DJM30FAPnNVdG29H+FlWEOEVToNCIa7P6w0vfWWk0Wr8upGRTwwxIjq4b6zWIQYOrIsBkLbtC/+
kaWORDU84fcTAzz94QhOdZSlwfDDImanLKqs0ZsSmYQrD4r6pfFdG8BKTax0yuci9g9tMJ8jxAdW
e4eRYoeNb0Ghp7ZdWtFRX46SJeDmpzUA7rMPS4EbCigizNUKJ5Np0ekupFKxCDU6EY3TG4dC+4pj
W12XDuNfXeyyUMqFRCxAQpv9+FpeLygZZlRHY5L0PQOh5bDGlpcFlCgnNClQtgznu2vym4HuIm/I
j9a2SOV2d5QdsTBReCbF6VOblN9SBiJk+T4nA0iMXiGkCgD9Y0KrOYiJSRH/7FFjtFZRYH3HRwAK
877Zy9Q7OytcKP24KL4ZvyEFRtQbnogkuJdGHPz4sSPW/vU5wM8bfya9yMJpyAYGMmUg5tIvdXX6
gfQyHKRUmoL3R+2D4o+rJcu4qPWJkXMcf56mCEuv6ALp+d+E3U9a2BY/zjcf2zYQkD23qjjBCbs0
nWvdEB4txrjeaV+XYYHI9IgwOvEwY7KCLDNXLeYZB28RacBzLHWP+u33BBfeTksQP5dIbr3sjql+
Pw4X/EBlMrCF4TIhwKokKZfRLCrrNSe9SeOsCHVa20FmNv7rJore0Z9w8J+3cJKa97AZ2xzNSxv7
3qoWQNi9njtjUkeYqYR5BzVT7I6HeHwvqzhYE/6peQodRI9Q1kG+BSPm5Mk4pOAm9BtdjhGxCcOY
mlbVTkbcnY58vCi0IU+nhP2i3fANSSMkAnBYdydFqYV/O16GBBy0Uc8eFO/IcZledfRdkEBLEfFY
Nf0HFk5G3VgV96Aox1ED4y1d8Z87Kb+R7hU6NkTe4NwE72t3/fFFoUBOxBB7VRXA/8ka3KpL7ALD
QsQ9x1wkst7Bbsiwd1G1DKvAIhLDOUyW6zny/+TEarcZT3byIo8uShw4nFz1KJS3czhTMWWWaj9L
i/YxiSZRtJz2DWJ7Pj9qq3/jRVoZG7IvqNjWNE0FRcSJaWAngQba24g8jflZLW+sp3hEMpex8oxL
zDwi+gDFt9eExcjZ3mN1O0i+TmKwwtaCTojJeq5bPyjO3K9144cbQ76FmcQYGl/BdCr4XBLLhzON
nUsHrK3YhHLEnsoDY0fibHVf6IjCh3IT+xJTe8osZD4Lay+/3KjvtJe58DYCLYHxBLFKZ5YVxEku
7mkRJS6ZzyRq1NXBGH35LF5PD7C3zgQVdWsBvorLDWDPKFZw8wwQTc8aUutVCrP5mQjqvdLqGmbl
ts5WeCBzmBGSXl8C/MHNHlJuE+T7qIUYt6+xN7WfeMfhpX5R8aBXr2qrmYrDDs2ShtEpsk0y/ZeI
xNt1PFNvBiCtSKxvwD10sqLCouunugIF4+80m2yKbJlMmpPxICffXHwmt6Rho1s/bQOBZa0nUs6w
FfR88Et67MQqRA0C8jioQ0lOt9+LzzmsnI5AUeDikRWiQv8ohf6PP0p/WK3twms321PAMBlJaWuU
UsT2rPjZWfIen2wg6vdL6ZwXKlI+EZxxAm9kI+5HOQ31M0a9Eom1Q8APS/yM5qZfIS9LP3ArVOBY
eKa7SIOcJ8sfa1mehIFCsnl/sVBVNcCPHoaj/M8263g++r6KalGh/tPr6YoNhXS4rAJ0lHHbqDnB
rAbye0hCB1zqfUzVcFzx6MI9BNPcsmju40k38fO6JoiQn5WlVOzHvpeNb+iKAqAe+teLYAQNQH5W
hyCgIV+Yh1kugtfQgxzDSDx6rz0ov53OZ/xR+sMV8PKDko2WSNRn6QeyfYO/UrZ9+k/1N8T3iDJj
/FDeWxuwI4zuEQ4DG9xbkM0x2xo0YZoFzXKcoCF+v/g9hSi5f6tvzcUhAM2wL+ydwG8nsBdZgy7a
bnTzhy9rzq0AslumRDYwty0Kyps8gjSlcyXwWnqhDyqfi2ngROn4hKdhWijbJhAuV/L4JVK2rue7
N53m6gMJzugjgftr9yZSa+IHwUtImH5C2M6NZWY2YRUlVbP7W7w+avhpLdxDbS/vIveSmPkzuPr+
BmfPIe3z6jNziCxKeU7bd8VPWT4I8UDRpBZa2lFdeFrAPAZsXBihVQ3yZ240vPEWFdzkWytir2E+
fmN0mYF03+S5G7+FKOZSEGMpSClF4EYYJaJE82OHOcz1s0MwjZeCCtBlQwK9YvZxgKcJbXeATp/O
OEf3U0VafhNUZsv3b+p8tf4r0srZ/LGhvgOhiO5ynEbeIHxCC/YFQuVgWP0IM76jlEo+Dij1xQDl
8QmpV8TLlbkg+mhxa1GvbbXpPmew7iZJpNGZ3Yzw1x0iRK3n96106yJUwdGNMj1DFo1oneE/qsLI
MF3fQvmtbctzNjc5JRobcftPyg/HxK94lC7Vf9L6hYBljmJ41ad/zHktB65JmU1TzR/Z+U2/L83k
IPX3H0gi541PZh1lfOFjNGsou4b6PubTXOJUPg7Vht+VBMk8zAetfVPETac+B+CAKqL05AZW5Ik6
i4JvL7nJ7hmD6J/Gg+Z2RJx31FjW8xYK6U31t/7u4hKMRBoKxLDAxrLPvpxlxf1FH2GbR2FaRIJc
EYuQ7Ga+El1aQvqd3N9owdomAzgCypvRyCvofZuHW8cbZE/GUr4sG7E0BZR+eXmb8bn7dYgxd6BV
GmTPdnTUQdPGbgmN9YBs4O/BAb4uXnXUXtHm/+DdDaoST3aoUkl2Wb8mjlvDBu8IbgaYWk9MibkX
hXE5/oq+NpbtL4UQD1bqr0iHFt/mGQ20exerjQ4wpStw++L28wWdhahmLxm6u0l3CR6jDLUOffhM
Be1nXvypoH/6FYX2cd9wzOcLejzNVXroj9KVwDxjCZ8oY28gK+zCYzHzTa3jYNT+0b1reipIvFG0
QawzYhrqpAdJr1EsLxbXhHH9HwVjbO8jeNI8rpWsqBRwO+Usunur+rHBeAyYBk1Sup5rfL+hWeDS
LRhVB8uHzATQ+BAFwPEOdlyW16XV98hkjoXMSEJN3J+SfMfCQYEIX6uHbE3MSO/lCfF1nJaaK9wh
+PmAP5dY2BOALUjsJtiO+0jBL+ss8Ho004O/GE0tXmHEVScdvJ2fjoLRpCuZIMbl7kZoCO6hnNEO
WsApZZCm9sFSj9y1UrbPyUX87lPvANnFSxBMAm9pDAiN85934Z/78nxd38cBF5hnsSbtz0KPAa6S
+c+5DS2mzHlLxLqNWFlj33br1xD0eqXKg/fU5/NoDTF3WDB6hlUmRcVLLNSCH5Iy+lmLon0cfjTw
PQRK1MBRnvxBFYMXX7Cnt8VLEK0mgcqgZZzNJYwo0NcsIyIKb4ZD4mpybf7m7CaFPPUEwKUmMkDH
8VUwR37PdOUtYxxYXDaLkiRTe8tesJhnIYvVNwUzXXNcIs0ruw5xtjEEZdfEaZG7AmcHQ0Jsbvor
RGkhObSTev71OcDUSUsuVw48mSykIpd4XXlUGbeQvMrP/BqHDcjbioEXaIOZxf2ar1LDS1zjIGfP
MyqENIa54DaE7tdtyZV70b/50PMkfbMRvCOZRDMAmMS3A3B/0VQRhIN7UdeLhIzezHX9Nc7daLpB
R80aGyvdBlWXQNIBkGYH3gOp7Jfm7/QxGgQcC/sbUamj6B6Xt9i+gS4DTwAyzY9tjFwSwnBZW89z
PFUH7n5QotPDNWMmCdxS6KkiPsOGVfmELJGkKF7nrXfRWHes7WneKhQRtiwj4md2vQVTgSLDc0eD
mA5Nh/WDzzehS73WrjbXYLsVZQVWZi7FsenoUOiYTx3qSNoqXbBSQI6DmRpjHVdTztsPuFcisEgo
J7HxQVEG1t0kd6oA9W0hrZ0rxliYb8N+0A9b33m7CANUJxuUaSbUdbiyYKcPBcGVmRzL1r+JMaj2
vYeQ/y/eaBDZwILtuGTWNPuuCD1xlD4VwroXECXO4OzJ7lRPegfH4HCuMKlzzqYAkD7gMy0nMAXD
9pUUFQNURg2S+gfQJJ+2WFte/B9xPIbHTPP+ZHU1G5HRP1MmZdDF/spfvxium8wz2HQsV7hPN6XD
TH++jgtZl0oHAyfqu94+sBxYYGEggydp5FaOkM3gSOuK2fzYLNf+t2HhKt1f1Um1bi5093fue7fQ
GO53yXj3+90Cv44tTWSJ9MED6rtkyJpa0i9nLFOs6i1TkbIdZFDuJb1u0VMyJliMK25c0nPjxupq
P03jNcn/c7HIFWDbx+E3pQabpi3X04f3qmpb3f9UHj4+uzM8iZFmPI5PVH9ICRjLebXqYCVO5uSE
V0F4d66n0xDB8d59E5LwYrj+sjoqZ4/GMYnXWGXyu4DrNElzR9ibABO3t6+TKAGeu7RsZ1ByyXHc
OiQj+4rG0bQn/+FGjmWZjthhz65+GV4jBxe58RbR4lT/1FmuXiNrCHjy1q1yVgJDTzYzHFftS4Gg
+E1CJVbAYeSZMbf6eg0zCbznjGzTkZk7Q22hcEimfPwAXrf5hADoSuvGijJPLIEwDais8cX9uS1+
bOQIxef+Eb1tyd88t1jCTvqI2fHetjfqtIC1cAwPWNNamdvRtNtvG20G3bupme4/dFXEdXRTpE7b
aShSx5Bv1FNxjYMnzsQ7C2OpdGQG39wifyR80mgi5JD4rpE82m8EVAKhP4l+n/YnCZ4wdLg3I+Qb
ipuFwzDofbGOCstKIBeXtZz8EusE4JBLV8gf2781tFXJQNUEzD8eOq5CK+fAHF+l/LkgfEgVLpWw
Vfn13ZNblZtD7wEJtja5rrv4/Nx9/Hf2kYSL++dxNfqBB53Yuef6LbBnMb83PFUh+qYEliOy+5tv
66TZYp2I0WAVKlx1CqunW7VxClptFW/S1gZ5jFSCcBDwpmB1a4omlblZa0yUbx951mtPtpTRorMp
iSFtB2DjWO+XVUtxqKv7Rv061qIyF3P5+wA/B3BphKe7b8ZI184P96yIuoFLbZR6xDUko4ifJqCw
r9UjBWAIC0Id5dRBbTA0HkRnWphfbr8WNyP6HiNUtVztJzPw4vIr25CU4dmghVDoeXx//l0ZCfRv
j10jlfJL1gZMhO7ext9bSX7CN+qOpEhyXEpmns4qIwGME1chN5utw1vR03eLiYKSwNFeHehDdIxc
WehCG3jUKiAAgmgUHShEIbKJLOPd6NYOfBjU9No9Ma2XSD7yRs9iCwV+7d/OE84nUea7rRe9kNJm
bFodJMq9zVsVnAxe2h1DLouTKqhii8HkpQ9uZUpmONR5RsmarTs47FqZm3aXspM3vVyivPX+UlCT
ii+cYuxEKwQOduWhu6h/2s63xeJc2sBGyQxKqfS3G/gbrOCjfBXArG07G4BG/W1t5SYY+PDy0WXo
EGohr0Z13xFEcgEoL2FCoYQ7EzGPn2siRsWV46KwEVqiwcMHq11RbvjZwcukxi34bxEkP+IJYJzd
XpsPIHuORK3dfdN9Pz9JozUGW2hakT5NOa7TvTGu3wwzSuEzUVdp5vNXXjmn+WEigUNdfTlnjVq5
1zHWIANT1BiD810Jzs2sJKbkiXrugnjpOaKTtU+SziHD88H62fCMDmNXcJP0ZUC3KOmyn4uMPz1H
p/TmOvxv8XnNLQym0zwBgTDDzi2LIhzK15erh623i4VfPgrKM+I98IX+X0/YGlfFwFuz5UbJK5kS
kVH17tIpZ1OAmxY5oN2jVUFB0IYwuRZ2fItxnUb9ktmrU+9cUAkS1DzL+b/ABgveA6ze2prLh818
eZzcP15mvBwKOSfUgimTp3VvKwEXbX1bhoGg31S5JepJUL/2QQpkh78B4SAMPtusGuJTpW89jpF8
xei4tMUM3qfayjNgSOfWb7Qypt9Xp9zAaHa6BYZbXrxclM1G5SROFbCB7ZWeh8roZ5DOXulym+Ra
fYkG3g1EHftPtYM09+MnN2dSUeNXDnIbIvRqrDUCFdKQIUkl+35gugCIgnZviuH6yolcO6o+HcL2
M0Xr0FfREPB1gvpyBbqL/UQYfBphzO9ZCennWrrZPlgtSVJvOYAlSfe7lr46EksGWylOFbvnKBOh
E7BBqcc6rAAdyoijSESaWkdTcqvxZ2YedZetqzL7AT/z8wZQoJ/TRObtqHohWXLH0x4jn8yYN4zD
LkSdgFsSZcDWHSk6FR93TlNCcAY0mjn2XIhplIKZPyo1hgR/V7y898sf+bSysqs0JILBEq0sp8sb
azjVRfGyxUBHNwf1j9mzRofVQ4S3TTtP3UO6N5PNjZxgQEpJcR1Iqgfb0x6GIHqIE0Ss9P6wgCvy
hr6w9ufM9KYhVc/6H1gyF15Kz04ULGfXjJmxkucrF0OAegdAAaJcukHq1cBeLccY5souVGiTpRV6
vyW1yJjXDJSExVL3P47IYNE3ihmpG6x3YE3XxaTvNi7Ubcirpa5UeiMl8LA+29NWMDNOOZjo/DvZ
zUccSskz8XJmkA7z9prCZIWfcLqc8/HXvMifdvGwULMNalcQyqVQBEYKJrMF8uB3N/36TUFK3HHx
PS8BH96x7qMDl+eGcEtq6JkXg6luY8fE31h3m2YfoA1pdHhfh9Qai42UVK0Ui8zqTqz8asVRwISW
0LY1ogGFqjKSLpaSYh9Xl1XrNPe1euzFVjHrW3bEdkInrigPZ0RoIej2mN7xuLdomj/EpB/h/T+L
+vI69wt3aNvBp+CwF4C/afgTao0EqQXME1+B+iS8zqJTTYLwI/QP10J0cOaLLWIHwMuR5dS4NepU
BjxcxEKfx5Q6s8xuj9vlKL8kdHIAklGWM0/c9XPbfTFpDmfENmM17acbPs6sy1sFCFs1RHNzAwOP
xBOYqNhI7B+Wc5eSB2GwPFjreKD0fdTJe1e0g9pq/Qa44ENOB2vO8JfhlAcCZ8jbdpCOtYvz4vrO
qHQOBx+7rBSHhXrdJfrLXiYMzaIvRax+BYgC0SH0LH4PKBUJt4MTWbE+owg1Q4fsLDFivxxq7ZzZ
f4nTKCUsX2x76Otbh9seznheaejr8oXGB8Lybntt9VqIYTF/N20kd30Q4IqrHQ8o80EY6bRShRao
t1WY2nCrqO9TomvBecCsAl4SFonYRCf/o19UBiVfYec1k/sNKRGLxoytZUbkNc8z3yZvXH63GS9Y
8yEkIHq6u/kr4HiAs7p4KUwwRVI6pwDxne1zHMNi59CAUzEkQa9sa7G+Fmem1aWLCqAj6lg7K14/
6z5nF3+KOziTvzYdp8fabg9tso+x6Hj7/qI/U/7kFC//fOEyHEPYmxyRrluDJKsxCtvWoa4y0X1P
PUDsPNLRzx2wrVvmNaUXcUUh6/Xtp8BdG6XwVuizNqKrd2B//dThGvXplgPIASxHWgohXkKzfBqw
dchrjr6jR9F8mdoXgj881ozsNuauNSsyk7Ba38hEMu8LFUTvktwRsIrJUDD6NmBTa+8CTNubrKiS
bxKAwFQYa5woI7VRbbDn3fwQOUBrG/X7+Jioz+HvgE4sDICHHOyOc860lyofKEd/XO16SfJkgiuv
dzwROv01FcC1LSEyQma2K6VVBXHcgsLU9h37AwQoFKpXjia/xD3ofTo7/3OUnAVGDf8ppjcqvTrJ
i9s8jgEX8wl1vA8gBAGX6EATaa9bafvLPA4AUCwj3L4RzdxnOkK2DQBmd0KbX3keqeUYDO6muwQc
PH6AO0ufb/YvhulFd3j5lQ1yxSTx/pS5SKeg0lQ1aCd+Uj8Eb0Pc9Be1fUCvuKxeZbyr3c6o87K5
4CwFj5hrVMMWDvEm68K2kRkl/Igv6MbfvCHtzPdz9LL+ZIlo+ZJn3VKYaX8X0/2xsAIMJVRMvZeI
+QvIpXSXitd8Y1EjwVvsL1w0HrX8BdppUJBONDtHGdH8LaXSGo9bseTTJnESjSliDwhTpiF1QLZc
pETz6aCqF8fHuwOhVUrU+8vL8tq4UnOfVLDBk47K0uYmZgVbZE7ebdlrwikuk3QZj6M0wakkc+oH
tUQg7ROxX9tRbMmk3qIYFqzCpmhlvPeV0NvoVfE8CnXyDxjDHoFZhxpfSk34I0nc0zPrIszgotN4
tB6yKHVejy/B7jlNe0GVIR3Vo9VWG1ubvq/z6uqZcVc0C2N6LBGCmBdBDmjooN2AMn5vIoYxYa5G
B0/oBUDAVKAQ8UvLBIFuGT33eq2QZxhkEviOArlnTE+eIqStv2jQrwoXJIu43evKnrd4MS5GDovU
MMLdxj1ORxxorT1n+IWXkDo5fCHtiyuY2ZlbxFJJnVuIQw43diDlGWqI0vHHNxDGcizy21YQUlaD
dDZKHDz2thGE11FehkUiEoh8kXEIblW20SLSOIMMpXE1yT5ydtzVa1dQClo95/IIrwARwoHjiDks
ViawZqh98Q5LR1gLlxorhBC46QdsJf67gkx4dubGHftdTCSmpRB1uM0On4Ihvho/D8jL9UJEuuIG
p/AfPCNXM8gUmQJNWmaaLmRWwW4S4prfTrnUcuqCmr6S7kUnaRkzLOhAXG4+0ov+4zvH7Y0gMeUI
Z1CpOXfHliXI3ng0CK4gQLwrtNblVan4klRCuYGNrH8sl0NcM6/VH/qzFiCSM9Vd1C5sRrXioKaq
M97TjeE9CchXaaLaI2S3yB4R7DjBLSwsnZwmJ915SyG9LatCaaxBn0QUzce6dCBkLlYgf2CXIprH
JFtW7rUznMgmZ2tbbnT+jSqCdXdyzjS9uICGhk4gPECDMnwGQ6+a1kxZoN6zV3zkS/hqJNBJChWD
MsnxbVMMFLh1g47JIP4AsECBG99fFhr523LzdVhFEI5jwXRcsytF+nGdaeocgZimV5jGeTA+DFtG
HjJucWq+P8JXcaPHmHuGY4yuVDkpXARXWJQ54rINEebP3zXvoq/KxKpmR2f81aP9VSvQjR+2MvrU
h+Tr8Y+rL0sM2qGWqVoBwlYwjV4SHfBvv+t3ogk6uP5XGrIfnHADjq8vocPowaux1d+e7HLFvtOv
pIo88Sv7xAEVLt7Tdf1I8VJSdLQMsYAJ8lxI4V0UUdMd9hFCyxItmXpY65q99kJmR6VjXACJMFjt
QfsGLT7Cq8vRyZNXGN0tTmJzqcBGJu82zx3BxKuxjO+8+BUWZnxOY/bVvvL0SW/pu9DulOXgbj45
VTKeTm0nXu/jFmQrnarXeI5KoZyZTBkFh17KA3dU6dgoiIz1FFI5FkRKJMKEZvkO9BwVTe7tnG8G
6UA00t3NvCuRJI5nRDASBeLbAbXjpbAbEw96HAmFYD8kilKUS7dkpMzRyr0de+fUB1jgmKao0I3j
MFVXj5KxicJC9dIP9vmbCAHwiMbyt3MmzxMfdd8r3gm/SgV8wipx5kD6VOfstKb1n/g1Mcts0EIp
ZiEzhoLFpLDTxbcFwOzIsHkhW3hTCtwWjHJ7xMNda1MenrGSBQe5ChWDmELoH7HZbWjwVE8PcSg0
VVYDCei1gzCvQw/2UGo3Cs2DVpXS3WVcJf1kzKhP55FCSXHLvBUK7/Tje+CXkz1r0rUjsgEEJysl
V8O4Qbfp4xySjx/X9U52P/pJX15bmu9AI/gFNFeE56dXMYOJWxEMMUVMrNzKdWVQ5vEHwj4+sT1X
1Kne/OS85w9l587OFPQ3bFexVZswi4qWfqasjeVFbfQCaF77pFVCCGJACNxUFJuAxTPsqEM3JCI3
/uSo0A4wod9Vu+GL1X8gBt8+jlp3hO0nRKp5KkNflQAvTuWJKaZqFkFjmdNzCs5hoeZU3fSYodYt
ghc5Wvu9jNxopyhLbwhRjCkTruIpKe4v9rIVDLQM2Lz4ds6FKFR8XC5lvul4X7jNVCyppQuY1CCU
WAA3LEkIzhA8fAp3Z4iGX9uHT8+QLw5fRw+yrC6frfmalGP0kpJM7LmMKN/YHz1qLaXYdPEQ6UaK
bKcXLVAD5qOJrSbl8R3eQ2MfH1Zf6UU8a4FsAAftU3WmMMLpQeLoDztmd/1ODa/qP/E92t2LMc58
DKQh681w3AR7Z3B53pcl0wV4/je51gOxtA4J8RWTdQaRHvGnNzLMn9Spe1CDQPeQQ6ES0hmrCEmc
B5OwPest8gMRYFnXLj1zTmFqqz4w6zclDHEgywyEPReURYLuDlVK40xWCWqQP4y0VJFiT2/gHbP1
WXABv6BE9KbWGtyOq9fFipVccpp2Kb/BliSmTneKTS898cIRLAPn/xUVjABjhakoHMH34rDz1YNE
NYjink33xhtuMDaGVq3Gx6QSgbWmP8FnYkwzEA9ih8GvH8Q4YhYG9V02tdT7EgSkzXLPgZlLwrOy
i74Od5P54H469m0Q6UvQhwtTin/lmA+X74BomjAQOtlNM8CgtIUY4JmU2Z4yjZ8qS293FUS1RFaR
hfe4uQqT9qrTGo7pxMm0rr1hTQGpUuERvL00Sl33YPnR9hqmIrvrmJwBNwnnQfaV6PBUYyLcOjRz
/KL5+sEpbI+la0GR0ooXwmfpslF8Hp8cAa3nY+o+rMYouk5N7a33lA3h6anjb75JxvP9TxpzFR3D
hDUGun1p4jM0BYWGbYvw8jbvDYIHkrAi2V0lqpA+x2QqolkyhxVi3CnHMOWB8Vau/LtVf5lH4JA9
QvX2pked0itbZeYQ+OlVDNMlvp3tfhWXa8XfOrobdaiLsUHmBipPp1LzcuqtU2zAmG1n59Nr/+XO
aue4KlIsDbopte2I4iIi87zCT8oRXKMvhLVr4l64Fd9fX8jnuZ4KCJz01RD1iqJmPcKh7stUy5Ho
IlhULiRmB7ONduOd988EtUqvvmwYvjgmG+w8TaeHFT+UqCgyP/Eed4g6zlabvTKhCxvCBK1ymu1g
xlPyCKgJuQBKBUx/eS4NBt5BNB9joYTgkRwfGFp0PoLSoV8dOtSpFH1rOzn363Jo5kI8n+DNok3C
RXUERNI0wyuHuuEi36jQeryBwQu+WDsmctx7uqAYxelNJSoj4CcIAgKsLZjzqKsGftIGqkSaxQ33
VONetDZyfMBB2MgeNmcE2ffUn0V7tovWCSFh34scxMOzjxpLOvoRuzGgA597t00unzV9yA7wgv6P
NJUtWeA7LQtdT9anMVHLTqEhLZMkG+/F9i73/gyxe1lvYDohu/rvLcAgdjhXavD82ml9IM6AXw8r
KPosTdyVuUH6YPxszvwbOiecDiFyjouGURPGyiogSrIYXPUZBeIzFiu09Fh6o2q8GCl2kxOHmoSd
c6MrkPeOr1rJbg616E0EQsTYNES/XYNeon3Frv9qo7n6B6iGcVn01Y/q4DKKJ1oq9Ufh4y5eTf8U
OgTEwIrOZ4WfBuYKfU6I//a82sM0ACXtClLWmhOxEO61QlQnzY2D2hrQ38fJ8N6WHi9g0njY7+Po
ReOZgMoPkHgy9+Nk+mHgatIAqS1snPW90kzZyyiV5ARff2uCBUsVMVPA5oWAuaxp19uQLGWxB88f
IA4DTeT5z0FAeTnqq2ol3E50i47TgZAURM6T6oyHA7QtCF5CjDuwxAiw5wjDETovgF8W19r0Mtf7
mPk5tECJDjgOCtV27Pnic3TxHSgQzofLgGCDMCqUgdJxSz1JlEQvprmvAfzNXvN6cMHzp4KzjzBG
vPLjKtQoPFz+pfr1HsZY7UJQFMIyY0HKovP+NmT4dBwW9uY2Vz7JZPbIFxcydWqVIE3YuniQrRNh
L1t6ltiiHkQXLj8UpHLA7FfSWxReIxqC4kP8HlCFIvNA2weUYwCq/Qhlt8yLPTXIMsI/InFcS2gv
p5Bvu5MgoT04uz9m9d8aDC4CIgM5Xs1r+/7UC7/tSE/zO5T+grevkr4ISdNL/9Wz5z4KeNUxIIHd
/Dgqz4xdZz+xR5U8bdH07jPwRPYFIEK25EMFbuBcnW2kcUWQdfExPiL2UKvIBNWwGlxZdzpsylgo
jSRFRLD3AvdN2nrGYxssSJzY0NDMbRyBFLRVkDaDvzku5s8MoIU+ZrHWO+4+ANavk/Agp/nYyh9e
AeHPaRhDscpRruPiEEQlsaTho26VZwlvFETU82siArGc5T3RmSDDGIzDWAxwLs1JjRAWNHwVXfv/
510g+RlF50LDq/MKehgxLu91q1fk4HWe0FTkBi9t7YRzMeKHNp26okY4OeA2TDZwMCOXsJz529h1
hnWH/n6VlzeS7CVjWgddV/ECerEfZS+8FKP6l+LAPQV4urhmh4Cx3/8XjO072qIw5nWuio9jahDT
7YKLNvV3UZdSFUQle/MAX8U84un04+JGlu3WcifBQSg6zLnKaxTAwGeZLP2+lM0PBrSknHhKGpEE
D0aTUgVfBn9Cj7PyiVddTF8vv4xuJb+23/Tm4UZQA3npdS3Fh2wrg368MQCea55LW4866QVkBJ44
B61EPD5cAXcPq/ciIyu+thGR/kHXcq2nnGEV7HOZ7f3taUfRYHeYMDOaoWh5mvP8wJK7tN59uBio
qvwq3+/1yt5AiC7utCKXHg9wT1FhWK08RD34lrSt/UIHZnP+6OyXU2NSxX8PDBBkoc31Ar2E2s8r
j5Y/JoE8RzTdmw0mlRjnOyRsUYGCjs4x36aVwd7sx9A3OBcqNHqFLoj2XMttYOE80Cop/LEL0Yaj
/EB0QChzJMkGYVsRxv5Ri1uopEdG/HzdbpXq1D5605fc5EMLXqiXTORzL1IZHJ1KDwPcqBZv+5fO
sfQ7YD+lRE/m89GTHH7QfCDnF7E4v2hrfCb93KaBIRSwoQit63ovV8fg1o4/6A7tNBwHsPI1QIXU
WSe2wxxgRqzsJmDMfhZXaRGLiHNlaDf4rfTvXXxJijfpFm3q4zcJUqGG4RwkKvPCwu3Q8rXFGDQT
qfOAyic+4w0QMLPTNiW3yl+OLn28P58nGUh8iarmzewl61PW7gKtTb9lC2C9s+EeIKx4A3twSt5k
uKaVz6f06xfX0qMrrkU9ocF3OCk2YXqJzNyCkUBtLlJEM26RJsT8Q2+Apab4G3x3DT7FrZeWGTUw
WFRMWdk80tlEMgoZPmjP7uR2Eq7R5p1q8LJ0rKhNnWs8EtdyxFvb/VnyqofLUPGjLrRNurrWLrnU
H1cnh+CvgIJms0ykepfiSwj4GEN6Bpj9kDLN7h/8de8OhUgIbXmGjS3p2PMt97/SSBLqO5CnlAaL
2AfzOlmu03ubdAsqQAwPFCYRXTXdtyLewsvsbJu69E4MZWn8H6w008SxTVdL4PfxYPhW105ZXM0+
mY1XMEAw1mD1nrEIvPcUaqrKGw/j9FuzUju3X3hEUOoTFyQ84GLSTQ6wyY7EaPIRoDNsu68MoDej
CHhC9wOkCnxK7eICuV9akH/Yxgvl1PiV3jqOBw2mbGW5E47bW226aJAjCvIajjvILCgTaAXyGAP9
F1zUXjfrM/RMHbLAzoGSq9cwxhNGYpdxlpxkRTpbqEI+H9aGfqP0NxHiL0eX0DZiDNT8rYRV6/e0
5lgerBGRzIylKAvJEiuQvB9hmY+W3e7ABwueRKHhbqD+RbMqUc6Fv1E3C1M9k1gKzkXcqGo9XOCa
CAuEh36vVQFQT4N7LNxV8831H8dZsm9/XceHYJorEOo+h0Q1NgjQV9rzoKN4c7UViZghWK2EklBi
f14XKsI8NGpCVmQUdXyDkCOJmBtxCabS+/hTmbX0ORVD/HdFovHUm+dQVRv5yiNB00kixMCxZfku
JlHY7iVWXgQ3WgqrDJ31xVTsqIrK86uKnYUSvNgc0baTB4HEIVmupFluCbr1K7jM3BgpspBWC2Lj
qmSo7fp15qsgk06ECCZByl62pbnVOKAFcRaOHw3LRDU/aGpizXrKlAjn/s5Jfx6yHhMkT3esMr4I
5zGRRHquCpfO/rGkX89Zcyt0ooEi0tFeHsQPLH5fSfN6Bu2nU14399RCXopPqj48uYk5No5J34mf
RpphuwM6suYhugnPWNS3edDnLpGeH/BtoHv2A50/jTpc63AfydrT/jHznVA5Svxjf2dPcYMn6phG
fFfDQFn012VYC8U8FbvramgJ+TRczuslyFG5WYYEIei15f0dgY+xCURieS/trFcYR10HJxk47rD4
q9QTuks25MnF4jXckx/9cLiSUU0vakam0DX7u6AMX02RJpWt+FS+JDxHaqX/kHAec6GczXmDAyAs
Lm5232YKxlQ8ghEkRI1PCaO2YdVuF2mkpz11cp6y+D++lvRgV0mDWYitHRUcJF44QeWJaFqDcCOi
1OT6TWpXhbYS7AfzIY/8RdtbjfZO4G9YMMVXAKAUZnVTue30QjajAo4J7RtA5DBo7WueYv2e60QH
6Gx2BTiSaDQ1t7Ry96Yrc17xWGEE+YKkGf2304PHrKlKw88DhVZXuEz6CfnZoO2iZy2UoOxVYpCj
7+Hfb9MzbBBCm0ID/aYAa0UK8UT7R9dvILiVhah4TdOKSrPHaC949SiHehMmHh2KjaWjRmkcCe6U
5PYI3zCKKzKcEzDssXjkk4JMweu1EQG1kvDdUN8cw7tlPtrVbCXPyB9hnAUdePrK2hBbk4uayeo5
UB1jj/2nB4b5qNJQN8lOKzurpieKJwro79dY19PB06ZV5Xg5ZizL/TphoImWj/b2kHi+QGSsQoJ6
lW8+oSB9OGRP1gufoHHXOfg78zHjtAJ3nUub92tDZucmoYTf/iJR5OGADr94nsqOQirLvE1UlEd1
K2U4kjMQipXFBmC5g2rKMmfNUy5IX6dc+OqaskXUZtdCbstZvC/8vmJBXBtyBT+c+Bwg/tam3sOe
wgx38YQgwRCeXh7cs10H6h7MleVBda8ajm+QW5faJAs3fSS6YjGjL8DFG7iCq509Z6kwZeVbIPig
UWxm+021EjsO1aIhf0LauC656RmW52Leq8EECA5icLhSh+iC2ecfxu+HbtiRrKub5CPRanWXSM7W
SEv0bfuEPTkFi91SxjZIxc7ybx0LOvMNg5SJRCJEDvHotZ+tnd0OkWVs39lJ75PIlgOsQsKMPE7T
Ko+heNJrlLd10drkj+X1CzdZ3eZ/ygT/7MrXLRxLZr8466rzNYMAnRLptIrJObbyedjBDjtNd+Yr
D04VAsDRtNCB67A+en3ToFjUlxfeo+C0tz9NMJe63b9oWtD91sxYGVDW4FRD7vmLtLYzBvhnoKZt
iI0ZHRk+CSGsmugdBUn0jeTP5B5eAeejks0slgScbs602WyzCFdngWFvuH/CfD7ZWrT5VZcWCLKX
8o8OuIq7Rzrd51Jur4/C7C1tcXt/dA19v0Z/4K341YJnTtToBirF9opkQG1N4qgiR2DGMwurRijn
NVDzKiMTO2eLOu8VW6FG3iVGB29aXNYR4caZAyiwBYj56pbshpJ4CTMtuXra6UrNESn7GbYwLqay
Hzh88TN7eus9eJDiQ+/4Xp1ZZEz33ziwBID2DFCv4Ry5A+KjRDCPlFP/HgjNY2w+bww9JUYBr/ap
Z0VoHyPzMom6MlLyi/u2cmfQ8iqFijMHPfS63yV2gdwbTy/Be4rYusxjHLe9oat/UgIaFcCIDpfQ
qlhdFFQ8+6fO7KeLOXhmAdpkN84eQMAkBBHSbsdVpxAbk1IYFEfcHnHE1pj9GRH8jlRT5KVQtCjX
OLoVD1Iwf7YwP0iMlRHp4URuz5z1XXNQOVN21V7+hcgfqz3c4pc3RGuNiLQZB6SnkJYbcjdiCYHJ
bQGzr3kig0yqb5jPo01cVBPpnr4/5Wd4bl8glktxzWiYMpt3LYO+ZD2syeHFjn2PbknVaYqnl3ye
yzFhdhTNnpi/pOX2RxC2CUa1fAuj3GKjRLS2tl8DCh2pXVxNZerz8jfII78CtWrqf1d7//sYsMAK
p+8NXS1WFvHkV5InGQR5aWVricKSpPZavKUqC2VUyOY1kJqUFY1PQeOWhBYxYMUELVf/QZnUo4D+
3o23ou2Jm9Zd9uvBq79Zn48du4BNhmEqeAhlC+C0e5ALWhzaHNqtCBGJZ2F+dyHbzRBI+aNKIQv5
SHRYttitRD/XkxlicSkbyoxEhArfBWn080XqPH0D9bHG1CdZeBn7SMcDPdZs7J3Ps8EGkf/hOIZ6
9yLV1DOjUuXdGQ0B1Zshux+LZmfdCh9ouw8xiYjhtx+AU6OMDDtvRL5hKPHYF0dPYoZRjOABMLB2
S7FtkZFegoQU7GJCNOD9eMz0E2xppZq6cWvLjfkLsHm/FT6zpWhqO7hxlEXSEfN0R7JOOYNP7VL8
s2WSquwbK4Ne4Wc4WAwnxh6KjdtQOS9+IV13xC2k/FoQZ/7aEvqNAqwC43s81UUmzXRrPS/AnJPW
fuAHkIoSpxXiBy/7PqIou/zBZJgl2lnGNew/hUr6KXiRRlKTuq5+8Pv8GlNaeHzNJYdVQe9c67lL
amfzb9LuGFBQVKw8AI24k2Yxtsg6V99kzDbMhSzCOIDcUVBMMZatnqXIwtpJK9ZnpurW9YomtPGO
BhHx4S1DLkp1Vd2i8u4ZZoTkyO0yZbB5G3MhuYRhlK9Z+gcxfxNQpLxOc9ECNg/vcepauSV4fxaf
i8YaPM72ZxbhiPhJwFNQrVMOFRju005YJpYv9kSCDM0qM6Z5bm68G19bkj7ObYzpojVZ6SWPQNps
nJ/tmcfioffCjx2Lo6cu/9T2Pa32sHGXoDFF+S9kk6uTksOuPXcfEbcGL5UVR/Z4EG29PiS3n2hw
hpm83GkWATA5+q5ZxYSKfQZV9ykZ460MHviFoQNXFHhYhVnrgxqhwxzFDVsqZx8vtp4A0ecK7Y8T
kGi7o3OKT6SkBqxG0tv2qAsoL1HlkGFaRqvTYhGQvJtDuRKwt/1VgtaClhjA/3CuN57T/Lrxpd40
lIcZcmLu0oRolF+dd3M3SYPYQOa9HWAmwS4IA32oFkzsMejjxr575qAucA139aedXlA+PRl3ZiDg
XPgkcik/9WbgyABGLt6xnBRUprrjHn+eMOYJwNulz9kBaxLw7UfAPuYGW6pbmnP6wZTzoLd+WaWm
Dcg4SIvOrDsBZlrmkRw4rGY6oEQe8PlGPAg6BbmZ9BQIDEVH1DtQYQFx3lcIVAFG4iREw92cJi29
sbVWGRpKQ6yhYsWipJPGYnKegooyKH8a4KagE8LhewZ5yzNHf6g+rIllua6EupAtLns9z47qNhDw
NmAWX82Hmg2nS6vXpa01R/U5j3jDQC/goI2TVwB1I0h+6zEfCeQGsmk+9MYV5MGQHEEkEVLKJROu
bVqMPpKrfZQ5C8Dbji+PXLp76Uwo4HtKseER01EmpIAwiPBMshUzwyQuTeoaEuQ+4LGJzVqqjsS/
ObRrRjL78pMpAMT6crvFQFd6cpLTTF9iqfivuT1F4wBiHyEVNPnquQff9PEPZFmiWoFVjhAYf/Pu
tU41DbJfbPlLrNAzdu2lzkn65pZlh6Kw5OQuyc4E3EpwZp+KjbQouBq410dbAjpaPOj3AFl9ZqWd
qjbE3TkzA/0A8QPXdZ/VIxhbD9lyy2tim4SMA1KkjwmW8+ZlEvnlBw5NFV3r7tLoSIZyx63xXovr
cbKI9IcUBInuWrrHZgDvOnIUM9q407zpA19EHjOrdCgrNFKFltfJZtb4V5ltiSsDF8AwzBcCVeht
2kGBnqP5Qp8rqv0Pk6b9PNRrTh8whNliPyHoeggiLdCReNqYR/zHX7gnS/ivqS/uqPz1ai9nn/lN
aiSXN1TDDTctDCXAIgVXBBTO3iNRx7B1djYpm+z/5xG4b5WrEhwssFzHPC4LbiuTE8YGf85L29+d
KVuFV6WT8tDNJtedqJhQ8u1VJZd0PPfSQLgcUUgN3RNcAOHSFqZTgxugvtP4n35NUjQpVQehWB2R
tmye4heN4N0KBbrfT9r9850u57o/dpGFKSYcg3pzVIMxtRbem74newKPYcgEk6Xb5O8GCu81KXRw
RK94yWaPNApHk/vsgEjypkXH8InfNKp3YcQ3N7WobzirpK3qqtqzh9R6TjKxo/KMp4lLeHiKAU5q
IzaJx2nG+fczDmBuFcj1n83WyDmlr75oZKgJuDlTbX8Az7qe16CrAu+QUPwNEWO/1Ehcx3W9Ayts
pvVM40BypwLg+6TeW5AB6rg8wizeVvBFuRKMRXpMRXxHMtYYKzKENdl0UJgvoD8JBpA/tUnae38+
ouisimSMe7tFqfM0QG577cIr/8EueNXNWLhBLxAQiUvnLmxVXuRJMwNSI8lxnhBfpC9DrnkC1i8J
ZBk9CcjR6ucdOUZUIlqlqmmySJFDmu8kuXWtqZUb6fd7HOmXmr6gRkjvSOtMTmCtXXRDIkO+Uawh
v7THskySx8lt6yUAjYUVv0IGH4KxkzMOz0Z1zrHyS/Tc8rjBRtYRfl0fRMg9JKWf8zsTvMpROWjG
ZvxRgG6KTiRYZAqBvvspvGntBTcL0xAwhTZiCD2nqUw86GOwjstRCfP3wc0YkRzhBM2FkCedzBgL
J0QRn/VtqRvKVtD1rOO9I0d7wgYez4ReWpozgmSNP2FvLNzqHNQ3tfGFSGWxFd+ClHttk9x3Ee3s
0zZxnCJzsAmQv0buHO9zmBBJ9mNLcgzlSjucKaFwzbSxgv/Ej3d/JwAjlINpNRHnvQjHd3NfaG7z
7RQDZEV3CEPOkYoIBqPiWHzOrFF46uMz3uqvKuO/ndMC2f0gWaRJOEQmqRbbDhtYXopk+raPAw3s
Lg0dPMowrnyiKhloqzpHmMvQasAzUEQDjyQFKzQjotlULhjiz8fC2Q2sbe7DwgIxfqSm/KgYC9Al
SF5/mYDnvcs/SdXf7S9asCtd59A4fvb4ykq5RX6m4pScyX2X6Z8grG7Um6eYrAzX/HlLz1zqRV7r
WBLV2lq1VGFh+POTvZU7/32vDC4OwVNGSGIha5O+DeKQCSh+u9Z/bQo2TpLMLv9R+nI7lz6Xou0r
2Xno2aS6ccFviFBkGgFL7znIG1ggO7NIFV8F7w423Q9QHLgEarxQ+FyGIHrlZZtfN9rXrViwsV74
rooF7YjLbIHZO7EyZqOFcIGci1LR+fr66mx0m44LlBJ5KwoGohvE5WVRv3+weMVX4zvdJa7CeuPb
1l7IBd4LDxN7rT7lXJCqPXK8XoCiZlEtXQ8V9p+eKr/OzHO945+7JshuR01fp2eK7/goIaEmTe8B
2oLQnQtzJuP/rSaZtA470bNq7l2Y3KhUZ8oCe1tDPBExtm2eW+wBPuaG8j0IfofrvtHRFXxoyvPn
CPbT+Rc9LIFTCxFczvZLaEdJ3kTRVyvepbl7tOSKByvuRt+NreEgmZoEQJMeV+YNJ4CJbd7g4LNs
Mq+GK9WD0hUFwr+lEg1ogbQkrlr9MpMj3n9ZkEae9h/BkyNtX4NFD09VY6Wb2eIODMonNkslYFo5
BtcozrRq/EGlwCJsf+DkrsuP9a079zormgTtr0nDI0QnsU2BivHDOAhJoaQBI4IJZD8TpBCZ0iRo
0kqGRjuFTrq56RJMxFFE4W0c47wHlIgOtjeTZiWvipoYNqOi7/enYJHtLsWYPjU27ORbhg5fbYnl
PLB3vym2FPkomcnCBdIbx2JJMecm/oXDrf7UG4jf/lMKqRb0wu6xW5vAwfXhCCNtPqM9lVnZEpAZ
zf8BCjt8y8F04TWOjxYxIWTl1u1x4NtJYI+vekJ+KAzAW1s4dWd/iUjXXPBjsmbUoioKjnaWBhBu
lHjd2vPfNha797Bxcrc7qZf7rCKBKMW5BTIUTO48Gc1Oe8FQvQ5uA4Sx88YBi83QqQkN0HaGlLPm
E0ZqPz1EvwvdGS+Bs7ZHCuiIM2fJz2dhA7tjXzEvArznI2U5AFGYUsgoNc9qG4OD+XRB8mn7u3AO
luDlyeBtmvNnyaeIaMo6gcGxcfAFZnN3weOyruaLgJbNbKcZ96f8zKz6HTJw8F7Upt2VpF899ULL
DJINfp5XF3PJ9dEivYBWioXsR6Iq/DvnzIibNdrCFaekINwVQwCtlKGYzdhV6HDMOl49U/vWPT/u
BeLhMODHXmVotdhdW0dGehO2iwmURKhRWiKPVu3QC51bKB4KP9t1NFIsNLYqCaV7wjbMloSm/LOa
la9jTx5AnPHevF8seek66ggwc2WBNxrf01Kta7/Rev5P9APEMiAi4GhW6fXpgq7goxIONsUEOCYd
SCETRkRm5KNYec1x+DVEcZJ5ZF/h1IlzXjrs23BU6iiV0gqCV3oVFDtJj0c9ZmXGQ3JrsOKLkvNi
vLkdVn4hYF1F4PM4ZVsLcxK04GZ8KCx7eJKm57D0YEAFz6Ml2SM4DYWKGXcBixIlMHf2A3oCH5Wl
W3UxSbXZnkV8bnpb9NUM5GVfx/RGoBeD7CtorWKX3s5fheBwC1dvVZBJk1lpsOrVtEtByAQLMA1r
+muDqwqs31eNvfVROgnMjUkp3Jjo94JkGn6xmqZc6GsVGAGPH/WCynM0kxUl84VxdtxUxEG3JczN
4PikXfDvlaswhP56tB/fMzVARDGRJbiMBhygQCw5E7MkEiDiSJcOkTyNebVr1NfrwZ/1Ac27rgLe
ajwLTIXFfGIySNHYAGX7XezE2tRpjSOtFpxRPqQTXJKQP5So3pE1jPSV6B5PRsDkonN2UJwr6cMj
woL+9wgCAwUXnsybfkOO3MAkhhppAI6wOpXKKhG7HePgA2TNRq5lrdMFpRLC66jNLC5QU8rshCVO
OFQr30Pg29xTn08lJY6rXmlaSmr4lM2btIMqWRyh6vjJqfw3qN/W1L/qltBfEYnaWi20qwjyfTy5
kU8NK6AqatHg7uRZPs0g8ulqQ7xKMa/RKUoStEwOFOj4lz52kiRSzcUFHIaLcP3jYq0QaTT2deOk
fXEx7nXRKfSsdnwPXJNw42tt8Du/B372Sby7wmM1Nez/D4vIzcbMk1jlM3VeI9RY80NN+q8iuKeH
CHArRrLVpBtHZG5lrRElEd8ZQoRZ00xpGTrWcrdyXG5G7F4LCgN6F875DPI5USZGVnpVg1S5DM/v
+s3h8kjDVCOq2Wb+tdarIdohPMcLmOe3h+FGig8SSzc/0kwi8o23H4QYYUzYCFWdICtPz44vA7Di
8DOmYTJ8HK1I5d9GDRzFCeJKIgRd/6xVp329t8Kqql18UnWQKWXHrkidkBeURDzZkCFr6v6bINPr
XNroX23msDzd2jRd8qq/TidjIraulkb1cslBCIHmxGC5u0UByzSt5X97li1ayzYnexbGdUYLtgd0
Z13ksC7kllUW2bITLWvfPKunRYCAyCy014LM2LR6MVJO8MTxraKplyJBC7/kjQnevz+3hP4AUgbw
XR+GUdm68GvxAYEi6+R90aIiGVa19ijhtIfmzb5C6kg9xOzjE99u5qhkvxvfdwJLGBqea33I0ij9
/8KNRwnqIvTS/ONGFP3Cdd0aBM5ixPnPVkbzPhUazKEJjd2KSgvBmqrbDCEmp4LPQ8EchEGLmyVH
Fe6GfqyoiDhpm/xpt7aPKq6kV6QQH76ToUrhw45WqO7I++rNOHoTXtyo7yivWDt39dcJA8U2WvDu
D3e+C2COQcGVTLkb+VI4/CgQWO3AuH7uK0myTc8EkpUuDDRHTFtitBkv3CcZp13D5+5spmpRV8bk
b6hnNbppSsX5+cd/8n0EOltgJeOdFQ8NEC7B8Q/L6uNXrnrSpd0J+BAG+cIF9aIOTu0S5BYKMWl6
eLfb0KCTFsLVUKaxMspWxn938NE92ynKz6AbQcKbCQOaN0+7wrbIS7Z7ggvbH1aW7oB6j8muHIE4
reYW+kJ1JVX5Dq82BZTKvyqSvGbi3tX1LisQbxdfnKAs1kQhC2N4d99zLl13agrQQ/w4sYG3nAai
+6YYccYTmhMO0HR9KNgpZPsS1KrSXNz7JGDrACz3z6fDfEbCozLRmDOgb3M47cX69xT6hSjocf4V
Qp5LFRGef7gQddN/0SM0u9N5clxgX/KkVC7wetLQekPy/WiONzJtrE4yn8EIHso8jWKFj4REVcD6
Q58pFHQbmHIwBKxGKbN7O/Y4CKKfIQIuT8PeAq/noFsUAaNN+4NsvoHqGx4wAcdN93XhAN88LmIR
5zwkzsEoXSZmNPRxg83LzLWQzlpP3xOMz67u2QMJKSSaNtpgcnuh2jPfdUzbiu/QTcMYNsIU4Y58
T3pKosQZx8RSpFozelAFSsStRzpNzY5r2YYcaEurkc0cOIXDd2gzJD7391kH1vuBLg+mJCT2bWm9
zKylEU9yIlDJZ9x80RJk5i8+o+Q1YeyisC54xf+b8GKwJOJ/s/PGVAP15nO5A538CadyH1KH9EHO
d+Pjqpgh7ThjfjQg3s8C3enIBeNIEn5gEJqcywVVW4JRpCFfk34A1K9IaOIAp7bbNjX0WE96sn7R
mC1vXqckofZoGPNkbB15t14u53LfFBdr7l5mpGBtIwztPw+RNi7Y9m0wRpT3hsT45x/LlvvmX16l
ive49HDW4OuQ0/gsafBLldDkltzFRUGrYLB/RSYAQN3sCXX+OZPbI1vFcTx+OnNevLTWtxWipBxf
32iQEN8SzoFghyYgtR7+gunLR3tuRoQaNPTsH7cTdxwfyfRIu9Wv0WTsCjnN+Ymjk+eNsbsoLrvG
5JrF8Zacv/bFoN0JYpoAdJhMVlPPHOGk8xh88OKxvJi0SLp0uhfSInX5tcM20UwK1nKiddFKgOg4
q3XqXxiWDyt/WYSoEB5f3norTULjkOi08InyMYXkrjpzeUVGpvb1z6uxMmhvr65uAIyz7jihYjJA
mHolv4UvwNlrGNkDrmYk5nuYHKv0CMNRLd67h09JHLtquYr/2sNUnU8suI/yb/htOqnBtAGyPlkm
BpzOxaom7Hq65gfFbV3kkubYG8lXTkxvnYr4E62QRc7lEp/owfWd1ZiTFqBQ01+87ROSzPQtdOOp
YAREJCKwRyLpXGrthz+oYW2QjYU0K5+CWbV/UMX/Zrb6v2lpgAeEx0OhtJp0E9ryVxUF3fpRL1R4
sMJj607FSRWi9fwM6mg7+kSYKnTIsc5YK+8tYfYdUyAXeSvBuGvkYvAw2OOTqrnt999P7KzPzD+D
XqJTbXRwnVJ49vTZxb2d0hwfGevdFGGCLeAJC935PAKkO/5ala7b2I8qDs71xaVAP3EXk4DntMnh
gqsVtLkZmelIush0yfRGyx7l7MGUFhQ4UJBgH2vIvNow9U3RYHWgdeBCzY4NXrzDU/8oPTKW5iaE
e6tzlXlSzt0P5o9Pv1dzM41W5D4eXDPavbHr7wyYRDPfcllRG1NoL4KGCySaswEvq/AUWj/if+/H
pYxJzTMV8PrDdsOwo2NQCw0+9TodOnOxXBDARqyXIekNjs8SeMb0+IibX7zB7y3qoCOQEUpSO9aM
OVFpogTV0R5izrmgqQ5XuP43yEjjL4jSEkINT59ZOlBwfaiOsluFuqV70fmoc1SstIzn4xYO/ITd
Df5LOvF9/RddqiDbOcLyahW2TrzeF6OfcfxPZIf/xbWM0Y7pxZyMjJ0TRpQDdTjor29HOIGzQu3E
8cL+8guqZWhfrt4w7D355EGB1jVf/SJGFRKIhZGtOSkrUjm8Xt1VvM8qyEu2GABnU6qjy+TV6gQc
4NlhP1HAcE6b5TqwHCnYYPxmxbuyATM2ztAoselh3hz34Jcz7LqQUeanOs+7Sx1G5ahUFHmuIRI3
OZDcPQI8N8LfFqg9JzSBMu50V27pUfIyC659MpTuulfwiw/N5myOYmpvRBHnaJMwhD7AGVquGOAd
daR6PPrvLDdgMWakldNHZ+c5f79Tim434iq2ihq52xhnhUeoEoQkJF59/0BfVN6Jpj32xS+qTNxV
o9dJn6ckzamKYHQNBDzYKfP7/JY0Jdk1CmZ0JHrJzJiVcP88FxnJm5BXL1I2IohVCcyYMRSQRYZv
2nIZkhmhYfudpZvp4ZKdmyXbReHR++wV0TbeXg8TOfztpp0sPXHRsRFhtFbiXznHi/PbYuKnpNjj
vE25NjW8z8c4VuuEk9/tuAlfyQwtYmTweS/99cuaagz7nj6zZRLBGI0uoLjRdw83UeugCk3Q1Fmv
8z0i1v4lfKVVUQdHIv1ocH42/fC0HY4m2FAMYNBqtKJcA7D/HP+qmkGnnOP2Q87KVwPXSnbHYUnL
S4isgMcZqm66LIi3hqwV7hrvvk2N7QRe0DJSwxCkF0yHbLgfu9DynUfeQ5SzGcSrwswwXubzbtZQ
DRj/X28POsbaVRJ1x7xNSVDPxkSGoLtvJS7ZsNxuHzwgBBh0aUmVMLUJBA6Q6vrh1gpFYfDYNTGM
7vuFByAEXGAsvlAmuKNhjEZIrKDdib564lJ2E8/h5JJXIAfosYHXzisHg2iBTWhG4bBfuFwGpfnS
aXdlFXblH2a4NpeVfWdxin5CK8f2Pbt/ZTJwY6qgd2yHfKhkG73KURd9fGmttaFHfFNfKrAGmivS
q5m7K1DoiMA/COvqnY/I75F5JqZIao+S8g+PIG8nEFhZ8UIx3l1Qpcpg74VPUu0glUJrI6tmn29L
YDzXXP3tC8oQMEfTNTHhiJPSJTppXQ2PU7Sn+bcORS5VPVOsx2GGAtSDqtvxEB0r/f11gZvnX4HA
F2uE25KSp9zSzYytzJCJbTFBq6eIeQ/a1vBZt8sB0nBsuaW4ENFHUiCmwU0PClWFVf+VoEj3BD8u
VTI3ZfCtjwRq6uDYR3Hr7ptCfNBcCCOa/grncQVyZfykZREHn0ymb0YuGThn8401ZHLRe14TDNIY
hngZlFlzZgN5jlUHk3x8KqI0ye1G6Je4wEAyytK1+o1MUz6RQb8Fcpc4+SiCjeF525cXoRlNdecB
MOKG5Wa3jMA1i2w48EcoEEuHwHLUuUePpg6A3BOkourp7qYaczxhSEwS8kuM36FeQD1QFDHKcJ95
RUm1AO6I08lt7STJiBotr4Z2sym579PSoKxIlZA6wkz3hef0ejfrQLCrtgoYjnChywc7hPUtRXD8
QFFIpGdmFDf8240WJZ2QjskcwkM/AwDucziGYLiJ/vnRHzE4AItc+9qV/WOKg54LANa2tP9MD9nm
x6XYsmUGR27BKwDR23zA5wLpgq0WdpaQ0G/O5TZJwWwshoJq641SXtmirbPmovjYn8NTN7kqaChW
OEu2t+Fog8A9gsBqteV03pX7mJPIcWacQFsr4Uir2ioMaf4DjOp9CLtR1xZ7qw9/PI2yd41I+IIW
/FXyZnPEGg03JRLyKvFDek+IlN4JEAgkypdycHVUBbQuDDKDHJd5nNVyUw9UCCQ2kJ49X6vxbwWF
KcbaotfSJDUL0mz7av9wmWVEppDrVLrrcZtwsqD8MHUHhgDE9Zt5VxoO0suL8jum3zh/1gz1J3pl
673oizi6xHY1ImIEs3I58A0JSr57baRXPJgEkajwD15Kk5Zd2D6+bv+2xev1ETQ+VKfITaq8Bzs/
Qw/5j45AG31rLkzPVh9nP7u9smKFso1IpJTbSmKcm4XY2ouI+34ZjQ/Y7onXQVuO6DzyXvypLDzw
c6GoafBnar1lRBKBZZnJBJnz/FnAKUQ0eiwu8JNMnYfC7SVjCPux+KYEeKPxL3XCVUXOAcMMcoMa
6uYv+vG1XPhITWVVXvyRunp6n4sZPXiUUM/Pab2Vz7oXwCxxb1K4xVCTGuLtvxBqMoSpgM0CZq39
ETOsRfq/53Jhbc4dQ+jJaNFxBFxdrJ1qQzjdyRNpn2DpxXpQsGm60d/ivU51DQRo/R1vN7g1yQE5
rGhBg/Je9DaoDlTyJbTESvo4OjqqWwEYjpMrs2MPPPNtJ3z/1+dF7vuZ22f28oEnIYmMdd+Nlx0/
zzjO2BYWqPdOcfkuWnxlHbc2t72B5Co7SSSfr5fIxxW43yzXxNQhQ9Ies9z6F7TPpY0+/Uet1cmk
RGIG6bD1/nKhl7V/V2uYM9yrsWAElQIOGrqph0sNCBuxecsRPxfrbepSyEWlv1XaNAc01d5+3xwP
FiHfltRzqzVCWfw/u6NRYorP4j8FF0AiOY0iBQVRzCzgiMtYo/5ikAdtkw4Fy/mcTAWg9cvb6WIc
TKwKJ23rVTxFyurWqbA5sji7/Yx8+b1Na2Jx0LNGNjn15wiowwBHtw2PYJGGQrq1g7vPCQBtL0/a
LHwiUk0vd6H/GgFeDxMhgJQafV2oxip2y/uR44yYfG6V7TCiIRfCDOr3R0mPNLhSRRPnXOiyfwJQ
0qmvhUiehtSCDpiBWq6rUYgRmr6FP+UlyxA+WG3ApD4esYnsIZrs3mi4hqKg7HEIr8pUrIyRfs4x
xZ8jxUrrf6prdRGXM5HWJrr23DeAQdriRGX0e7j1qWpR/5+n5/dilg04NqOaGCYYzFotS/Zbatc7
AxyntAOkoweO+yMaPsQLUuAG426bMwG5JHRAkDVBb2tfoEaZbsoeGW21+flszSvCEc91trnYz9DF
Cfxb/6u59No+dov4483JzcA/o3VqJo1i1MAeXPpcPr5c6CjhK9RBga1YzKcl0jgieFvpsXrCRQF9
UsZ0MdehMAtiQgYT9OMFNR53dHp7/rhS0NF+00F8crGM7MWAqCdkZuwX5WKu2bbkQtKFzdWS8iS0
kmLYO3UlIrJzQQI9+wKis+vQzngrRYclbBhE6wm61llXfTDC1aVJXP71tEdW4bjQ+8ttGZjOwP0S
LrwQwBJBPl0KmYQPkuqLAkiEwOCqjT7rAj1rLKHEr2aaUsOXnlcMwmM/rfXMIXIiTYeESk2vYOJe
5d0jXkyIhzyMvQ4fUSCkl9J5YNADFK1kXXkcpEJTEUWf8r2TEQ2KWIwzDBLxrdMstuR/OBv/gnbW
qrIxzvGj+VUoCttuX3txP4v/3bKucUixCbv3wVRC80INJBOIQVgeXDRk4FMbUDjX1vNeBEknuZ5z
6S9eR3CTb8z313ZRfa+jtWdVdE76qbNs3shO8LBbwi5rxCimOFqVn9BUiRhYCL4lSAMaXrEEShS0
my4Rp4QdNn1Aak/ZYCiSyc+U5JNQj/Ou+W8iqAQnma271s6w5W0iY+0mPYP1UEq3WlF/WvsV7FG+
MKaqMqThgIRwt2Y56Vm4ajYFZCBR7X5bVr846i+be4iECdcONXsqP7kaDSFQO9Sfytld9Z8LbqJe
DanH/kvCuEEC/4M2vm9WKiv7ReWXz5A0MAhfEDt/yREtUheQZbej8dWdW5Z96FAyrQK0znY+VhPD
Txfn9hriYpMF/AQI3YP0HcPWzPmyGq+rR+ANr6up0QcQ9oDXscfGf2DPZmFwUugV9EBx4Bm8Bxk+
p1idC+fc6VjjHrUi8n7VYwt8PutJP323BUA+v8EAhYLfU2RChQ7Vaw1S0Fuazn/nS6VbW6LBro1I
ODL7iwIxmR5KhfqL+FdEOnnkNCcEF5KiOneEu+b2a9oexboVCwTYuOQr2qK/qXJ++T3dQSsu8+fm
mtGk3gIFME1cUzp4T2Q6gj7cZRzH543MsDGxRKw/Zmgg7rqBnuDucDc+WXtgPS786o+gmA8WFKjv
lrxFm3nrOuB5ihM+5+vTT6qwLnfvuxdcrzRP2GGB85jcg3kihzwDNjI9ABwG/Ddef1S8khP5BwaY
nTjxfxISIUQ4VYQajMbcygbht1rCrTF1N48cH7j94KZ6/mZrdvg1mosj06LM1K0HynRv509peCfr
DMpSqUtlAndyuGHaNVW811OB8FYSKw2iDnhT25YuCzzlpJ+zslJq4RgbK7FX/QFEJUyh+g+MSjnW
FpnyzC981DLQdgrcXtn1Sh1Mq4mQDR0+bgUVpYDEep7S44Rcl+E6w+s2WqIUqh3RRU4+QHr6lyHe
lq/P9p5SNz/4pE5EuS+Zy/wqwCMIUX53dy5Mnpr/ZM/2QeiJl5vyTrcBwq1eDLNyiY3zGepCwP+d
vFxI0eBLTIPCxkAj4pzNJ2QJaEjaFXAtzodLloNFA3FaVrxFZ3Ov2fxgFsEezxl3FFqTsKipmrYb
N5kA8gGoBOHx2bpN76Qq2woBEiQgx1dAhiNiWnhAup4/DceMJgmOo76peshL7A0FfrUJKNHsdpg7
x3GQUG5h6HqKHOkQU1axAX3YzQEQoLM1coW6wRwVUfP3uNLfBpXntfVC3S/FgmIbFHawuBJ0mDfF
gJjZn6/+bmOfjHusmNieN3X4JAkJLDwR0hdhWweqMwCduwDK7fikwTd3jxDZDMrHd93XXpWrPgcM
nNYAXf6BCbGVujLivjOGtwK84lMu25VHbph8o/GCy73UhEtwU7HiBDrf9KlsmQapPjfOXIRQG/bC
wm8kZOTRzOlxqyVzzL/3GjMX/8XrtrvGa6DLpcsQWIJ5+hJams8qYrhOhJozO54LdleoCLN1GFE5
9KLUjwzKTzFF3RGr7sFopSn2izMcWrcsnBlnQ6K48ZNwW0Xhj5sBs3IpvrPCqVB0jGhTg14rA36T
SGjPJc6RmcKjPhSJh8v1odScp+LbHyw1WiBGXowh8V4m6VYgQg0h/QDTT/SCnEzuVeqM3mpWNSQw
iFmNa1qdYqpTR6LUZh0gBUs1kntPk8jt7hwkUFhQZ9AXezeazoZXAXCRxIGdaeFk8a0XGUzOoqLg
xUhOlYO1Ogj4h65NeYgCbUK4kMt1iP7HY0JghCtJNltIbY8lKMoADIPVzkgH1psPkvaK6SoJarbw
mfKAWtMUpD4nDWA2RiRpBEQjTgTpXzz8pk0siNVDvNFX+qDiudIGPNr10R0FYOrHIPrT0Yfkdzuq
0RwrXRQF0kHYX04PeXekFuMRWA6ENTrqQtCJMkpb7z8Ek2ZnMuC3aOumLEgnw5c9iWJmLID1/3fT
SPYhIisAkKznEaPKuoX/gfjr+JBirs2r56T+AoFoaFh24dprRJdyr+EupE+XjGN0HtENPU+KtWPt
JXBH1/wEA8PQnUXRDeA/5FsiSurglewRba3zJR7HPDULLVz6ZcKLS/KIuDpsDZQA8GvKJuPE9pEm
p1iHvnWPOr86rbPn2Yf/DkAsNR4RKr4Kz0UGNa6Pzl/QzZ6flBH4WmojwczIgocVZ4HENVJrINWy
gXhQzKDZNcCcGcoax38DVHguFxfMOfyw7qIqvBq+7yBp/jo+w49r4+x2ULWCLE7Te+EVdtHJBB5m
ym9pmfA+dw6qSGG+5zstw5hs9MYzDRHfJFeqkTADIEwk4AJG5Rl7WrVEpSfpfsWirjKAxXzuiOO9
hkZ1iLXBzjdhW1jEGnKI6JvyzU05dXoK+sDrYEcZT7mYRGvxeDmAAEMnJD8gj3Fk4h8iYo7sUvN7
9VndI5TqDjbm+su9WaUWf6eRlmB4Yv0XFjdTC3jffOroobRTgtPx3lLbVpQdoZeAlSMhRBzHqr8R
Me+n1OQAIfuWGrSxIa2CgIDRGC6sUEPVMZqkp5o3FLUtaX0MdsVhcZDj5cdDcZIj3KogUxRoGnaL
GATUAloF5K+8a/RdR51gw6nKEo+7peRBTgXXba9B9L3kMOBDb+sjbDA/5VgumPY2mrdZEWnoTcub
idmjm3M3bV41NlZZ8EbTH2UkXNK1HnXfBQsDE5vfFkmhERGaj/wO5yVliR4AvoamYm5FTjUfNh4x
hVkciYaRllFpsQtmXI6vgYCF254M6YtDNY9zNgf1mQI4HYkI0YcOLvnYMQJIw1rzs+0QKUc9Ex91
VUbDLhRc3ClrvofZFdIiY09sAcZLW4LAWgJpslsa/+0A5Mqu56dYYXTvbsITlE//VxvbokWLdwpO
r6pFFS62/JEchLk8TiQB3I9W6a3GMgCCtyrl2bsB0XuZvjNU00zngcMm6dU3VxAQiy+dGXEzx+xO
YG4tl7WAP3JYwV1s2l55pPXBk5QOOafxNGPlTPO0+89/eZOrpFkenOlpixLJ9D2SNIO2KPtsG+g1
YUGDTZ/FLpYpXCpxwBQhvuVvCVLtjiqhYiHG8SbZD48YBF9G2GF8HUhaYlJHXCGgRa3T/M4FLUZa
ZnxMXR19p4G/XArSg3ZvVN3siTK+jdkGqfuo4pthurq40KDkiU1S2mrJ8EtNIuUfSaxxaHnvUxZq
+zBGy+kTBO8LJWMnlpwit8mBDskDRKUiuMh1PV2K9Ea9c3KZTHkcS+IK+RHiBK2/gt/NSc9wGHWB
JfoptUneYxqWQcPaLbDsK9GgVi6t7EwgMxPd8xQwDMeLtNivTbBCyi88AjaY/vegLZ7iJGpDqNXk
yfTht+SMO+/onQ0eOKsGHU0QhaMbLPnj4fWHGHKZCY5cWnDD/GN9bh0ZerXz1YbFUxSk2siMwXXZ
uP+xLFKat/q3VL/86vV0bk5fLBoKxU7T4/+ZX6zSbUkW1veCBMV+36czuoBUAIYEQdNnaBLdGmL3
pzbQ7UD0j1EJF6KFmxeAmHCbxSYM1rbWMvvGHCH6e+tUqf+giQmA3coaB3Ho6F0bbRsib84UqJL5
IFoY8JOLr1m/f8aEV6EuCL/2u+TgJE/KbyjRgLIouBpfK8o/0C3hcmooBMrPpCYF4pE6DLxJM5qq
N8rjMNPoXE6Da3nPnklfSd7ihyophPqWHaLvgLcaN9PsMo2tT8308uoVZ6weaX8MnHkjY4YswtG1
LeVUAj38zYsNSe2DRsGWiWTcwDn4mbYkb8MudDQ2dTaufGzt60yn6qjsr7AoXJR7rcDtQEP2omLh
IDBrQbc/AG7TpVu0B5TSs7MeZ6+Zp+w3G//j9TB7+e1qGWybr152h3L0oirta2HUHNIX4W61SIdE
3jgdStN4zIEXAx1kfXUf03MaIkK5kZbbXuwiWcv8l/bzIwl7EHG/qKRcNWf1vqmj6l9f6UpjMjdj
qV9YT8jmla1VaNxdMJewLg3g9TZZHowCqJYz1Z/QPBdwYzi6El4UBhHjCsqGm7OF4H7CgEWKqHB2
TqOjeNCz76H1MsNX+ZyCRxj8xPYD5J4tA4z/Eac9ToFczzdex4iNQo0ET9PlHyLY1Lv6V5Fq0uLh
ZhYjNoZ9zrYoqgJs4zmIvXHF+5pUYCDzCKkb0qYastX3ououQ3R4Jbhb1ZZ1MK9a38Ii88Iqr/ra
SP9qeo0nCyiOG6iObpJVUEEi+qAFREgPBEnhARHyZpmphaDsC0T54InLmWDLDQUJcS8Zg9NxZPWr
qS1Z6dr69GOz1ZKqmgNUXt7FnUVx/MWqjjhyxbdimv+trhPC+QdCRDbp2JzAsJUs+a9PBDpTa5lo
xKP0KQOGd5CjXVRWYHXm6L5Cis62/3OqOVrrekMbxvqH54p4q4ba1UoAif4NUy+B4xA6tIjyFTZM
168C1soVdknTgIDQc/M24KDfosP8in+BshXp8Ee/0PUFknvM9TRrVIdFQKJBE2Zg+PT7UHGVFaqt
78g41qOwf/v6H9lebGi8VCqaRj0JV2t6a7FsJJBgDcFctg3CxPETygus5SrpY1hUG4ZiH13WTwOI
eTfslOALnhz7cBR9M23hy5br123gZ06vkx544ZH2MJ1DKygDVy/BM1KUQVB8dUzlJoieYXK3Qsxd
qvfrJKfnTcwf7myPEGoNaLWUCbRSqRZFKUTnqJ0IJ/rf1DSrJiihzgV1MIF6kYZgi8SXZ5mDkEUq
8BCY0aMXUnDEkSTrGNttuFSOmPoiD2uM/PvArM3ezn4SZ75s30TWXjrVbIj+GmYmulXY3utZwxJZ
911zB020uVtrOnQHmOb1HBfz9Tfja4jckXOS2vbD8+Gb6AF7GPVl6HUp99m1rMzelmZFH7jjga9u
SxNWHS3MQ2ZeB4brWH9bvAd1QimFVqW1dTiiDB/bFOT1XuDWTGIzhSkXM1pDd0qpq2I0oABPjZOy
Kf2iEdnVM48jf6nVsGCV0JuCrjfTSgGD3FxQ3vGUBRlVjhyC5lKfXR9tvyNQq+FVdG3VzsXKq0JN
138+dxEdB8yFAq2HbJ30dp4DO5XFhEfsZjexd9d6pUbgg3T8gmsikqIOLD+z8ZO4IyKoxbbBnhm5
ScGMoneTxvVUJ07MTeXrjaPeHoE+c++/Fdn0XKlV/oVPXMj3rFJbUxOhQDUjh9DuLxTp7Y88WPCV
Ywui6KuKWz2u0r/aLsSVXPUtlADAgqwZSYqnSrfSnXutOOeZCMJo6p8hTIYe+k19K2cmHnnBqlA3
tRa4T1PXQcmHOGdRzlFN4JSeko7VT0I8IltLYro/0tm2ZFSq8HcVVP4GsaQi2nur+sedqFXjNDsB
TwEybHgf160u2J8kTkmLWloECeUzFny4938GMMm1pso1GsrNEBI5OlGfqvRJNHwOsYYMwm5tujCw
piz63hSaTcxyXLI6uJVyPMHyE06n/q9Yi3BoLV7kIeyDTLBhfz4siY5lD9P+tyiAbsyYkvrx9/Mw
kykpSFp0sQv5LOkc57cPN6K6rKz5kTYyjyCEq1ncDMgQ6upkKmIDtp0CCCSSMMNpZV1qI5llTSbW
3882xlYp08/TxMdvZLYBFbUNPcrpSMUWOd00USkEbYkIz7EIgsi7JrDZx+udu6I2r2e0uQX8+ddb
jAyVdfEuyqizTaoyPAvYkWGQleKL1mDKvTlQ45JQYRdZi3uslO6s32+bu9kyzhrGT4WVzgIKfSTF
DQ+sfcA1mkW9ufBwfZWkxBQmYBZMTbgpa4wm4+i5Zh2AtYSzd7FCsPVy+hoFbLrmkoZK73Hc5O6b
hwQh9jA224W3DDne7xQ9ha58DsnHNcEPBaICJVdDXN2UvDpOH26QrwqiKIVj4NVffKIUVTRqi8Ci
wsT0dAR46h0MtS1YsMBqWqOWem5aw0xZM6icGSXvHXyLvyTNd1HoUJm2RM+6VMVXnpACn0qjYE0Q
QiOyarcnCeXU5wH6ktLGj0bQV8vrZvLetOD6jMgVmnOMXtsziyMiut0KbQ7l5HpxrozYW6INXRif
SXEvwg3MtuhQt3GwmDJDBOEZLHsK+bK18TOyzpAvpvupuMAm24DM2LaO/koTWy3W7L7NoPYxV8FZ
EVFyy2zf+AUcNJQudnXplP1ezLEebVo8hHa9Gl1xjRgznmqxBe/TtEhDdNuVl0hVTB25i+3g4Ka7
bALkrmKnQGXwOkAqOvUMwEjPMXLzJ2P64mDKXGTogt2sgP1OzGy3pB/xIrBkHRtsxyoX82+rCrtl
GrMvXpmBHJ16E46ay/TZA3M2EF/o++W11BNaJDOG/qDzni+QCzRxQypWo7d1kmok2cmax+ER7DNN
lcuF+/io5k+7qawlCQQkb8gEk48O2KRsJ5srEMKkJ4dJOsrj8yLMJsVitTciUmdeaIlEAX5Q3Y3h
XuTdI518+2oKFC+CYOxviHIONfA6j2ie9aWbCXGMr+dSZXUQldoDXHmLbppjBI2Yp5Gu/hrgvF8A
d8+WJ2RtxZQrSCvUAElrFY6CtHQdmNZd5iamg8r+GDDwWEZQ2w9srZ2Dq+zG4I8HG0TUyFC6khjf
oDxs5mrMlO6XYC8fydN+hbu7QJI4shNgXZVe36dr5uiU/QuddmtnnTt1VSdEKlBp6GXPtZpHp9es
XGPR7S7JXuhfbkwERnNoi0IEWUl7G+bzHDESFqjYK96N9/xXBSh9P+A4HLfoPG0tO2DyUeJY5AMf
58fv8zcqj0ztKDiweKyvrEuFR9cPfuleULwuGNcQyo2sD20ptRYKHIAi4m1CluRlQCaMvq9W0V1j
hD43Jq8ZWuewgNpS8nt19FDj7qa/4f1VcHJIX9f32WLIo4OoMEb62G3TtZEXMWlRgxCO8QDZ3jUl
I3iPq9+nY9o77DQLuEFSxTVcZPe0aPMmIghg4OoOt8wNIjpSh/mvm0uhj5HCbY0WThqrY9himNE4
2gZV/PHLBF+ut1IIqzquMmNWUSTDpTfQxz5QqElWNVLBt1opvWJJb/YahQN0K4qRudMXs7b0lLxX
/au+H3AyUdTpKsofeBGpwSKWn8JWHciGUoNr5rb2wEIlEYwpDHArmq9r1Omz6XA8mB4sd+BYdSHB
u02nZ5fU6JQBBLmeSaPTGSEyBTVpKdFagf7uG75/SwiY6ibLnF2UeFHtlJepAX3Tf7N6kddy7ALS
6ttbUFby2nOYr0dg/8l1ZV51hx89qtC4qLk+LJwmV2vqiUyaNi93iorRy3zD2TSf3V1+qTtX+J1o
0RTqa32wUT+LzAasAPUxz/LeF+cK63ZfLepkcpTQydMtv807XX44jQrqJazQFIHnr05kXU85Jdim
Ns5e7jpuPf4VWRUHMjDyBxePIhIKHCt3RZtaenRBtfskM8GjbK5nXoWFhgNR4wM5NVYzih8aiMTN
+NN3W5qNGiHMcqsnLaNZf9QHQVY8kYEsdx5ne/PSlhAtUUPcGQTJkH8NlzdN97oWzZxY7vB+CKLc
5exlDE+nhjjrkSCakN4Xw4dSfBcFysHjQZg7kHWn2N9hqTs0pMBEC2zmpXTEtY/KTc5qztAF5fGq
P7HvupkNC8MaAYNK0+jCrDbzGOpE0geq4xw4E+VO0ggwakMBqkr11GZ15yjwzBeCFG91/nRhAoHh
WCyiSlwnSa0JRAoWVb6BnBD4xjBt9j0tgAINRraiNkWjCrSa3C+FkiHNahZDfNWIZN05B/TVArzQ
bxfuH5e9EbgZz3yixPtidtcPrEvgubWCMzcXeh3kB0iPNox1kc19H08UyNE6AqW0bJoTg0X6v9v7
ZtlIFsEXdW8RJo0qWMS77O3RhongFxI3psfUxr3iCAz/ZgSQ9pHvhSyXpsfnVjTVFQ0PNYoLxJ0S
5PCWUKT0pLQGYpvEhFNLSBjsu4BtXhQ42QnrghbIl1ue4XPFaMgvrnp137b+d64eHU+0sR3SR9YK
SMoDA0oNTguRkbnePgA+2otDMRJqz/0SKUUhJfmVvInuD5x11EIeFHsSurN5hj8Jmg/DY0aMl5J8
uK8E4JkyslcSvFcowY+eAvS2VMpWLEw/9aH2zRmuo7bpAYwgH/XNCJe8Q92dLm/PFBG69JfwC/3e
8TUkEg1bT6xIakF0iIlOrdnvL/HrITkLVNB4bK6PU9tFrJ6D88ugQfq0OcNp3yEpdFTwUwx7Ziq1
4PErhgTVMQfah6Fran7cCSgdasldVeFYzxm66m8c0G3p45Ke80wOgNphBPZ7+60PFNMnxHw7TD6j
U0fPS50bkXOG9s3T+nqQe4gGjGqe967rrDasmaQ3tDrt8C1ep5/6/pUaimj/EiFdO9jacVHM3J0r
xOzFkbBEOLQ3NHTydWfiauy8i30rbHYQJxTNUX9RC6FYdYv5ejXXOvAyUHyEEkMNArQMv8g3mnji
J1oFW2D8oqeqseS9+ODFCOUvU4remVl+UoGFaboR7UKm6CfCcTLsQOWGNb1ezTJAV990INhGmiaF
ejzyf2b1CzM5FSK8q2HCbe53eT+5wQ87F7ZFKlB8LzwM5SS8JE4fQgghQ2wfxSf6so/BMENQ9W+y
BOulNj7hr1LBuBZDNhElICluu/I/5VjeP9JWmHPDbRZFt6qBrb/xgg4Dxdnxut7bhsGI94VS2nOI
nmDyM9TuXM4Az21cymLLtKgVoBVW6wfQ+BX07/Cyo0eb2XweeOeUNkwBpi9T+/ezxzOPTx1ljXIr
WtCrb+ExWqCVHTl1toACYy7IV7stCLpLwo8gCUytAm9JX1NwEDMSGipW5ljdtLe6rotHZaX5aq21
RF6IDkXqm0x4qN5jnnayebzCZPHTPUSBopKF77/nKPr8HGnLeJkGIiRQ3rN7va+TXWqh0puZrPj6
RyrHSKit/CX9HprPVZ6+fA3zmnv+vxZyptafPDogYCTzllmKm/zh9dAnv/dzDdPygE22pTmYu4R+
12JQWFlaSy+NBQtA6MwaAJIC5ZV2/nal2g/qlvs5konSwwHqu5NcXE4vvXhf8ZXwp8ht/zCQ3/iI
7NRp47g/IxVFPXrRCNJEkR5yfsjkWSpXlR22s0ZgRF7h8gF6uYkOyWLo8K4FO4fvTtpTWOdi7jrY
cTKiKfR+sRGGUsoh++C0tvOd/VtYv///DrLtrFYXk6J1gKXEe6l6TDHQSt11zgon2IDeCN2haCY/
5GxD0hEkaQVF5mv4SQWj4D4GOex1GiTI7q2aA1DjSRYlUp7iDyjs03ZuCA+5dkEZ/K1Gdi44qfAI
XWRl1U4XoFDZ6rq/lJU53h64WHsOTNFvMvzIFv1/nOKRMy+3UPKisk5pj1LVDICrVPyEsc3zNGUC
cswuldipgvFIL4mD0Omt8z7Ro3VDq6baCArh8PZLec5yn3Gkwl0NePOFz1/A2QCxbWCo9xc27Nts
BVhkwuaJ/9yezz/BnK2XSXOTqVjnYc7JCrVA4rpY5yFaqnKgKR2PIXmVjdCKY1vYHdFWakeAD2B8
8IVBWIOkv0RD1VbcgTAi40DxghZlrJzKLKmxe+OWiRQJn41HBQ5XNoUASPI2Ibny//U4fG2cWtau
jXJ7hYcCbwnCldNhG4xgyC+JTHrHNGkSNNt5hogyOix11lETZKr4s+DQgFpzyqIKtGedIw3pFKIe
F39I93TJyTz2xKYwt1xtqfzXtTwb9qyXX+W4wZeKewtbLbG2Wap3nFTQNubmXn7D4wZnkd8TTvj8
0kIXC/2OwAC2MUakB6AZONS7CM068yNCzgW4TclTobMA+sDL8XoObUUDndWW4bVR6G90JSryW6NK
FXmxhQwp6Z8GwmQ1M0e6otoDjMtCQNpZsGSoWXkAxjrv7jgi7P53YJO5jFU5dDJTYFUpiyva/dQw
jkZRxXn9JU8yt/AP8PDndjAHCfeivNEor47dfDcZBeiIYy57Uk1qnHx3vYCq+qQa3B9wb/f+Ojjl
IDtjWbwYuHFUH2FQWcP6Cz1zMnTPO9yH02fr6I/6RL6enIjnH8bc1jSqy+k8G3O8qzazOsFb9P31
KeAZGqU4uLsP+nGas7bMjm+au4qZ2wFI9dhFF3eFDztnbsxH8rG59Q5Tm49dzZEUhk4zH06phk7k
/p9pgFdXQ9kTDRbeXgBABgiGm4Par0edFyBwnY29F1+0S7oy9gorja9jhHLuBiWkCu7/s6i2wkIa
F9hgQlhSx9m0zPEChwG1WBtQ3Dt7l+5iaVS5R6MzwWj00BaIJ2oTnKrCNozH/SFnIVw67x+hJcv9
qHVn4ls1u6TsR7e/Wkq504sOXB+1L82XkNDWWObxRUpvWEd/618k5dryT5lqtXYEeKZIvyLgoy39
0AXJfR6h/DbLELkSPu5Yo0mfNIPoiy7raYNCkKPNHFkEMASNyF5QPTdjX4mj37PgcsZSzP4dTM0h
STW29ovkIXsCu237UHBztIUWS7gC3v8OMVYHkhnL1k7NKfjsrZ90nr/OcKY1U8yuSxG0iBT5OH6S
m8wYTaFgah6af2VmF7KzhE8Fh8GbJa5Y1fnGU0jq35R4qGHzVHioM+O4oVFGG8qxP8JJbiR/rTCr
C7CG4RMCs4GwNRjfkkEUfVWSBc6G5T+kz8Xrh9gnB6xylwT+Swx5nceRHaBwQYkHI/ZzpOYoNbhn
JXoEgoAHa4BEWK3kj0v6e9NBFcJ9pXypfnLhONyj9bw190Fb2IfhWrSRkg0Z5jpt4/CNMFxUhymp
9LOoh29qnCuyk+K6EMx8nhnWrjkdZrNJBzBgSW53lfwRun5cBxsetfPEKd8VnQIPM/r56TtWNjQ3
IbD4TzjTdlxvAJck1IpmL1pVTZaujrhMXqwJazQNJBUWEXUKdBlyLaEeooT2qE4HygHAYZyvV1Jz
fCCy5+0L51ynsvfBGy1NkRcvyuqKcliT7s0nwqOM43YSRti5xwjQfcmob2yRCALj4nh7zNHW4ojM
OShYSDZB+C0EpzuMxRmhg1JszZXM0HW2G8urX8tyiFtS3i7JUGI2nSVLU9Nd2vMgTcOAE1xKKdzy
6E16hLcHmWzJ3UGVvyMtj7nCwz3VTjVCJKTp93nePJx+EDt0QUj4hgUz2mv0hX2gPf4pDAHintHR
aduanv7VHwS1+pTnLg1IVmU0+l6hTUfaXi+KR6r9eI+bGV2Bn0vSNRRk0pii4Nd9aOsc0cqQ8Jz+
X443dQTyS54D4IjTI3Sd21mo1dtqXVhJo1H69Bzrl9rsWsx5zujRSQhWjU/R2T+GSipNCDwe2Im/
bTAeJ/5YDGzKlDPDC8XTVTcIwRHDDFsIBih0HCV8kAiickbMUeO2+5GsyUY1WWvKHhHyFfV6zA9v
sO/kXXrH/WrRS/OAc+uQbF7JqEfWe1chC60/bwwomqQ2JhUB43Cw0zlU9Cc6MyaBkpSv3lGrC0fU
TcuZsALa9urPZK4ouHxTkrOwNZAl/OchCTdWsv/QfMYUUOty0dAUAA67Zom+7h17iMXb4VXx3meu
Y1JihxTTJ6darXK26+memPWcDAL77whnwWav7SQTdrUzcede8VA1TJ7PLrzwjuIHhBI+m+PSJPUG
BA1L+9OOEOIONqAE2S6MrAAEMNyGoQJpG7G5kdB5pfjrTFKQroHaBaxHfWcK2AhDcZxE92QV84TR
KMHJymSRuT1yyk/ciTSMQDSvAomvU2YRzo21Hge1pQcP5eimoQR4wslYWKm1vPmrQbbLe8Rhm21q
IuV/c9zQ4JnjKGz1i68AuxKu3/nixs2z0FQPqMg91H3Hc+hLPzWlVL45jUrAX+LyXUqjfLWNFto1
4zVOfGGCR27XXn/qYeEUNN7kLshu/2t6Z91OILTJkLidNPZe57mXry/AEoORAhjL1/3tdyAtwGmj
DbISNO+csOEQoy9piASoj95ul5N+NzOBSSMg4L+LY2KKfKULP6grdNQkjVqHW2bUJ6uvOSS4s9nz
ZFesK2TrLVu5JBuGTUNgxey65NNOseFn1Ne+R+eFmkhYmSEjhiDrOtQPeAihoGiNxToWNoJoi0Q9
UzJMwjFRvI1vVcPelWA0CTv72Qx40nQpOH0YYnqLxshHB4ggjgKTn1oNgF92Prq96KE2jqROCH0/
jyGelFFDHTNoGG121plnL9lTz1dN/bpeAY0jPsGeQIvYMe27LQdNyhSUsHogpq/o+LLtCkOBKp4v
mn103cHZ4Pyp6T8ryfq5N+JcxHw7NqMiz+8Pkng7SoMCjlyRB2/IOEKHXHNzMGoca3REE1TuaQrM
gjaAGPrG3jfZNK9z4wXnJK0Tki68kFQXmzWgpA3bnopx7WEHXEMoezUC0OyWd2IHkarrvdtnZqQT
8Y0Xjf3C5FTajx7ahzl6ZzlBBV0pUBLwNtnsZl79E6b8EFE2DnUdSGaqDAY5pH6Uw2Ktx5jwF+4R
jrdSrqiygkOWP1Wcs/Y5NOvwlPhpfAsu/nCFwQE0KOwis8HCucm17h5u41KMKRqdXIYVLPVaZUnW
dFQb+qzkrrlKHDfhSlwBPPwRqZQRE6Gk1MZ9rpaBXMXdMy3wt+y7JID34u8+OrKkolLzYRhUt40A
AYaPbdn+3xNI/Idj7Nu81CfxQf00LFHFlzkIHhyyrsNP2K5gejTlDF6gq2Vmi2WHrDons/Kq+/i8
VTJp7CJUsk1a9sVfYTjQr5SIvbLJbwNCwpI/sfdRl3+0z3GAm3l5D47WNeQwk8a8mdSA5mBR9+eh
c5XWX2Ut2sD3er5btOI1H5O4oVWtOxIUpMl3/zunr1MUAfNG3NBNZPCd6ik90wUXGbljFAlg9NuI
AlLTo6fieAeKoCJ6CX4SC1Noa7HBQAsm+z9cb58m5njlYCD5kYIr9mx2STYtEGeo29BXkxvOIMNJ
eY1qLq60o/8Tm27gVwBpa+qq7n7h4cbyEMEoxyu+U5KrcCaB+ZG+iTFtAO9Xodhtvi4DrNvzNvee
MfRO+b5RyN3ZMFvHm2hmsFeXBDdQribx+SScOTZoYp0gH80P2iZpSkTyhj/lBBhV2afEpaP5eXSu
bW/Vpa9sPEbpaVOLICY4xRRXplqnzNJ6Yo/YRYs4xGiCLwb3hOI54/OThubGlnmZPRBER6Osrf+U
lE5SIEpCf8gjWq7n+esZTXBlxgECJ0CiuUzhT/l+EmqNDJbQa9wby4HLf6zY5jNKoxycVirICeXD
+UGxXyWK7tyJsgX9pWOClqoYLn+08osZ5Uuoifo0agWszzQhxEEo4i/gztZJfi/Q+5T9YcdDhrZQ
/Ywd5UJ02W3bFaL3mfjw8nDJzVH0SQmAyYcHIvlL3EKv0vUUx9POOe3kTn4JXxXboRU38HxOkOLe
gD6E4Q/0FYZjXBSJpOG8yGx3K6n3OkbhoEEnz1FtJRCfOgBcab1BWDVqzTaLrcItCuBuddRxLkP1
HEiZilYT+Fmo01kn57rto8FyXyzR5Lt4A7Z/RSH97zN5bGqnlTDoG4mFB5yx82nM+7V3QBJF6mGm
VXto3l5wj1bydZ2dmjbiA1VCtmBrPUn0MZGxY+ZlmeHMelD75Ol/MCGhNjz8taq71fxTu2YanCMT
fgsQlrKJUmNtxMR7jS0R2QYSeTOk1IeCf+JMuEgb2MFmQHr7xAuE9ZQH3hjgsFbbgvgcQcSbeqGg
fsHtZU0SGxQdkjaNez+2ZttzmCViSDGexQE7CGFsMs0/2FD9XCcXeOTWjk6vPxe6UWShaoOJ6p7o
FoySuGx/nl5pwfUYFZx7cZk028yXeU/7ItaXpYvlP8zpuZ74qB9OrRlpP4Lc3RGu8DQzxbBRwdqg
5fbfmOfhsvMnKpqhbVd1FgwGx3nVzNd0tGPv9dPmeZQG7v5PbLF//ANksoj/6JqKeOgrLkYhs9Mq
uUUbgJjwPETljklJSrD7MORVv9+CPD3X5+/how5DOSbm/RdG5gMyNj9SCJxVICDQjRvpeaNvdFAx
yLwZTeP8bktiYTs9rweXoqXUyB/e0pe9mZdGZDms9R2sxxXrh7U3vmH42c25x0E/rW04gxfuNba/
3IEuBZr9YI/1ifv+jZZjbDnyMNQUyjk67607v0KAya4KcpDXPyuRKFFC35PpDC5HGYBAp8X4PvzA
y8rp/7vZMod0v0lBUTo4Hf38XoBlOM8xA/E48QX4eOPR2+FFDJnfEGR19sPsA2L38ZiSZNwZciqe
Bvsm2ZFtiaHW6s3MER+04B/DFhP+1QejQt2c7jh9grfmEDQxTwQY5+NgxWt6TXodxybas4GhNVdZ
f/JA+0W3sDdD9nzcB/1xjkrtx9VQMTjZNN5c3vkl+z6TzZGUCMdeLpDi9SN/51ZhfReOgeXTCa3E
hubSRF/hiFHCMYKACiklzVrkhPe9kQYGLBYqgTFe3RvxZ8Zr/tJhs9N5J8S3Zs72eL3H6yKmbETN
l3g2V5wMS6FOm4Rqrzu/JcNE7EhRlVHKLFIRxW6HL3FHl3my1pKmEqasGV/Sbnow4uMqkfq1tA1I
2dWmIfUcWatM9c3I+6abLrm5uaOB/3O1eUQ8SUWf8zHayf5FSCdUSeaD0G4J5PiniLQbs7s/ccLa
GJi05e54PjBYEKNozCWZPGlBhwR8+oKQHqEClSZUjiYtIRUCJO8PIKpCEC0vZP9+Aanx1rW7gBEr
YXYmB8w8uM9Amw8QLMEgRe6xxNfGyVXIgPr57uP88T34ehu2FjeqngSRAnOrmFq3wvLbwjnxTf0F
vCXz76J1opGfvMYp1WYO4ccxzSgqdVnSQzNp1i/wO5XDFWVqN+bwRlQC4eKoWJsI/69nzqVJNBpU
9M1lEE0aG0eJUAcqM2GAKzPG6CM/6NAk3/u0jGywuECacFs8jrNTqDcULfyrGkUMxLrogxSPw3WB
pJoAybkSFUX5EAg/YwJE0OC4l1ZEIfaj+cU6uOKnrrL3KKcaHcyxfpg3rBW51kde9DLNRnY4MD+p
rNjwqY/zj3tQ8zEMnhH719OQYqJut11SPMguptEc2qmw7wMmjHnEatXhXTxhAK12rMr8Yay9tMk5
bmAxSEACUcEIvzLl5srSlZJVMCmv5jvmc+C/LvuAOkkdfpg9y/LF8Z0jYSU5A/FQARJAas+yL0LQ
+qm5r0IFCZI/yAppzLW5dbn0y/n0v1rgnBA6ZfauAoFdZfMVtm5NzSOwPMG91EemHnJ53TPjl8Un
dmOVkfRj1AhIJUZ/gNrNOk764HsJS0y9LB5b7eKkNDIYoEjC6MAaIbBPkzKOEATe6JvT3iJVfR1y
pu11pYWj5Mq8UzZIlF1V1/JLlnM79swBRSPvIo+8tScGR8Z1AOYXh3rC1yTf5RDLNw5+Vta8dEkD
BZg5WZlW+mHc6ITv5jBjFR0/0fhnxknzNlhtm+XFXpcygb0qBoaydZRGGtGRyHiOnwa1nZL0E3n3
FelQutibzH+zC3/yRGeRv6Kfx3HpGppkRNzn3Tkbl3X+WaiF45PLbUIVbnYRmDl3wsFtem75rCmP
Jatk0d2XUeH+opCj9t3j23W623d6OTYTIRKGrlj0PbfIEJGfAHl9LBSnV6N/DV1YzEYOuxiW+ZhR
iAqpFTA1eB8U5rYPr/x2WQR/j3x4iOWpaSxVBWt/FOryWLpmfv/oeXguxX9IZipDAu51Hun1nwud
t/wE9eJwu2N06QPuE3BvC1vhbqKu+6rb2hl0F8XIae0bv4a0OTpT1Q6Nv/tB7tVIsZV+5wQ4kiML
ScpUFLiJMwFttMp//QefN1QnW/SdllqxRaB6w91WKBX7YkIOkmBJ1gNGxcsaMQ1MTmmeONqHkBnk
71SiCoI+WtxWlCpe4fLGxLe0RualQxFwn+eDXganHpPZkWL4jZJydUjF5gEAiJ1iVlqLDZew57wr
/fnk327Kn39Qlznw52csbkqUvE1/yyOdp/Ehit452vWATNhXmv85Fxx0L/c6KK3a8QHmo/BgIvzs
mxF1mMHjWzyd2XaiqZSOhbrtPTR2XvG0qAUYCWp7oEvckrbEjU4Rz77ADCX9Bx1J1U7amS56QAzw
71IoE7AYQo+eB6XkYNnMYPmgl2bVlhNxB3W0r9TlWGIa1EztbGoEbRXAUNmWuIBrB3CK3IeORlpE
Le/QvYJlcN0dbQoueIYEADbcMq/cRT3i8SZ2lUgmBCJetwM9a7JCB9k4Vkv63MJBkvW/OYb0VqVZ
6hvIZR4qYYfjsRf3WapwXtbrOqDmjF6wJ6jHuRDergovvImkx3on/YH3FGlo5PrlJJABBLVqlhiL
tDbKbpPDx6w1cNfYbJ96nXJT84D2CF4XAtnLTUPggwwqJmXGAtGZfS4v2TLodUQOsudwa670hQA1
v61yxieJAbMbYQndF0sr0P3/AJ64ygakk/kGuzJUMXO2Iop99fi7TWYe9Q5HjKlXr/V3xu7/GqJe
IdDcVt1/e4LndcnRw8o/iI4auMRaJuzrM/XoNvdyXWDU28okRc3xS830qM9Tty3e6Yuuqp6Hr4z0
PkCAAjPBxz/ELc3nDsLv4YvYyfMj3pfcR6e5/gF5YxeKA4MpLu+cQnY29ZjAN8jy3TifyNIREWVu
0hvdC4tea6vhHOUtu15uCMaoA/DRN7gkMYWet+IrNtOom+qwB7jsxHxWUz8VvrH6Vj1aw4o2lWWa
0mePHEkTublY/f8Pn8kseuTQEEAjRe7Fxlwv1QvNDmVqEUyxG9cweR032jPmNMBuaWYYcd4tL8Nf
0cy5yz4QiiSVvzqfPuLhr8yswKsSKCHZAw34K3kHck4gg1lPA2gwcjQmoA6u3MmtuUyfwlT6gcnW
bBX9sh38u1/IIqjBzk31MmJa78ibuatUZfLDW9I43Te9mdmUEd1WESFaLD55f5vMLSj2VxRmunPZ
eP2KGuWtoyeJHjSHcLb4+RQOofFI8kKcPe+NwH7Yrf36AfTPyecDCWWrAJaMLAIjYi1T4JibA6Je
wKAMiYzm4W3DtCSqaRlKtcgmTC/BchQcA7EJ6TVNXkTSXTsI4rVko+HCOTmtnig9wQrMGwKd+WC7
S/Qzr3voHqRtcAu1Ee9AtziTBSKYlh5pUeXpB+cViEluUPmEXLI9znON37JTu6E3eesCyZdLpB1p
ketOGNLePK+X7qrHf2H2lktj4qvcS887Rl1GBXIQW44oH1Uqq7B+9eQy0t3O0UzQ/lLvuAlKSaUI
kSdozyKiTt0hj+eq073FTvxl5GzfvXbrRPrNB3kSarBgVmIbxqo+XG/AU44PsGvBpUqQR6WGFIXS
XuakzZ2XEQpP9MYR9uKhuvquJj8uMiozW8Xyd1NfKqBT/UtRqtXuqytHln8F5iqIjkoALlezwymD
mHmXENteFZZc8efJb2FRfibFO4f8TnXtmH/tLsmcm7ze5UVbejxlaOpVqUOpMsyM0irbxUFmEk9m
IN9JS+MNBFtjjgk3nbHzi2AO0YSDxvX7pyYxmbToBj/RMaQ/bVSWVt23ufAlG7EM9z8m/aj1uC5p
emgqJOLuOTfEs5A/xEkFeZ87U6Qc+6DLlDKDZXmqAZbgmfKQr3Upo63bSon665Sye/FTYSg1fWvG
sZvCK3WCUT8GQK4bSV9WywwV5e2YF6tvX3whMKcV3t+iQG8fljekhRtUKE6oF6Ot574cHbG2WnoB
S+XpGLOv4qXLUrXTSm6NR6U9/+/B2Yl5sJz8ZRVmBIyXFJ0+kWFqycfgZca7CCYN3ehZef4rRR1Z
x5/vYe2AlDhn9alji8t9Nrgxk+pC+UhehEiwTDDeSs9Gp2VrF7hE9eA9JBUNd/S9iu4wTSXOCib6
13pW/WPMHYTR4VbXe91XRzr4zNUv4uckhRlqTgwX18GSBAHgEFQo0BEMI5hMWjjjlqR6r45keJne
iUTc5jaKvm3UiTLoP9P4yJccxMSGL42gs7DWRCRgrpSyH/NxKYzhK9nCmVlBrb3TAq56DAiuE+N8
m3xmcFwMO/rRp95o7Qn3QbVKZiv2MPyqqNCTZmrqJZNC/nQSmeSgsVWHAZXpQHLqA35pGlYbrE8q
msk2DYUJckxeHPhZ2kbam2O9xKusfAwh79iB1IrlWbF8+KaZjr4U89UyjKV6uUYytk/cPbj6JHIJ
tEMyfBNCzQljph6xlSUklSFw+63dP/f3YdNIwegU5i7fU3x8Y7GV9kWYdal6a14Ix/V1VvxU3i36
34MjK7w/J6QhobYom0D3Xs7+umrDVJ0PQnZdDgqllTmbUR7sGXXNiJTSMSK5pAAf0idApFQ2eZbs
Nv6ttHqAAMaP9pQykHIOrZONkwzPAe0EXfw8fo30vqxYe13FiJ2eJHk2W891ydZIzBci9Q2yhCpq
DkQit/iVFEsupVj0302qmacdYM/kNVwjV3T6LOvp5ALGuAgXHGRIdL2q/VezIZ/lbfG27Zpo66+n
EuLRBCMsL6Fov9C9t0RMFmlIf0/6zD3Zfyc3KXNKxTgm2j2uVa+BMQe20FQZ/XNsSLWbWMgu8wro
vqZXP0ylT6Fz95w9Vm+NmspWingXElruk3PEGCIR71Oe9HoKthf5XWq5967tEV+RD1alp8Pns9KB
SCQqzMPeOEdmcHq1Wcmu8w4juPN/Dxc/vn8risqbVJPKonVGXY0cRxkBquo+bcdtD48GLKHiTl4N
mWZ6gWpwmDaRepgzWritvlQ10wZfcYu6Huw1pmEaTn8m0ZFWrUUITo4DVpWpiDW+SesiOO+kY6rn
eRb9fZK7SajyMsjVeyUMqOB1fAtwMWVzoSyRv6MwOXzAyxnhEm9S7d6oFSvg8CutZcIwD9vE+1Pv
qNM4W9v83V32rsnjuIiBL4YEsov+++3mixjOUHSQatVNdvlvDdHVbZWqMibKwQHJxGLLArqtt8Yv
C8YvxxjLpnhZ/RI4471bSt77LpBDB+16qK/C1RE7Lpschk9kDhdjrFwkqqpH+7D8gMj7rrR6dQWG
bioVnP7yRF5fskkLJ3ARoziPupW/2JeF9xWPX8QUDnjaG87xC5M0stkxPzxWb4u9Zwl5sOvcWGzD
0mQh5R3htt0GWu1uIAG3q8MXnw2mSAuPAEd9ub0SNHd0+QFRrC5pDVsfjtfGQqMb9ClaCgDjqpTq
z4WnJYC0KVvCuPqwBEufOwFWhjXG+noAcgtZHhEXOI+f1MldiynFVPRSq1VZTGxuByozLs8wEFSt
cfnbM7O8dqZzlQt241M5hkKdoDFZO2h7u9DgO4X04emyd1l49r9h5BwtXC5aAYzL5rTc4VsxC/8M
nSVH0hFwtI45SZ9OetEtKIMbm1ec2ee9AdJuNZxFgtIkw90NW6lk0bc62kHU9+yrYFeplSApYfSr
Vy1dJXQR6c/8LF/YEZer7U/GNOSMfjdbjmg0fHxW3azkkASXGeL3taqDAheAzkta2xN+RrTjS7CR
Uu2WKXtg2j2lfKmm0rbwX80uRont69bim60ro/3TwKlu7TClZBcIYBdYRtfs/jCq9V3eKiDAESqm
CPa/gqN9h4wOuanTZIH7XqiEB8ddTNJFoNRsB+2x7fbmgSVFtxqBNLAhSlhRLZiD1Afkj42ARTXw
mFrw+ed2QmJlCkinwWBtc7ikK9baIm0rmQUivTXWvy6w1BLColMhOfvOKE36QZfUgZH2GxBmwMLj
Nz+PvW9CAPIwBTbtEb+cE9ShOrlaAkoelo6o861S4UOmgqwLfnsZohTAUpGaPPOu6cvtIAOi/s1X
znATiEJo7DoC5E9Iiz9BzfIlroRMVH+KB1GwXn3ir9XYYTyiYOB4rqk5pxKNB24q/4Ouhs7FbJx2
JUxb7loN8zPnHSZvJ3MbC6xWLLmR1fE9AFNke6lTT/2PQCIbkldo5jSOJAQODBPFsxE5ZosJU+Y2
aFcy8MRJyuqrbpGwPiG8uiItC+1DwxdHDdyUDewOt5fl6M58VrZrzCn7xo5oweWmYlM+vjE/NGUK
suLf/E6cDB+5tQ5cDl00bNSvJzKp1k9AMgmUAil/K92EzVAs6eSoIjOztPGRxPxKs2dSgB+09bFG
blJjzljRzkkx4nuyhWm5aKzc8/pt4oG0lg7q4WxpHtdquDbeTrUhHytwpvISwMK9R8aABizmkVB/
8tzQ+xkKDBLBjErlnTug8wkzj4GmSr7LrtQA75AFpjDho3ANxkhZjGyvZNS8qPcrUXDreNqr1pTA
MyOJVV4UI1dyAqtqUzoTWXoLaSB8ATrUMUb5PdlWl1xD+g0ZJBLgmdRj6kTbNrIz4VZArWnirKka
GTlYn4KneWpAvG5bez4Pvwec49mhrRutgGZu7l/jfDZXr1dcemnDncCKriAC1m8F3Zn6W040X2HM
YMVi3F1v/QrUHerMAz0qHyNEUdbJUClD3rQlI4ukWqpxtSS5IEEOmVZaVydkwELcIFRU4kMl4mqp
ZJ8WgREMt1/Ryb7eLOKFQ7Lu4UCcIh0x98Ql/l5aWTennlOduxW/UrK/xDFN28MOoeHtt4mxSZh5
akM55AZz6l4R5ZReObSHE04mI45ff1a7aQwHo8mZ1jhpEYESKu1usWE99AbsvJl/7ak3BLFRLiO6
3LC+31xs6BiWfsJtnIaOOqAOMl/QYkUcslKxVsad8pg2X3gnEXdGwb1lxeAd5/eX9JOVhA8WDdyT
pcAVR02tyW5UN0ScqRFSusUtB4fj6JT0xB+dl4As4+j3NIdRbxMYw1QNfEHVRZZK3G0RZxzlrry+
5XpQxAiKOcT1nVxG0TLNCbAq4GxbVgaf1Bha/qpagw92VaJELAKH1xMIXQqRzWC1Tll2GH/yvaOw
DT6SKJHR18RKNt/2B47cSIHTRLFR3QGWMYYWv0bpsOShDWRYz1dmAzxZhUG2xB1ht8vM1eyAY4SS
e48F0C1L+G6GrzYPcgs+Kg+lU4ihFf1PZEswpdOdlHwXT3+hQ+52QbhQe+hImPKcdbvgY3J/50Sh
ANFPuzA+UMPcsYDruWScgUyzjMnA5yH+L2iFkbVm9WDAfGCMqW0HMCA9QxgJ9n/lh23JdbkhCE7p
vI2n8S4KgeaBM0Ojg0Co1/DPd+Muk7Ksy9sJ1QRTaqAJpt5K8twNlQMDIGndJ9UOgTLHz2PtQz7B
Kjnzef+swbH9vJdVCVPx2oCIyv0rZddL4N8O8sLf2EG3iV7UTGKn+xCCN6WNf2P8KXzvlFkGh+2K
uuKMrEmNKLh8AGrI9r7EUjuPRB4quqSsk+j2yEGBySLUWiei7IdfhOZVEBU4T4VKs8hO7of/LLHF
KA9QQEUMKg7ag6q8lnYQIUSdS+vBX79zhuppKew2hX1GfZf7fTFulx7wUiU3q7ns4YvOejqDEs3/
SHg7kQVKE6ZPW+3QqdAf0KprWUw5aa3vJ2rflhEHOnZF+5YYRiAOAW2+wllg6Kdn6i+yGQ/dzoMS
L6O1AO1baNev4SIpISRvMQQBO0axwaX7SbEq4gpLzg/N2jbUTxDI5FYFfLjcFFuEO+qDu/OnzZ6i
U3PvNiGCPn7s4Q++5bATHg7wiAXfcGrOjYZ4BpvV/BvRKYspHQd09bOZO1rYhNGMKhWD+Hir7Cup
wZp21kEfhJ7mk7Z7EZmkyqP+FGA6043y1NWCPf8A/cATWE33fWPJN96O7ctcHM3yT2tvsEmLOkKY
4/Xb0G978YXMMLimjLdBUJ8YOBEa5EYSTbjtjhK91NKGhjbHl91Onr2aCYcLE+DW9P3i5h6NvB1J
EbwZAf/LA41YT25LYvdN4QhgsRyweIT/71sRlTZBTL7iDcXyYfGe0dRc1GKavgWIzbWTmXx2HqFQ
RL9ociLoXWk3pnWLjJmWCZqNaPwRqAcMpToUSEL0VJ03cepIJ1PPrgMFTdFlLjDsgDt55lWEOIjZ
nR0U8XreouB3wec/21/BRNg8kwPEjk2HuWS9huWUn+t3YhVZyJB4oqaUdMVnK2VyQCiqQgirl+/S
uMbe1Q1FaL/vJXhZTOB6jWCnf45RNTc5qS/s+4Lk5UKYLek4iBpex97FpEXa3p//p3JsL2OkI9hy
IfyeKyFB38MkHR5fDPDlIRgWPxp435i1wPaLcKZ/npLM8qe60gRf1vIck43WxKiP4doqLon3NqWE
K6YSh7HEbRJFpmXBGW/3J2KT7idAqOTEXjS7+QxtwaO/efUAk202AN9rsO78B8g2BifWAt/vXsJ9
qIa4NMUH2mkbIJWoiqShbcBMowX5ealf3imjSWl32jJxP8g3SGWlMuIou5T5dcI17NRFTp8bx6kK
12sFQKe8e698G0URTT0jdONjjDpyM2iun5e0MK5NkFrmPlq3Z9PcP4YNA1L/Za3KGuc7t9Hpvpxw
BbUGf/rJ/s+HYGSSFGYLtTuinHoyWKGT6EDbdLcnDGYGRRseA2THgeNrbY6WWj9oTGkAHfIbLAvs
7OxMGsMD2oiqGVWWjujnUxW7J+E6Pnu4Lg9wWj/y03a/mvaoSexi0lwgxA8ZWjCxS0Xs4mUp0UqR
FD5T1v2es+XXhodBnnAW2eOJDQ2upvd384qr+Gba7AzVpfa3nanK1/7wDrjaQcAIy1gC3DuI573S
IsAuR4AzdeWfjau81ai3EbRBLBRs3HWEvcctlu/V+T6zwaTbT7w2SATfnIslzEVFXNFxlwCDWE3I
UF3c0+5NgiIsmmzkbR8z+eKRyByDE0yE23JMPLA24lrkoa3eEoa2sIr70gFDC4iQ738XYYQqK/R6
AyKSmjo/vIUb5zCLfBEdb5TFJ8owJ516lyLZZgyyriHoQGqeZaUkAfoZ1rSHLsbJTKgUAqByIlWf
7pIWXkzsHs4wl036SvaesqQjwhTfZKEVS25ONrbcnf37T/0FapolR1xwllP6C5dbTDYRBehbqoXl
+5AQAz5idZzFc98sUQSfzX3uJvGkmN+7l8l3m1O986NbLiWA9F5oCJCLyLnBsXMi1TFJMva74hnn
Bhx2XSqRwikYbZK2iVL6suHxvyy1LL26ESL1Oh3JoQaQCVyI6SF9LcToyhO7eszytrXTY+SuM50Z
UyilimUKCEZNqL0H2K8KQBbkH6nQuNf/haGzjIQPmam60gX/EuVEg8G5LopDLI2vQWhW7zITmdAC
Ow49+tZUNG8smXsXG9WKHHKu65JoPfPoKazLr5XCky5YwuJmAZ0pJ8JqHAZDXMBwihBWVD8S/DSW
+cZpwQKVWQOf+NwrG9jGbePmbA9vUNSIZUyxPCoGdKWiILVb7T6WVrAD8kWHs5cBuYlssJ7Z3d3Y
gKDzsxNbGbIYWZg1ZuyjCkeypSUN8LSP6yYt4SLmOpaZVJqTMyj5GolkUfG7WE4H9WAY9kwsx4ha
DZmvqQbP1WjmfioTsxbShq6w+Sz/WLOqc/KfTkyDdRcOHfFrmLi/N/zt/0OwQq1Daq4mWJjkzHUd
GufbUQnvM0shnxm8rzzwhXWWTAUdI2niRm7MAgjavUVkpFAb24V7sdExgzPaUZbqtfBHyrJRGRds
hhXtICI2QN5QmLlnjWwUqZBS0yzHY81CFGvpXlcCeVifO6jEiGHaUvV8S3Kv7xEZ7En7mR1iI5wQ
bX/fb4TT98lrOG10alxzxF9AHJslaRjpN153JnP1i7EnkS/NK0Cfl8N0MEg7z0X6kQSjJL97a9bL
FFzxOSwEuXe/tllMxLWFFW2x+UTWMpRc28vLb/NQQz8j2WYzc2WsT+aXeX+6tj8cteg4pdsxVFwO
Rbu/dfdYYDsQ9SalwrHGPSi/pEwfPQI0LS9GYA4O53QiVzFIdjVQeS99NSLYfOFVZakNzm7qditl
HmXZbWIX+xtvh33q07XEmoDt0K4jZEj2PXJHMUqOm2ujOnvTwRAqkyKJR9hiylcfaW6i3XPkK4uk
qUn9vJv6vAiXYDgLOJwhHj8KGjuDFUXZ9WaO+Mizijk1q9lQQ0oj7agjzJpzLoMjRKcpUMdkWBN4
Z2BiQdLRGlNP9a8ywPV+8sOFZQvBsORDbRHbnrGeDX7V0Z3LTYj/0Q2HcWvkiODtd86DbBtO2bb8
UcVsk0mKdub35Bu8rQaCQKl2cpobpVgFngvAFfcJir6CHZAup6V8mC1O2o7Iy/SzaMDIGUo7mbMb
hPFuoCGmueJkMtmel0IY0pM89Uhts42diZhatR3+HSnRnp9KffpwHcfFMhbSiHv2CbUJ+qoIlk/g
Hut4Ys2NMtEIlPQqhIsL7ZSnJDoHv75rrL3Nq429/ha9a/BjHRNmGBvrXlcz0PDc4/w7GYbMVlII
WHyvEj2XbCMKN+p1KKsHyr+VwMgpiDAvDlRQj0oWuZwYAK4AjZ+QndraQ/g6E/2XhmNJKcUpb9Ib
XabVh1ta37CT5qXwCzKvftSLktnDvfUW5KYSy5KMYCjtzA94ldbB0JAyDE6jytc39OMBEaOOOX1j
ZT5GFN5BcKaF3bgK1hS1numkK+hrpKahqlQTB7wKF0pN/Bak8EG5V80U80j4UxIL3c3a7XzOXiTW
mBr0WGHN8UgLt0q/eIpZ6OAbJfO2IjuS8vNAL2UyIrSmO5r8PXFXC/pyXWMV9kO3qJrGNLMNh1O6
0XhT+ur6hjkGAlYWSCN/cP/PlOMRMj/KPjaggSdCg3Xynn6DF4/khWGMtzJknISp7QZpT77HYTv8
Q9oFYqWsqLoqicmsZGy3e5qolo9kOsqjT1QFYBq1cSQocYplm4xfPedll6ZELnlnT5czR9ngjZQx
epenG4Am3XuUnhiomws947dJZ6Gb/Wfg3XGwUFL1RCWNScjIDIg4ajv8wcy0Xzp42Y4LuzjjwgHu
ISdmg3CudARDrwrHxKpIfmneYpkBmniSbri8XL7qTh0uQzESwowKWuzCoE30jBX7prRCoyoFCgCi
qAUU17WQWEZcyt7C7ioub/mTc5GvGsYFc6KqhRZbn6q1VfAh7CDf/HCzktWZy7KI2ptCHdICrj0M
EN4SaEG7MYJbsNd2cuU+/2F1OvOJ8SBwUt2mTMPEQLfW5Zq6u/d3YTq0n3pJERY1WmeYOibJfXR5
ysDQqIb/cZFcNVJ3wZiiMiYTFmf4kRXNU+5kDGeq7BZBk9UaOgC0O4ukEIePSVLk/UwiAQa4gInV
1Sua/ADwpUWB1xc8tSnXxzeGT9QrKMSoIaoyjKYzDW1Ijcbtg9K4OmUfu8ReTw2I6/LDTXB5f06p
lTB12dL8qcJFOee/WsjU/4t9oW5tS02auJirD1/Z7i1lYO6zYY8axP5769c7YiYuitD200KTcP5t
fYQg6LxHrPgXW7qkidjFcBD/MBEUynKM1T5oeIZF3GmhMEukSWjLnDo+lXTOWZFvueNHc167yu4j
ZtVTaTHSDp3lfb1Tjiu+2RVm5fZlnFcuBULFAawyHDydCUQvXpHmV5sYbYe1+N5pwXv7E8uFE13B
g5B2TU0sCq4heZuJmmZvgGuHwIMHcCHuHfhAcU1awkEk3XPGiTZaqaSQqfohrJ05g//AhfcDMkph
U+CO8lCNFkE/mA2llowAMSg+Zn5/DAbTVwm0onqepAshZIMe05YG5LXIueRj3thihxPlAu6wieOx
8OLZTtWWF/gmfPQEO8ckaPPgRejDyyUY048YDKiCt+Bt/FybPw4b+m7ixqoplcjYNPQc9rAdQTbV
gmPr+S5XHf4HffBids/de31zTfHgl94mFNhlT9exiSSZHDL7U5XbMspe2eyGOdGGQaa+1XNocq9E
/sWPakwJyc9DwZGFMaS4XiygVSa9aUotFhyJNuyv1gaO5Gu5zw5Sj5J+7Xdbu58GyoIReeXiutnM
yQk+B7XGQ5JfekHwU3pW5ZkxP+YCosLnVePNXcXIAmwGPbNaHTemeF0buMRPBDxwxrFt1ll77OOP
BkRRGgzsEorppkBUdn8/E0NQm4gPnZagFPxsqMdnbjiQ/zO18Aqaqgw0P/A++0vRlPhb3N4O5Rmj
kn/wufZPWrv7E4vqBwkh9BUIRAPsMNrisRXt6eK0j11o2m9uRcMCN8mwqdg+fTOVmHrvlz7+wfmX
gdyh8vtPJpyjk14FSiWGoiYOlY2i8/4AmqGLchhSvMHCyPwyrVgCX23ROqFb4uKwICKf52p3Ll1N
eOWD4JKoMLOA7w++rp4y4RJ8YQr84T+T5AtBGZkGyi9jLDJDf34CKc3G1UDernbYOcNqTScwOQs1
l0i5LyQOK58MPdCNijguVyBqm4HArwk/1ts0OKTzPdiZ8c3iDQfHLJRATXmLomj2glMiTTk5AHPu
uJ1tTnZsN8NAB8ICUa5fbrEYLAwb/kKyeIks13WnlAIGMdHSHY6Bm7Qbk8ZQBM90B/hPLKEgMucn
O1EWlqhWunoDqI6dz+qQXvteHXvCIpg/7T1qpPYpSn0qAOnRMgBZY6neiyXdshqwQZitfViycpiV
CEEx7PuLxqj/S4wim2evW3LvCKRGbomIun2Zg9p3GdHjGTtC7dbFOSxbOCzdjydKnxR1Gjn6+yJI
I4DGiWl7c4+kLeqHKdIqIzwtZ7Rq0mscrsDvMzHHB2TqGKBSgwp06BvRtYYzREO3aJE9Nu0jzVWZ
K6geyekwtvK0jbq9N0b3bneg3kCY4JBuMLsfR7cbZvjr3CcTPclaZWU6kRyFiRuw5JQ3FZyrVmTo
QIyeS395+mnpBb9dF+PkJVLPyzLbPKavuQD1GXUhT9Y8QiORKCNtFQxyWUyEBTPb9WrTI2jh4/Z1
rxVxHpuKyaGOH60WaXtH6ZBdEY/7omeJPl2BZ1717sfqCMCsf0qsbW2fyV/OeY0O9ZEpWT1wdYuz
VQZZzfcCFE4nUUG4Rp0KBPfEiSp+5ID/8TBnVOXAqww2n7LxAicdoEvPf3RuzgrZaZSHiBKXKDNA
I1pki5+KwQLwPVEGxBXLsKGbjkCN5OlZVPwXDbAVoMwrCeNC/nsaLHRYIV/NoFy+lje6Vc4A+Lf0
yp8IqY3jypBOrBn5W2yg65I95KoTFGo6lT08Vda376zizJe15AnYURZMwToV4XoR3WvDzIrkq0Ll
WXWyCJw8E/vainK2uoOfgCWqSfsB24pc/odIKqwFiy+AAF/FYBV5z/jFmG5k7Ckod3XW3JGkYYDe
SlRL5ZXR55R7i0Z9Ig3EUCyyKuRCeOfiye0b4RmwVmeeyHrnMz/rnC1vER3lHOBkhutxhrzRtgc2
+AwwaCSH822RRrfByFbszI0QZ5CUbiFx1riPZ+OgREL+uiSxtIlcgApevyDvBNQFy7WoTdNhNew9
y3dHnnPJ4igGSSQrpoq0FWra67OiFalrUBd8+CXi8luOCO8LlpHSlp482Ld4NJIoOo+HN9XMVG+d
xHlTj1wLXplfuSSfe/nXM8ITLHRQYLhcbQT56jM6wdEV44/sf/wWrfzZcZ5itwIbA/Rni7wRybOh
J/5hydXTcObwQC6K+LbhkVfM1TCa7A2CDhx3ZA3t7eLU+P9ITibxHKLpWQsrUY09BCWmfdb/C/ZJ
Wmie/2maPsvLLhTrBsx8KhiuR4D7VDLUq1gfkJLS6kQOrMCEddyDYorTWxWnrkr74tD9E3y6RlTb
jfJFMpzUQfdBvZ0bfAm6QVbvReptAYLtgQkbFCDbyq1N+38E8sWM0airFjjbpFQFFvA4pIpfxifK
c7l8MWnu/3lsGX7dO/fbgoyL1l3OCKnMfuJ6yVSuYP7OYpjlGimILDDk3EvqMNQwOvVS0Onnhh6A
11PQPhv6q+VJ+THkBt1QoBWRK83Wl9OQ2h8ZdeF9QTa/t13fENXCI+ULoDWPSfLZbXrbgANAhmJd
kN+8UYpk1AajN5mNUEXI6jnb4d4DXVPKQKHE/LKj3FhZmz8s6mGjhbc4xywiwLWkbMFeoWwEmy46
hL7n0lU1eupPDkAVOdLJokCFmsZkgv+QpQYxFX0xNBoHoXzUbHWJyJZWphzeYvEY6sr4YVeC1eGw
/bAsUSJzETYwLRcuIWLpLj+oOpjCbm3/HyfKmAcKDa9hPv75BDpk3cHJ/Gs3ZlSgxxkhjLu/B08L
V3jyna2A3H9NtR0xrcw9ZI9HI2gDoCdGIQVU0akrO2CewhJg8/+KLbSGCcrfSbbg0TVT0YbaQoDq
nePZutjHAZALIVMVQeLs8xXfK3+D1Tu3a/iwcxcr6Wi5n72grxdFML43tCVDFIECfHcj4R3dKNJo
B0qWTIUoa5wwyauZSh7xrx0cSAbFsVLp7OHXF820dr4GIxnXjPcBdK0I1frG5YREcSi9VIRPn07H
v98UGlNxS7PEHEaoMxGdpIiRt9u/WqKSuVRvgtVgwcxMX7dht1LcoulpNkuSl8CsdNfEBIaWiemk
4uE0WujPRjFDniqyMJ7WEwUlDfYQUYHsqvTUvpdGM4rI10Qm0QwpvVU6do85jz23wkmuJjRaoJWC
hAB+Xi5lx60/3b5H5vF4gXGA8L7jZ1SQ6Xy7j8i93cfkEprFRf34bLiS9NrvXSbOVjaQ4Wvo1kwe
BJl6wpg3JfKUHuzcOLtACOmUf0PzUAkPqbJMpk5pva/cnV6+JlwLweG50KFKMyrvxHyyVOiqsh0s
XvkP70CBxBVK2fHcE7i53Y93bOOG5kf7sNqTziVFkn6YUeAHr/PVmcBfapyjppdyMIJqDFc9tl5O
8RW4oXd//QIAgQVKvh1jFkQzsTwNjS9uOD8z2FT8Px046GtjR4JPqZQX1v+ONmIqA5UMFNXh0139
sU5l5k5PHpModVpvfoF+nSpVpCqhtPFbMq8zBqykzHH9ttvGB3efkImvlsB7Txn57WdyyK5Ox+Fo
wr7fG2693SFKdzpZ6lMhlUQeYD7ABoIiwYYa4DSH354153fxCIb0K552tDUYVpAuvPk3J4SfNxCh
WUSlK2AcX29yOevNIJKfUpBeF3rb+EVscYBitCwLeITDkfiXDYlJBSY8Ts4EOrVQ0lduvwfrZ8ut
IViPd9Bfv05ZSKtMjNy8X8EobKDmv7bJmwzCf8GtQNlVUQqbkS413i00LqmhgHNLVX5q7MgDDSGr
XPPf3eKyBP7lMbSf/q3B+aT3Tv8sqZEWp2gHGhfuIxteO4Yhtcnk0fFm6y8s/M3RpIggHoD22V98
mYTZvGNSl1RXNNPtQ+7uuHgd2UQeLRKsNLSV9l/cKnALBUpCFYMa2KJM98xjxO9kr7KFAa1d0TkD
2VhVp/WZUFke+sdIT9W15rk7qsgHMVZa2UNPi2QcImOBq7K8xAKK+YUy74dlxeKKHN1vhDGzQSAp
kr4rqmo7lo7uJ3LJdIK8DTngvBovU6Fl8mC+uQ6/PiPPQzfHylZpUTEqmLf+y7W5etGXbBtoRus2
BCRyyj9TDs8JNV8QPCuRsv4qIwLia2nijsED+97IIZLTVxkbbSn48NaJZm+8tCp+DfoBFfWnqU+A
46Oa4UP9IlFCT5MExKFlQWq0mkKwkBemPFF16rVr9RqrfiBqJshUXCM3XucyOr2T7L0378D7cVfo
WeI3IbuQz8rSAw0181kgkQHBawGc9noH+93SHK5awJeu6naX15UZU1BijAOfsrDwqCoXawgm2dCy
RRXHIE3dMEvZQRZ6SDoCDprRqfo+W2izFlyvDLSrnrUKkHyFXEHkiSHKkNDm1yqkHCnTf921+9G7
+nXPt1o0K2Egz0HdLZzcwGIWLMccEiO209RIzbAdTMGkUcveNlA1uuOkaAllvJfEXlUpMxB/VXhY
AIo+kjwncFHKvB7fsEnvKoJ18QDRkwGL8zjGBjPZjOcJFD8aNHVoyA0FM28PgYIjG3XwJMfFYMfn
U+Oui/3ql9T76aMgoAE2S24gyMVWn3ccq6sjv/7m2QPq/CGEmg5Q3gjj/NIeC9Jmb5A1lBC3XfSy
t5gz7EIpwkMdKb9XN5u+ChR3ARDih5ugei7dPyurGKb91pNrRTJ2npXh4W0KyMgqrJ7Y19KWf5m0
q33b7HebmXbueFBWjt2uonA8eemU8F8MVEtuwD6UboWzFucWXoQ7opIwRJFkYV/QCJ07M/mEmBGg
hQnA9n65+uzD4wJDWKGVOxjE4hlx1aYeCAl/1oIUX2ao8dDkFfp+HEqSDd2Yad/AIo9S6g6055oq
0XB33ApHaaGnNqpGRIc1eovn2a7lDcyHupZBzcUzdBMDITyO5Vr7S2Heqpe19imisdWXXwaYaQLQ
mTAf+VpUba84X3DnmvWurif1UIzxSDQiVnk65JZYWNboLbGFfaRi8pwd8oXcmPBA4Nk5ISWLud/7
PI3n97uHLiAXH73p9C60bOqU/cOq3Z3bgdyAkyWa5TzSqSO01pyhxuF84iqsIbR06HcQogNoj+Ef
CqO+rq7rn/TwKtTe8Q9k4flhzJ7DvRV2CdK7OK8eJiC2dNwFOda8xjgYkafTqxqbb3gctMVgnEh2
tWqxREWjnS0ZsB4uYbH3wsuJDNyPFsEma8stMXeAveskHjjZ9Olc5JZUPKa7Z1NifOb1dG4k7K1H
9IREgOAhUykbbSL1syV1U+SCYc4Rylafgpif4hqxQ3ey3SDXlyyP4YgMLsGe9TrCbS2u1jsl1WJG
XC8yvIW/KYp6VvEZrNsS5wx484ZyI1XjHUIeXzR03/r2FkmHWPFnA0LogwGGXxgj0O3+XAIGPhED
Zt40hYi3xpmqEPlf7ACH3kmlD3TjWbRT0ks3Y4aIkCJlm77Su2eaQ5rsrA4V+0r8RCkoDqNeFypq
qt/oLcZSG5SFHXt7G9OaAGNZPpBdMZCeMfWamJd1449rKMazbcBqsSBKY+zuygHf/LTE0/3osMeW
oJssvgUmbQCGfP6bWP7zKvhdQCsVnM9kMvBN6TPhie9AAnk0J6w9l6qcA4ebMIXc3CGHIbLkPu2o
3eIa84aXucTx1IWppqLSBo3ZXpNMZrIlPw3TgRAOutKNUNoC1lfLUvwEwBuQ7dzsX+GSMva1zwDl
uBx243ZMow7wKAKiaoNuM+teSUNB09vP2oV1n11ySq5jkrpu6zTVvpiZLIBAya/DDWF6ZZOE0UPj
gY6qtFlj3I/hXS/fFEi6q8l+nfJb0w/TaHNRSH0eYlFsf7Kl4hzCaM7nzHp8T2ZpIyjtI7AzgjGc
vGySUlBCGAgV4HA5oJykBMqILt2m0HvyXeO4RCyt6HOpqeqpsuG5sDViD8CWWy4/EIdJYdAiZeek
/Bezf/nR24Xh/BpdXATnUQ3tHe+fb0PMk+EF5AAsvzasq/OKzGo/YW/VjE1tav7kQcrRbpL5oVbx
uOjqqW9lhvtj7/FtzjUALr7KKuJKtFuAwPaAUN98fYXwMWYVypvPCtVpMPy1kD86L73+jQ4VI12o
YC/Zct3Ot+d5o6HiZ1azXDM//wLTKD1ujq8XaCw7f+sx5dP/OnQoDMMgdCrRlm4hwVRsAq3pESqB
kDcYETrR3SnMnjz5+qTlNBu5NheP5f0DRNy2V4fGMgXwMLnZ3TZy79Rg2dNrUFpMmTL72YwXnIUK
78Z5OFAl6R6iUYnu5D7jd37zDA05b1OPIibz1sBC9gZMW1k8TOmxOwpD9oW77eEMRRJ2IpGZZu2X
TBz1Saga2NBqJcJdDfSurcokXZ0QIt0yWF6q/ycKfZZCEMUzaHIa8RDpzlmpDTY2xnB7jRwOcq70
J2mkHWPjf8tc8/Bll5kRHPF7PtuCnAUTOrHGWHC9iRJFLKSB74MLABTxprxkQnZjLAF3Ji9HX7jQ
+l1gVXmBhBZcU34IIrHSL65OdWu/gniSE+kyNRICzvgvb8sILEukkOiKDyw+ZW1xHTssajziYS0c
C4D4p52N3X57cSAIveuu/Zu6iZm5eYiuDfWijCLRcm37xvDZBHH0tecIi5qENutBiI4Nm8C2g7vD
+wKVU8Wf41rtNf5p5RcXKbOWaKdyy+/xFMhhd5oR6eFdM4f+RkB4RDlYPckNAF/z4DKoRlN0urpD
6bfs2tRBbHRsJ7AJqeDxR1epiR6NlAmQx5q2tMr8k5hzjrLj0EZ6WTYaC/82YObNxydvVJaXVkG4
93s3Hur/7sCTEMTVL9TiaOubiqdWkNTzb6m8w5Unyjml5gi9/egFolxvk2TO83D7Ee8rk8W9Ult3
4c4PSBh5u7g/fZeFzu42zU1Vrl+oIFgY0CqUkaM1QI1AgyjJLC8ts0AiD+T4JM9YGhYBtN1FGNkd
4SK1oI51x2ek99SevzRvtfXskK6yiyh4zN5dNScdEZi+FmiE9wWjwyxqL3Tsl32xzguLbXhuqGiI
jF3WPFxhNE2DUSu9hYhwPsrlEAnU1R07A8X0hLXXOUQY5AI734aIlvVokRZP5iyCRttGTIibs2Kc
aQFo+0aiu2YSox5mrVMAKK0fQH7zPITKnkYmRoY3xq0JzrnH4Kv8mutw57YtrmvrEuQ7JlPNid7h
QcKlFXqYz55dc+5eEr6+gIEV0iS/4bK4RKsrrMKI4pHxq4etC/bLnkYAKC1vhQOEGAceB+HyEE9a
wBCnB34DvnGHD2Lhd0wIcc/qdjoew4hnSYO+r2xKPgPqFAbcgmH/4NqsYpD6RB94lv5RUXx/E6ib
pfxYXL8VAjFD9P7gFXAu385ufbmFEHIwni6YF7PpXmSfNfVBjoFymda4HIuEptls/h8uHPXFKNrk
9sWOq3poJ7Q44l4esNuFSCCCf4kYAcF1lap8XjpT+dc6VLiOlf/rFGiitvXkx9CzOqinBAJfvK3e
ykJKn1CGgyZcm23iTivU3BUOeQ7uhA/+yyBGG3L/IVmNbU0tJ7iJ9pvVypFK+FsYlalsKiHxZNO0
xcsCl9h0NN2LmKqHhndedieskQ5Po3zGLr4JKvywL9+uf3J7r0zt8Hd+NRkB5mkUkDCm/GoBtkSZ
sa5jrEU2CMhLNaG0VRyIIkTiEh/dZ3VXwr0+NLhgDbeMy/KBtdrTwHvwLwhAEQNYT1Xa/PBCnmlA
ln848IQSkfeiDo99o6qEofLENBaZ/s3F7WyaxaTK3jKR2QA/GDvPtH5j/o8b90WcDGDq0p+QORbM
FzlB4wj6lFYJO/Sqhdw3RkBkeD2fd4PGiv68MOFZULi1A7OuUabA9glBJ3zT8PskyXk2aaBb6ikX
16VLqs+RbtQsVc7V+Cfs9fzC7AwuY8a1nX1iU80zb1QheQkBpV/58GnayQrUTtYFOdaRo8/AzLg1
ZS0+XTNcbRIsy5HNeeTi9Hn8J0TDOAdgKrpc4hTFQvvaBsq0bpPWB+f23B59OclbY+5ZqajwN6gR
BjcD7LPGXioi1fxHviha6DHtVuI9/K96LJ/84xE8U5ePj51+vlGWFoHqzy6xIFb7MJa7ZhwzZjRM
ndrNW2ED7B1oEk42xsApsGMmU3vN8lTiSSHfjBzzfw+MnJyvkOndDDRpFR51Wf1fBOyk2a+SP3S9
QCkBTG6Wg23gG0/zpw9yoH7VgkcUGfkU4ZfIOL35i3YqkU2ZrL4WG1XDQXza9BynAwWqroYpPkPA
HWn+g+36PFG+mhOLNyQboyhGYVtGlS+PXSu3MQhDiRVEtMinHADmbz39lWPwYZxG/zGWRs1MWIW7
GCBTeJ1qw60+ED6UqbVm1jSsl46i4Nr1Zzpu1FALW2BLpjoSHZ4QrasmLnE8ltuQEfkRWfV5vZ0o
cP+HpCuKujtFTB4NYAU7GCV+KmVfUxGvEN5uSSo/hWSJ9ksDSrTJYonOEy56ve2Ads+lfH5PpfDp
wItdQWSbAr8LPqGaOlpDwQ6shiR5XRwl1ri8puevJstHLXy97xNjDBxRS7I7S7I2VAUB+RQHYuhs
qsU0wxHa3MzNURKRio7K6LFKF7lel9VF5fVxwTG4LTTwuABr2kv8ghsIUomBV9N9XomWaiodfEOZ
BDgxzWTe0/15uwD46IBjuGj+MrpnZhz43+6Wb4sMhOOu5qgLi18XyLyLyIbHVr7gu/5TQIVCBL7b
pbBnbUlsfywaEa9jPuedJdVW974Fqb8sXa4/bvvaEjEqXt5MHZSa8Sd7zEiXDPwNbemkwOfRk4V3
boo2RjirS0vL+UHFDegRZ9hysXPLHzWVHbBwM4XvkQGrd8vDZOPs4avelniozltQMhAahZBj7u1N
B7dNcTO8fku5Lg76E8+PI0pD6B0BDIAYdCGSviYQrVDjTpXxbgkvyQDFKIHlgniJ6LKWia3wDMg4
fN/PECY1A1v9mhfYMTGMzldjt8AWtvxUnnT9oacS042bmHQbqx8kXs0FUT3IKllxInrbcevJ2t8n
nHw71p/56UkIc1iYH2M6Vd0B78pLd+OloN8CyhHg/032eRDy2uLSUhF8tzqxPfnGX6U9QC7cYcyJ
6/4fQrlgzxQ24JHLfDKmSq5EfyZhgklnh6AAuxSDe3pELyBi+UGR1oka6PjcZsdq7a5sxA9v/frt
dec4ShQNN6npqGKn3z7ah0LprRfcxg4bk7Lpg5ZMzix/JsHSh8iG2rapjkXD1KkQ75A3QbhU+ZwL
fjb3l1ZRPWSamDeF8USP1FTfCsVUi2Pab/Av3W+u8ackOSWv+81f4YBgu91yYcJDQ1xoUf6fF6jH
XJC7LtnNTitLgjpmMzAb2elpsz/6nY3utGkARKQz1nQf0GOLfPlwgIcO+HBYE7Llg7u39N1PIpD0
lgNcmCKRLbAbZD0FfrVzp6GJqKNYQMCnYL7grYGuTVJnZi7GytgC1/aqKknkJDo0bwC8lJTrz/YY
vn5AIfWRSzvZSAQ45PlltAOmFvuYNPA5tapvzLLKg/9lFTNrGxCa5hSEkxz3672MtZ6FuV1sjoef
bpftme7RY68cfGaUecyPbEQjxAdLOEHeiLs0RRtkR9Ym2CF7jZUNfmtxLtw9HAf2KgUxD0DzYs/C
v7eyT8PaXFQm7gj7M3hkqRY9IzgUGImZia4oLiqTqjcjOwdLYWdukh0YoKsBoigzW+ldhvx3Tw/M
qK7pkGZG+ctPW+C3ldH09CEF7rvspiBBsdd9PB7OWyznkWJhZFVgy04qXj+2kneztNbXgT3MkV5o
fTAmkgNY6i078RWgvrERIYl11SGjmA0/CbQZUo/URCmC+ptN3NZ3kQI55uU9f8qm4tYiQCZVUGO8
Dq3X5axa1GiHr8UV2APdXgwFofteegoqybyHZY89YXZ3Xn/p4oBxVXWTTXfMRveooisqkGWB5HpQ
q0W/T4jJJ2UVFNvgfp4wQ/WojopLDXpeNqw9d/63jRP2Dk1cVYvZfQMuTjXr0ZiQIF9jIMsnpl8P
Cjm9OsdOWFzVrWrGNUnbaTT5h01ngu8z2z7UfD9oO1XxzUIR0ldGA4w6dt2BgyXEfMzGM2oWlxwD
eERmL1X0kry9h95eIYaXIngnihFD3DkDrRvVNCjIQHqPVAl3tDLPtyMTPxmdXhKihlFIBH+VhjBk
6SZgo9UQ/d/qCoP7BcF8qvf5Hmd9VRNsF5qkDmwJg5hYhLJT9DmQeEPePMKnvboFe7p3x/peNNyi
REWxoLiLkpakZ61mLmy+SGJCgJ4QcklTNgDp2bu49aXegtuGh8dUU+lCeEJjcyjxNCOGltUSjE8P
4eR9XGyUleydCY3ls2E0gXkNgzslHLemDA8y9+pkUzgs0oOPBanDYZlDB8SmLv20Va/ZcjpRPSEL
SreBa+tWuZY1fRxI/LbsevPz3nDNe6rFeQLgViiw4MiKkiE0cpXbjJtGGy3+Ck7S0GdlFO2wpYdV
YynNbq4BsI1C6KJ4DMFX45ZOIC5Ybu40ty2BOWTCGr2eoLI3r0yv8WZvJCEGFN+Fjdq26QzHZPf3
awBPRnDgOvz9F15DKsHsh9sbab14r8G2vR99f4yfWH7UIvGv7T9ho6qnIJkHfNnNXOh6RUJZQfDo
Z0gZ5XAUOeWDVtJp/TMbRxgWWYIk8dmpUPZtV33WT/bqHB7f1n4l7lzra7VwJd+/y3Co1j77pTlW
5PVeTEMmMfqU55wI04618tW1LufaI0pg1KIEV9BpdA9aSzDKHpPGI8zftDhMRvt7B7gTfTBzXp9t
fjLYYucTFkJW9vZWtBqSdWC85/ov2rW7FoWX7eFAtfqcjweKGBDdlrTMhkqOnWBnrdseWX/XO16e
PVocqkOoE8UQUu34A1OAnZIFxn3Llw/X//qOuzezmHje1zDU3M6pXybXdlZ4ZwuZVi/VoZa6EuIP
xvyIg7L8ogKwI2RK3GYAQ/NTQLm4ccpjmHH90FvBnds3IOhUXDLQYRZ92r8fO+jBLB8Ym84g08Db
OmujSFDifCkGLygeteeGqGKyVN+VRXZoqKHfCK1gFI/iGA58renhpyo2Bau7noWMKNwAcJCJmQhu
4BSwtAq4L+35FNSbMWhtupUFCXT2xSBbcYLIGDoVlAlCNOM/+9cskv0r/RJ6Kjum45x53FZEBuj2
gf/U1E07tlPyA9QJFnzbqa9dk/WF//qItf/y8ruLgK8xqEBDCKRuBppZmtDx0wOgkHXjS8VjiziE
SPIT/7FoC6Mm5yUCfCO6EyytwR0OJiJ2Nw+XTzB/NDyj7+AA27TQ72lJirPYhG3zgxzFzLghm0MD
wn0w6A1vDumuz10uCrKzkemyOxi8ofK7PkCQ02XAkEUKUbL9bt2fK4eZLrdp4r/LwL2mRwllMJ5I
HR1M0C70c8G3GuUjRHxGNAah/7VkDMYbtDB/hSgqP27vHuYuBm/ki/4igV1QcRKExEvzG7iNr3fb
XY2+Gk1N/1ULQSP0TE3khAeFOBJUG2kFu5vplzM/NnWeweRPGYgjWBWPl2e3YxiqmphyvwMrCVym
+E3G6GFMCl36+pQgZVwvz1ryJNsre4DQsy0zyxGVNHfgizKDVMUx2dhHz/5ACP9fn/LqXRw1yCI/
bGvvx4zB/7oqt8tmTk7WFRUYVrEktUUkoGLi80lGxt+BGqLJd1eldO5ZGZN0IF54ud+DVAFgeuS3
/HsPww+mz00WjXztH/v13bzjfSpjvFELjjfN2XGBKzjyByOSyL7RvCtHEmQxDY+Vio8nTDU2eja4
GxMJjG4t0pn+V3PzYuRQcQUABBfeLzgnMaqMmdsEMSMIHyfmdJiUIinBNmBChLqEGk8bcB8shO4S
U7y5BeNePZP6/mrZoU704jfvYjYpcycUphKHssPYEGtNHA3CLj6i4hKJ3mWQ785gxSLyfCsQiy6j
fm/7BYgLKb765BMexVx4AVR3H3/jz4HKcYLV/2PRBmuvCaGcXHY+k0DcVP44SdZm76rZg50B3JB7
9+s5m0yVWs7k+TjAyGKa1AMoKzYkGWh4n9CAiLbCqFLsGgVpVog2+gIEZVC9knO/hJw7Kd8Cu57L
7hrXcZwey3pKOYZEM2o5jEaUOHdCfefzX/JogwWIB2mBTYuE4ATa+AwxUrrHOxKDleCAbLq33I8K
6cGFCJt7a3eMuKfcYDn0wL9VXcvJgg2ImGLKRCD1epULykR79BPEEGX3A98jOe/LpmS42A21V095
ULJwMbUQdvm/oqAWKUX8kVW8l1z1DNdg8ls1t/Hm7nkGej++VpSbhnEjWLbp8jK8uoYsHiCuXJVI
Cb16kzOo1vuMin1PqQUkDGY/bfh3if3BqgPE7oA4x0cai0QThucdHGh6cjs7V5fAPQ6dkujDoJqK
J479G1+gdOJ+sOob0YGWwCH+2s7iRx7RfdxTGmMzgoDJvZMthWjWP+6ql05s9ylftwFP18zGIg+C
9h5FidmRX26Yx0Iru4eGS/nKhoN4weLPSBsXBKbNbblUZCe/GIvvAu7A3SZAKuYXpvMKYy8zA88J
wqa2NGT5pybtR3p+4uCL1R8FoyZ5o5FCehLckxsSFGxlo+Vdo+ky50hU6xXYkDl/gGQdPXDXPmBh
ywWumxQtx5ruEdy1MCE6KrgD1sBR+ep9KC6bbrxDWZhtOIuROdBelN7GTKt8YS4/tyEIquc6u5yG
S64Em6I44Jnn+Xk1azaHZZMbdiUuyw9ZUIaetf+ekCl5RQ+AxNiOAuj+ADirbO8xs2GaoqOzzuOa
ybehbU+g6NV9fH8loDBb5vaQIP2gk9HUjRzfSa2HGkn07sJiBIpHnYVmywOJV81icnh5F9BYW7Pd
eytpIqWgkvaqSO3pKI4AsJAKR5/E/4SCOZMNex2pr8kq5Ox4jpcmq1+FEcSTi8lQl9L3BkPVlvbB
63dQQn2UskymlLus/pIo9b5fMh6OTc2qPJqvia5vGqODpetgZIjRpf9pdqh/EitRtC1deYMFj7i/
zh5QlcVQGzv51Z61GYEO3MQdBqLgXS3UjrU5pbcU33CpqD6WthwIsKCUOJV6StZHhoOk1RxQKHOx
9qoNNyz7tWw4pxnqX50liLhB5SK0kGcU51zuHK0VWnzXpiCdZ2H8PKxWW3y+SmS7jqSA9Yv6ZKH+
KOZ5X2oLLoWMtp/EHT5HmdRr4HlXn1sJ0diWE5a7X3IALelqDrn1977saIyeRa59Au7ZBsbdM44G
QgRbbxEmD4y6eXezRrNkollOsNC1AYi1S6oWCHc58MQWYQ9iQ//vgISRuHEKwe4uBj/Db/dVzThh
AV0LA4YIJ7lzHN8rYSqL4pnHyw7v6Bl1GMGjQkAROT7CXJS+F6K3994QDucfyQIDVBfE9Fix6J/X
Z7VX8tY5bVgqoHyItY6op/IqXCCmP0XDfcOu/JXiarA9BCehxxKjxp0HQrifmvVcrW9viMt8hqIs
yg2rqggTElNoolLgd5aM1IKaFHQAkleoyAmTI5OVjHmM8Uog/8Ej2AnKWvciszUw771kwJQEnkzG
io5Q8fvCD53RBB8PBUJhrKGGBHXkWHwXJV5jhLlP7FCzlrSrITp9SVggePC+gqqWm89+xujsL9iC
DOGgNxRjOFkrGleMTsMKkb8+qXaklk+uj+D0wanaC48lJUzCB590L4R/XRsZ6HpofWA9oCSDqOY2
e4yv3kTCbfFvn+HD5tKyWcnMO+d3eSltEk7Gc2d9mtHOHyJb1p9tYWohMEx95o4+l/YiDEuLOt2x
GC8HH+sSTYIxQxnYwJD4Tz7BQJL8PbY30N60uzg6U4I5AWjuhAEc5xMuFwohdEHXGOEOvM2l0pe2
dyR/Q/oCPLyMzKI6pWzIQpAIcG5bcXZeMFSlCE/tBS31DhMY+DPTjjWn+6+rLRg7FR9Bsy5eQYWf
3qODGVzgJfc5vhpYIAtR6ubNfftdYkVVGwFeCWEjhF54X6JyXii6S0dXfE5fmJ/BAcpL3fCm2EOX
us2YWYkKalc+pSGgFjRWK0S8MrceAGDd5x0CDYZ9EzmuXdNnmQui6h6TnKjBCVDsKax9EC+JXXkF
FgpoDtlYQRmH+47jOBCWOaGPByy+woALj5Pq/2niB9FupnelaKUK8383c5kWD98wwJwtoE4zlkGr
Q0ip6teTJf+P50Hr2B0DCbpluaRw2E+uWNx9kYr8gCA/mhZdqc53U2QV+V4Sr9Oqsp45SOmE/IzV
L5b8L7Go0ztXDGIpw/56/hG62/N2B8YdmPDYdVIorOxVmv1F0nqVGFbFfV5D4FxqzE/i2is4VAXF
3BAp7VBBTjqhLKo6Hbs9Dmvb3JxOhn+HK48QrJna+Ix3xD7HfKDltOb1afcPVo5lEFPo5/5F9GUA
CeJQsQa6Lx+1xcGjcObWf+3XFXOFijvq3U6YqGFv5jpx1IVCJ0MVrVBSdWm/EVdQ1QqVqKGMh3WM
BE1Ts5cUvOdul3iTyCcHGe41Txh0pYPHeh2Zj4KeUVtCOoFvdWranDmli9f0N3cVZbkGVmOPi8Rl
PyeUEkKkgwUZEwdTRi9lCzhEkeC9QzcgC0gGCzHwEMPA5I9So3V4lEgmsPQz0iiBJf2VsaGf0WfW
iSBrlrGD2F0bZup4TDsN5rQA85+afmg3OMcw0uKJJMSpMKeyLFFt8DNENi8jmrnoGt8YI/8oxq/Z
Gg31ACcK62qRWhF1U7+WfKEwc0bPyDRUwL16QCKN+o10FPGiNhQOVNiWCvKwUTnLlphk1mG8xinw
+bv7YJkr04QvZylfmEaNNdMS4pZaWEt59/2arVbzLlBbVR5xbwBJp3gDycrQG9Mo+OqHEktDfvqM
jGw+rcNtlehhFLGNrqePf38+gRJcwYbQTZzzrfz/EXwfT9ExF22ULnAUgMkMgMn/Ap9qVCLGq0XT
A6j/EXJueEDfiBuYzVAu4voYWoVgb1elBYXTbm76NGAont/P/TtZR/SkM1l1in7UpuzgOtPncqgl
JWzrB3vLjzvJseQqGGP5ouEdKkjTIQQ1y1XJLGeX1STNveOJtciVjgDiMOF2WbZArbq2f23eodVk
29udrf4i9klI4fw9p4gQgCUNtSX8nqUJothrwpleM7BtW+cJRWu3C8r0SoI7W6ySkicAso+MLTiL
Ig4yaqrfboQUyuEi4imKrTZ8kXqSjfsrahRy9psft2EAmzb9C9HDdCOdJTcedEzj0A6K6YGKVM8R
KgU9T0XqLc8D8pmKWPyxvdVhvtfS1o+LNpPnhGtD4sbKMhEs8nR3//9x1h3anwSxpOBux36Ku5sH
81ZX1/jz41iSDwNOswqvKuEw0IShVNBkd103K0V6ZmtMmvKPnHQPSgz2bQCBdYVhTB2xJfuHe2G2
+6kaCBN0aSEneRhYfMcEOAiMJmpwOjslR5OXeqA9FNelMbjIB8OeAfmQ15/HgJ9af40X93O77dKp
JLIeV4r2TXdpETHk3554cKwtZed/G9jLdcUVaA08ZWnPYA87m2cwUncI6OREr0WdVyXsmVLd9Xtj
JtbbCBGLDkaib9TvHLDcrdGZBI5Z/25DopNE3eFrFCBpyYcdHpppBK7q2MWZSJTONYxSmXEC3uDM
NyIuYWunFFg0CPNCV8awN4IPiJQvBfgQPtF+tRXEAoKfkv7Hu4HlyPrmeY2/S/C5XPXXrGp/aZk6
vQZ9w4VsK3G6JjJzH/jQiy7+eICzB76w0CZcXst0v/yDjp8ext60FVwW1DqDm/ghb3ZV7lAd33pI
9YW2TCmNXUwLsOVQ1cGkX5LeBZymthtGi4zWJN1JNdA+2EDQgZTeP2g7/h1Cnr7n3/he2isC42x+
hpNhctygT/Tl244a0TgACMy5bU4dxFT4b/UUJ4u9Tlb75+4H91i120d8AqQWT9Duo4iFrsm85LNI
jo2En9FfTMgHqzEgNilCufs+yHk9XJiN/gLemjqdps5oaEB4FKczLBwn9oydcg4pk+lxMpzoqdUT
BHzn4/P/3oZUhRrPoKCaXbNCIVInDXXpaF8VWH2ijZ/Fg2Eq2m1EDWuxMaKryQE/4PjigiLTlVr2
xlCgRWdIxM6MFa+3X/ZAuAA9Q9aqa8elZ3RcwqYdsuVTTFRzBXEJ1qHeR/yGKR06m+Ot/y5V3JTZ
vKttVAO/IeJbylClEOrC0H6evQCx1wPpyw8gk+MhxkdE2C0SfLva0IxjFSbBN1ayeRUQHIbFyUCy
1Ydgj2taD/SlgL7SvlOohbtKYKu5DrfJIfkDXfiaiza9SgyL+KrfdG8nJL2iZWiZts9rBavIZvdc
xFwMy9xvBvZb9cAEkYyBxvendyOrseoFRmj2EwzL4crYcexmnyP2KS+8KpSDVDTq8HhbVzyoqlD5
Hy9GrFfsuIkuTtKwsbAZVj6Y3T5CrAvcRQOw/9tPYHkfAgJMse8Mm4gKkOM2WOqBOlPJlsJUdWlN
QXobyjl8l4YUZzlIUULyW5S8tgScfmkolIQ2kzjlW6ZJk33CVWzmU8nWWbPvUK3CBOL8K035QcdM
W9wmXq4YdJMDhAqWu8k9Y+4FsLASq7fhUpiKXXMzUdUeKfQMKjI+Pv9OpO0ysGoq+oWbd9/vUL+E
iTuDCdi8t68EJFR5yuUhyRjfrMlklc2bcSROfAcE5wSt4pvN9rvxuBaIGCqzCKSDiVZdjZAKB06J
TrmF9XKh7G79IpUmA0LIZmX3u+Fxw7y8RF1cu9N1ptxUuSKxHb8BExeID5XzRVL5nKWFDmUiwYVH
BY4lfsPdUJ4UZGNARlIsTR4K7MmmlciRNYiuHhO3aMHk44u/aGFHxSYlB0q1FrfTANE7/mtpWMza
3jev9LUGD+Gr/Rso+CBtB6TP2h/+REoG0fXfSoWTj0MkhngexWYYvXMh7lQQ5WlFTzOBl4yJy2p0
zm5kXyCMc1tL/0NkzfGzslAcJ1GaFotS2xJOG3N+2SPIlGxKOkQhXW/UvhzjrOZ4WXGeWgbwvWr8
K9YT4XNYjiYYh99VRPWR81aweDVHISSLZKLwJHfnSDWURybx4HZ8QQbmBNOfntFtWSOvn7AmAYhF
OxnfLIHmHFOd03SO+zMzC583Mo96+WF+xRVZLE40DudaOa3QgbMkFUoT4ggXdbZqZVzQnL6kXN21
7yu7QOrAe1BuV08TC8fInPMoTQKWc6bABh/FEMxBH7b/CX4y0k7JcOegu1vlnY+VA8FypOrBdwH6
uf3Z2isZLqbSsucdZ6NNyLobxsTNo0IYll1TVyyNi3cOfDt8tmh0d7krPPAZlJhaXKE3lOnwxAZt
gmCjL3Pn82rS0/bvyZMRHCbwfEiAIA6lPKZcO0nGA404PmGGFLgUknYW5vW+ElMypHIGZkIh3W50
oli1eRleAjswYFiIa73Biq/5ZJzEdhD0J5qSmkNWbRtLCaUnjTB6P/nmVr+fT2il2wfKk/1unkp7
y5F/QTi/Cu64ObgoBQ8mNNpLW6FcuOencupQPBeiuh3EerTTljb82jUjeZ7zlk2QY6XfuwAmb66j
1xFjnv3fj0WJHfob83lSIyMbgSv7Kdp1ufX8oV7MLlQj3z06yKQ5eOXxmzus53bI2XSd1Wpnbe8H
5a+Q9X8SucAmGQB6TuCA+ieyoDzk5nfN3s+uCNMDuZ0KEAKayHCxvp0ZvJLEXgm20Y6YnqusHKAx
j1o7O7jvcFazyIvzhiMX/jRk4vMB83rI5jCcsr6O9EkYSJ83NM4Mr8q0ZNiyjpc+Ni3QDodoiE/V
cEHvDRr6T8ZZOGjsMjcSt5Jb0B8NsEph0ZBeCA8ZlChJEmS4qPogLBExjC6gQk2EIwGaZeYtA+h+
OJTdbyuuvR7vdtxvXpyZaKP1piXB4Dzw2E9aCjCDR8FDhSwHWAgURC5vmv27rGNM/PwHQsVUx76I
Eie8xSJd1aY5KnqAzEypRRcfi/ENOCsRehYhHo46hw1d4IVVg921GxsYrNQiANQheLZpij26cDha
GhmyXQf8zKPLinvDsdc2Uu4SymeXUVllJXbSGO9RkplSI6HUoRAOurzhj3IM4pNowHBgU8BXYSjM
ENXJbUzRPWR0kfYUos15MYKQHDHLPqccsSSU/waDwJnRkY1eu0Ps6dh/7+wN49YwYJYRsJdoVPu+
i8JfeXLm9zSdJtiJogMPCiQQ070x2lXYxeKFnY9YDwD66MFodv1EGGVQc5wAQq6Iu2vD8FmyFXWa
/TR+o6M5FskQlcoC4O0lkCY1b9SlznAC5OC55AE7BKPAa2RVQBVkaBjIqmZwxPw+EX0EME2KKAq7
7vBbxPlBLwdey/WFmpjdZAdCry8jEYe//s6sAAT5XVcySrcUB5BPhA8eZHYD6y6fE1m09qwxvhCy
OIVF3fVS5bCdHVStQPcdZJyaaNkx1mkhkuI45T0w8tazVqDX7V/R8sLTk0Hom3fo50K5+WTx6Mak
XqixAc2sG8y/uDjtQZ5HtnHVnurOq65tqpDTGlI7s4JHNJ+7gthJeq2vjBGS1FhF/fi/SfZApHUF
me0k0pmE64bzCGNFMckTsfeo+yANY/1ysfHOTcbRTftVe8n4+DW6tKfVsr0YAal3vEaUaGKhM0nm
Sh7p4OUGbFZft+jKFdoxhxXIY3doGWEsrxqjkamYmbwlL30GRX5iKy4vS0mJYBkrE30AkfcJBP2R
QkNmLYHSj2bSQquHDXaJZ6oNyTMX1wiTsbdnG5FaGOC74tFZ9dfWwjU7Yz/tKGW2WT1SgG1DvmQo
de39CaiO0OnkK0C5TlEVRVhdCVBq/WWe4GBtEj1lYgBi4eHKIRdimaGsXdY2ExpM2E0o4Za2nQzS
fX27T+sX2KgVxKgYGIONQm9+SEDvRLbIpckPB4T7HiLb5pgATPLcf514tICLfxcr+ljoWV7ooAFu
2vKMUAosCTJrmtitlnUgPCo3jX7YpzeCB/uVIgIGNLZbw9EvoeqkS4CMfwbyPE4D5+ioh2fq/UBa
65S63YDxcV4sZW0zV9CyE9CIhFPpeMXWLfy60EWnmLqCGAEhSwBThdPaJ4vZpioWp4qWfUzUgjHb
htUa1LGt55mCX2gP8TK7jXQRh6izE3GlE/s5iP6dHwT9gmNWc+HVRQC6c2dHL+LKB/N9cj9AJtFF
Jts+rDnyVnJyX9ntPJTXd1DDgfeqeT6YXkiQkpaTC6A9mtVjYvKKwz9CZWE8t3MGFJlHisuBP4dZ
3/RoP7g/QBlL2V3PrMLC9yWJhP3WqNNCCNwolHu9Vqdoft1uHv/6AUTb2h28hytGwYdzs4TmpyXg
PN3bQvEcRenicVUmLQVIduTBNXjrr9/bCmzepMS15J7mC5REbRLEI9KBl/mDGARUWVUdTNnftppY
BkqrXaGQhtSPb8l+9t2hKJoKAL3Od9l4yX7IABqTICPJg9sg+p29hPa9/uquHjwHYtwXJLfAzUrj
F27/4NQfI2Msq8NeOvRTNqU3Xsbl1dpYgzCcA11OQAOUEpmGV/iN16LW8dOctD2zd6h6b/h/ACOb
U6wXhu3GqmFAmIujwIZ++jM36mAzV3R0tNfP7Us7Zn/tG6gZxXyh1OHpK0JVlKaUpKh3+XBbucl1
Ms8lt2eOaEIcFacn8cHN9u4gTECtTHx7+JKICnN9e2rOyl7EDp+6o6F2k87kZA+CgvN+osMgwUlw
QPjL9xzpFNazBfrC+pLhIxQyvQVUExMhWnlHrcAtjJ4hdY+PxRlXQ+un26JNK3IHBgRbew1gg64y
EY68elc0Vq+vWeChtunXfBQA6ERkyVTEYf6MvwUnM74A6mWDEHEJ8VvQvRgmP6AGnVaCu8L6po7J
U43h6ef3P69rqQI9aIt/KQjBA6v/j6H5T6i2Fx7Rhgz5OlmIO9wyBzsUEQLYwONg1JtQrbQWsj38
JMTxIwIsoD+PdaaCr4QafW7WZ7+3uqK1qM8EBGSS2qfIYg6ig47xtDc/BCEdCFplaaBnrhwcihkv
czJeJqcaWECpVKaPPXmKWzwq4b3xJyorfjDLdikw11YonQgfPvx2OEVyQMswPZcLg1Eg7xJBuJz3
p6DGlxMf4qeEy6U0REoELzQZbAVfUB6rvMoOfO8LawztAaeot8skOMrvwoHL6YI6QhJInDy/koPm
Nz56uWa/A3o5n7++fPRYC8jk7b07plPWQvz1Xiq7FgX+F6J1p+P81h/WV9L8atss3fy4yVnUhBVV
CZW1JzdCC0d1hLA63zYo9g+DZhU+OAEMxjrs7zew36VvGn9buTFp7CfiQLsg/LYXFOKfmGgWRF7I
ePKaGD0xoiZKA1+EC8ORGmQC68IZYToPlaQGAavx6Fqh7cBjOHU1w2n3+0+hTd/WWVf6Ig6yT/K3
WdLRqNx72zSHgpRxRqusKB2AiGatCONXFeJt9B1HFhHL28oeO5to7/jt2CtmlxtnwHSC5bjCwD6X
VcJMjpZN+Uth6RgnTQr++y8I3Nn2rtdO0xH38UvON27D6ADlT1kVoTUseU+G8v4pqbuJJfN5UoZx
efXV0m4euZgk4nhzDGvFFoyiLtN6V8kotGQMRc0JEHgOH/gYevjovb9BNOotEuK8W2+8i5dxSuVL
wRC8avUtJPe0xS0oQfPYSvTRoCZNtCEODOlswSkA/yApNtyadS2cTCHW08jjGdB7xvtwwR5JFTC2
+DYS7ozYI3wt2QQ21CgeFzBZ4yGtDNRwssbyXWQkHhwRG07FkicEwueOhNBH5suOoaE15XY9g+Y+
X8Bt+ZXQhC1DM1ec8A9uAruDXw0Mr7KGyrgxu2N/Zx4qUrpBtoz5NSBkJzdNhaAYwWMNH8H+Pf2g
w6uydlFW7892OJTUsqcBPeDXaQPlaw0mDRnedSI23cfb21V2Bnm0tj958jXkA1oEWFnfmdTu27RJ
p0vbUJIufqMmnqzCKfNWtzeRGY5sIYcP+9litKjzsRRSpAHg5xDHajuHnYa+fjq6/PizNnwe0djz
ukYP9AAnD0cL7MUFbtSvaTOVQr7i47hyvlOI8+KAdR9GnzQRwxGazVmVkC5Elf0jHhh3usmPvkPS
CaNnV4Px0hnDkfYgJKj524u/Ka9At9zIgw9WB7ldjV1BEe40xDD0gEf/CMgf+OWkhcrfeZZ/FDAv
1z/dKl3V5VPtl2E10JKr/5HB6hB23kRimIwB7nYvNQfNQyvFWuerQIc2CijyHgdN6iLZkdVFDLlM
FZ4G6rswtlWM37Qx9IkVNOGy5OptN7OA4sjB8AYnT2DRrdcmZjgojBtwsAAwxWxRGIcrxNndZOu0
pHVJ4v4SsgbDptq1eeXaSkHmlg5xYIPTAz1YQlaaradiFb9vDOKLV054Byt5QKPbOSmeV3bIR+Mz
zCHX5LHgq+4Vo3tgwZkDA/zn+GPwScWn7jY/2G639+5ovdX0a/T2nyvRcG3/whljrcjAm/SJJ3ZL
UFWgSwwwRrcrKWcBGapnWoeHTNjqUwe+n+8ebw7wxBtbUFysDXrK8OYU5mRbbMpW60Qioap0KVPT
RAD6uZIhRxHv3iWGnp9LBYuc2E2ApMk2+1Vh8KZMSixv4la9bqu/FHgbDuYdMLUMbD/wX7+ZEFjC
W+F/3H+HZ5tQmDu6CLxJ6a5EWJbsJphOikYCXaPeKhqq5rtMsw0Wwa24xfIG3jjKJmrTYd4OaT+5
FkI/MOSihSClrjv10ShdfZ9rtY8fckibXv1uj+6HizhwCcY6wfgZC+3efrl3vVjvBuxO5BszyXl5
JOAlO79VZHfuXo+iNzYAcpkIZ+tswVHu2+SGF2QwwloeTr3bgeBv5CshDYTxikR97jgHRa0wwC57
tZxsPIdDX8Z40IhFjwk7Nu/8Ut5lKCbr5Qnl+M49wZy/bLvIQFp3mt5LQsHNIH9+YpUTOJ4to9N6
ylCvxUbyJjAy5NOdropoTAsFgTvxZ+sE7aOTHX1pushejA2nVHkqXGbbfo12Pa8XTUkecyIaudru
pBmy9OP0pxx0uJcOrgVvsJQUlGlvm2M3UDpzc9FcXFJ4LMVRafJXKX/jurIl6VZN0SUwBptZrw55
5YKTmfowlLYDu+saLy5Nu2j1QljpyxL846zzYsBzI8qCe1GS1plOmuSYXVGVHj/gzs71rEwMJLUa
WJWPWKAGM5V85BdTEnVF2xRdhmAYxRoD/dG+5Y1HO3Lm+9Mfc58uQvaxUjKQaGSG+XDiOGq4ixnq
F7HbbduGm49moossVXutDtdq+3niz5HNfaega9FGIVZG6VwpLRg+1fyNP6b6R0AMkw3nKkFHVNVi
zOcVf8BNyzDSCRxDVhfo6v2j/NJkGl8pWLCB6G/FgQKOfmPphA9qCyt7F2Q5ewv4wobj5zZSRceA
HMp6crt0zPkBGdEmXN4doug7wOv0IJ/AwByeMvE9jc6KlvSgBPV2y4sC+wPMz7pw2yxl7+MOQeeY
SyOCNspT37GHhsgqgQce3BNA6KV+DEXtAhIuBMp0zDwYHQDaO8P+RljzUFRhrOA4ai8nkiuh0U4+
2wRyamtZfSbAhPlu+6H7RYVKTQlJUTUrJ4lKUOTC5+BydLTCdJwUqSUYLnZHvxjGAXM5aiWLWTXr
MdPTslph9E+4AsV4aaIzgMDvybOVJ7VD78q4hQ+pO2InMZGxN7vqQKkM0plZ+08eQDuUjNqoXCo0
lPTkZnR5qxjzAgHZCjhWDPR+gpW3Ehxv/0oIdgFrCQH4fSNjPRTvbUclB8hus0v5Z9K1Nhwbym5D
E+2ntzgAP5aBkrz8lXEH+2sngHnVMjYTwWptp66snNbhKKaw9HcZiqd1LoIorrgmEaFnHwav7ecC
51vweb3l+sheuV1b2EJwd5W+FyYHU5ImecCKBCZlyPPwwFzmibGiBlZUk5X5l9JqMa5CMkDnroi2
qJT457nzrHqf5SXUwf2Ia+7PQO/oKYepxF1Lc0bpG6P/VJhGZIZwwtsQl4SMYjyRA0vfzeBtsrO+
/SsXxbxGBiI/prlCSVLAPv39LyaZdsrkkeOBGRlWIzJiMG2lBIvNJ1EELyEWxLV5SVoBMG1UL3gl
Km8u5tjEVkp+EOgsTBbTEi8hjUDg/Ng7fd/lmGWU0sToholw1CHVuHlhQxf3x5ZXrhrrFTpIgOA+
Ia7hk/jCC993v3LJlRWrukFcWjYeWOW4g1xh7GPurNy2gb55rdrM94D+9I7CAcdgl6PmalQF8AIj
4CIt3d71sKX2vN58I2Af4R+Z41qtdj5IcI+fjP2jF7onz8FOeIhC6d9ESQTBrAMIpaGOHPe3XjIh
sGtKuOuHabrIKmjSw7N2+jOrrNikQ45h7doIlXOfjP8FfJVRM3P3iILCcpR4bmKhIV/3A6lZPqVD
hrLmjkTrNk+aHi0xKTQMd0iCwMBqxBRzYxs2HPfVCOFILeub/r06Ic52jiuBOl8cGMOIcjD1bhkW
6SQXrlRDm/Q7AtFctYm13pS97kR05v+EBeaDPBi5EcyNTZfRAyafnHVn4mfKDixLPHZHO7dvLVKP
LIndrnjPR2NbRHRES3hUV8BAri6/UkYTbx2O99FnKe1L/f0o9WfOCdcQRPyrHe7lHjq39jZM5u61
Fq5IXw15aI8sj/lUraaTxEhYGMX9H6QAbCDEWqedidK4WvuXz5Q1nojYSZ3YDBVMLKQuphIpkUZ6
iiCHSHfVpLAf07mtZWD+Q/teSQEn/I7bew1e2+SFDBHDtC9r/HJTJtf3I8EYcg0LNsJJjra1hl0/
7oVvhZWXhQJiJ89j+JWCPIjyGCDlED7H7HqF/DZKcJkziK7VOv91YuWjT94oD9EwCNx3BSP2yGJ/
n0f0dnqj1qxbWZRu20/LaLvxilsLT+S0bHq6Y6QS4qlHguU+iWRHFsT4xXDCjkFNihhftW2soEHE
fzPIKxGsz25EK/c3HkCidM9Oz/rexahllf88BSC+uVclozpjWjDNYJZ5RYpeOuo81ecIKT3CvHNx
HYIoz1z3H2YMfVIl46ZpTqxgx8MW4OSLFc6on83/4APxWmtrCW67YxMk39z8K8OrKvbzqR0LSG73
hAGxjzylUuOmRo8GZcZClLo/24/zOqbAN7PFGtfUgvJLGlkURT7iQCzMpsGT1pARV5n2/v/qFuUK
9i7qsfSQRs3x/0vy57TY4Of0JWIrV8bQlXlWsdgJckW/bIeWdl5fwBwzSWYe1+82ug6C07F3w7Wh
sWBKgrLI2FJHxjx38OsUjDu9ywZUXZoXULJmMRCmYc79feJHT9EWAO84AnBrBS37Inhpnjt9XOvd
I2HqhFkdKhGwUiWN4XT7L0gGq3jFX9FupLdgySlGq59en332oi/KKRCwkIeFUd5EF9wBXIqgTvOJ
TWcEseAJHdKwUzmCy8JNgu3ZIK/fNOxQ0wOQXEsSPGQslnPYBNI4yhNyg6N18pDwzjemx8FBo4LX
I1ccG7KVKMZtiGl2i3+Pf12ozU3WhQub70h7n1MN77EdjdZoz6kpJAVWvvP/iRV9EKJ2mBLXtVpR
OKrt3koS1t2I9B2nqT9O4A1y/l/XqNjOf5jDlQxbiRZune/tTzSFjxhEFXO4zPz1JGrdslx/++f0
3lSLu5emSTfHN+altvTq8Tct9RYcOU976zaB8OIIv+/AMAoTgtTTEZUuXcZY9KRikeZz+cXAQIRK
Vz5ibx3IyUlzKvsF3wtVzstbczFrFMIXDILezMY84+q1C3FP9qq+ZW2dmiBybqhcL9Ippt7giA3e
4rsVKmc0e7W7lhbf9/uAkgbR7q9WLD415y1XaXGtsjkXk4pICk+MMFKKjhJ5N2WYywsCT5wiKU5m
cuJi5oipVhvh+B093i8GoJoKe1EyVVi3C//8xIKoCSVUQsgUOBhfmIn70+Hh3wtTmOgW6nL/56Vn
TPwn8DNRwdWU06kGjBgAJHD4qhKUfIKSVj+MLM7bfL2ZC8ijtc3tIc0h5KJCF8WBLgk2BOTz6ICr
2HmxvJ3+x/XNbPIbs4bg1zrVxtJmfR5zPpCQnQwVOdFOdV0GBloE1VYnzyIe5PRC10wcenqq99FV
nUzQbmKS4de4v7q4UNcGa+ctSYiMiIgTt4E16KxRMho8MFoq+YI6djOo+Npjxbs8s+/ST+CTGt7E
IxJUnTQDOmsDMM2uu8K+KAF0jIo+2uA/lcFQv3ezdR9dcQA5Abpl6KUx1FhGkqEJOSAgWl2RAYal
t52tnHLur+Wj7zgybzU1R/6LVW7GNU/wsvQQr4FAhrpgrHcnOk58EB34VLCyUVsY3SDIkrTyIGh/
S2NnPDQvHEmkFfeBmWk2rWOnVrXLcWfHASFfQdfhv/U/6/MQahdBIUHp6DNKVgYEo56MxYvavXEU
PaC5l7KwW8r3aa95UCMGia38H3mMjcqUjYWNdKDbMyFSv57m3IOuwDVILiGjfduZ0BBxNOZGF0gy
cwFrc90ndHM0HHvbE0Pgl9gyErsD7eq/nDeVajS+9u1CK0Mc6k9Es+ykRxD36BWpfQfGMuttn9UF
8/rR3NGbAL/Vw/bV8fo62vSC7It2T4qAZ76t+4/TqoEeC+7KktNTFX89x8A6jL6OkPNkaW+QyicJ
RMX70byK0O5aBCj0iiLv17wIiVUGoNy2RggtKXM2Z8WMOIhy3fCUhXtmwrT5fl373YgawRX7bJt/
A3blgyhyH+nTcRQ+7+mZt/XYbnnKDaFWQTV6wHane7EJq83Z4huJX0X99SCPADQzHjesUw9ON5Uf
YNDOYBv8l5/2hJ/d/KnC9erNxCpMALxu4h5P1BKJymApbucudjssrEsFkYVSIPsGe1R/EsTD1RVa
NQA2h5Jyckr19sUlr3j6nJwh1S0X6KyVQT5HEWtx1LHz8FDTfzmimpbMADykRxbcof8PAB/OY8LC
7AYje9ix+IKQ+27VW6vHxRdlpvP4vACHNoJVV/dmQMxPnK1awTuomVZIfU97KWJ2UnmTXYz61oSw
sNl9+t0G+dl5qJ+bBmPvndDtHcIldv9cvZsdd6XmYQDRPCQl/H5tM+DJ8WK/mylo8oKZ7dGV3FrS
Xf6nYsaxUY74IqnBvH6PS468U2PkO887ROj+6mMSHJigSn4BnqtBgYwqAsfa0iab9jd8bG5qw99c
vOLUzZLzWQ0Ckc22vvapGOHlZUHG0tXZmyN3qEQifaXpZM0MHp/VLibFg97sorSiwPRvW/Xr+a3R
zEo7krjpAfk/bvJbZRLxS1oBakd/aQxdG8mlI/K7vV/VNOVpwJl2/aAq2v5Zn2B9PuVrLkkRg2xd
2wBhOHxi7PBaBFR/+6jFjTvFwAtxdPS2lWK80Z4OUAc5mRCkPPIuj4PbnfRp6THaqyle4sJKUEXU
XBimkBraQzdoA3I5SuZfwywy19nmc+8TTT8DfvodyGoy0DCb/L4GxYd9jZalTxVr1nUSqnwKXZ6P
1cClWVTkPcIN/d9lL0aiQAplkNce4vIKUFh+eVR7+39zaguRuzMcHkhgM2a7ieahfNvNoKH8zyJw
Pwu1p369WqAF4DJ0omtwQEmflOvG4UXkT5sruKrKUxY+qJEc6lkQSxm6BCV2Vv2De+wj+/gWZcMt
EuhSr6SD2IZ2pwXXDzSPkqSkyF6Xu01JG7+46JiZIbsgMI4muTf89EsOOyNtOb0j/6AcH2Vfid4n
asauLY7xWL/1Z+mNvSWZZJ0gQ/OAVqbfSXz695NofY+cVibN74V1SEHPGbbJT/Z4ZhKahhlQZFTW
sYHBk1npFbzNZZnQtmZek+P4YpMYVQ7Hip/I7cfOpgzz9uCzcQRcnFo7qFngpGVxMv/shYDYCzKy
dXZ1x3Zot5RGf4AwMl2aOPBNhIbpein78hqqkhSeNdeYGapRy58xtdp6N9ZQk0Gj4vpVg0F64eTl
viMaygSdbiZPyqE97kRFsqMifTs6guJhq28TB7ptKKKMQuNyuX2bS/uuCr+zglzo5RvNiH8ZcPfM
3hvjLIeEWtOd+s+x2FXRhv+WhzSvcfrbbR3qDHwsW7rKkcEca99NDH/vfTf4oEWKz9O7tuyIm0qx
rw438l6xTjTrqVcJNEJk1jmk4zYc/G+t0BonS8D/8ORClBUQY+127YOvgskwc0oqhTUAn0RaW4A/
oW38Ojjz/5Rl5DybuFRGMvzOkdeO+wklkCliDQOet3mqqh0LAZwkljOXXVPWYWBn1+ru3L70VPSv
DHUeIgzKyQfW6CD6hB9golwIq7SO2asH6quO3uzAMnSUZy0FQVk+HYD1fWFunH3XRV99aTXCTu/F
zfF0bj0bljTqbuXbecj8pxsC96HLo7i31RrKQx745O+TOXycSyu7Xi/2/+Uwa7IoDNOwb6T03NvP
O1hO8aXAep6e+UsNu3RHystzneU9c+jhK0UZGdW9g8pI/lHgq0UyKgCiDAcmnor0xDutnNHs5Rlg
4JaPf/Oy7ZB55gfw4o22OBd9yT1qwBulPznjS0dylrKbi1t/5RwjF7CdFaywLp1DVlt4TlEZBNdQ
uNVCzqtvFQWy0cU7qu13vA6w5tI9OCvWtmenFE2f2kgxvRaG51wSkZH9d8MlGgo3wjDglPJR1rev
HQd43zAAUoNJonPAZ5ciwQEkw889M+ufqY8gDTUedQuTREqPP1T+0tkAV4oyI9gEF7r5gqV5kkQV
Rhv3gs1HlohfY50H5jNvRmNV8so8Fb9BtY2joHAnM7vakd7DUqNfIcaOLhCGGx4ZdJ18R92N54Ov
PE3OsYxQjN6CAIWhJlGyZJMc/rbPpWLtbhFtpRUTl0uivo+kpISXhbPNXhRoa6oiVHsSupZuRNcv
j45Ed3vBvypuUTrMwqpy5KFHGk5T0d1FqAG6DMpZHB2mOJyrVDUwcgjw2PRAo+LL5nbFBL/RDRpq
8aCa2rAtd6nTUPwqrJEVkFeumUOPE7BVSTzuKcL9YcM445MKGlLlpkARMgzHh5hgvjUDnbDetQPP
lsAEi3DKk0L/3DAQ0iK8LDxYOvIxAzXtj6J0vTIjCHPGrTDQzSPkvEAEjF4HnEGiZM6WLnnmkM/O
4NpJZDTcG9VgwYsn99eh6Kc8Mlr8s3J444U5dxN+jdpwV3COJfAB6ClmYAIFyyLeHwycVmLC4uNZ
H/APncnEVXN/i1zbyTTcoJV6dIgWjrCcYagXLfm9SLAwMJhvjg+HDDFK5FErsEZhKZ3LaBQ4sddd
eBKjuf+rSP8gXQmrXV7gFm385nn+uNldsBM6PhgMjZgCtqh3ugrEvmW8hdwptWrU577rvLuSUTCF
Hnvdf+vgPQlOI43GQ9sKgoUVlcoq7bn8zi8wKNlFKa0la8fwAP1k7qHHc1ffONjzrI5qXkjoOTf1
DWsjfwEKuQ9a5ols9DqDpuU2X/w7VKd/eb5yPtNDDLV7yz64WhBoPRa+ESAGo+7nvuTISztg3vc0
kF1N897DVCMM9i9LrvDofXFRQquRe4lT2QV2Ck1I/ThkfThmXLwsR8n3/EjH4V79+v5o0pbbk6EO
UQfHKuUPsfYvpDIpYhPA7Kq3CGIdIs0PkCIWnghviUsBnvgHfXAtiGztQNC5JKFAs8QEkHRwvgBd
liwg+kwEQO1JWbd3xUOUXGTWXr8dY4bo2/W6+43u6RcBT8VlSimrq771G7OvslqwsUdLiuNqSlXV
y5FJdHVsQJvYUhlpSoHwb8ZL+IUORHOLwP+Kr3jhg+d2iOLVVyJkhINMip2Afo3jrURZkUaremU+
Im8o3hgBWhkZ2R8oGx5V9VVJlCsGMQDaRY3ylrwsbFiQTgMQw0CY+EgYRrUPjGMtNoReV50XsCvK
t98DE2rf8Q07O2u6eti6IwQzX7WT1aY0QYU2AIwziEfKcBgGJ6WeCmebQQnqFOsQJOCmvsrMiLCM
pEFWB5J1OWHyxdZx0XnnynA3mWK7kaZxYonwApZ4ZZdniul0boJ8FGawV1PjvTiiszWzK854z+pX
4mJzOxBusaOY55TKRriEEGv54IJgx0jmd1mA3jvgsk2Tqyvvdpy82+bOzLgWCWMHpUeaVr5KUEAP
1RHbA6Fjbej0SOaD/ghFYZJhHEJ0yODgY8yUU64/aXtRxYzoUeddIzuoAyCdi7sEESMu3LEKzsRy
yrIlAlxuecPBvIZgB/+WtToxAph+x4cgOZMlKvkjzvLxvr3NxDRrjM+0CYPBpDMrgSDOOCiGkIl1
zArL4Wp5vXcioZjH00AbzMeRKl97bA05dwxafLHEJ6nicDmdodduIfJRmMNgZ7GJpK+tCEIJBd1X
u7JQlMwDOEvxrRD9tIx2QClcgwpJnXUcTlZ4DvWJZ/XLTPwaAq/JDP3Z/2Ria46+X9bizkdly7ao
fE9YulN6pcr+ZOZg6LsUGIHRqSVvJHBbrT30lE9SZm7HzwAQ/ZvRVLX8Wz2SoP8TzhfQkZg7dwnQ
7xPMG1w+x2gkBVLqSnVmLQa0Mp/IdI1SZ6R5qO8fHMc46FcuVmAqH0Y7xJI3qXKKGTANwVW/miK8
Kj33J/QuLYud6aCNTSL1QRU3JV5TvgKC7B+HIsgkCAUAAQhSiYWGEY2nINWFS1m/3HTeBxMsVrf4
V8B3HZ83WMarEjL15OXE+t2w2MGOQrkVJmRH8RLNMVJjRqDEmR80yXnx/7DV1NZmhzZLXm4CW5AJ
4J8BGDwXuKhuvyNJqNd3uSAIIaU6j2a7FN0+W5RezTeUXdEWhf7Ks6iUqnVGIXO2N7VpyTIAcqMs
bMUu4ZxGXv79qrX/rgzoFz7xkMP5VXE5OwXo4V0MYZnnlnbN9oL7AtxWvib3AP4ByHX977yfb4lS
a/R+cz3BY0kR4MmPIOPPebj0q+zODJ+1A4OirAhtReLL4DKngVkiWvLSPl4XYLcySH0VA4jvcNrB
iiKV4qI5wCvu+O9tM/nhJNqyiRfU8bPBaUlLYI76HeNXCrP4zma7qH7nBn2mqh2lfrBLYtD1xapy
LyfJQUJcDrb/61z5gwsdcUVIfi9br3IjNDu7Qn0QAXoYExBgskBnSdCUYDftcXAb9L+O1J0aQBXm
dVBWnrfEz5tTVoCWNFB7A+k/k7B7yddpNIB1Eqq10rID8fr87o8kQcoUi+5uezKsAQ5LciWdZ5jh
UPwsdmPilnyn9k0ROxV4aTUPq/PLKNBr5Gzqbqg/zadGT6N/1K5oDsANyaH0YPxY5jAKbXrzCmmf
xumUwWHTsKEquGW0mMpGkj+i9CQC1JPp2XM45dTqwyw5V9TzOiUJ7e5xr6yTKgifA3CMEDy1jWx+
3iI/b/wAQipnqkbrUp2H/P3ibA3Vl5K09Tgil3G38FAKLgOvVeSbS7KCAdxaHg94MRzqFgjCiEz/
jv4wMjVUoN8FxEVzsenb0AjUH8ENu4ANSVHgf8swNk3Y8+049Qp2dDuV1QuP4q3P89CrGwSlH6Fr
bAnQbe/c1lv54j+hfkGy2SAgu6sZgJ4G+ZJ3aQvdT+XZUdH9RvCVRlWfFzeYvIu6GHqTzce4N7D1
Vs63jf3M0Z5SHFfwxAZOqdWIf9dmQgmc+YPCgll8uczrQSZw6u3W3e3WgbjCu1UUbWYFQuKYlzhy
8F2VadrqdrfZMZGvmuJUkmRc2iHPdMaXg6Xqy587jTp7moI3E9jEg3XmGmuUc81cBf+es3omOB9D
EAGWX0AH6TnLBZMihZ3ifKz+IAB9+0jXtyF3i1pUxuWp/kyff7QSWPDm3ALvJgFKvfnToaFwft+t
o+MgGb6rdjJUNnhaF6ZkSSoI/z11k11uxBQKhi3ByIgslaz7OI2kshTQZuX+bA2zeoiCOrvJNYQM
ZWsB4GeG+7gNfG5V/PYrXgS0EJjbnLxWR+yjCqVoumvSu+WrSHdkRSgXx8+iN/fka/t4LCCxtNl5
jQFbdjZUGMKXZbk6trZdxlRSdv9pq05cBNyPQIwlD9UWKCh3Au0Apyjf1UfKuNoD8LrlW/u0rhQm
44RfdKgb/YopMxdeGZfQslnbM23m2PzOpFRWPgr8JPAfrZebpWunrQduvz9d/WXWneXufOR5y6Gj
Mnjy5XYhQFI59o+lE5A5lap/x3LZeTqLJ7ZMD2bThXURXufHhLXZPrpKJbCpAg5DUcb5CUHVvN8/
GYrhmvi9w5mzYAKUNRv19CnUrYVKVo+p6ebEuEl/7U6kvueF5+unAEJdlZYHVGIJYmzqM/Bycmep
Wk1T5QMf6sJj8FTXMl2rBeCBbMEes5kEbTEjBPsVjYrSj7ZWOVLqeR8Vp4gIAxSndEeG2BPdnSAq
B4tE7SJ27fCbC9ED+Sgklvt2QzhtBWCfFZ1Z2L8KlMmnE5LgM+i6xlIbG7OHQ+a/zsaq95CsoOCV
/EBiADMF7F7Qp1HyPAR0Nk/ZhOMcR5jPOa+5ZoUrHyPUqi4ASgYhwj44QBiH4QY8FfAHfVdyHUcQ
GJFjwR87EEug2ET7YbwRIjOz8H+D+wCt4+7p0NMVu8DEK+SvoXi5rCqCcVF4chjJN+IcxKO/RLn1
uWIfnU5+ADOcEdlqw2zlkgLi2bjD95BYIV8EtZU8UGlbtPrccmfU59N+jr5Qw6/sxAsC9WatXIRu
s+2WhaTmcewEat5dfFxW22W63Ht9CFsNOOYUnTXTpPbJxV401KYBAyg2XLbUobs7f44fK1vX18Lp
WeT0MQVcelUpHh8wYUWIC+T3e76a6fcbxU4In0dvEWOlDAftQWEUKbZ4aBlQy0gL0hF5NLH573jS
JC/l3l01aZsJ0HjvotzVi+SeKjZMbQB3HRQArkf9k4VcqihYI38AVOfIaUHfA+A2EHTeNe1zKkKZ
oYaaZiI3DJScrdkWkAXFKaVzFahIwtNWan0y4a8O+SLIGVELqJ+QIcD4HlLy9dWtdZhh9bCpkX3r
EuBlFinFeu63ikoEaneJp5QLJS+E6hTC8+Cm5Y9Wds1YegQL9o9ajRlSL7+YiTvDWZYRkDEPqNUK
beksgfboc9bffeaW12I6JcsX0TRr1y4M2umMSdwEq62jBNw2Bl6j/bz2PQz2bSj1+9M+DiwUzq32
lqSyhzFcSAYCkxSShu/Fc3gNh9dkmF2+gRRZ/iXEPxtCbowOBSwMZqB8ZiMK0rELUszkV76rTxd3
Lcgfx0zMJ4qa62v0Jv2oQdP73cAD6+BAtaEAk7M1t5GV9mq6rAoEnb7bbGTWd042khtsP/G7MR5w
kgTZs4U1Wf9U3iCl1mGKQZIBH+401UTK91JzlNjB+QcMXZXDevB+hAGmYfyIiceiqJwjxbnAxYMP
8EOGTMmDSYti5gx0xCLi+3YmJpzHLskdBtRzi2p/H0oBxjSBqGOOlCojezyUSPDOGjb+hxPahhDP
J0UiiEfX7TiDy9/D/tfw1oyit4Ie6EVesdRnmpspEx39OohY1BpK06LF5VIvLqmIh1VWJLWJyI2q
U4zp5x1/hiLKY58wyZ9hsvmLZkmLa4MEpTpaVNKnVyJIMidJNsTt6PFE7f+jbPVcFlpsTsAzjJ+s
mUAwK18foGNPU8DcrYNA/3lEzrAYa8uf1+kFzvqz5bJn4uCT/HE7yLww7PNT6FBaoyXcA0AkQerx
DiN5etS/P9/ED+G1g8rDoZrkfnYtsCqHAI3mOyGAez70ptanWayKYF+00hWhd1GCNJW5ez0+jJ7x
abCr31xO+7aGgdGL/2OAkNCpzpv9sDL+bRsOh23bIN6GOSogvxOKGHpnF1d9ziWH98uboBbHxeLh
PnCktnmOsLMe1kY7jS7/HQC2hA5HeQFmVmMDAkh9grgzmDk+lDcLC4X5o84Q4KQBPz0M2T/fuAAv
BkM7FNgAyad+nriH+Dk2dKW0Zj2Py9R+beKvsuQweVkE8wlBM6nCgFNqPjqHBdWObtI229lI8Pve
mqW8vQIx0pUoPI7dZA6RbUqaNfQKQEJ9w4Bg8QMCGlRxiNTn4dg5e2sbbuglJKjt3+p5okAzUkel
MBvYgjmt02YXPoWjvzfTALFe96UR5pyuvjPRJKI/aYQhCUgoKnfVTYAPK/9cxKikrqKCnjjGgH1Z
9wlT+m815bEloxTgLDMA45A7cDsNxaWelrZH28UOz/V4YhH/Skm31hk5lXw1ZpJ5loirjiPKOWyN
Rkl5qaWoSIAiYv7kQ/JymUiDp5vGLfbd4W88p0aqia088/oa95qTh7MV5Y4/pYoXJe8ZxNow+hbT
aNd7EmQP3p+GhjvMlBgm/EH103syTKGBlSY1WuKf2eQsqx8Bse4Ks9g3IfMbQ1WJgurYktzrB64Z
L+zIvPWGLslsanNRwBsOT/FHTgLd9YDKpHw59uccM89OKwbFWTLZQa0g9wQRnk05/pZJsp1gqPSJ
rAAuAmXUB5RAeYeIiZHeUPqy4YXQY/5PTIRJVIEFcImVJGvAlhIkKGaVFZu9ulw/obyNoGyrBSHW
0uIfWnCho5OuXeTtnfLXUjD56mBCuj9+6PDCt2OaMlEIWPxEnPsQSbR3vT2hRuTp7EOtcMo4TOh+
pJe5oUGMT87AX8TN9pIj5m0geAuviRYOThvHoTr9SiH+BTg6DFgg7w9l7j8vvvIXW1aCvlsvpcQn
6Z7Bw7R2u8RhplZjVmL824sIhlVR7sQehLeSNubPe39+bkkP/qY+2DbbmfCbuiYAqdt7X7rh4f3x
uIf/fFEO8q95WTVF4uvh6IErWWGRdM7Enml4d3hG/Id5BTVuBI9g9kho8oTny6R4GlMBnjh3MSpM
itVnMKv2Rs/O3NcdlAVJUvc88GSfIG4Tl7bFM3Hi/DFsQSZM9oT4mtWRijbFJJs8JjYEhZtp0s/D
D6YEz1fToU4R7ROTAjYUKXVjjf9VfLNXUIbYrcIIbie4YCVKnw0O+obbPH0UXDMRZr8NgMgMDHKA
P6w0Uj8jnVHWUcH22XklfsAR19kjIWvtzptvvrx1QKnncW3zlS0/tVdIwvFOLYJfWz6TQoCKNzOP
P77E5uFz6mNHvk+0yx84ySnakDMWvphba9VmxcDfRteS1Bpx9vZ7LHbCPk4rIe9/JUiUCQyt76CY
SOdZCHygOSwAdGzone5+l2f18G8kNEqwy0FresC5ARMEwF25dRdSs9DzTuWR3ZKKZJcFkUBkfCSm
9umH8akkvlj1w5sl79SwdTMYzGfSUvDAHIFFUgZzGXJgEeL9T9MbkB2S4ifOuxHl/d5jCD5PI+xC
2ZNTPnQbxN7mZ72cgE9kQqyy4LvGq2LuNlbF6FWVvFw9UCcCyUHRSrCvJAJHt+30j31zTxLvDEf1
3T6dW+aGwBozQRNEubhfwhVfF4wpiR02haYKhJRvEtAPQ+qsFmS2aiKSiO+fyMKF3UIOvf/YoA/i
U6tim9CAzNEUfDSU6PBD4boYm1kDSmeOy2rb76TR2FeUXkKZTkmGszJuw9N7po+ssgM4RuOBYAMW
uXDnMJMxJylJIixWuIdiP8YkxZd36Oy3p7AzBx86gHL4us5EgDf2iyRykqsYz6uQbE2Jk4IcZ7jy
xklIgvowo8ITZMdcK2r6z+fUxQ5Mro8+1R47FyIdBYAHPgcsPaavZdJ4vypQ3Bc/XisPY8br5ERr
f5lTPEqE0vh2CTebHepko446GZtNvsjJ1dIRBp5wJk8m6a5ynfZLoYQ42+1QPakwCksLwq1woSb+
bf/Qi2Cbn4WsCVBKc+hKw60KETToVj4vKFlMBBhPgxUMgg4Dzc0VneDRHNacGii7db/EOtkOa7OA
Sg1LIRgXzQjHnRNgref9daxwJBfoXJQIuLN27G6jXkrlVH2Yq/QDUfJomSlhRnmvM16LllpgkibL
p41+2b4Ro9BKNd9l8EbFTi5qcgTZb7r6K+QSluZQ5kk1LAp4+Qz8WKAeE+AG32+gwl5GPFPHomgm
xi1fWhVjY6vo5AZXdxhlbfHPNTcHHnZGPHa5diWvYUdpgz4sMUrl/VsN/F/HhMmV9A9TjrmY9wCd
kUj3kP1mvMgywps+Dzp6enApMgd02rKz2tKTvLLkfcofUT9V2cCt59ws9pRZZsmanbW8QZ4/Vge5
Y8DTu3KX2cBEUKbTKpSqffUNK9VFinqYbpsysMlZAFKN4rGuJvVLeySYDxuXFdojDI/J57LVZLcX
uIkJVtIst8LoNLcijVsB49138gc9//2Nhi3UUgx0A1HeM5fbX1EceB7NGwLiiZ9JmY59Jou6DPk4
0ykzjImH5GYBGbn8ogjuXXiI6V/V3mpUT3+qI4HO7AtZkRolzZMy1TM0Oe56fYjZL3QRaDlF4zbS
t0pIdKxoc2DfLnQKxFMdMp3IbzZ6HxMTbjP60clZ9kueRxvRnI2naEY6tbncr5bXcQixtHGTij3R
MhIb4jKNoptisLPRGn2xDjHvjbxQTLLTsP2bv8RZaUOwySXfArjpo/img06qPTdAORPk8iW5GTAv
9G+32ZA8v2C8Ni8x3bYvkQM7F6fLn7DQVRwHF8W3JxQAUGjrYmGfLrv1zhBwXrv/tfixKyvBu57J
633sBNP0cjDnuuTZvAI1OtKVKHPciuUj6EkKxxnFHRAbA7GMj2n4GXLqnqC3Ggc61C6Ugxv8+zbJ
DWN6bbncofoiSea7AVan2SlCm32AFeHNWi1GHfTEEFPUgIOp/fiC9NPxpKC56Cczh40DNiqXbL0m
VnJxncs5rbSoa13hOjA/9xYxTQEd7vwLjgySH3Suo1GuFKmCCUezEPYf37S7mNIyaPIkPaBigMla
veSU5PeZZdpTUVmGNqHBhwhk57hTkbjiJZ/QFsB2LQYArcSjHLdGuJf1dSoQnKjBblxXmoCwFZ+p
hzv9vFZ78fiDLrxRbLkt6B/3TgINzWHaEu1xwBj3elAUlzjIfXJSQQeT5zqs5rIfWlyy90aca9Hs
CEDl5uB3agLTo1OXTq8aFOONslWbyl5voOcVsJ2jlE0J6g2xljZTCZfGHArB5IxflhzvZGsyCbqk
bCDqeud1sYUMPE1Nm/sbN4RrYvPsvPfQj9JTXLJjKMte4n20E8q/lrZOCJ3pPB6vTz06ZN1MVDwa
904yFczexOWituu97t/RcSRFRn792qbu0R+1SETnbWHSmlRgUx0ELVO6hSqAdh34C2+WykTrOBzJ
oRCC8Jy47b+CcnujdbBOUyd7SbqzBM+Esmxn6bsIQc30y2/C403MubcN7n9Ed1xPHk2LhF540pZv
4EX/phj7Mr1QA/I6bvhm3bi5UR7hqbkasSxwAxFWuhFJd46mYIey+5/te6p4HlMAaCnWD94VKDAa
/QJWQk7u6qLNfsLPSW/bUWt043fM7onhy3U5D0so0d7iQJVAJmC7/gruqKqIflj9z7w6gwULk8ro
X0cj1EjlrvP51IrMGG07djJT9XVorvxdM8YWcKTaEZsksj+1rLd1A6+/5m29wb7uJiiVmj2u/ofM
UYyKXsxY76o9qyX68MVHA8sNnjNrGRi0YgCf7xCj5eymPhJ0wlx2PfsyqvWcnaaT5eBdZ6Jl910J
uwYf9DbI047QQskLxNKRXMlrlpUj1fYAYk6hbZ6f0q5TzoxfsaAPQNkl0zfShQV1oAmKGUMOTz6W
WzVgDkj60LT63q61/Jr6sFE8U8nuEF11+jURvVnSnW15PrommwPylJp/1BKv/acWvMJ0IVcNgg2i
q8gAmcUXd4UV23C+rHy8weNghXvcn11piX3M7GXZ57tw1pVkGUdcx6AS8MB7s5BO51VsBJJNgoWr
5qUIlkztOmEcV9zRZDP0ZFbw1gdf3J8UxzBQvYJJq1q6LxaW5gcmcaaVlYOHlo+whEnL+Bthr/X3
UIOlCgYK7PothK7e6p1EW4AXOrwY3BE+5wqtxYGtzc5IKOes33mvHFGGMvbaTNG0K/nPk0NkzKpG
d1Z44qPhkb6qEb0TbrnDC2itkE14zxrdJKoy7+27OtsdUrFcXZjatFZNEMbDu4wDnxCvK+WI2Ndz
dRqVV0QlfbHwc+fzf5bGVgjBsqxm4gD/qCuqaBu9rh0IUUSCzoxv0PxtSN61yugLgFbIFlntHimD
JODOnAc+wM+7vpBv+cPuw5Tq+ukkNxC/Zx9cwTGhBBu8jTR1uZNS7ASuHvCCeE0XzNvRoeIgdy2c
Ct5noSHUfYusJjZHlpFZI+/Qo6LTihwYLAYja5nAlPBZ2b7YogzCsbv44uxzcKj8yiVVi0Fi8s+2
OusdWQmGB80mZeO1XN7NOHmwEQ0NGQyMcormtEeKCE0gG7AJXaHgmZIWUJOQP1puB98aXoAZ561C
lj/Dl136qFypFal6h2858Ew+nnv4L3TSLglfuQWYQJ9SlBx53U0ZhXxWUwb3D1rtNrtcGosdnvdb
yaTuMhNRUVNcL4r3pc1i7sb8x/I+9cf7ojNcJSPbG/LXSKA5I5C+B6u0fyIf+RaMg3yVgnWWXOS4
0pdUPDKg/XUV3ih88X3cOJ6j2Xc17D7jUqy/hAQPahBb+DRAm84FUTa1g8kfqFTKwXOnjG8eN+h/
D/H4HeklTGe/oYvUnqFwgXBxQEI2qnW9RDd5wdM3e8e657kHLFXSDYgAWrHuH8vtcnsr1NeTTh+8
jmKlX4Og+dm650RgQDsa3xaK8CHtE8fFOYOAsEfNJgfb3RiSBGRYmQKFgz6PbX2ywpA0FhwYXEt7
OjKIf2T8G15iTDz9jnJnu8qy6klrtDvKMvfn6Yt3tAs3BQVPWoYHJoAy2YAmWJzCmT+4fVG+2t9t
vLbYVNbC8ezWaDca77qrZmX8WwKmxmCTtY/H5dhnGhZDpp79C7Digv6/1RLj2xmLt+AnY8E0nS8C
gwQlgDOHrVPUM8cAXrsj14zVxV18FlHVRP3QBWv/U6kl4fzKczrkQ+DI6ri2u1N+5FSzGHYsORz2
+T7Ed/al0dbTXkfHrUUv0nKUHy7W3NwE3ExObMvvL/yiIe8FNcTGIpC5fzL+rKJmmZ3i0+JYPik4
yiyK6qKOxZA7CKaEvBPhmmuN7xaJOaQEhy8Yx7LBdB3NG22K0aKK+VNaYEQD8sjwKDoeH+KodAhQ
N8jUpEBigEPtnkAtTOSTdaXA5sIvOSMo7uDGowpOz66FiVo5Lapv8JKp/vPU7fiskjd+HQuE8W/i
yuqKnSlErzoXcEB1IvYMlkop/QQ17AYJ/Xqs9QMtGEgXRl+LwaTA8pD67Ra/SBU6se1kUN6HbWuw
2327gQtid35mMBG2dOq88LvmYiTmltICswMtYo2qIzJ96OdyAL+deXaE8f2v+7VbcrO3W9+tqzGX
8CD1j4mi3e9r99mDafhY1AXYb52ZDAtOIlBU1df6tD4B8J1VpHMwEcF16Qt8q4afPk9vJ4j+8aFe
3BeJrjrTYBQa/rkzwT6mYZBI/cg0mWEq7uYroiW3iTYi4HAcZKKb5GQzJnvartWuepavHSA7mXGA
+pzdogexTIK8nHsvX7Qek9VyJwLkHr4z3xfbMb/E6RhR4vZ4W3O6XpppLz2Jke3dHJwyUzZz0Df1
xvwemhUnTpg5IYcrvWJXb7rBqlEfI2pbjJ6vOarUYRoGgfKHNTM6GivZnAcFlOnwXJI6GPwiJ0D/
sgvhnysDCK9RrczmuwkhMf0qIkJt1rZ7NKbJ62qvpoRZcyZYbOz4npqTWze6wZOi8oTLVx1c
`protect end_protected
