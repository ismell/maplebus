`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Zv2Hd4g9AlOUWNT0BfhzHBMEWHoqPF2fnLmeI6LnbAHXElIF5FlcuuWoA+A5ku715GjIsik+aFg1
18/R6u212A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lh0Kpqb55zsN+U0q46rGqvJJvdX8NRcCVyfRm2Y8gB9JM5COpuiYl/t5cy0ckyBBUbM+InUn5i9u
aysPsWpEH/a6TCFLLot5JOQ42xwdQhK2YpSvHF+Jud1RnJRXF2uuBQPuz/wsbJRinAA5MO1O+MK6
kKyjgHRTykoZa4fWjoo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YV1jz/FUblAxpL6DA0Nu68JH/UQobISC1N7gTb8V1JuwEhk2ID5nESpHZgtkocebrR/Ibk14TefX
FTiToLip43yq8pYmIR1RBJRKQ8TkNCFM67HB+R7j0oINTK4d4tJlsJBYFYM5WKILhzid/npd5cfZ
e14YTmANKL4IU2TaaytqO2jL3G++8gPBWFXH6wwl0rEJgz678oqtVodWUpj02Fqui5bLpVJt9vty
gq+Z2eRqWNVClhi1Qp5mrRFJPpdEOdaOO2iqWZPxaL05Ctg6ITtYWEEb511TryT7ApPEk80ij6Zo
DmBn2t1kVK2RGHWZeCL9rSu/YDepcfhKC8fkmA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fnNzo5b3rCZfiK7RWo0OHmDS7fgv0LGfWYMnkT4/wqu01vEeUaqSFYirsBrEUTeIW8xz75l99fG1
gPQc2fbGAXBEMFgUTjapsC3Ayli9XZ2gNThgZcuYnd4qCpV1eFddPZPMskkd6oBHQVGpYox3mwlm
X+7eml9aXdb9dTFWmxA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SPIIGBg6z+n+uSLCPFmxHCsS5hoTQBwvF0gEvvuGPs5MwN4PoUBbktxix5ABXiI9w2Ipjk6OQOCP
3XXf6uaW7OEaimjbE+J36xtjqhVW3P6TNS/DoSzqfxwQhMznZSm7mxZsKYLJ+jwo3/1WKud737PU
shOmPHhrJlbkdmiavUsuvZ0Gfb9XZTt79DgmjNYiLD41l0moM9OJ0cxILvRMHzVgNKykBEuI+7gB
pyuO1KnZeuPz9tGwNygC0TqqFCg9Ql9K7a/nHf3ZhotV4sNdy8+Ta4TWkVafvsqbmqtOXeBI6pRf
pXv8NS3vp4Dwh4qfVLWUVXdgACUP2SbEBgOUZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28928)
`protect data_block
KUCJWKWAEVLyYbov6wvxhM9DuDgHPGWxWK4VxaP7BluJEfbjycKgXKIVDLDWotb39rxlWNTa0221
80qBQ2Lqyqi95ibWclxRY0XyjZBXklyfrXH3CQbzpQVX6M+8h2OrB+TS/bIzuT76gm9M0ZvXfoGh
iVX+Oopgyuq6YYjZTfsVSDJPYujXG+cS4fa5NEwGTxHFstTCkujDdvahsgVYZYTvwfGYHttfpe9/
dtkRpFW3y94rBoi/lQgSh5EfSW0bIl18lsGXZ9CRk7/vmFLNpnbgAeYdRsbMYyLPUMbdtE/mkBt0
oQybztcs8j0BU8+3y2fddbILgAeAPAp70mUfSjUyv0x7m2gJ/eEVflRNDDi5MYY2oE3dCg6F1TJu
+0miLZMpUX5BsJZFspeQBwrBnMGzjQnoMQ96TIoHe2mWNkHL8l0BYu15nNtDDEA6gLt+YIHNcpuJ
KmKuoJV9Ely9r6vTk33OET2Sf6mFihQ5bq1kM528Fe8PC+5II80DySHqm7q/+WBWN6azQ/Rdm6d0
zjJxleVzI8npnzHVAPNBfWc9D3m7dDw90WHC5hrAyEHafn0bLwOvYzrpxQegMx9cNXaM5qLEgGMV
424BIo6vbpquY2EOFvJbX+8Xgx5MnYwx1drHjpc+eHmhzSfEVuBFD1jmwG6R9AnIOzaShviW7BDU
NGR7AFp06xYt1sIwIIgRzqP+ExpDFSJBh3PVQ7CYoLTX8nOkWw6wcEM2V/UmrAlH3t2AG2K5jW13
LH5pFrv62Vhl2MZ5XSHi+Mp6JMoj7GyJgXSrVoNjqMN8D40Q0C0Mto9kjXDzz0lCz6HhKGn5D3iS
Uuu2RDB7c/IUl+bFiOxBe3FSkm2IoIhkuqfJyDGzaCb8np+5dPo8Z3unXmyRFvsT0FJ03EgzWI/n
SiZUyt1P46VPRM4FvEtMexUw2K+Dq/2MRT3q+NE8L9YhPY2tf1QI3GzbdoFuWTzECIiagrZtECMj
oS+TY8uXcsNnM8Lcoq+I2Evw53t7B158k+bO4eSs0HKPE6KCoKbpQAEx3T8toP4bra3fSMJQMQhF
H0T7V4Izz00PC8oZP4yf4b7XlKVQxSvbl40uMDYFLz0bZegtFL/kl3XQByRftuio9aqC222M0u0g
mVbmcjIHAv0lt8OUGYae3SnCt7Znz+6vLGf5kVDFxlFcWoln/lJHBSNavlam8sqxkjkam6bPZXdt
zX+fPPhmq9c6ChdkWDx4cmrWmFOtn147W1/9tt8PxbHSenUzxd54fWTH6YgnAq8D6kiJoQULUgy2
/c72BPcR7ipqRsm0huDrOgz85D4aTEpmwdQAN5qR7Sstr1ws+ooqSEikIxtynvWptPfnGB6iHy5H
MyihygP5AHm5Vv29N3ctCQsOnjvw6B0NJETNlwueqcRoXN9Qw0a/73VnUiAwZBpi4cL0l28n3Wso
0/kCicQTS4FDuiTREDAQlpDLrttin4/4fhMwJt28XpJCAUs0qNuZCj0a5MHD7G5iVOcCCuon3FFt
prBkwTs7LexiNBM+qADK6AsQqRMJSzt8X9YnSoOFFrGGoH6VTFPoWUnlFhexdUX/AFEU00QuUYoT
7qmAEip8O115XwhqgHB8j+2LHbY5zLBP749AK5Gvzd6SMtVatb8c0nTyF0ign7P1Y5ou8xnm8Fft
tZabFQ2uzmJY5efnqi+Old3/hYK9kfoxkAnraN/KNPrJi/tEEvMCg5J6yE10k6dE7BO8j4/8Rclp
eKFGRf2AHwbkR0a2XK3poSA7OPAvFNqHMZBBN2qZOH+0Hr5GoIa5v8SzkWRUEqZlerWytuqqz5Az
kffEf96A4PjJKlE6JeS29yhkEGzeimWexp7Oy5gKj+wDOfRNWtOc3agMBAG6+Vk5PTjiPyTE9hYd
iV7D1fEM6aKWsIKkZPzX5HERU9VZ1REfKaNLiybKdg9HiwZMs1N+SJG1bauixfO6+oBoT7oAcAdS
MjBeB7Jfcp3ok8sFC1UYLxZWG+KAmQAxhb31n6ksPVG1Gi7vwzreAT4mMX9DHslabJyojEoaHEpX
AsKFE7BdefcFgUCCBCF39maqBsRGATPTkhscSjSwccQ2joTDcv4MB6SaILdvgiTfreMOTdpomCOD
8dVwMDkHmJjTfhgBbWrQJBywjXHg98XHKdAFntT1TcNsTVra1mGt0GC/7mes/qAGZDX+YhLXMRXj
7+EPubRStLGFwT9Pmf9jgqXFEBV2v9QM0im0V1oJ9NoV/7Lh9unNXjMpMKLZgnSeQ7GA2VK/H/B3
uigurNjq1/f0XNIUjl5RYRzaKqT5m+D1bRewGQXkzdZlM9yu/ykdyqn/N3Ur0XeKXAphGnrmHj/S
lFuwiImHGe0vgeKzIdAyAJXlHx3AYvrmU2L7mamFnEg0DU1b5gFSW8Ov0XAGk9OnWmQMWoEwEXSy
IwjMYznnvvLK/9Pdxyn039mokhZD50E3q2XGY222CoZi7ii0TzJcHRPjqecseIzFdy02JGqCQ19+
hCOzi2uqwNMYba42Q6g6zZbAKHxwJr8KQBDcY1dJitY5t1x5aXV4+jxjkCw37y3oEIz8DP/nXjEm
UziW+j+4jer9mP0UDwme2GhdvvNpeWgBlMU5TZZSAMBgyHsqFbsm9zZ5kPZ7yqgx5zZ71rY3YK4R
ZL+2oHgxoMDQDtWxS6Okihemgxv+3zjcKg9y/qooF/JVRRTKIBbR9+N5twNUvAZZxZx+hCBrDVQn
Q67pRTLxQ+o0G9X+CcYPncgVPZHxOGNWPfuXXD3KnbleLU0qUwdB67z6pm9wzZd21PkuQIw84Exb
kSR1LoUzHTK+2FH9DI5i/2r16R1TYct3epp/pJHlTf6lAyYxyBSMDBScMLyPQxEzjtftvSTjf9eF
Vs3dWqpghl32kEopRyWddPOEd0Zo6Ad5+rHJWIu9rC1NOTfRsuS2qzjfswFpihYV1ZHZNC2VfkyZ
jAnfGRW5kctT33O5lh0JRESG3EbGEGO60HafHVRJvPYMzAva2+3wIV2jpm1IYZFqF/67JB9wup/Q
R+mGUok5NQZCzVf28fr6GXloFnFSTMzGANeEHAa7vcPhp46bBtwruIz+0Li1yS2+HOlLF85BwiJo
g9KmNRx+7MJib++O4de7VRd+NVdSkTvYJEnSSHKheZN376pfqB4v5G1hiR/RfqozKGRDGTHXQMDt
GM6IgJSrQflWjAEAMaNwuX/eZ7nk1m3qimbi3ixwJu8UFwDD3rghMteRKOIDej8w+mvCJDOvL5l2
vwLOqaK4hQfRlm2QMrVrhIgxnjhtcGovmk8WRceIZBSmOCXJUJ8FkIOdmX0/1AHya4L6hv4rLRnj
O9l01CTxGqB8Dj3wqOuY8N7GtVQi8waVt/qrT62beaqO7bKGxvO77wMI1qub0cPT9LwCgNzil4ur
O51DBQe9pw/EuGBKEpVfUs/UPMs1ZYHuWYXY6t6I+M+XVcc5Z6YJ1ZS+DFh0eXKMwe2ZnS+I0E1j
PFOTnOSvE6eo6EMulk/yEGRUtVuiB14hHWVQZgjWOF4Ja8Q58iLh5YwQ9TDOzyACEixpuq4tTS2c
bzvA7bD1XXx6MVM3E2qXr/ATUJ3NZDWnpdwr/+bCImyi97Win+uagGaYI9bAo8XJzEKKi2ISTm0v
HcAJM1RjZ6ArKXe6zdEUPt9z6hFLuv+EjAjWixH2qaLzM+BSPhwIiGQ9cDSLULFudT0BQgn7NxrL
lKC/5W85YUloZoYWVQSEivknI0Jh7178PfMHP6N8pvU/pW6RZn9AcxH4Zt2ANJuf6eBjzJx/dkug
Du2zZXzo1im38wmtGT9sHOH3WiKujTbrmrSIGu/CeRlSJjtVbuomdOVvCoSX0om0ta0YYlQVQbS7
SyLHzCWzR8kmX3yhT4wetpycvlS3AIpl9m+rSOYbnW+KNC1hKLyf9sdHiuMz+ggM7GGR13Kf225m
GIzthc9ShW4bf1a7hQAgxL++kpUodYC7O9XG/VFYaO1pcco+pkIxDFa7HRm1kxi2canOoIg/Zjin
Olfh5b8H/nfuMcMWEW6iFmzA36z6RlWyTNqEzbZBooTxqxkfdzZYCMNaGV0EtVzuaxVqHDcVSJ91
GjsIE3febR/rmRP/y06xlJclpXeeYoEFusej3ULJ0WoHTVJpKwaiYfAiy3KCjtsOribe7XevaItJ
CU/H3Qlm/JbNVYMy2LtNdsqjfFj6ItJNkTFt0iEy7VhsHKPsYvtYeSShALkLDpTjb8rxjSvij/22
UtSloyCn7he2A04Iut54X2M10eDs+vvbekOZEg05XoWalRiIhxeaK68qQ18apOj1Xn7aWGjEQTWr
z62NG0KPFLHOFfM7NeGN/RP6FqgYJInmmayxZ8dGTbCTppHpv6S4O5e9OuWtVQhdvPu1Rj1gcz7i
UvCIGXfm4Mg2tul79m06aTNkgYCOT6yi1WWhKIKgISdUO6BH738Uyd9xvBZjp6s++wmNVPzbaxNE
ludQDUBCRd0pszYiQS1K2mcc2/+ARBQQizKysQvwVHY78N+ZcwqnwIca6spmLe1he75u7nb8IxTp
PwFlB42DH33ouUGTW0yzSYbdKi8HabZuq/47aHVsGxc+U526iwR4qQSPDF1NKqqD2PdfEjf/Oe3u
wFKtuIz8fqZ3D+QaGI9SqJx8oWK/Ecyuy862lOjqIYEy31GkSCCfMsj4g5lEeJdIFQ4idAiHY4Im
J5qHJZns9NkzC0DMaJITGZiF6LK4Ep8BH7yjBLTcy1DMzxyCpqogin2d7aejIAtFoRMx5WLkGijU
dN6+RBLOE6XbgNnNOUnU2JkEKGBehooch1/nNao29mQyz1psrfLmjf0dtnntWuptbMcmhRioP9O9
htzTqNNQzNW+YFTiJjPfMSpsOcnCcAWM83fYaavlaVmMmTPjOHnuJedCmUvvhIw6zyc2YS98DXz4
eGKmBSTOmVLmTcMbvS5hBTEKlJmHBGqyrr74GQgyyf/s6SOQQHhZ34VEqqVoJCMrqockGYFARoes
06ylddBAujcpZzHq/CBxa20nxcj86qxpVVKT7A9GulAtqq3sERtc0mi/WW6r0aYM2SFxeR1cyAFf
nNK5mNGieGxY5AkP60W7d4qFo7jyIMhmbKh6sObYNIoQ4NxaDt+5aKKR83Sd/Aget6uJGVA3AydZ
dLSiX2AWI/DECjIQHPixNeS9z2X/93TQOLJeKZwpH5/tZMDabhUGJ1qqxVwfizwJ0xr14Su7WvIp
w1Xe/+p/ZUPdtfyUTFhknNhAsRhvolOrrrLrqdOD5xEVzyVJMHn4uTpM6daAIdGlsD4C1Yxs33UA
OXGcblimOTISihgCiUCnQu+bsNe20u3X+NbtwyPU+XdzHdu/95tnslbShbBT4Z0LPPzxfQkVBm/N
ijIGJiQEXfdlEZLIwGzvo96iR4oJ3dFzzcYJAmulBS+WXSgjgfYYTUBEPG3OywRVuf62OlgBhlww
Due6kZAHyIFY3d67RaZ6LTCZGLSmhjATZNR8UAiqEQgdibEnwc214NXM0KYHDDi/E+9B1jT8H9jL
EDdLuJvoYdegjDPl1UDiI77jZ5ywntZIECjavId1872lpgC4hGSE7YmaGas9WgKeUW4DTYfIflD0
5HWHGfr75yVQOBieOxoC6PgsMKIJrwd84AQNgvFqA/6WmXNzkqKB5QqimWfDUnT3AAJVuHTv4ziM
SfuV6UdgkzcQ2TPdnbuzNJoYeLV6M0iwaU9UT2oG3WlPXRUxIQhGgVy8PoCBnKXCf5Y9ON6rf1h8
JOb0HU6YEcu+FNqyHRPmsNeSE/unlDOcWtNfxkdwmzihsT1Cj5l+qPK4VBrNbQ8Txr7TIwjqbfhL
HdB4/OPB6IZDQacjyD52duNdrsv4VrTLqWcQjSHLkRADZV86q+TCFX9ou0Z1tJdweNuRWD981/Mf
mndhLeTXffirc8MGRsXSbaveS+wkQkksjPF5/Go91v15Jjr7UpPClm5vHf32ZmzDcdc8Wg/5j5RY
yP1IieZvkl2l69CJ5eRk+pwcDTiNZ8ohtp//wBt7cx2dvv373Z/+Mw3hR0CYCoNW2ReyhZpS2HKd
kM/KF3Fhk0KeKIDK5pqCF8+Iv8qQNKZL8jq0J0DXcz+2+YJHo9TurAVblJbVGQYGq2zPuV/az7pw
p8NtRB7jgukxciSaVV5p/lYxbKUEZ+g3+WBCSawl9SCdY69H/1p+N+g4Uvm8eMgkCZln0AJSWAxi
F4B47LiJXoDhrG0YzJPOC1TZNUHQI7O3Nz5Kg1kmiOSsboQuFGkerJy8f91NDo7BYTO0tBxJGfiO
gsMKU7RkYE9ZW/bDHMlzPadEL+PRqcIzhYRxZ6RKJGy9oSNIddUh72b2DbhuxtQRPJ/4vv2oH4jh
2jlK2vlykN95l3bm6aq6cnmvne06fn+xuI7We0/LkRwbPC13ORHp9xJOdKKqPpWU37N7DcBAVrjB
xfI8iuaDENgWrRA4bnZ1HFvjcY7IkDRuAGcoEc5bbPy2mHAk+t52NRd7VCCIzNH1aeeprwF+rgzz
Lt38bldn2VsfxJ/cyOMx3qO6gbu331osojTJzudCD+kHE+UY2pKuGnyl4Ibk30KdENlsinFzxnvH
rB4Fy/l77iM4A+Qh5MGS7hSJqLAWswWvwUvSdmwfjWRaHSz7a8mqXe//tDIn+NCF7l+mymYqSsS8
f0kiV1CQ/WQkz27s0R1GA3RiEOjkuhjEtk2bb663E89abZS9zboDVD4sJUDTv5QDbPSgpBQz8qag
C3svu/uwt4MttUaN2vZbqK5Eqk3vUwZzuLV14U+Q6zFDoZzRJY1iUrrDfebruq/GWS4CjJhv3bqv
6+uA+l5hRZcnyq7Yfi3Ej8Ii7CaxEcU62BX/uMGdDH7tQqRI74Ca04zsvi2nZd38v+5+g6pGJ5Jd
F1aJvXrStRfpalgElPn57T1ZkX6stFdfqonBDjnurOd66RBMHO6dJOnYNfchZl4QfzAB9o39fVPG
jdBWXWi9+fHZnU4rCreMV0X30VEr+RM6DxvRXxqBWCG5gtjOnhSKE6ujKGlwdmrlkji//sGPCGtH
FIyWbh6bfN9KyswuUDuC0acvGUrQoq9RCeS1MFPPteCwnK6WbYkGG5KqHJ4bAgIjtU1gE9XBoTav
TFexDFojYL3/D+S/JDiCcO32lvgVh00OBJSB8OnFUN5Mgx9b1FYy3kJN8Qy3zqpzml1j3pbC+F0X
hleQ8iBh/rI4bJfimFmt144l32JYuB2hW3YuGVt6TzYQ8wTGFP9X57j84NWNCQ4XnMRkOP2mOyJM
LLESn1gjrY1rtIT06xts65PY50qyCYoS0kfvGlMTEHlcYFFrDTO4rIfPsonrJ6w6LyH2EobEpfGx
3b/IsM7KEs0W4m9pnGwfz1NUZyUwlBxuQPVD+BJA2Qmn9eWOiX8OZ8IVLJAzNTddrD4Wx83vguei
l39IRWHoBZPn2Ba+HtUloXtvmgFFcSRBL+ExljTA8Gmxxvl6XShViXA0pvHVz/JdvSP9xpXoXJGp
9YEdmfoBYvfhuIc0gDQ7z2IIdKpPohxGl6POKCApveYjIYqCly096GfYKzxBBuj59YoSXPNAbWN7
fl4Pbmd6CaCZosZ7OX0ecTL3sQq+PR/Gu0ZvKuF/XqUomX9yvO21I4G6vzdU2yNAibOthxpx9V5S
fyeNBIfFVPi92e+2KtbkEL/R9H4AdE8LSbAuFRqcl7gFRTfm+Jftb0fTQThC0YbbWr6PSZQkWsai
TbUOsicW7vxFtYC97h1XN7aht0t/W0C7c+TXq6o4/dvfZ3SoB3iZQIaDa8k0Dxfy6CW6EjveSxxi
pJ/Pz5iwgACF1WFj1RW23bpApYkPnAMHdhETRimMcePPo46CJDg5UJcFpReQi3OSg9p7VW/1K1SI
hHVmqUCIh/C+p/FbqxG+X3tGkFiW5deD6tPKu4XXY/shAJDF8lRf1gv+gI/60MIO/obPyzzpFge/
LZUyPjNAAkXRRq+Z/H028EPIWxexKtwwMKigUzGIlZz3nDayIFH3Rd0Jfx6HosJtXup5uiHzls5U
g+MtSkjahdbV6b4AxwAWqvJ49w0R9ZLCmu3YQJ+BgQXmzy9RTmLrmrj8cfme863L8YmvbQwafnMG
GuPxjO+gYe4jvnqAdB3A5XPwHrIqTcJdNZdVwcg5GP8/lcsiRAYFbzE97gfP7nbWQRRScFu+zpRk
4i99Dt9sAHVb+b0Iv6YiWNilDxgo+oLioQ92GYqBUvX8P2upAzYH6lJyfbPadNox/ZFpguDlsZ49
JYeC5bU5CWiNoh7NOggZmRHj4Tt1SmCtLdO7n7kKcGrSSYhM5rMXGDOnjxYDxOk3vn2+v7e4zjZ8
wlarbrNhrMNbxoYZ7UY+5TX7PQoqPm8tp8a7SYbnPdbX1tiTC2lqizC8Ol1swA4Ld/BzSySSX8Bc
LKilL7YRc9OZnQ+HyEsdGP4PzW6NWyFoa2+xn6fw7d1fia/WduVm6z7JJnQoAWjLe9Fet2+3NNrO
ejGgwb2S3WJwetTrnFwYncOxrQsqBqLhEByG4qjApdvNhtlEUG6UTwyky2KaNfk1G+MmR7VZ7Yqz
EQAhd4SROzfi7ZC+0dd11SThUonJDYy6Ur1xflC/xnT/PhU2D1+Q1fPUZZW27Juw8ZrD/s9OU58M
a1Ku0bFf52HNbkltyvwvG+j62w/IDkyHJuCSNADwD2I3THoJlSpy+Vi1tyAjeXvJt+hhK0Sdj5SJ
+NXAWzegYJMd48DLAhVA33bVtLtjZOn+bKficw8smr+Nj5MrD1RgDVVCbRn4uOos/9G1LYzAHi7/
wKj0+zg08NpuVK0Wfqy7H8L2oj8UDZE20ZH2Uko1yNNMmA1e9plIl/lX53lwR+4BCdHAljQF7sHG
Z0hfti//az3A4s4NhQDTkJ2Uy3Nju7QzGVja0l/YKTlP727EYVsY7Vy6e55E9/Df2Ns3m7IQ3oAI
Pv7a07MQ7Gb1a3g+6b77LUAkZf/JHU3QKo9Bk2nvCQJVFLEZaoflfE4DqtGGCpP+Cgt6Il70Jr32
Z5XbG0UyFTIUk1Ksno0I6cR4Ox1z5u107rKsngoUbGlOLyDA5w9fMw9bXow1QImLS785r4MmgmKS
/4d8BxqEs/TwOlu33q45UfnvYK0po+ThEWBITTEAoMIe/CPtPIrZZa5Szt8SmnQ9ekMVlT7RJoaS
+bi4ZI+PTI15p38kJORvvZ4OMtZCTjV0Kz5XGWowLtZXgSAO6oct+r4rPz2h7Z+YVkm7xGPtCA2d
lInyOP2H4ZS1n6NdtjOMiormpMIQ0XO8wNKplGwUxJj/pNXjj/Sw9Z6khvocdGE9jL6JNa4UrJP9
fg5+YIe0FQ8i7Qe8TGdRo4mtSqVn9i77RdHGMYDsJQ8aen9lFu0GYQlWU6O0q6lHmZ7S2mDCJpSE
kr09rNyfZbuJtlw5TwS9xcbN80N7t2Xr8lEdd5OsgboahSreqd59P5dyKlvvIoIPUIK60RpQflyD
HSCo/IXUs3eiTJ6UkmeaAmR/VVCcCyYSELKcKOYWZXFrbr22jGuGGSMKlkGawUIfFm2kLMw+GKsj
j/bkWz6LTz40/CurcyCwBM0ZX2QTWps0LW1fizv3or/1aRt/JkvmNdtjUxPVVtJQUDaJPZzstTg1
KI4W1eeE6VXcwi9woLhKNNMyV9tqgWdBlNHEEDzWgONGGvp4Iu4cW91wX6K2oHX7oB87ur7KiiG5
KuIG0ZP+zdafj/sRxX8qSF5qRl0953nCns1IKVaESHCb00inLDIGn2YlDjMhq1jcNt1V+oefD270
Ywgsel3Lym5rBboLP4ziDNyPsxb8f9FEt33KnGhsKEeeTzytnEN4cV1gYPyqVkLfNQN8RgvlnUHU
p88aR/7T5E/NT61/WaDb27oc3GuaiML9neUyIAZlWhaQaiiqepUP3KPosZfRTzd3SI8SjRR25hUi
xbTmZD/g0y179fRlpJcgjmzCGTEz4RxzILJbLVPAptwPiS81kggdRNAPwuvcbVJ+qhGWg70iIai4
O5/3OjpGp9mFgVfRl9ObekiKMXiYcY9Uhhv9nIbmD87Kk7IjFqbZQqh4GtXX5sGtZFTXj2VhRyew
/umHnsuZMTSNUyjethO090KMH1ZRdGYShZ5ZEuAmd1ES0dhtE3UHbinZ2Az3o/KTs2ocPVOflVA/
sIppnI//zLWmCgv9RuZt/ocGIS6r3lFwLtUDnCoUan1IvIiWd+ZQFaoRgos69paR3MGJeEVNaO1j
HbU4vH9EMgANtuQx0ax84X6F1/MfNp864zIabtDMNkwh7iivagnLcsxkV+IZtD4pewoM5hP/MVzq
bGiUkDmZanZfg/6290w6554TJthJ3s33rfE9QPc5ktF7wqKNrAJfr1dV23bBJnG6NWxopv8i7Y9t
XE2NQuM1clFIyb2GiZY3q7tlYXnsq9HO9XncRcoOvdvpDedR7pgdjyR73FcBDlMNMeYp6aEe1zjz
7xpu8x5eSsuRHWdgqHOwm7m63n/c84t238nV+CyQU/AaNN0/pLuapfZ/lZoxF0rWPOKl6zlI1tlA
ZmjT/l6sKdYPe5+PfC+we33f4Nc9TylU2AMlvyR7SaWLQhNz/0Qxwunpi622pHldHaGCbXjfMzNN
LnEVaVTWoUmgjU+pMXlzJAGkRXl31WAxbKnnkLpQElzBmDIDaIgseOrshY5oXK+rCqryMwrVsNpK
y8qxhLJZ3Klo9ixBWpvjdoPj6rSGwAdFBoRHMIm5Bl2yk5efKjHDZ3Rr31QBPtTCMSwh3T7Rh8Qf
iALHzwmh2PT8XwzMj3oAZkawlcDHNHchG445oQ0Bdmim+OiyGBKL/zj1le2jOqBflENaVxmRZlLm
LQ2jjFNv2RbIbD12REDpn5/tzW9OtiLxRdQbGYkZIsNc5XPBJ5iSMSRXdyZ+WBPI7VDy/4piNXhF
pO9Ui08OmfPqFxe2r+bn3LrKiL7TuDrFxSy6TEWOWZJZTGqs3ukzR9MmjkomiQMZQsuK8CriPIy2
HGXE7tM4YZzQ4y1lW7y1U8HYj4b+2jU89u2VYxQkxeEL/0RrHHyWyg5NQmHxb9ikC9pz5rX7Z1+C
OSAQkYOvBeKlHhUyTJQxh+U+BAG9WpccUHnLLPygBlO8TVej+54WmIRguMrG9Vmk9Un8fu900ks2
dln/eQI4lH35LkHIUv4R5/zBRFw3fYBBGKIZZijskY7l3ZX79DlAzPS7xCqwzbZn+z6Y/YFaRIOS
bxzObI0sv6fQocJaxJDXtdPcKZ+LdmfAhthRMqrIy4u1B4UBXBJKGfKyvonYjAGE+nu5sYpKWguX
KMA0J0tSxoDZq0xbwfC6u2ZftS75sAIkYsqbVh2iPvOv3ELHoTkVBlA5MzjIzEHlGm52/ZAf30HA
W6syOBOL1s0wXLIJkwQFJkqAwZ2pgNsm+mgfoJhyB6SCJxNw6oPsuvMAFgevc/eyNEHxCFp6abrl
DcwAKsZbaxTARQkdhkdy39l1lRsRuLU5EHiEi7OUSsmYmv/0AQ3DcQIjBGuhfo9BN9J6LcmoHksH
lbG2R7kO0Vswzmmb9MVpc7vg4T80dKzlMb/CcjkRZQzynEQdreUfPKbtksdOudqONY9N3FQmDGZa
AynepChK+hLYQZmDDrXL0uFtqXcxI+I6TMZtaLca9fvLXZPkCty+rCoybD8nAYkoF7ir9Uor2gny
iRoBdhB+OYXx77fX+NJc2LxTH/upZtRnSwvfqfL7tpul3rbzbx1Tu2oM3MklMwV04PHdb5p7brzU
ZnW6E8pdT0mRPvYUGPHMpEe/51yCF+Wm64y40b3MyOB6MtK4ka/U/ySmdjdvMzxqQB0d9m92hV7E
EmLeM4fJ7UgKSG7xcDx0q6/Ws/7AcnvjmFIxIlW5Om578wfHPfGMTeIE6tOpSKtzw3iRCjFgEGjB
kibrC1H/W3bk0voEkj3YpmWYMyV3ATWnjcoAbL3t66CGEtzaxfyLSq77FlT6sN2HiI/r5quSb3FM
2YyGBmIcnks6jKyN/aE+UT7shzxIYcZyrMtlPE1hlIAsru09eGXOEAfwHb7jjCBPTwGydGT28dPt
m9zDSixlxAdaWkD5zoS4QDn9Dgn9XnNsZDUZwd9T/OPJUMOmyQ1U2mVt/cSiwUkJn3aG7D2VBdE5
hMwrGLpNDRuOva1l+L1vcLGdrczgszbqawVMcm8uHIF6rHz6iPRUVUJNhBpuCyFCdB0NPKFs2wga
VaEoKMqgrjuNPXKt2lu1kyhxJq739snDfQNWHb+wnNXdvu16vEDz81wNghZlRzeVttRxBgIFfDzk
J79VgxzWRZm8cVyQmSvyTT+v20TNlAZn1gz2jr/1zoMjzSmGIiszG0Yewz+TZBmTxyqWTyafuUvx
WKuE9uyTrA1xkH6iXZGPMYIVUhMPfHPh8B5tIJHd7bvUSF4KXziH5w2dvAdAvmD/EKt3scABjG3m
LCTnUshhLcwLG8NGecGdlBDCXccw38Qd6IASKK1LBnssBapXDAc4jQK6chDitKrTYeBRVw1J/Yje
ns94TM5Mcf+Ld5gjpzYls3K71vBzwYtaV4Jk1tNrX7pEioW+a+lvJk4aeTfnbCDPsPOQGkMQRzBq
CRDE5wMNg6c8MRzMJ7eOrXL/kuw7RIv/T9ksQHFWg+5TdpdMtlxLjaYpBWIxIHJJpml+EIKLGcYX
uklNwzMqmb/QsU0x6nCjPYhfU5QslFmYRr3+kirYnwuP6UYq4UATC8WuFlPAoWunm+Emm6c8G659
BW+LZ/ksudD6Fpt19LwM1+4lhwUWY+KlwwROHOB0TGmjxSe33nt39VtmGpOtcAr9VeWlUo2FntCZ
bD5D3Zw3sC8Y46fmrNDjH7vvmopLj8mSDuQ4DNzfTHLHk4jqMFHMHmprsKTFMOL6B9wzRp6O4cat
ktFzNWZzGDn+fbfkMMrizAt/n5iKJj3CnhQ4fIjPIrTwfEm/7hBhPDVlsZQFSFaRv40K0UA2XgHe
PV63p++NpLri27IJFZxMlwLyacyvWFbikXnbkQkTalmnSJFNCYANfp8ucmmWgIsrrRo3PfFb6ob6
9hmqjriEOi6fxFnD8wln56D7vbq1tdIK9IN3Vz7snVMaADqW6UVtZ08kR8VxZGcRODEeHqtGesXx
QcI7cd5+8UXSW0e7eS3NYOJStt2R9j29Gv+Svq0lhFNjDQtDvCYatA4zKSr5kRnz4G0CGDRObIP6
v5l9kvD7pXWSQZ3ZIafglFuKfpD1zYNsSHMqmMfYAqS9A75af1gGF2eFWO0rkgxTmcwD22W2C1/T
O9/vCBe4zjgNqFad0u9hkUK90jC1Zmrn2qnGw3i6jnYMNu3ToA1XQVofGlLE/hsxosRcMKk0Y3Ps
CF6u9d48nRwctaSgJWi/mhpVqJh4bZQ/Fnnq6rod6idmV1uYA97dVWs2mS78cRHUJ1S9XXcGavFM
5GaDSRRkKCGJP/wsuoWmrUMg+RJl1c70ZuCB0GtWOAT6EAN1F6lx+kBWlyCnVV4uExmopLVSZ5x/
bmDgF8ooIM+8hIz9EJK28HGEl95E0THy6TxvSwrgDm5mbsxJqVZUhIKsJSCQA53DbbtIBh7/7iam
y7cLz0EGxPukiidJLAUgfZ8L5lNL+hkSHBrxMhDy3uSga73xtCanesurRf/4QxkIpcQclMnhFbju
xssuHVh4NeenLWf8VFzvjXF6TUHrWye54JhkuKkfAfU1MX4VkwrInxRB+8VMyfvWgwIcBwox6mB6
LHwOF7D/Iwb6FfYcv6mkeQDjYr1dX9Sq3bW3iBZNoJFt7T90dbH8ilzJXOsdFw3AeSpTWhKBBrOq
NCrKKHNIpDTlaVzQzP+CHgBkf+UMRK3tJRu963dvpLLnc0C5kt2+A4lniAWignj/Xr+89V1XwWDi
Erqu1z6nyhEkVeF5h/oHF1ACQw/b6V5hCqSTTDoEKHFDar5fNTlSOuYX/qd4NQQ1Qv74xGAZqg3k
VZqLGgt+bNgZijzvHgtW1X1XCfCRYgZyZOqHNkErrFWRsytST6HukimulVczmecCYrNI2LW1cO0V
XP3BEw5jQ7IwHT1DnyhnoOSN4kHq1cnSujD6oh+wtlhYj7elqLOM00tMa2ApQxZJArDvvI8eQvfl
yW5W2wfzL5hv5hQda3Zec8vkusrkPCgX1ZApf4MkwcE69ybyQt7u/2CO0JuMtiNai7pY4d2/7R4N
M7NeJ+gXk7XEfo/emtX1/uq10AfFysBIeF81CdYKWxTvsNcvMxkNNZS/jJqdGCcAJP8EHjrxy8SY
HCYxn3NCCKXks1f1Sd1rcqt56EX2vSoly1LNMA5V2PjMlkM6KQGGyPAcKJiMeU0yWn8FY7uIokTF
4Re5QF65r+CSVtOV7VmzTUcxvPuE2t1xZz6uEfaa1/qIzvPydL9pGcUsFWAhIGFF3bg6x8fViA4f
WXQ2kn8wgdxxldPPdzuFotvwC1vtjRw2NXrLx8rtQ8cmLzqC4bO8cSOhwaAkf8X4OPqd2BxtKEIH
Vf8NZR7QwMddgRK+AezbMvZeKKgZEEFZKVhjlSLdHf3Q48EwSO9/206oJsFYqNptbBLOMlzZa7nC
Uy9rz3hEpjZNk9tbA0hBWj3G/lJ8VYnKpzkGYQzlfZ6aiTI0EPMRrtU95M2n78wOks0jItpmFc9i
CAM93D6YwXNai1Ly2FbuhtQuuWMhBodvhX5ZCfNESFghybaC8Sh/nVv3ymZz9Bd3TgD+W2hPYIKK
4SJkXbHGGOGcF3q5gxhAw9dck5EopQp6im04WkUB4T0+9D8vGCwC63K2SZENCQElgBwizl383eeI
/t0e+hRY8I/tE1fCZ7qoytAQtwxGCozhu4y3LjkhpzsEbVB5ug68/PQAD1zhz10o10PVWMpUR2W+
tFIB1VL6WXy3CwD+QEwc8F60r7HMMG/jZrN9wEC+2xR7axqX6feCbSBoaAnxVpxKhbpt9e/bdUyG
fzupHZed+zMTIK23QNmg7f4S9JEvBkXk4wmkbxRdttmyG8NwYnaNmCJhDIEAbuY9vT/tO3BISW3F
QssTImDLggsAkRoIzhYM0JHD0lUeoWr1Dh2YMSPm6k5/IWVLfEupNCXzrxrdk/udH0Qrqg6kEcjs
GU0PEym7LWH3D+PX4Hu3VAe0gP04J16rpOxjLwLeyUTmNcjMx40KZNHYhcoiiVuxehQISTDUkkqe
v8WkrhIiqt1rtdvZsLX5Zti5oPO+GYckivf43+dxhMxEwK2igQ7RAL9xDfwD+1cs9vcfXXQ/W7N0
5o53sNfKMoa4Nx0sNFA5R1Ak1hXY6/YIkvhotOj6RAqFtfOC+9VbK/09+7EloKKIhLxMgMTQQXcZ
XJ4YZc8ExTO9LfYrifAHloCSRlYZe10e1yb5Kcz157BUJuPWMbYOYpbK5amGrQ6H2jfXfR+5XHxn
ZAP9qt3bHOMlBP/Wad8sRmgln3nXqwzuHUu2JcsvTAHnfaF2eHaoZfMuS2fx9LKqnFuIou2qCi0i
E24gFcOdKKNabuzq5OWGg215qX3SGWH/TN3zO9/VudFJp8X/Q0+ncr+1DN5BTjmTPU+xgyH8PWkr
UJ+lc5C1sn6q82PRK18F2wFBLfNtqJwux9lJkkmoECjfb4olYkHUlcciOePy4ozFJOZn1rLAT/ho
WIoags74SHqJr26zgmj3wcDJI59s2Z7YlRY8ltYgpvP9wFd+avsvlRPmO8UboPxx86nPBPNrsuJq
/IJhg8SqpPY6prqK2j1GLDQ647BNJgreVQdZTV+lFhwhtzvkdcb95XKeIDLNZANm+9t81tBbMLqz
kNWzYwbnMmnQTyLpHb4vrL0hMBiblbTvcubfVGTGSIrg1b+Roe/+fJh2cfzOx74N8Gx1aFKnJSp/
zz14abC4Y7ZUDmMTyNG+9AmWyj2xgCVecomDE6ypSpD7gZMtbiZVshXPtX5Yo2syEW4YlYofZrTO
gC4hdVLh4aVasEMJejY3rt2lvwTK+BougMIe2JeBGQWkx/6iE2iPfW8XZp+MQHUM4Fqg7AsJ1R5G
SoAdS9oIPegLlOJNT2TphQd3jN23r2ObuPXBDnLkupyt/OYJqn5rxDk6GfvC/XofC7/3qBV0UA4U
gsI3bRVvPYIaZ4ofjoH+SnK9g3mpLv9ExdfyRtSm7srTaE75tRuX8JyxHFUe3KEyp8yf8YQY1iGK
ixSm19UvioZ8Afl2ccBvGYi40yTJVtLSKASG5WdnEfBSgMSTh39511jLszl6dPsKvxfUdIGRHxwy
Elq+Pea69n+WytUL3zEQUhV3dKFNxQkPQThgl1IMECBgwSn9jDqP1baiqavUxkHSpL6DCCRPJU8l
bUT+2hOu8TyyJjCZbZHxwv7pN/K2rXFF6UUGOGfpYjJ1p8sn+jGC5kBTITcr/5A2sQe8RXnL364+
J1JkAOLgBRK83REkaRJnm5KSOk3ZPk/m5QsSyUQzVJC1QhKHfEuhQIqDl16x5BU4Vh/BWytXCQXa
Bit+93wN3q8WiDglspjDnYoluGGbBebdmEtG72bfwjCG8BYm4xDrz/k/mo/aXOTRoDoOg7FtNMyc
P/Szx/tu01UZ6y+feew12QXbrexXJ8A+GC/CHjTpQ+N/RZiVbGZdrcDcep09gSiDekleH4SB62iK
fTROaF5YTWZdFZtMZpLHm1cRE2/JagRGPUGjAujTTjeZRtTm3l2OgCVilYOV+DuwS3H4Plh5Wyjh
bL7u3SrTemqa6o5yBsJpBHsZSdSDsbIxj76X+cpUUqrZyKb4Uq6lsjE/rCP/e1utLLiHPS53ajeC
LmufXSrt+kGVv/fJQb6PudlpjpTEkZnr8VI3xc4ZKTXC/O+MO0UEHBEfoGZsCqWUKsSSEk1veJS+
YCgzLiyEh1eE8Asz4yj3Ff3ek0WlI8qfjymMWKqkQKx3iUyTU3xC410XRZ7OQk0Z0wOTP57BKoYO
oOqe5FhRBT4wDxj346T0Coq9UJjS7Bg5K6G3cA+qEgEF3IDhmUOORp8wVvLgPhw1QMQ+WXIhn2zg
Z0edUm58SBWe2uNmJwKb0p0DhKfS66z9ix3qly39zOVuSMjsDwNO4/InGUpGqACaBIiPE/po8iG4
nKOJJjUql9KfP2d3LoC0a1M84fVsucylgMDbz7WIIlEb7//fVs2k7gubTpkokvUrwopQRNP+SW8/
tjRZW22Fp5hRwp1KiLauetqLH3kITHjE/tvZcoZk0ZzvyTrhcaEXDipOsV1Pa5Z2wIywtc+GkhHC
TkcxKSWqi0rfEoDqTg9Jy55gtEYtV7/qDVk9KojKkrXRSndZzdXt96N4zbuO2yS2DI8+OvtPiA4/
VY/TUf1mA/EXGxrjQtKD1YBL9z6xwm2uoGV+cwpnjTT1oySJuA49vAZCuw8PxPQAptFzuGFlnq7A
8652+5pVnxtdgA1HYQ7bTRRXA3FcN5sw2G6CcLTcSFVHSKDfF34+FLAQtnEvwaFwxR+ySY/5dco/
8bySG/RdUm2QM+QwQBC4Zcncz27Af/bzUAIN/KkGb87LGpGqJu7iN/f5C2HM3buzC/ZauL/MaNYw
8O1MPGGdLKG/ZPJmeolzbV3Ca9AJac2NSJ6odP6sjFN5+tJbxYfWVekCJmu35gwmO1EGI7NcybKv
7rpHout1Ps4ZSuV5A1E9dTb2KV7Dv5Z1Q2lU4Oo7C0VJteM5oBmpyhjopAhpXgrL+wFfmV4UQLbe
w3cAqkrZa6g7FIyPfUOcuYd05KZ+c5JoRfPF+eprjFxCXjgFjrgjt+Uvc0qKvyA7A9So+I2IAY9L
2AY6SLN1z0hD7Y/DhqxqB7O9Cyp3mBrLpwSFZ9Ax2pGj2wOIK4vuPkOO/SCbVadOvc3W+1btHgj0
IXjIBMuF/YUpLHxa8SvNOPGLbBKjnml3KVCegy+ld/3re2sUdk2NkD8cVOi/e5vR/jL8tHby09xC
iCqpRwlItQjPB9Zfm/G4b1PsydxgiYmOduH+NN/VJP56U/U6eY7N9cSQZrJuHFfIvHnxD2OEv7hm
vcrm80IA2geVK+wNkG4amr+HXx56eF/aIvx3QVHzwy+IH5YJ1aH0R4IkRehi/2fY0Ks1ZgSOdGDV
T26WIUs2XWN4I3lAbgljlT/jSZ3QBTr/afiBTAorpflkTKpzhbkOJHZuirYHLcV8FbA5slM2FRry
vCebkOnIMq7MJrXx/eYdYyAkCvEHE2kpcHND+w8f6nVwxwZ7P4QkwaFhIJPuEWi5Bp5C+iOMhJ05
qwzKa+soP+4E6svn+im9eSTgWGuoZ3jTuhNpEiModAmWTo7TG1SJT7u5tuMMDPdFBIH2NHVTEVgs
Ag2h0feOIsOyIkF2OQwk2khK0z1kEL0VLVxAguc+dk6BDy8AqQkJd8Vcjli2Gh+Q0XPuzQE428u4
DGHi5yfzfYfRj2o40al2c5SaPufE/uyqFm6+n+cwNhnNvUOZ7px6gFkae/hhVdwqSnbPMgOQSTRH
cMIK6TvAM5LSWGqm05FhQKIhHKLSHVjNXIOrZb5q2Gx5r8o+9iYKkt0gdtNZ3ejH4Xb+onwbMIir
NNKMeuXiOhJ0argfIUFVpCEHMF4dTl1+scdGdQ07M+m74lNh9qoVtWrzmWpk3jkNaAMtsmfR5wUA
QYjy2iln7RXnYmUd1xOLjjFJjAjjtM1bJgtzivoRuu5GyXJgK8TkcLym0EAarzgJCSRm9TAh4JJs
BvbQ+gU4dAjSsN6yEt/xqVkMto1E4JQcxwTGGa3oQ7sQ985KktZh4iPEBKPpJtSVXyfX+edMkmjO
DtIQub4pBhxy2Etfxn0Cxmc/4fT0tN5ryNH9b0f4O+hqvLNQLKg205/vZq4/VIPQ9Wxb0X6+rXoI
Hufc/MDjIW3gfNkzGY9aE58amP12WXdTOcl59TUHlXSG0GbxBU+xZ21chnD6Y9pgDvlagvGqP1Pd
tSsz8CY8OIkI+iXd71oIQ43A1ND1zGsd5uDZ92PC4zj38GzQP4jtu7pbzfI9UWiMQEQKSQkJilGJ
ARcvusZCdvOze0zRODbc6/qbaRPynjBVrCHjNWv3cENe9v999Ha50HdWLIbF7DIEiAMW8nah+OBO
O6ODMkVIwWU5AWJMk4fhRV1ASG264aGdtBXgBdOFss4s7kEc3wgYIOpFy7kh5jTfMoZHK+iYYAFE
fncKr4f3lmCysNboeDpqacytxQNo+KMStfwO2roJvMbMJS3anAw06G3zL3s04WDCJUNv0Zoi44Yk
SOIKCYFh9SFMHIegq2P+1bCaaRfKIzph/0SZtIH1BedzzFrWnaTIGk62Ep+dZugE6ZLeTceBwyo/
TS40oQ2OogvNpN8et52T7krJD7UsZS3q2+U2XV/FcITa64Kjtw+dZ/RIgEutPKv2Lqg4Y1mPvV1e
oE5sxnQC66QG/q5fBtyA+wjj6anxbT4Elw/MwAgZpgXcDqLlScT2FA99dRQ8o8PDE5vb1SmmywjL
AZJm2+67M4Nef9u8cevduHT/uKNxZBb1uck8yXDj0T4JX6O23VIUFLifKVb/z0c/VBMVB0/2s4fD
VlbYh5XkdZNufpfoCAIH+2MzdmAQSMjb0w2JlG5cqnzPNbkuuOUFESvl0th6Hf6uKt2Dgimw/KTz
kg6YKX7u46PmwcCYk9izmfysDL6z75+HPr6w72GeIZ0Jcx2oYQkq+yHkUL0pncGoXGUEl9GEwkFC
oSm1FGHIJ5rfx/FAU7kS5azp0Jrn3E1wiRU3GFp4Zb9ibK/ll24Ws9xXj57RG31Tik2tIuBMW2WL
3HWerqTLa5owjmPsdvnxKJWAN1kI0Yvx1pdpcZXlZfq77JBo3vBB4bzA8B28TYOLf8ALlX+XTXoW
eNHPt6jboFalTeg4CTcMo9xqINgCs53VEyXRVakUIQ/Sj+rBxYF2WGfZGvINj5686lRjwHKuvRDe
XK7qmReEhpZas9S8xWSwbhjKlyUjATiMMowO1j73ANbXqEQ27/pSvYsbqxSKRKhkAXkRGoTDCZsJ
C8kyXe9jL3UN0h578/+0mlIwnYqhLz1UVkdy6xlPW4x/Lhz7ldiMzjjReJr6kB+X37Zw1EBUhEXS
34zuOtPKLSwJhKD0XebATlnzosfrjCrFIAI2g9hrrB3xGeC4xYzeacmKbZGqiL04qVtxtNRcJqwr
FWrWB9bNlOzYmkcL7jBj5ZKjPviHJmx/CJzhFVbRuayWK+xnJjgF8VojvbEKIDLEJotA883m9oR7
Ltq2oRB5MLz166ewYzYXFugxUDIPSG7/639oOeZWZOoJ7JaUUeQtaIqyKoOXRgpp1vLZ1x2o2jDW
GdUL18djw8CHIso8KhSVQsC5D7BzwN22B4Ihni66yhJJ16ir7bnbUGwEmEFZ6LKrJ1FQn7PhK0ES
+tuGbhR9VUxvPxChkiv333ffBnEbN2avb/cHRhL0nuKKemM7wzB5LCRaRFogREH190fKlxiGEGOL
UKJnltbRgbq9EgYNXf4ZAV7oQldxOZ0KhEa5OjIqO6zUN1S6b4N7d+VU3o2IGGmkz243o2a8jy2Q
kAIGYtNd/V72jVbAJaHSjrhZUUowRlToKT31LXOfqVHVPHRMXImRg/ZgbSfzWBf/R2aNLRcJw2yt
SRuDcZq4dSJ8wPRpFAyBvzfJeCbTbykUjIknoe0V0erAfvcVj3kwLGqlPU9li6qisRnpjB2deXeq
BLfu4/4LAd/44dOIqnriICUgdhe1BCfh6CPTX7H7X5YSwk3JAGm1/GH6yLlJRHGIYxM154VV9j5c
DYHMSxPYXmmbMtD6U+6hJDR4SXoQ6LIYqAEPO1fTcHX4zphIIjLUMPVr3cTh+DXfzxiiDpjzP3su
s1bYEbFjyEao6pLil3w5TQB6feFdqcxDS4MFxsdH1WaNRPSXlAY7TQmcsJFjczFWrWYf7TvN+SrE
Ha9ipmOBZDK3knom7ctf4XkQ1oPGhhHJ4g6EIovNXqXPSNICp4rnjWLaIpdVRwJWOT0fZr+rUUhI
ZVFhe3uRguV+rVtFlkOhed4lusLzA6G5kCbZVUaYx6/OkLMUndyU4752+7lbHMq0q65pq8DBIVV1
2pqiNLiN8f7wGWAaBKwkDXK/u92DI0XWshwhrqSpSsO7TkLElKfarTmLEejwqNkCI38H8SEHOBU6
d/Au0BZW4+Olne4l8NhEN1kWu0TMZwk2OWJvGMMe+DXF9K0Vz4UuuXbHbH1lKbUgR9XXIB5OgC9w
L/znvsoIGJptI9yuX5JH77RQgQRStQMFLoUn7uJEeF65zHxGJV74vDHEzNqRotXVUg6z4u/p/9Mq
p9G35q34Vre1+v0C5yUuPhBlSuKG+3iX2hl98FMaUrQZplL7mL3GoWINC6DFJT0qiyIzMuSL3KKm
l1Uv8z3RcmNVIdnMNWWrDofcPbknzEsyi6KKOWRWv7CpTW5a5DAeiTBon8JKy1JGAdB8oKK4vkym
GhTjF5XmCmpbEotjym3OxhjBUUBhIr6UwynJ9Akg+He33H8xDsqUQKB92mERizcKTMHZvFBGc9Gy
A+Mtn0lp2HlEABdLpJcxGi4A489VCyCtCqNh/i6y0+61wXOwPczUzjJhutPrv7tES1jElGOWaU3y
dGO5yvfq85ebTLH6fUomNYSjeIisJet72FjcNAEY3okY4IanLugfOaXLe3aMey+Sfj97r/zH9/oa
DiTJAdACTQAaVUJ0AvAxGHuR8Jbzcy1anB4IvvWEfMfizMOUl/HEXJPHRgXLTudRX8/C0LpBLumB
Xq/dyxl7TC/nEpKLcKfNIdQ9bjxqtcV2qCRpyw+VFVaixo1jhtEMs6etor3wx/gdAk/5U6nGeCha
qtQt94gZrOtrmAU7kqCv4lDoIcrhasqNm2p6yu18z8lnw5fiiY8rG8n0PyJROtf/XYWba3u/IDYi
rakovvaSfZFvZUCt3h0kbNmvT4nd1TNzilXrC8NvsnM9sUVmMyykjM+QJOFWynNdFs45Sqy1ChGq
Ojl+7kaj2J06xSkcCkZme0wcTajd04vz+RaNwVNPjIFxIzEa3Lfk/EeeVv36MDkG6OilZhkEXsAK
k120juK7y5ypvnBwi1ACrsJ/8CUjWY0xz58LxhKgNBXpoYci0pDomslCWpavYZDY6Rnw5oK5aL+d
hxIRvg1QSv1o8yfU4s4JFhpBXAaBU5ZOPVm9daF1JhUB/skXqOinjX3GUtFesFTqylcRAG3Uu7Pa
QRugAEWUHuc1jIygUva7ePqbVTWMpD59W72e4Bcf9Ai6ZqmAhJ8aJwSuqK9Ci6MuWCPIOu7mFH9x
xVTO+4NctLX7BlsCNYayWgCkszPvhNOb0cKaa0gfRgKjrE9adiuzbpIE0HB56+VUVxbhU2um1Xkv
EhITVjtGyK5Lw+45+fuNH+RkmWKuwbQUddJjNNXojdDRHXdQQYvr+e83d4kfqZT+j+/kNLf+rGjQ
/N6yiZJUQkOMoSUlUrnHesS659q2YpYpRU36TwTAnadsunIlj1vra5Ud6gzixH4pulRLs+fQYwk3
DmkobsHfWveJA0n0sqNoxv0WBRn6NJoyo5Pk5SfBgXxPYSfiFwlc4NdRa4eHuyWORARtsyFO+zK2
EFj8x2EVR7PSA4r8LOIUTwUbxV5Cn9ahRRCwImetXy3b7RD8MEE754pEp8tNHI0b4KlZnXp3f9xX
7Wn67SPHExomth7hsxG2o54uVqNjgGLx7TGtYs5o0eSke1chNWP3JRys7eXVs3EGat7OHW7F1/ST
yFTfsNALG9qjfTapufXnbX9Y5HmmEN8qe38SSRpX81LxmRBuYuXETuI1t4+y2cfWl2zci3TFZKDL
KNwNgiYfLusrxDSda80J0KPkYobxzYE06kFaPfvIdgQioheFnn2y6Xh30WWjSsb9HhH2g/xgoBpu
MtE1XDomU0620n1JGTwO7Y/zEA9z/eFwyzzMfZpFzBHw0UAc006pjWY+S8q8f+F1zs4OB1XZK5hJ
ZDtKnaDyNIWB67luRgQ/jcrv8VAdta6PGtfZSkwb5vBkg51NvKgehUSX+tPcvIjW4BRKiHXXtIcK
AkPUSxdqmZaNuku/uPDYSoytlg/JcW3cZ5lJrIaHNj9iV9TlS12fZryb2ubBuEcyc4ckKe2K+p2z
VqMujSb8kFgnn0OjJRimU1JSokuB6xO9WdJxiQb7r5zQuVzZF80/T66ZH5Ca1cGW0UL+GjI1I82P
iwmnwpqc5UNGOfl3eezHgHKZ7HD9wvnsFV0e+OKZ1nmUqwHVvNo/UxFTddcD8zhEPNRWWFIuR6Sh
fhREMjyHjKt4SCxdi4oGOF8hKXmHP16WtRbd1IFZT4ME7S4AeTBT1b7qGPoFbdWMIVoMsTN82p9R
Cq+XONl4UM17+t4jgZ1wCGlTbO/DoQJ2VonRuDJYQR/A9UsNd1FnLt3Yf9Ugqvzq98p7Za/s0bRE
QM8yaJcq05I+eix5oAwRNNAFV60xwmrVm96iAkwdS0VSpc5njOlIiI5X/PU3Gt0+y/3n8jPXJifO
eciOHJjaUj+cDs9eo5KcUSha2Hkafzqk6WflAg1ADtI5BkhBwkIt+IjqAaWJctuKfV0AnWKoEnHq
K1TCm72yONTa2kiV9CnpJQxJmP9H2LOAsjN9k24mdcDJLcg1fsHepvtDXgSYJ1T9Teih58SuKaqN
zHZPiFQZWJsKtr3ZYQVUDka1dseMIy9gefXlE7Aulx2XCFsSnoePXP6t5jqRE3Ln5wjNQetbRA4a
rIQcTnArbh+f9C1ZCxEuCQT+btQ27kADjQih3GLE8oL4xX5K8N8K0Bau0Kl21inveEnsmddxq+3/
MteMTOrQaFEvODYrYW53wq2cVXgoeShAxmKB0baVVunY6YSnfDO0NM3riqMoDnvpM2bA6akbvccD
hmwLuN8KCJPoKIqcWp7bH6OZwJ7V4hhRpF25CwdJWkPXnCdbKfh51b/c+okVJeTG88gygjE/9CtC
la77W71l5ic7annI/znwFsVaaE042nnEuiQX4LsMRxD1/zenyvN54PZ7mb2K3l0vXNVsKsTXnwGZ
JD7CROkpY8463I5jKBvU+D35+AIcT3BsdsMNdL+wL+jt5LyppA/XDRExMys5OLe1NCMgkrckmoii
KE/l1rN2oJKgqiwPTLc3ABHzKGUoWV6nNHyxBeFML8JuinbwgW3yMZXwFR+HPyD58Rd/PdP+0wgj
ZKzBkdVBko1PA5qKzo+ADRqZZdw2utDlAFqUxBW77kEzq8IEmTpFJIc32EH8H5pfXDcPJcYKFq5e
USVI32/Xu0O46CFrs+UBcbp1+Xw+M7ItH9tGaztAgjqAKpJV/nyr8KHPkBm6ihQRKdBesi5nbHuE
CRM6sLVek2ZeI0UjHl1rESps+Jk1sT4mPGziw+3CklxI0uB2HNdbRXjSqNWHkL1gn3kCRbSPLP6k
fH2AlzebK+0C3jQ4EBu/TKgF3t9n5He066jgbDLyFEy3Q0ufcoEUqsfHnsnxNugaiN5YIzL0UYQ4
fnW/WeKWY1rcAg+jOwxoUnYOcWT+1S8jHDb6SxTa8rinzqh0nxo4UUJPSQLIDniGZ0uAEieaL4+z
UfaHKHY4td8/Wn0UDTzFnumzAoYEosDn0DkDzg2WhCgN/Kgz/ZfibueL2X+Rna1FyNFAKKygxNsq
xLmD/Rrr/NGIBN9LqIQfAAijS5jGi3JOJubkRKaA8z3do7SkFwc2Tn6k9ZvuOh13b8PyAp+E0VoH
UaNqcuY918lFA+9LFG26ZND2PvbQRj80UfpOvbfn8jax6if0EJ/qaUnO/s5ahhmMCeWEQF+TmQ3v
kv7Al3Yo7uQNXBotgxVgj9jdb8Tfn/zAcFtk12Mr7H4IpxCkesQn25L14TQuR8RC2QRPE8SBZTTN
OtXGXXixwp5Q1aLA3fn24GcrftY2I/lEcW0L4A4WMh4BqdJSTDySIPyTflWBo0BvqSvQBFapYfGn
n11XMxnTqa1RycZtlXbDQf+sF2Z7sWFxYUvW7NNiWdrrvknHzoK4mkQ9Z2/gxiC0N0CEDQwFt37V
rMs/AmRsp3Ewn8vcrvk6s4tDpLIAIzMLTA8/11sBsXt36zmhwbO0vObtLazOl41u0VBPabDeM+QS
b6tq5Ny+gKcHeE7+dZC0GJoToV7TDbYtnYjmN4hXGYfOJcAn5d0VNxbQWG27OvaoHkUVFee/8Vit
S3vden5eE8smxIM/wxuddhLTkteDb5YVzyN+QktwFMoFYcsHh7xQKSG3j95uN3zTkwHT1O1NxT+q
mVibX930a1ljn/tYDkqcMLyj6zIPoNbHrECOYTezlsaRrQIiaTEr+Sy2eVJicC+C+pslit7VrNwU
fjTmjXDcW+vSX1gZn7vSLJtjPMrz7UBq5VQe5OxZ4xMtezbwWaYZQX5Sy7ZWswWUSbr2BNfI4M49
DTGZB8fN6q5lH469CRgmSAG/kBLpXcnG8ZUDc/U5UJ2UJLzyEZCiWRQNE5c2sX7QFso5qPbBq6r+
mZelz+PsiGPS+QnnNrodQ/A10l/MAjqyy2KM9NqPIeCd6pcwXQgiWVCE7IcnTqdJh6NFoI26B9Bt
5Nuzy5E/+Fccatb6rc5cmMAfFVvfLAE44FJTrKSNDFLvCBrxiuW20kuZpGuQZH4PVPK6GmfM4+yW
gaJYHhGLzJXl09pf2ZNAgWUYeH4+TCoqX+lQmC0n8PerHkELL+50nQkau5wBvmcl5Zm16uw/sq3A
bd9oYhZeiLX8Z5A6M2xlJrFSgTVrTnEvFAjZdQUb+W68PiiXQXdlVxKQTLU+hlfOjIF5kssJ+Inp
HXNsB6iwoNbHHA/8ga3kAn86bNZgna/47XJZKy9LsnjF0O7oEo74PrqJoHmNqkBm0gxf/8OcecpW
vRre/21PARreTxG2A8+po1NXP7463V5SYYn3s8FDiuwpB/nJAnFXoIXAWG83RNlPZvXYF8KwpcBS
Ww5XkSrmYOXlzSpBVG3Dle13vcTRFdLTp+t8phxg+6fHPDw+77/1UBMC29r4hKSErTCVED5qsCvf
tDwoTUk1Lo6vGNwPJ+wSsuZIEjFCb9QMSEq0H65k7BjxVpoy88U15BH5C4GuBWyNcHU4Cf64dtVp
mpiQFNjyAHvuXo+2N4hy31tO9o4de5X36xdwkZrPBkxkzmz3Q9A2VDJh6t+k8G9cqqLvMEsDYC5o
hhFb6DlsN3adXtWkT1usw0RLNOFHLnlO29Fb5AdTfnF1x6ZD8CgAKWHVrwZ1OtQtUQP//z12FHrK
5YQ59ZfBnDxTwJ4PYlVq6MCBw+d8vswnx+tycBm4CUI+hf9RSYAclrzl8mDFJENbn0cPzC6oFpd0
5GRKC/TeatqkWvwSDJZ+blcxOs5rEWo8BKilNzAvYh35HmANKzkfWJ9h7rih0G503/A+/3KK8KCl
UfKKIW1EoKHe+g3ZFmNun/HwNS87h0/e6jtPUmllyXBgIKAMT9ydRdemJ4VcuncOrUROkqZ10mSJ
7vb5lSp6R3PKdlwpz8nQ2ubHcwEjlzlXbBeUJvxBDySX23KKmhZexJLMkbWO3GZkqW5FumU5igza
up3uxJGyGlY5Qwege9VsaI6w+uTdHkppust4aMtAUV+tw2FckQluhYWLgw1QkyPAaS/9NkhZX9BK
z7NlQQ0L5e11OHceEF0s76JGyfH+Z3jljvBn0KQ5NzkhvaNHRZzUhh3bsDQh+1Xe1UqVsZDjg2O7
G1vzMlSv5JGKxuOOaGcGDyOuWDenKmmRgkRAhsr+tQMbK/qLVw1EPMdUpwW0zSMX61VibBE/ABTM
K6zCXmhxLojbwZNosVrbjkbw0wLHGQ0PiFWOkkbYc4VY2lVOt859g7DwA0oD3AcCd8iW3xWRoYTh
clRpWQKLivpTDNQqynIHHgJgcIN7yJnqRG/G1EgcKShOvOwRsv3kpiV5TNMrVksZX1Q+0yrerOoE
1OnWza5xlBAiDP5uLMy+7rJhP4+Pem5zNXkK7AON4TYrA2mG8E5SOmSO/y+aced5q5zPZOoGm5ZE
fQS5K30ARsmXsgEpTl+uNms+TmCycQQdAEsMYYu0l9zClCII4CE+PufvNzIPEE5CR5VKxsn8aRhD
EKMX4dFDZ9yII2q/KA6hWLCwD4wEH9OULsRHyMyzbDEdvr8VcoNNwRjkqrcvlsAfcZj9k6L0aqbx
pOHEXDcOzP7yl6WEy/9PRB3dylhXqIkJog0968lXBjYwzKferlotLuUms74crYRYhEgtH/fPmy4V
i+MUUdA7OIlzRQ71kNjySL983iJjMsfUlvywLTee9Q9E9uFFgqspiM3gMZu4p6EvLOdDzSsnWq47
eA6sSIYoOQjEHkGMR3Ybg6aFn+hKkcyv35RB5PmvU4TuvnYIWktoV6n8ch5b3fi36QlJhXVbGg5x
hJmrjUJ1TnqNeteSxvZCc0T00whoN0+r1N5sGdXfomGv6NgNtRqnwXoeugB5Uyu3lw9L6+zlL6Mp
mUh1aVxl1QHm27bC1QenBfyuzt5Eitv2e/bhBcAz6BHh5bex0p77ARSiYyjxO0WfRHY8s1AW6DJm
V3+hNoqdgPdCjDVk8SrMmevpGFT1bU/5eE71/ZM3P3J/1+O/VgR7EPfzR35ff4cMIl6fZ0YS90Ye
XoE4HhBdycC+/ko+rLSESnMGmqWcm1Fx/nw6RqM2uVGUxpFEAuUDjN8raj+mKAoRlnYB9HeZuFEt
KJJth6Xfdc7eD5hK2BeB/wTW4t3eWh8kp09Jfa/3gGePmPz78JyjalWUdgwew4R7ktiT2m8l7XIF
ezxC3bbGvGayC/1ELoAp+OAt+qy6HZc3w9QGrX8b6Ohm/YcFYSDC4FuY7WzcvSCX2mxNwz2rZFhK
wBCnjqYwQWy3ZwcrR6FEeYvWy7tJXZpIIsMclcUmMbNHu/lTnne7Hhlliic/gUzgwtzlqFrglmdE
5lFsRl0xShTzJ9EbQW/c1aRWihzHUjXMHdSxx7vK8+we0QGWMzcRsW5qXHV2qEQ3aZ0tiQB2qqq2
QGi0P66taKQWBRrXrXtPreqD0HELlXSJlneekU+pZ283/25aVwyE+ojyqg0ZPgwl2GRbxlKn17RY
JYdvfWAxjrSUD+rRB+K3C8mWBozO7BE6u9ZHYvOqRgahzwOyWS4naMT0/jg6YFjPaPtr0VCGlzOj
wf8flJP5rKpYpfxxSoQVu1wyhwO4CEwGdoUXqzqZSpO9nJtzRrPMajyfGbBEaxLFdoEvrKhVwU4O
rTeCN9OiRUWfTfQOxTKXsxh1tS987J8zCDW0mJyaZhkj/AelDT7imzWaAF/DYf/ugute1BGNn3Oo
bagVISxF335BuRfO/GaKdViDoVNHzJkggUONuJwXQBge5IGq283NNmbGQUkcjVFOTxivlGIkm6wx
LOvBAWAv9Z/6BVg5bTL4rp2+ZvvtQ0aSEI3+QYABW/z8ba/Q+gzI3TubzSpsvZgJFNWoj1soF3xY
6x5+diCM0FhnaRl+L/dksSaRvGwWfgDmqmoZ6fYSzV3f7K3FXmT/9AUOC1k0kWuCREJJ781ToRK2
JYlyQC1Xj4ZzpeRNSQh//CNBUCnFA3uAlKxvlCQqzOQSHdCDiyEuWEB2xMVP1MPrmmXjeCIMDWZD
4FsLLmaWKhKGi/lfoxF9awP1xnHO0NCoZ81xOu0Y6YWtjt8VDdN5Qi75//yIkwwRFyPaUXtVuhbS
NmsxFIKZbT2BB22xqp9JzJWqq3KexMDxe0GKgbpKVYvf0T+LXnl2gi9lVxkvW+AgiGrkb/Bos/Km
GKhZ+i5LLEqc5nk0JaS6BB0nBJ3YkXfTzRiYnmSA6aqolpu/bMRg++YhrSaBNJ3jiOjdAUPQkMMf
ZT7RirC3IeMkEu1/CCIx49JXtCChXDvwcjW1pLlPYzMMPSbI+npLF3hknBPxbOVhf769shs+tRZ3
bUeI4wARJYEKcfeC+YwQXPGMzG8c2BNjVyuI5/1wMweKF4wMoIpW5ft93Sjt9Jy1Pk7mlx/eqnHj
eGQE3JLyfTkJ6tbtQ3ySCEsW+qKyDNETjSUJOeSwVjlk2UIoJa/QmZ40T1FKQTvwNYSG4jLwIVnE
eFIjtigaZXjbZPgX3FR+Mu/zzCz1IPNQ4mVuC4XnhOLqly6v+rtSBKE0tDRzwn1ge1SmlM4zYkV1
geQxuytpBu3gf99I+gSu1yV765qb8egeIYp7Kop2hGD2pViHDLDd6xBd8zc3Giu1GWljlRey0SWz
sf0Ci6DzkAbE3LNsjCNqgGN0m9etMHTaO7pyr3HxVhvq+QpaXijdTYSy3dPIqpe8hpdO3mX1bjMR
gEulTi6eqfW93cEYpEaxEJXrTCnBadu8vD06k6Vk+2a3DDdH94PaUIWoVBic7OrDB4wps74Qpi6T
LGPny0dpmnUz5pjM12ePXpxawiD9anaEc1vsS+Sy40aNvRgsl0umVYXp6ZJqjOGzc8bnNc3px+2q
AGmv2ccRwkOX4dTLC/HTAfVN9EcXWmNOTHkaAFWQ01WyoYQUYQAXA7mMCt4I3q7SNw/T67T+NVsF
Ksl1ukSUTbPn5ED9NiYxLIxgSE468BRuKivV09Ay+CFggxaQQoQdTrCU4zPz1QEAFu/035ZQjovC
MwrRzxChuP9IJyif5tvbQnSSkUvlG1e+kWadb4V1+IjDy/ucjSSDWN4BnqQusm9zXe4zQL1E4n3i
0f8yP7TP9QWrv2j5XMQW69SF1stI0DOHIhEvuTmMlAqILXqKMXL8FHqs3Hi+Ug/xzcXGqlZ7u+K/
9KCTo4bK1gklflbE3/Y+mkSHIFCOow6lbwVOs0C0BY58Gk1VNXMt9SOZV82Do8ooIvcG+awHEJCW
D5RJ93fy4jL4BxQ3+E4+4cwWftfJnmRwuVXSFFZF86zp9sHsff4L4S0/Jj+q1EjCGMicuwhhH4cS
X38HM78R9nPeLKXSvEemhBZqJSS9rqYxi2jiVJ7RF0w/KaJlaJyH8Rnchg40qnGIpPGjy66II9ts
ZcNVA8c6JdZMP/8XOqB6YcleGW5TlJO5tVbGAF5ovkOwPTE3+j9XJCPGIOdyyyWSUDe6352j2e+R
MhMcmpEP5H74wwDt7vnGwPmjrBa28NLOSxaQOR6boL1UZ8g9TNnGLM9MYu/niavDdlNKuN5pYBpk
ApIYT0L4jXACYuRlYoct7AapPMhzSmEPKksOH8iNZCWyooBID/sXlMydOSZq2OcXMtgT56vR8RbG
ZIA92BJiwOSp4Oynio6EHV/AINsJrVgFKdNVaGxZqX48VI8VFIMiG1KTlyoHTu8nRRuLy4ocmiKC
BA9NakuFnzJ5u0Ey15xZzIsmW/36fMkiiAtwVi23vpPkRsAXKGyp+om/Fo3qbLH6I0861C6/qIkj
rEDpNVUu9RNP/fPsSaXeMfcx1W8XWydPl1dtN7Sm1GS7ozHNza4k9J2nE2/77lk42bJH1mZavv7k
N7pCyAOam4y66BDe4DZisB0nH7Yg1Fn0VQxe9Xtq6G/MeHiVYDK3xeM62ilWccpRcuHkhKCiZvry
MuPQP+KhglAEJZYG/8/kuV+HBoevJUqfP9elFaZn2QdLi6nbEbkk3OCN4JqIg9ete7dcf2A5j3vV
JXHnmlloFpTNgVU6ZdPh5odobehDvKW5EwowKeRwhvWfnC/PF1bNksEd11i5aekIWFEZr9lsmaWX
1YO956FeWIvzOz7UAW/FvjNgQQccumh6fAAXXeyxN23l3gH/8pFX6tmjLWfl282OGyIqWtAJ4oBE
buA4V6cljIOz8lt3Z1JQy7rtvhxK2p2ngeNQF/hjnPSF6vLt3OjQ700VNworz7YsMhzGgpkcKtZ6
AwACJiHDp42cTYpwW2eE13BfcdvzIWTg0ieZO0qI/Dy2mTR8fChJwgcmzVydV516jiqLyl1Wtmra
oPme2SVRS8m/TypwbIqIQEYxT9yYMkIcmni9kTEcc/m8BLmBZucUdBuf2OAuHS/sqGQB8c2P8KsC
AluYmLDtffA1Y7I9UC4AAhQpJWDN7DWcksixpnoGqXW2SCXdMy5T287e0qyW/7etiIr8huA1yR26
xA/UdGoxdYiP0MIFX6ywPaTDkiCXX4oHw45McennIAq0jAZa28uetki0L6zqZ99+XPxyySHeQPRk
ovUo9C6LdBog8iCC0nEsfGf2M5tT7qOM2D45EeTGQwXqBA5loksmy4E8Zq0pfP1xNS3AVh+B5t+m
n7CdFrPa7aBpZ1zFSVnuqo2EEM5dNnwD3YkeNshih3DZUog3zO2EEGqUpCMX+kb/82olNyXnF37l
5skwTjsq87D/2Qm7yFtspVXZ/dwW26B5cLqWBe9+eET7COeU2eb2RcpXFsKtKWiaEPLpTb+p17P8
aCd7S3YVbHruaIuipmUHGEDOi0mXbGZcwpM8EIGl866oe3vGAX+qxSysrWazRLX/NXMW/B6p2BpG
UBBDgTBAa56tNIt1c9Xb3p542L9sXUxsMV1FywUUrq0HN94Hyqw+rewMJq0WQ7qHXDgPmdASOLaG
jrd8aLAyPPc9SHKUwfzHoG4xOD5WbG6fdr1YBnmzr5WQkQ3CjWHg53YKfFohpox3n4tDrmyenX9g
1qKRv6XY0BsGKSsdmes/zu21fH3+opWH7m+WYBb61nEvNT4qTkFHtN9zE0CMBAaXPuhcAfTsxocl
mtYamboSvpd6zaf+M6elgdlxLmZLFUUtwO/f5M88BLlKaf7R20Qf8gmAYcHc4BvO7Wu5TNWg17QZ
W+uZMafvv5JHwFgnN4eOPq8Vv2vvA6inP5iKxym2WlWaLbUS5VyfELUClM5TsoRhBG8/Q6RZpCa9
K+XSZHibix8GxNdjUm4HJ6noTXpvThLafmQeg1rVIMXgN5AxiV5jCaVhu3XAfyUKHRpHsaxbHed7
/zxMlnb7gsdwtv+//XfN1K3+ziSgbDK1jqBxOuWZEhYvANj2Q8jFXabJ9Ib9axIdEXZfUoS2dTxu
jlj6uiq4aXJfNdh2C/A+upj9hFEquIRBpfrDjnqQvCT2WGU10oYt/QeJByNVswtlnlu8fs/K6BmL
3Cu389qqEKxYv88jNGbmEkF0pO2grP3SDpKo4JLA0MisXG9Ys09ip1SyyOZgK2r76cb+ynQ0dOdJ
vbn0Q7fqeuEVzhCy4pvvdwvqYSlwWV95Ae9I1kq1GNks8GfOTwL6G8GZ0CT0mz0tBsxKSEnmOwzE
6iX+5/+gjsU3sYpAuRBdbnhJwCE2rMqwH+V/v+mzbRAj5ybYayo3nv592LOIy2E0ac7YdwHYjgiI
Om4W69ZyybaS9t0Y0XzHABLfW9q2Eec3EkGmZ3pF8VB1SIxbnKUvB7/B8MqJWFaaiIMdyfrBBCiQ
M7JEnXD4GHJaptvqljEYhizdWgyUmfaNqY5RLL5/MXZ+HzrFQ4K29pMXot/vwTAAJzMyNNTD7e4/
EBEGZ040Qik2C4aISRlHKANd7Tjov5Ge6v4enjczvmX5CvEdfyQdV7q/5BKmyDsDVid2nGYhtjWJ
Pnz1zfGoB1EzGkUf5hSdhNOqmpF/+EZgmGhmJ+SauM+qrLHW/PBrrKBHNVY1OX0S+WU1rfwjGFAN
YWuTZU5JrM1LIGvDlrLpOHCRH0zSEWrNQuluqhyh/q0XJ6wX59eu2aBYZ7DccG9krKRdQ9ZNJCjk
tQUZ4BVdCBavYOVsYCUUP88Mhv31//I2IM10mnfhZVPd3UbY8G7HrQHFLeU5+MSAV+tjhSenw8iX
4ntKXINu45cWz6iiLCDTNoqCQgDXncgx1y11PxXN3Lsf4p/xgMxaeNKu/lDzM6X45w4YI3foHvzu
A9bGsu1aFDQx4ihkoPi39rOASD5JSQMVcWKTsNBwznHGR2ay3sGGsQn6788JNR/sz1IWsPqeQi8j
bKqQeD0Sljdp7pOsWeHR9JqhRoS7fqySL4veC1zBLv83InYr+boLlWWi5FuoUXREWo1FW8AWtE5a
43Pr63Cq521fkFpENcjkhzJii3H8Jz10t+HNnWaFtdG2fwkLP4hdtZlGUvDpC94dWEg1bKRXEOSj
BId2gnAIE+HoA4OBaKUOfiuRdPQpDzRF0BT63vx5YK1RErLUt9L9Ac+N9/Horigmr5XD5omhE1bm
37KvbCg0MqNrQWxkt+/ge79NHYvxFRriHSTdzA64i8dCHseEZvuQhCfLPPUSqnDTuNGYDIEkDpbr
Fs5zqe5EqdRJVT2d6tyKU+LWjXdVEkuu4xUqmLAP/PSBpg94GQ+PIvNZJyxoI2yl0rhtsqXERlwm
pjhKvhb7js39tqU6IlDMWlIS9PfmCgtmIEuCskzjkHgupCPn4cuxF/NcsyXobDbS8appdGaXmwfu
gHqd5lQHvMXQ232CDoh2pfjk31XNfvqqpG2LV9HRpZnjLvyFYKVxW3CB56E7zZVe4RL/19t7xajZ
M5/3PC4zoi10pN1biIcYmm97F/3XJCayMZ6GSzdK2wf3yIJfMrxLCTdBjZevVtpiwI+ec1rJN9zB
fxSfyDwX0/GnjwhnZV100WCLRco3zPg+87TjaoCekHCNTUpqPE2MvBEiUXrOo4vahdH5kn+BYyIM
ubXeump0r6dBlf4orOAtSYv7XI553EqWs+wQpZykO2HvzlcDkya/bwayxmc7p5H/w+iYNxPQT8JR
YYIeL4VCzdx8UmbINhBD7u7M7XqgIk4z1sRek22PjLJ4mNqdXuStb/kXlZysVgikETBdiautiNNy
2V7+cdhTVgAQzsW5Xrd1UyAkcCa6KNDr8SAflQKekWDd0Qn5gH2bHCD4LIuby1etPdJD5Pe/PgM8
1v76TjpMJPBLQi6l3ciOkiisfkJk5OoW/Q+tZ40vzudVOruf3dRjpiO+nfCwGlSNEuT+ewdrgw0n
HjFR8OC2O+SHz4GrP7JFmCc/gl2IDRP8aKPW245Vp4SrmknRf6hi9AM9uD9Re0iYHmtUnl9kUaUf
GZVzqEVGmw6DJqaXPuF4P7K/UG7o56e5WK/zh3nLQ3P01wJNU/7lvreN5EH1Qh27x1lO575jcKOl
+pIb6OGEEavCYq15e0A5D6u/SExK0X37rxVKp6UoBHPe2u+ytlapFfrKx7sOWdZ/a0000ssL9lUG
hWgIh5Q1bVPk3xWctTM+BN3kh3pHfnrOAvSh6eTUzrQNBj5PO0WHuFbk3VY913+ggON0oUbGKBiZ
eeyGxU1I95HSaIGrKsr3RNHYB8dNLeXHlDrhZXA1Edtjk1w8aBqFp2tv5n91DI5WHkLQLtT7Q1Y1
PpJgNwPwtz16nCWYZhrcwo7K6SUy6sN4DHjxRSL+HmMmUqm48GY3EmMUDRXFBr2kX5GFlxjaVTlo
Mx7rMrqunFJrpBidyPhGDSLNiMiEvH0dcL4CeLoxEV+ZszZcCd+kwxBFQ1r4fRp0GUXlNuyyR6ue
jkx85iKcOEhZR7WRZoWvKn8UQdAQH7R0/gwQKRNaOpr7bwO0QRZJukqNFCd1UGt0T2vzhAQ4MYUh
8f1jfekpGHyUtNbVpGB8ZHOCygXUutaVZVBB/nAj+u9rcbWqgUoiEz64s9fdcrS5v0tEg8gbBUCY
hv6NRsPiQmspQZrCHzmiOZtcC78UkF5ENQqDywc+4Jue/S3nSN92+S39p39CRKQ9KfjqCCujbESE
YQ/uzonwDipNE7rmQyZlp8Q9c7nKd8bo40YCqtZC8ufq8p91MNU2iMiDaBT9E8HN7khk36qV+LSy
Xbky9YTrTFQjv+JVu5oDnl5HpD8YeBDBcEj/4RVdJPqVyuHZccufFG6bl6mS5FUWNEilDmTrezba
B4qW1Mue2v8RZz0GSjNiAqGRtFh/Z5usBdWII5HCmrQpjLehCz4J34d9+Xuo02bYXTEZAiGEoE37
R1X0bSpj4U1zb3fLswuU0unP+zw4VnDzO15VWObj2ZFYqQn4esLIsSduyPqRII9Q3H7BvGlEGAbP
ko/jvpaf3EMirvdEDmM5yqjJieGrRMqU+NWt5neObcxx1UXBfwt/qlX3ICUWgCJZnpW9fZTvAx6W
OQvZwUJB14CQIlTdjzF1Ejo2BpevI7bE6bEw4jFQKboG1Y7/hxuaau48DNpG801SSWLSxBGvieB+
LLcvV3vsjIC/ePAWUmIO8gyxFFsa28RkL3pHR7BGO3QLaAFCLQ2gUbRJy4Rk32lujPinBT4mHVHW
LNxQqRfAuvT+82ZPt4eHyBwGrGYMO5CETn/cThJRSErMQ9WANPylY5CmGEdZaecM9QgLW40THbOY
seDloCrFgFDubUtaR90mtDfy4H1hK9aDojs5Y0ADB79kaJuTV1F9XWhYjakh89uPD0lv8NVhutU1
/RHHT10kXmLx15WOJIJGBMN1UkbP+X1w+8bhFF8HyrKo3TdB4tr8CYRWmZScEoPcPBxfympPk696
1cpFrFfutyqCQZgTTL8QwOndt3dRfkV9F3m4ps0lFQNtaXz/sG71Tp56YPrNoeZe/sdqqWGnONht
0QaZezfH8Oc5jA6JvR9QUl4FlE65o5t3hv6g96mQ1/GFTqySjZ7hCrZRlEhblOanMZNI79AW9vw9
yJbAugJCTgNgPDbVJabjmj1Snt9ODjNMytP3/PGvQc2cAXu/PiNLUFMr/tMBXNe2+Ixpn+UeXJJs
zQkqe+VlQtX+j+dUAADSiG+O5dyW1fC79nzUuGezmtGeyckQC0ArDOvB75xNMGBOivZrIZf83Qqg
axcnj3k/mr5tqo7i1yiy7Be625AYuNNXsA9IL5nLE1oi2QCVQJ95jTXul1cFkGPOJwO7rUwpWB1G
Bf0YsyFI+L7v1VoxeWVbz1xmeWsMwkJUKemHVmp/W9+g6v80PukmQCwQP4AMYW9bdLNNb1RAGn6K
nHL//b3HIwbpiWlVd6bxKPI2/DJh7T5a6GHumpMzu9k4/p8gJON/WFAenMlSJqviZ8y3QD0WduIf
s5BhmxlVDqqM+kYYgWbepClTmnNvh680y49RLlHXHfxCjf+0qLeJXsMghPHlkKWu83Eji/2NDFex
sv7VGwlAZuJWBnqCbhncJwkYLaSxWQv37pD8TfKRyHaP6uFVmNBbrLOxCF3lfj7Do0ly+1ZJ/md4
Old3OEL8EZ9aAlgO9BuGee3oQ5pkoFcINN169A9xV4vgQlNA1leB8ZbGp/oFsUfa5jFGFFm9vihP
xzOladkxrKjQEANCAsDnw17Gb+ZU4QJsnNYqxw+FS22ubu3zW6457dCUewxN8O8nwK1e2HP95KXZ
l77HlcLieX8sB3rvUd8BGSzDPHPE8UiNj0wQVmG3+Q2kukIZ8s8d2Szif3zBeSTixAiHh6UDBGgc
9sPFs6J1Xcu9s9wMoHiHr0N5Hh2XPmtrMlFE1Kq9ho8In3FtvSOywujrM8KcENOTzjFJv7obMzzU
QyvlHZri4alJm2RCWikOD7q38DfuV6ifvIAys0OE6uUaU6VzgIigBNTek7B5M3kvHD/PG6fbFmOK
VOLRtvhLsX1Fp75RXOeCSTFdABZ6r1D1QKpY8tOOhAN88Tc91AgXH/sgRcilWu3BVPX/zILOj1Cq
O384kzuAvNGfl5v6+oKaIkxu+ZftuTKmXU/72zzcJXQlNVaisJ7AeD8iszkS+IZECcXZpL1UPYQG
D60UT92A98WaJpTWbXgYGR1px++A/GyXQihubPiycGheGKNSQifeQOfBcKeaAwzef70J1R19SSmE
zAhBdcOmEGMQiZeCWe/MYCYlE8JIQV6oRXHh+huUHjFNpChttXmPaXoU5ZhgmKekpHzsOgJD8R6v
ir8Bu+42uF30COpj0DULBXy6+9tYBCnbeufxhxk9xcNmC1iWV5tcjgpatNUHhtjk8gP5S1BN0HFD
TW785s9nyacfveUG1jZ3OqOS8+hXw0YhaFA7K3CEeYoRHlAoXeP6w1xWhxWFq5oVSNtYgm25/nCs
T4ltLfHoHouCqzrx8A1YMPK02Ik4tBWkLoAL4SY/q6c823TDOvbDU2K/bwU2DXdWFfeg0NQekLaf
CC8cKIherbZZ+kkALKSKopjAfZP5wi61QqsH0PsrrpNdOeo8M5mPnYmPi8qfPwlEIagCVs4MX/Ha
9tNpWZZUeATw8FWst/wNZAJRpC+/DFctrVFkX2sAvqJSA98s4ZExVNusXredMF99WJYQfqek3Osn
aUwZKAAMrWRjw02ZeazeCUcQLS1jtXy87jHhZNqNurgt65NutS4tFVguXQuVmhUapnK3Ql0BjNmS
bI+9p+e0U9TjNAGhXCSF9rF8jse5fYAY5T9T4mAfMsm5enzkGxpe3ZUhSIVP+0skTXi+thbuzx/r
inCxnTnWVLIVlzOG5fMCqequJgZGgUOudewecaHRJEz0RKCGjq+ETFv2MD70cV2zmLNMbjsS9zpl
myRv1uErBXZd6bLqqSb65fRXG0EwHGzz++V1L6GiWsZpqY2V4BNbQlYw3BDmA5Dry3WkaTHmquaE
EmZCW5It7MfEcQSLBe/Pys9cLzPwP5OZTtwiGUvvvqEK3LkJJrxM3Em3Ypsd7Bl9eos7EGrN88LI
IbwAF0kXki5qu+x2R+FU66idOKZw0OouolgPeiFwz03a4oen6KpW+6TPvQozMIp3FtWS6gqH3zG4
svIleH0Qh0S+7mukjonQ/I/HH1MDWDSYqH3oDD+B+to8d/l4ph1m7+fDBsM0I77XsuuMdr6jR9RP
8hkcrON1/yUODfdgsGHXaSZmdLx/JRKUpwZr7zix5DZLMdQ9z+C64WjtuDhlyBg+IawTSOgRbLhw
4Td/zVyv61w0cSg79WSRqIH60/FMmR/PnqYjWCE+oA16VgmTQGf0VsHDRkir4AlQnIZrfm+aN7bg
vKnrWean1koQ2rAD9QPv0Ih16gyTcL5kTktO4IOTTf+eAZNidcm73/Ya/DYZVgBBJA81wjWomFEv
lyudGpDOX4z3saRJIl/xSlE+grchltYKoCK8L7k9CoO9wzDkB4emZKeGfCW/fJHcPJ2eDUhlwsng
VWJC9ijDz7hRq/EDC4Xa7QOSyF8UNokoXxtna/LwYqcQkJQ/16L5ir9LQhyO8F6SlyAxepHHTSa0
PSHcpkXsxs1/z57AGTkb/5jrOjcRM+kh/tu/Uv2OjmKDzQHCZNHN7t8khNK2rejsDddjDxW6UNcv
IuILJfF0LX8p9qYzrhC1Q4XrJUvMIZPM1sy84soBfUSeVIsTADKMV7fb5YXqJ08c4q6LISlTGosg
VUNqrWGIyAQkUh0tFbqOgJaIAJUi/hDcQdCF/KflCA+4y7m+mC8zAOW/l2FdMuvvm+2EdwsvruWS
bg93nUwNYEwrvlZtzhFTSepI6YKOm/SAimhHsyGEXYfVA06CxNVxrOI3omeLcw0rz6ht/agA5z2U
rLNmq0a7BwEy7H8RKvzTuRLku8QrPSx/RvKYBNp821gNcjSAykwAYVE1P4EBsFUC/qiljfFqq/kG
eGNLfWm2E2a66XH22GRO209PEEc/IsNa1qJelabDOrYa2lcOwGyDz2zYqZ4wmetsM2RwRS2298vG
GM3ucekKjuYy7duL5A7UxkQaPiVm/bkraR1GenD78WyRnOFEVlWEGLsMtOlnUP5+TQ1gJSGBpnVo
0BVlKcJYWmba+LNx6StuSwZBqXYvxrYUgAuarM0=
`protect end_protected
