`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W8BTxozyUsN2F6BjwRpQ42E+TujraEVKRNxlVQMmjMjEwSUb+2s/9r7M9+9lqZchtUOesX9+piND
1wcCUUCy7Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oI/LTdi3eVpOco6HQnYXoyfPCEuo/LfAXbvrO0tV9YGGwVCn2CUNzYl3JN7CQL/xe4pLyAKZQaMj
HAa2pW7ncGmkLUidKmMK24fK1s6TXopE8cF7YxREGtgRC7aJOibofX9Ogcrru41CTCbdJgWCFHos
suR57vjMoIlgGJQ4W7c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bHl/QJUYlA/ScW0xSwRrs5EF1Jk46e66BBLINgQIFTDiS6wQLsM9W8ubvHql8w7h3EDwrvDybQzy
bgO51YsncDymBOShwtuoUUI1xKcF4+HxMrP26tcJwdDWr1DOjPZJvhn+yTssqx46K+ZLZY5JJ5kL
+JFdyogxAsyJ8pZHJi6KSceHjqKYqpSgRbG60TFe5iewx7soVGPJiYWNbvWKstrZFPmvUZRYceLp
JWJp83yJPrfuuIklMGOwXkZaqsHkjQNeeJuVyNH2M5mDpERHSk5ZK0EKbynVWx9OeUJTwN1JK5xk
xNdmB9KGoUNCXmPLRfgUmpjGp367VWZGqvrSDg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nJ45HTbnUaxsP5OcIUbGi+R3kyoohlxuB1IwzMnBuG9f6vydAS5bqyYwD/Axcx17UOHXWIZB/ZZT
t1oa80cuA7F0vNHqRo3ONsL4Us1WlC/zQJTR3G9zx4GZ7dbXyb44eoGMOS2vIFErztGt/M1M+09+
rrKNXvcUFD261fFA/nU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dyvaUtYZ9xilQ/zyjGw7jv/udjaIjl41Kz3OxJOVoVlSEnWNI/m9jMn9f4aHC/GbxsI2xkNakKFQ
EGOxvB0qNsnGrES16l4WuuaWrtg360YLYOHvWQRh/iauBb5c/JAN1fb0TQyX+7f/z0CPAg+5L3h/
ubYn0iWaxt8JG+6Y4I8ADgM8N6CzGq/8lJw4/3f6SxioSiORIzpzSiEdLNUAHWBLaigVvMK3vkhH
RoB0pQzlaI5PDkpi7SlefyeEcA9L37TBBo4O34g8jrraNDwjdJt3rXgOtZKAYLZoxx4L2OMqQf91
kxAEfmTV81CWBR7YiAWk+slie1cpyqBSlBiEGg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30848)
`protect data_block
KV1RooykKxUVVP22XhI6BYdwHEwv1s/Fayg/EvsgOFSdLJ38EL1wvzQij2QAUYLIOzcj+DfnCpBf
Uvf5izii8DlunQsARQB5UKzYZLAdyNBLGgl62o8c45tDeFnZBkbu1JNrwJ/J8njeD1u2FTNKpTlA
yThrUdrdICtyCr6uziUR/3NGcklzKNnx9xaD6Uuslx3975UmOYdjGvLbUDt4tOle0hHIqFUBnSE9
XHhJyNH2yAMdw1yoQu2rx+pP3MTPsA+4DRzLgv+CCvAEm1+2NsDm3ksPb4X4M6Fnq/tYxmDu/SNL
G0FGOkmcVun+ui78cI5HDCKU8sE2GM/IjKEBbMISkGDSZMNUsmRNP8rJDAjEhjdq+mG0nes3eXC0
RVmEAiI/W83fXVJjHFtiADPFaCUV8XOeCvdKwuVA0YFLEXzHqjjWP6xWf22Iqn9zSdWOzrNbV6GK
hvgTFQH9ISMKHqG+3NNV73xW1zA/6N60BACUpu4Y3Uf2IsbSBoWeU90EjBV+sJSaA/hsqqdcJ8ki
RnqYdBcrJ1k/HRIF8qmD0SAfepKmqHwUzI926opuQ2TIucOOAEOFtDXWANdrTGnwYsYnWOVq/NqY
PYlWwC2fEUUc3idjMpEfW7vk74TCXOqk+uqrdXRo76PVE2vvBAJwXdDdPfGI/mNqte0JM8HCyxPG
rrvQ1G4KpxwB1kETZlVpqFblDMxXavZJUtx2t1HLTo+lAut0i9jwHXUUbUoCWRSh4wgnUwzIuxIj
/4hqspQIRyW4rJg1wgA/6wiuDHZqRON9FJjCgDsfuXBWL99hqVqzTuCdWQ2qcCPq8ZuvBZHMqzru
6XarPp6XTJuYRWP6kgCJ2eY1UUKQA0f2QEz4FoLtCHzTqbgZuou6IHxxoj1hRWcWn0FuhgCibrGT
jxn9iOyPra98562L+ZyJoEw7HsCgowRltIWqxKlpiqolJ6w4FnH2MW10nPsraBQ1rSJzZ3PLEPWG
pRdRHBicF1jBrNeXQ1nuUUSgcBfHMbHVoXjSjZ4FE089QBTOHl2aYA1heDdDMQUaq2vk8EDpPuR0
CPjHDFlQJ2T5eWlpPeuRFclqzZSFZZBNG2Llh29PoWWisS+FAXuWmKrHe5K7URA06cl+1+dof99n
Exl96GgN97/fXCQiy1tRyauxolAVhkO1Ytm9qRWowAJyQCJnITFlrYvG4UwqcLoX6ZqIp9NFPGZU
lWG90jNJep1UjtHVf3z6ey4SNtd8TqSPYZx9IQVJYXQk1jD5uzU9X0TO2rQREc2xHviHUS6QSKTW
DXc4272oqo8VXw+TmzgQuNVAszCPTDMMhBQ25mw+Lft2iCnzjOvu9zzBwS0awkzs72c2GaKtR+wB
X8Fko8xrycHlmo6d6/hzDkUe6H6Hrsil51jp2w6/SU8wHesSgEJfeDzXzeBEyUKz/AkMjjxFkrNv
BKffimb4QxomCpbDizFlhbN3/iV1K7+acOCNyICPrpdAF44Z3JmutVLCu0+tZJojAFrMk4c7jei9
LhMDpNrV9BoYtIc2nPOsot0iM0AFI8vHmh6OmtNteLkV0Oy5SIlcOLcwFhLoCPzcYYFsOA2+ztYL
4wemKjeNgGdxnS5IKVAz/67gy0JYK6t5MT5U1Sz4QLtwXRVwIl2cnzbKCGFyq7PYpXiUk+xR6HP3
D6mYkc1yqcbEe1QNZTh59CvgBcsjPTbFlX36h8jKnolNGaPTWIPc6uq1LGVYK6i/lsCm5Jlz3zBi
KkxIA6XM4p7DqB5EzrbF1wc0S7vr1nAQcMqNb2MaqV2lhipBwC7h1gosRjVMiFpK/ETB1oBHY9ix
HyMVk6RWfNJ8htyT3y8fXpiP6a+btexSyGfXU53o28z5675cmhlghA5VDi1abUgSGJ+e3ObpGh8g
aLxrTk7xG4hArl2XL/6Mf/EBq7oYgIL01MXTMtkop0FnNTyx7A+gc1PUXQ5NxnCMDNJhYD0DaLkV
PDlXXr5gHAfNhYW9zPUOJHE898NLqpMQPnyBO4cBxalcnnbRXKT5C4c6Oc1RnoH+FHSKyLcG4C6o
cfzKCBEHcH1x2K/cHCYbwEiDI1RJOnM9sBskOTuI9/M0mDoWSML4uVaYFO+GF7T7eSJ7DWeJ0EtW
JoWX5eWmcaxb+/tobbyjm/fUo4Xy6UxlSaoQy9aNjkw+2rX8zsXEsnQYLzjwdxmSf2uVcbzhYa1C
NjHQ+vynqwGnIVMe56J5SN3kOKwVjCw2B+g/HJmF+4GkrU2artd0V9DQ1v15j8pK0Z7yNpNO6gOn
Xw+XesS+OxKW6f7nEf8UgxzHOf2JzIggLCvRKbCBJyqd/q77B1pa96eApLMqwMdvlOMMxGSlPNpM
1pRP/nhWOZixDxdkIvf1W0K4wRJJ3nOfKrZZ0FPn8KKiVX2Zw8dtVUc4S6x2GX98rr5F8TlIAr5q
cr7ZbGHCWJS3hJ1kHFttW6MO/cTHULZZYTGW8qHxFW/wqoclsQnbsEHl7lJqIL2C7lCZ6A7rd1Kp
fQ6uFX3UU4AscNnbjXWnnSnODj0VBqXeDKBBHOFaOHBxwzb0OGIjkjV1zwtUlBz1+0dPCzZZGobW
93LV6ZxTR44EdBrpCvPFoDKLAR14oHgf/2lybIysoFpHAS9DuA5VQ+daVEJojx6ul65cX0FKKrSJ
62K/is7K+3MPc6EAlq/RQnFc9HJbBmd5uvxUxW9k5ZVPXPPmrqRb9M8XRWn22pUpl4Z8CK+QM+w3
S8uvw1FhYspPFMY2pyWA9sT9Jd42VNnpwpBIqSXYVBh4l5lSEIaQYDaembmUNT2/UbVsRfmLEbWp
PI31NfxIG7Qczovoiu1s2CeaA59Qau32hzBOs6PiBCF4b1Ts839hKw9qOjbTozLQTURkBxQcvhk9
4uXwsZg1nrF3dZ62fip7dDZiwHdnxWMucQuDK2ji6qpU9hb9ud2s5MivZvM1c1BVRaRG3WNKzlte
g/VlYO0G6UbxSgjo8k82TipQhho/3dw7xf2MWqjoolzTR98JpSFDta4laGK+m5UC5zZJK2/pEbnv
NCIH05L7Lox2Hhgd0m7wZRElaKiu8jkCAD43ROHzfgyjqUYCq3x5mMeuIhwIVoyQbfXgPWfLRp+A
1+CAVrGfn8mf1TS4Pf0yzsMFUhTJdfz1n4s0NOROzN1Mk37GVdGMQf6bpUTUfVu567rHXtedM/Yj
m+MvdGmOXlHj0qlaOIh/oX2cXj9b6zP7VqLAvgqdu6BaG+e83NwPayVaDIMppjNs6QOQ3k/HaBF9
G7h0btk3j/wbXAFL/wTYeifkf99z7ctJtxicuNab8acglGiezsyb9bYTpbzSEfezRDv8t3tSpOmQ
sA0RVF1on0JcwwR5YQ8QXLfNNjGeZu559zwjeydGt/KlZqVJ5B0UfvK5fU3alGYPUEdjJ+n+Yewk
sfCnV1ljjRd2FtBQtylJ+tKrUbltlTqH80g22Atvy0DG6MuDt1Je3pCk55v3e+T+mTLJ7iWlfVIc
9VFh/XYqvu4JX/WpsWRbTuJn+3AnIvoGZ6XE06FlwR9WwC6uwTMTAuU2BsRC4JM6aYhYDlfsfIRB
N0NNpiwyen9Rewg0j3N6YvF8drfikheaJVaVAeEiPyWHOy1nRcdzpTMTDgvLKeO4uSp3TlKg2UnK
aNf0LEGyAl0qD9KukTV4gGM/y4qT2pyvYGlqtSdGUrP2vDdqAKiRVTbAMbX/pq4dQnhQX8/w32d3
VoCTRSnwXUegjxWdEU5dDF3MOKYMFAShiTOz0zb0ZaH8W+kQFXhyMvBGq46Avns6GV4HumDjEiQM
kvhWaJcgmFEwWj0kvlDZ+qFo4t7BCXINUc/1HoRizIBz5fZcwCVLDlXSMJBVWWeaPEDotXQATBXs
rfMsDsnCnrOiNgAVd+XM/ye1MfxKJQJ+5KZZof4kO0pG/Jk21JMYY36SH8mbwqkf0Ztmb8k6gEqn
KGM87Omt2FC5UQiRKo3EKBGx41Ru2nKO3QJ3VIBofDGbU+kdSgHwOxdqTQFqyDrWj/4k+kvML3J4
Y9+/I/fp+TT87ZcDpcc1tIil3y1fNFWhsqLh05TJgvhozk3z73psTnCwuD9PlSwbD/rRGcCFojjg
W8Thw0tW2ITb5/b4LuDfydycfYqQRw0Ojw+k1qIodNTQtZfbMRUKDF+Mnc3W8rJ0rzdWRk3DVp+m
pY1yOuKf2Ym3Hqirqi/r0hcIyHzOVIqGaplkzOBX6MBxAa/tokXBrw7s/6YpuqaqLRKjOarAB+dg
VXxoCAXQMXHXYVTLrjX9HZcdKtbx6FgfyFfMnqMTd6ffFuq+7jnxuldig5SUD84gRLx8MAgF9MpL
VQ2U5DUOSIRJjGYmy/W1IVGcSXUCDSoBnUUlUzH/wYAexaxtzS2R8EutpToZQAZ9dZcVw5tBeXAH
kTiDxeYhOTrHnHTvKf9oyJHIWLsrPknriv+sSsHmeLhR2AHGTKHPM4AF1TedlsfJM/E/nQaRxP9O
YcYtOb5FZFQbEi3dg6dNYB/3vbOVfv4lOBOOvj6sIzPg+h+eywjpLXBS+chSHMreeM66wE1iMxqR
huaDWS3ATZgfhNoSXOLrT+3I7S1g7HTopNXUXpy0/JTjKIX+XXxfyF20QQe8D/keRydINdNfMeVB
GpPv13zoctZMZYObxN/cFXJ2dU7t9WT40yBviS0IsrSiDxP/ZyCBKPihP6heycO3l7i2mXhQN14k
djp6H+3sBxecsL+kaZ/56/rd/gX/9kcHfQ/33U4eCrzUrn4uynMaKapbvOuPMp7921JmxsvpwRg0
oi63lME7toFIj8RLL2uJNBlOmgD0j6KovslbI27Vw3uZ6874d7q2ltVgR9+meyw9QNE+gq8xSpoi
3ltTVNPf1UnTCFoWn+2IF/D5ycghRuK9XhuWp4Q0I+P1gdnJFDlgKyKfmVHhyHSGTRt4zovBXBxQ
a8hAe4SI3PKPo0Y0ZdhRu4ex+gv9oauy8CAyuEFY0QxBf1SQORMp+L6IACT0w04cfvOcKXMQ6aUl
Y1mKQjyy/tqQD6dnB6MhD9SMUF6ALOSO4laSDngWvXsEUlS9PpsFRWYXx1nQFnz7TWkRCVcaFjMf
gwHnZVi0WbfX0kvaRaYzkTFs7MHHEV0/ORXkBifHI0/3MofrA+NCr0VJCx4FYSBHrctO2EyXYcnm
FVu5LdK75+p1MPkQ/TciT/mgDPLiwstEAGBnDlHOyMUwjea77so8uCh+e3BqeYO2ZGmhYWF5wjfM
40akdQD3/e9hvAnhzk8vGrE6eRdschHhVw+fPv9Ksuw/zWAE2rvTvoK2rGWWdGnPtSUfEwHmTLez
5IHI3oMAylVttlKXz5L6YGh2aY/W8KpCcm2aacvMq9Big91hKo8IJiQKYP2o43z76GdqU8GF/Els
XbPnj4QAcNb1pWsnQ5KTyzB2DKe77rZK7p7CeRiFFa3WCxZDENovS+VBVR7r1IO2QTWq+OJ+i3wV
ndNae5WPKym+AOj8eMZBYkpMASCJWcTVkbXDOSG5DFtucOMnsywlGujXZfPHnVov8WaM9fj8TGoz
SHSNsCMPRMXb4rPE7+sF+61V9C+Y0K1+NUq3Sxlu9z2SU/vOAsHxPyQROGwySf2VbbCzCWs0aSPg
6l/fKqe4pTO7uIUADjRLplI1fQbrDZDuse+Nw1gT8+M9aqn1vKOmFFTMtr0zRQUd0hxoweQpjfjE
HirzD81RMGIgpG4B+aqvu8gQrAI4iaiDK9YZBkAhXvAy3UZiwal8wyFxc+y3KAt/nZaCUrPtiHO6
hCKzMXXA15NJGd9P8/8zypIp2BL2kHRw9LsPxXJhYvX8e/2mrhzVUcDIlnLOMj3R0B/x4CpEGTye
fD5OEjD8tqIhBQNHMeMxxgwofex+UhrXlzwiqLV/OLFjDriCOc489t9KEzAeFiDXA1SVO+I/2J4B
lLfi196UQATgWVr9exksHFSxUqvwNT1p40R35DEzQMm51SZLz83h961L5JUAet4BDK/JGmYr2l4G
5gjQ4/HMC8d4rgbs3FQBI6CPhAqqhkNMrje+FFmn4OCsqFWqlemfuJO8bsggWU1q6ea7/plD859I
15uoE1wPZtt6+5v1cmyU61vhdNWdoWR0YIIFD9SezMVUILrA4C72nSu9liWBgcdJTPt1x6N07ZaF
27/bNu8/b2IuwLBbu1swGd6aUQiV+D9VI2XNRuMRfK9Po5EfWKOmQasT1u4stengVrAMEqLdN4gV
C21koMol5zf0deF+RVAYSO1uTxlpEa4YN9JANlPkbk3hvG8SiL0JCiuyhemHRurQWMNI3JVrE3rw
frknRzmtCTjdW3aa4H16fM/lUwzNidJeqaEQRokeI4dmaq2v0RWP4f273dxD2nyZ0dtIXlVwQnhC
S4wZeAmY/UQQpu/wcL4+f73Un7cqPJAzR4i43sKDNV/Et1vXK6f/ScrUnidwIZgC4pLkcJKCTDYi
sYVSzQ43MTXVsYPPtX2gh+SriyX94S76ekUSEJKi7JmRvl58yBGlikdleqlR66Dpg6KmUekcI/V/
Ze1lCFi6H1+rmVjfq9zYxRj6S0RjnYwr4WPqVow41JcKJ20Os5lnkBM5hPwEUO7H0iJ28iPzQel3
xy3Y4FIh1v0vkyAGA+VryJmlEW+C0O7urbPQr0oMCD4bJTVGnyHNDfe1Tdc0aYwo87KNCMV2eGvC
atksv18Wx69huYefQwiJwjwF5itZ9U+mUzNTJyoPwvSVfDzpKoc99BUUig5R8uScLuztKCp5YXtf
jxivKd8lvFm9aE9U56Ghti/RbohYiP7c4vTkbuSJlQgmJ4ntPvTe1ONQNMDa8UhXCs0+HtCczPRv
XHH6mMHvIzjjJ0CWmO3xAd5PKd2YT197uPS8jNHVBnX3oJjuGNAvq36ORsc2OU7Rc8fJqY3IUF7w
kA4ZyWVRBR5+L/9+DVAMbtR/BBNjIhqGwxNRc0K4+hzDl0VDCCIcOO8Q+rQO50XYUP8QK6DZBAgB
vs0Zx/0mHrJxsta/Uyp2Ae5IttK7cezbvjVMj0G2X0/lInJ92YhWlfrbCkjUGCtiSIYDb0/bDAWM
Zs4h6PX5HB1EH7kEt3dfgD4xVg5JOHb4eQd5amnj6qqLxhDEN8vbFD3mEFwgNSVmMZMmTcajs9MO
vYrWu1Yn/SVa+I0L9JQ35HegRaOom+muyxCD3KjeuIh6y2ZIShEsaXamqjpMT53yOh93jYDi491X
stjdTizKZoB55usi1sEuB00jtLbvFCrZW6Hy+UvzRR5ksBi5PxryurU98SoqbWyOogQRR4FTyNmV
e4yT5nZ/m5kOAiRJ6AJw66WfArK/g0A9P0rp3ExUjLhr1Ar0ZkgU91ItjGuWQSwObXHXXNoi8OmR
TQcp15zasrVBl0DCW6fD1yVvSjTg1ENVZxUoU0apb6zIv89CdXsdq26Tb7ijFaMJ531Ns29gyWeq
IT4pzJndezXi3Ow+mrwA/h+d4TGVfCcN27e6jP8ThuwyixmDNDKacUzk6HUKB30PNvyPa2BXzYC5
gLlLkUTQtQ0l5PnA6+/Qf/e58L5G2YZxHkT0YYRT/B3QtnrisJ5CyQY14JlO4GjDMlPNgvTUTutw
ydkh7pHNt/pQVZIU2VcoBxZ68x5yNeSi/mLvJjXvG3VuswyNuw4EavJ/Jcm4XxIva6a6TM1tKfTl
2h+WzrbUCRQ01wd/nWzjnLkMWrbuHqjLodzrX6+Nso22qeD6aY7iKzkjcmaHDHHALYnZFjXZtKyx
chF7XbqqD0gsPGryCbZVcUp6LGzi9h1BksLMMYLGtD6kyylJ+mb4511IBsjSNIZdWPZQK/yMaLs2
kiHaVdJRuTkTu9vAByW5cVjsL0FktnGnr+XFLcpLilTmS2+blH4thWrqw3WQa0fEA94t35Ax22Af
p9WJ3HfEgziSaFT9C7xC/uYjNDGoxqdBtepvyU6WJhr1TCE5Ej6c2W0xkqUHddWpHhVBxOpfyNw4
GVUcq4MHIardLtiqO9DMF9SaQp/kVOIi7TFjYybD2oQs05AIiEyy3ATzOn5lZ46s04IgPRkBYN2T
QWtw6F7MdW8p4p4Ox/vxcXEUZFw2JaAC04RS5l82cJtyF43pPs9iAodylprrIYsurIhPeZnsvGeH
bQu1VngQLt1l4TTPgxXMYKHrT7ZcnMYSEDToOvRlyt2kuz9Tthm21TN8ZIe+ndtq6TT5r585wNzN
kfPTW1qHK67HFVosRVIhl9HpS8t06LdKwpmGbCv3L0wFcDHbKDnRvCw94GrOrizY4salRo+Qjuvz
w9nnBvYZyjNbzZYHOZ21yfXneCULWHT0vQgHPC1mbZApM6J8pOmosgGUlshOxzN1vmAv4A457ZMV
DUy9VRds3XJl1mqEqWluXb0vWE10WGED/83ZskFIyZ6iliy/oMhQN7uTMZxf55M1xvdzA5XiUSqm
RUHB5/Y8vsGwNLeq5FzNt4jxOzn9aQMEd20t01GoC1oHwDHL1ltigF9YvjPBL18n4OA6QSpW4bt1
f2UJ9EC+s6WusDOTV0Q0c6h69qNFLqSe1BhdLzf72E2AbyEkmgCpkCEaT02C+nabUeB/29K5JPkl
Hd1mtBr51NRzxRW/nyKX4Z8m5zPwYCzsbSsdDyQBUYfERUdRScoFdavEKzRLdctMWmmGhg+rQvN4
B8WNJoBC8H3PQb4rUsiEIMxeWHyLnF1HN+EUr+hhFlKAiPwn15zrtd3z0UWtuJoXkuuC+qALAbwj
4FBaKQRpqRwRhhu+SVAZNJDKqekE8Pew2Nr2tUXYqXNpb4frtcwOlYwmrMX/IEWdSRImddDv6/pI
PUt1GC33gRXr+nsP/z574CVguo/Gbn7Rx7yfEeDGhKkig1Eabn/2yuNNVA4eJi8wrYcskJlRmQ6g
sbkgOBJ2Q1HDonqoCodLIuCReT+oRRDHwFENq3iz4GL0BEHGrL1Rt5Vt52R4BQqzAqfRL+BTcTEV
fGB2ksEoH8RBI1p2eZ6yHGB2xPSbsUFzc3c7XHWtd03yzjoli2+vD5Xk3xCThmI2dqlv4v5GHgc+
SY1F6DQVOJqMKYYEorFP+OhaXe/hnGhcJFiuuQeCdy004PglAmFTN8nDgm2iVTUU0pTuOVQ5a6OY
T2lr3MoYhqIwbDXwLfOgJg54TQf+60RJ5/L2z5DtZhYROFJs1MrUk8ChMVfVym4drUvrjEnL9SQ5
Ll8T+yayL+EuYlcdtdyDDwF3AqRBnqH1CDvEwO+f5hU86htfkQ/1lTgVC2dP+lRXYt1TQ4jb5D0a
XuvV//Wjm44FjFNIHcO7tjfu0ddHvIr/8xH2dGpJczK+M0vLYy7TjEqh/wIvm9wcm6PAxMViU6fs
eYShQsztZ3yzD+L2Z/rIJqGeIgl6OE/HcI+J7VETQmvjI6QmtJ7gZ7mbMfHkZpUesvDsEAFlfiBG
wmdM0RDMT7XNynmGzOq26ZTb9JkLaXS/bb7EHNjLj4EKT+zkOq0uS0VenIhDScnw2XePFRUPSpMQ
xJrtnb4rperm2S8eKBhp7IBO60EYNCMCydls0IS2E56O7Gl6LOsi3yhrSDlhb3qZUeZcZU7EZVId
7s2Iqb19YI4UktYB+YMnts67S3eTIBosoXP0C2jsLzJTCQdjZcX8/ZcWVWNP1ezLSdp++i2/efM9
ZmtwXHGONHgw5WwagKapjmpZPr/u/mpDhEws4qsEvV84e1Fey8FciKasG6sHQHM4HYP+zhRNvtgf
QBuGv06lNYOdhWbqrY4VLAcYzVmA/VETu/Sc1UiEUJtuIRlmhhHri3FzxQWdxTdpyWZ7fCOEtlQY
irUIOmsHtmCnp/1Enez56GQOQfaDYrivuyDCH0PIFJ/tOkD8Yx826DXN4anED8tjDXOAL158qQdQ
MKpKTYiIGy5E7p8gmAa+GqQJVrv9M/4pEtJ1aNwq+AmOOXaXcEO+ZbPK/XccEwsYpcZ6SciHbL9p
eKSpl6tk+nVtuM8Wadl9NFk6gV6Grka3LvdS7p/+FxypH9CEeedFD2dcHqUDtcSgE8YDHM5qDDTB
yWi3gAWpJmS3eHgDsmTenTJXvtVAm8/OnYlSAaaJ8DJUBJnCQg+Lc20AscM776tFuUZxarlX1miS
GdvQvhUUNQTiDQOOeZhviXTO8l4SGHR8z4xWqxosqsaz4xmnKnNcreL50IOzRFx/qP5wZprEyZpe
JV00FlLLKrLW5x167awZ+6lFn0aO9rgMIUgY5PAtRQRvQ+zc9aKGdG+J5tKLwM6QDQCCE6jh/ARl
zf9Vrf9S8xTXDYVzjF4RC7Q1DAcb0oJDj3fx4Q/gXjxWXYJBrUc5d3dWWi8esO7TVn5NhoVC0tLc
zpA/9B5ZEJpqdjKgp4bvTG2sJ6/zMU1ffeuddJ/xHJViQcaXVEVZIaPEC7zPbRgKCjg0aft0h+m3
0EN2RLwZbLtGnrBQb6RVFGyBhmHGpTNIXTeNlgq+Y/pilyu62IAQAo75mXR1+pI7gPrTkkSfWh+j
oZF81L8as3fBm46LtwFPxZCEILZ4rS5ctTIS7aoA7BtZg/Kjr2UYwP5djjoeDeMjTAGnDfO3JYvQ
RKkgAuBw80iD12I51tSg8xZHgc/0S+mqIham7QgKloJsoklhotIiqlJ+vqmbE2nqjzL8XT56sHtC
eNnvoB0L+/vGoE8Nn9C1Jku2yAiQgo2l6QKxdr3h9l6TIeaQd8ROZPspEpfJ5766DZ120o1pN/cY
AC3l0tcacLnPytQ8ms45NPt3Gxe1CrZ7UMPk1+KihQjKV3lDiN+ER7rEsLrkji8h+LNXGSPSD+/m
WDeZ7MVRIuud4mi9HkSOcgE/CclNXEJP6X6AdRLMeHDcNJPz5uJoGTdbXKB7iYjEBJYQxB9u6zq5
jqM1UbxrZnpuCTeZqSeH3WpOSQ+7kmE2vziOSPnwWqDK/e3KXJ2glkw+dp9Kt+DF6u9Pog3rexWu
3UIGjjWDgdrU4l0jcM1JEspqddlmyru9BYdyZ0lauhGOHltP1I5dT6Ktp0VBXfiWnQuaZje8JYG6
gGH+/7zG0JqmJhHwl5Vbw35f62KZ8RrV/XJtcvmLDANtf1t1xk0o93NmvbKlerfwcZDIAfLgMA5p
XV5oDZwpxMMveuQanAMfB1rkmgFHcfzXM5fAzhJQNo6Z/OA/11VA4zYs6zQ40SEJDXjfvaYGhWRv
n0CGH/tGOTtOGamligxGJLbMy6Fl28C9RGBaCy3grUSFc/AqzNhjjbmPO0vIRmv4YeCyIk76nhaJ
FTssnZpKBunplXhtNs3TQYT8RnEQFCkFUFOIF8QKgLnw3J2N994cvheCxcMjVBkpm6aVmEtWpiz6
cZitWPOC0WTYoxS2YMTb108rct1hyUgFxiAJoEW/4JAtUhvQsFAZkcVOp45yIoRHjDeGMRkkI+g4
7JFicXyojIUj4RnbthXsSPOExCX8HnYpBu3l6ABI1Fe0lrcIZDVs6NaGIOvyEVLR6yBo/Q2YTyuh
vP1uJeQi4f8At5Bq37w8KORCvxB/MQAPyY3sf9GasWNU0AxL96/jaJQyMFhuXbS5l9cqL80TKU13
URBB3XoawQrAib0zUfa38mkL8g5rL2vAKI8eOEVUQZYbP73C79pqOjRmCWRseFtyh17+lrNjRGH3
aO8DlnYok1m8bHR8a7qErTUhUN0Ds1Z1VARzTxTZz2HifmMwDQy4LvddonRCV1htlreF+4SJjnVL
PY9xLHiqRLUTwS8JDZt6JEytFNq6dJw15v+y1uaC1yZU8n/G+cwrCyou9e6NXUoTmc4Q3k5YzWFN
01tPzV71lTc4t4d4jllYEkW/9O0n7UYmJgG5fIvb0975DNLfJu1tl/4XQZf9NyJCTk/f+7s3bGRh
6EgVz4SZ9licOHzxT4AiGbL2L+FAJcqG6WPVvcbYyjW+WqIlZhTS2lKEESq75YrlvTH9C2g+CdkK
1Q4sNy2V7K/IrYC2b0/RBYOR+OAnohZdbri3AF8otQsuaIbIwwSaKvfI7zXkVi0n4dHAd3ufP0Dc
oWOk2nLlgqQB01bRrKGnqqB9QJJViOhvIC3rMxrrSH0jjq1X6LFpPiPEQ77L1oPJYC94zT62m72O
ROllxCgaOTVHflPlNXD4yeth5EKGwumE0zF7UszLt8ZNHKuNXsVW0/zkh7UOdWX/pwUK1BpJUXHH
IUMJtgqBywZZBVgP0G6bj5AyTJTyiJVDazlCXVDrBlGcGD/lt3pCefpX5IyPU3ZaLfdLHzGblHgD
erJTWju2ValOzUIt/U2SysP0SMGoeEs3yO39kfDnQMYMlH1401RL3SWeoZ3sno5305L5ifO8J0OR
ILkogAe0ek/Mpv5VPXfHh7PUTBis8iW1rDDRfe+7gQAaC/BPGQX6XhWFh1ifsfVYDjiibFrFf7aY
Mph/GIYLvGU3LjVVNGly4myZBWAnRVcTNcNtyjSVDAOz/xXxwWLsCveZOezzZ2Ws8wiaxIX9o8Mn
qIMpIUz2XMtEyp6pAABouZmkmHF3qgd45xTfl5NYQWGsD0VIRnxSljIeKH8538ndBd65jjs/uyk3
OxRkAeuos1ExlrmM5YD+eB8KRRYVIB/gmSnpoigmsE4Bwy+BF+agb1Y2atAgB+jWU2k7EV30K11K
7EfMsK72oPgISz3vb/XfS8bcyEx3bcjpf5qTsZC4uk0X5sGm+mCNLq9HW+hKCrQQOUA+ktoPKPlZ
+aor1m++zCsH3txsQSiNRUy4m25UJ/T/9Hc+Z2wez/Lqs+B6PSCDgVoCmhu5anqoyPNtMJ7F/rfL
pBnRc9Ltvr5HpUMwfyk5oGRTXisRHS8bw9k3Irj7ZVytByiyx6BhSAFST7UkzADZlRxzvm6Qfxvw
QLeKYGQoZas9r8ZrdP0hFf/FsgDHAfpAl8Djk/0esVHSbfbXQps3v81i1v53J3vgirdfkA0KFu9/
xgW8kyfLmJ61uBwt59c7IsS2s7WRLcFlnrxAgT+NdOvBIoNAE9AykKfiqLEHM1tUIbo7PD98HNLy
DUrhvpa6n++9RCfL28tjfBDpPKI23mBpgN1aRVjDrN8F46HM5OCQivdXyHsjice7Pn+D3TSLm/Hz
sk0vb2SWBCqDvG3F4NZ9Ee5BVsxHJGO0eJl5tKNBiE/LJewmCW0op7jTsysb1UDmWtLCo43tP/WR
FbSKqFMCXooc1VwY4ZsPBQD7wJdX6qAf/OoxKP/WC7NPKwj5YYNptgBYEh4IW7Qf5oFidax/X/Ng
zQvOg6Srrj9wMR8VFoSiTimMye889eeT1GHNmAn2hlsgtTLHkyUL6gejADfAAGEbCzNMwI7m9D5Z
/sGEp8PD5Xf6m2NC/KT5oNQqIJT21pw/c+TjZPgbVWbt0hxBkv6kXtlYigK7VdABUYwSQiMcYI0J
K84pat/R3+3K5WQfqMV0TerI+nXxjJSpGeVrhrwlf9+NIp+1icbuativgwuZ797cO0CJ8SB7BJgy
kqjd+Ejh12qIm+LMrJ7HbR4yh3MJaZHwkHcf8xcHWVVAc3DcG5aSkHPPGyl7lfAx1Ihdv0cCrSNf
9hWSNm8RZZO1AK/RfEA6iY8hiK/muPgK8VKWt8Q+Quk0Jey7Ixm2HmwUPiQ76Pj3rmEhMiVF3oP8
sW6LYie9HGtfogKg7ek2jfwnRfAtC3mypuoagu+9T84y3t2+PJJqOUkrgG3Z7c0XdRrTJRwj/wTd
SMTkRPcVfqS8KdqX9s+vBBYftXQsa/jmUp2Ih3e+zcEcsze/Q1a6RKwnjQhb0CG+mtHFRVZgiH70
dPGYGa5tYJN40KfToeyAbCJ2jbbSWc7q/cI4u6BVqWE6Df1WDx9YzbpN0+Gh8z7KlhUvBdLAUovP
Q8E2J7chW6b/zCg8IRmaHYrZKcahtJJVo5ESpOlJvICXLWw9TTSi9WUSvgGCMrzlSwsZCpkDwBPl
jtRDfwQxIYCoc9w7vxZ/p3FWd+DsbTnto2NJ691rBwIgVid1Ek8YhBJSYhfUFa8ImAS06pA9ogMS
AKdGllXzvqmo2NxgnLw52Zx8xkShZ6x1cU4cutz6FX4lYWVVbqBLZesbvNANkuN00ausF7nvKmVG
Zm6g5KOut40ycmrewHrg8qT6yRqKdkNvTzO9s5lN1ZMBMMoHa6afCsgwaYc332y0SsR3BZp3/Yvn
zxAAG7jJkTexW6SAIMkHSiErbukDWopfGwIVkpCYAX7/rTIDaFzbmfajma8QpUlYw00BpuU0/7N4
DYRiBCTEe8SJl/3Qt30XHi66iDJOQnRQTLvmnGPlRykyfq3W1uuEUwnO5AtxJQXF54mJ2FDQVZmf
1Cv5dozwa+oFniEgdSSK3GE/zzvFuUd12oZio/LN6UBu4OPASOxZJNO3EY7YWR8O+8mew/HGzyTL
gPzGeHf7NP0+zq7Q/G5AYOfTK3ZDH3xFZ/zGUm/+F6oTTfDRDRpDec5vwwX1dlQ4YLQK0GILtye8
hhCnibu/H2KMXPvLcKG/94k17VgUpV5utwanmmKJkofX6uSk46zmI3ixFgBAj5X0NKN4SewLKjMy
EkR+70LPKyojlQCzU/Ru0LzND6wtO4CgwiqkwCp5g4WZcL+c5/HNEP/3uQR2w3AXYZGAejNxrmps
eEsbs2K5I2qp5q/oxiG+zkrg1qRPgTvrFpRQXtJBU3FYwhEe0/HOCGjroAj56PqC0I9/wdIUaNd1
s3Vy1uJQHHU7MhJ49FGE7OVdVDgpm+vcu/svfNArMu8lD/CkTBEqxYjuYk+FmaFJGoTuoy669N5F
+qdOWBoYnMk94lnwZmo3pwNudB25hoMw1NMy5aojVWfpo8OFcgUgpa2lFx3rHn1otX+sO4cy58mj
RvVsMBOC3yCF9BH0TLtGaJqDnVt6+XpMTnDI22AJ21QXB5ZsBoi1LaXHPZbqW8pCDJMTejg0oZz0
5+pqQVWUs37b8mku0USN2/aj/K22oq3TtguPvGH4E4qVmWy6PYSaZQz+qOkyMzJ2Ux00EfBOSDHY
/q6x0TUph4ESqCU6IzozsYulsUIa7GvoCYt5SSWgXrkqt0MhTwRC0BEIzmgVGvzG2aIOcZ5+mo78
Ijawl9K1evWFFenskl8171tAtV+hZuBc2KK3s7fc2D1m1gvhJelfUTMPmJqgHptG0n0UdTmu9LNC
yLvNSt9W3zQuLyKOnX4ZgYXeOtI4IcABkriRJybM2wEeFQtE7IQ3olnE7Qp1ygLID03b7im9kynL
GhhW5yqgR7Pd604gzQ+EBGeRheOQhVe5ngcI8reUf8LOtBXmnwE8+dIDw2L8gatatlicwHloqgdw
/eDnFn7gN6GfntQ4KkCnLAvdG2ufZVqeQUHybVOYOJJccMc/OpjLnPJhmZAZSroOlg3mDGO4/Cgi
0ZMpWoQb6EjzHnQodr0xhKCGoshehEyTv5w44ooyGVjUqSUhcF0LN/nvv2zK0U1nvXjNUYYiY1Bq
Gzw3ZvGYrLXXtEKKVLSghIscXPKCxf8aEE7LcSFIZi6awWRiUG0Nj1IzDMyT7tX3TfWnF4oS0CUN
vpDLzOzwbMaTKleClA3/gRY4f1Ar7dpaaAdZ6s9Y2p/xUCGcAUprDuZa67444U4lHHTE3V4hcT3Z
NejwRV1JrgADrShQQsEAktJ3KL9nIZztp5DLV2iyMxVkZgI4hkstoOBNlJuON7ZqXYhnqVmC3DOU
Q+cqiCdnQVbyf6jnIlutTH+d5DKCsg+gb8RoIv9sA3sbm+oyt97Vof79+htgeEAn+056s8lARU2U
bcJSstMggBMx9HWNbCM+FrxwhOjHRk/O0NLjCmAvthF7xNBLLu4GAYeFVaE5jrTsm2ArupPJk82h
pZju0KFVCc8tXZoKOCNxBu5Q46dkk50gBP3ScdZZvouQRzf1jcTuZqsDcv3XqpNsOCKjYq9XK8e2
HhkKv1D6zGEZ2yplIpHheDMHJT87aLJdlagGXZ9z9fBvSKSvCBbbkmfHwDNiz08XYxdZS3wK2bjf
Lg+cd3DO3f6g1dyBv4y/YibHVpDwLCvVl8qw8JFlE0RPpr6buVTI2C5F2LGYU07P5vARdu/zO11b
MZxHxfR9u1GindjcoQXoGyT5gCn6sZeBznY7L1Kq3R2+3eOiQ9rHF8TQJCGdO+Ezk10rwOrM5FDR
Kpjl7sopSTJMcZVl/numv2NQWd7kPNqlGwJPMiynYLs/gYzWFItdt/yftr7B2JNo4UjZ2JbhzksV
PCV2creR6QHCjSahs65g4b8tESXjJD1ldzH3wrHOKmvF34o2SXkTkGOclJQAh/Rwrpb0Salg54ZL
rQ5L9Y7IaK1oFLj5YE2N4UCWGHdDJoPGSCdG6sCgpVuIHbvxRWR2z2V8NT0EUgq+oOHoUkIVkPTZ
dxKso/xFojNnQCzTPVQ23LxnrfUBventyo3m6eRk4Xb8Ri8bPslFeqoZJEwanUbc/QN7i+vRZjN5
cpaluk5jKlxtVw0Bw0iuHN9ydEmmjFNwPg7PqBpHb4xLy9ZkxgeQlagUZRfTW7fNR+ys2JWF/5Wr
O+h6+wI5bgnpC7lGoibC5QZ9GlCTRKFCUvW0nS9bVrwro4J4dyZYOgvVyFwkxtI0CmnPBNS1IlO7
uxOX5mVwNbXCCUIXrhTSFjNxRoIPmSxF31WmZawSwhu57U6mCcp3ryd4b2JdgPz7YNKVT9HuG4Yt
ZvY68Z7noD2UGkbXsT0CaoXsk+dLx/nc5lokTMNd/a94r18bNwjoeF5JhRJOUTTmDG99JGeygGE8
7gLUeUp5QGlBXyBt3THi/WIhWWFI5rQBuYsUEEPjqZSKnmTakvdnvnDsBoWwQL5b8jN8+/wragk/
ipXHXirVW3kVU81xjmre92UIOoiHVBkzQLc4xFdPkD3ruvgJMYIVOruDeZspki+WJ4UKKK/S25D9
Td+E4567JrFv0PA1H0ARNuABOopG1M+tkN+Tk4MAdLu0kjSs2ECWqYvj5i7qThdwKc5u5pM0sxbC
15tpRuSt1TCSlf3gpQnNvGTC8LeO21Kz6cwGQnA5fJakbpj/j9DismcfXQgor2wFFE1o+u/02L2z
2DZOrVT8j/tpkg2PbHUFJZOth+m5YBqh0cAr7N/OrwTloM1pi8Ah/qUVbfFvDutqwCVkxb9YsdqJ
4KfnRcm0W1Eo1MpdbB7YihG8wK3St8dgDh6GmIy0AuUoOHlRZFOx2wBM/6nThs+moHGmxrXY1Wh5
Jt+nsagdiwBozkOW5Jai5IKsML/ihL2QLnKCQrU8qUzAUY/vbv7xHLqoJMilll6p9qhoElB2XPgM
M8DeploBRcTzUbwG6HfPneiwTXrJsTl0vFIIqR8/fy9dZ3KO4V1GjluFZJ5m/ctnDE94jNKxSRYS
/vGZWJuUHhX+6MkF/gV6WRqko9y7FkSTG1EZkZ/UqahDC1T5+wZD//vXmQwx4nhHabqjODkicStA
TQC/JTUttbqLFV/LATqmr55reqLm+hTLi1Qj4CB115XidaN32TSP9SOv3V3XBKoq/82TPlmWvvy+
9E74BUjqawz5bQnJ6BH6nmwE2AF+NfK82vQRmN6PJpPMT8rwewt1krh5WS9xGwP1+Uy5i5FhiVhp
RnVrJJKnlGEXwl/fJIf7ESuPDa+sJytxzWfy/GT0xHDGAMLltr8994D9CrEiMAd2w1ZRMwZYm+rP
aIOXc+Om9fEMHQ6KY0EyRbASyBgIyX5vP6sTUWjvhztrPnkK54OfrMocLK0FDLyc1RDTGKQ/jncW
Tvws3cqNxXnMApxxaJMLX3PVJHs+rdxBPqJawNrtVSa61d+9DGY0zwTM2Qeb1pUWtsCZ1VpRvdD6
+Qvyewnyb+EDXFvQBOXEzj3JKY7DNuIFA2favVEdRPqoBQrCId7OqR4HO/TF5jVpGUeDrsXnhY+m
v0afUav1YGxy6R5E3BwHj8ee02X2m2KmGz17K09xkQYb+z+8jIZvwjyH4Dy+0/90XrhfIc8nUvYc
ZLyhSSMqKZVE0xUuu+wsfHxk/l7Mtbf/IAdHj7p1oti6SVnMsqGdlVbhwz4222ZQ/MCV3XA/01yl
dkcUYRA2Q2vnf0OeVkKgKbla9Yac12OlKFKFa3MceG0p5Jto5AjJiYQUx797pLM5svS2GN/+X/SL
5DEJlrZce8gMQpmwdU8JGdWWHJrf3fWSQQBgiIYdhpLEOswQnfQl8fLEFamcooTaPIScaALb43F6
ZriVAC8TGCSEk/zaJkA9lxTBjMYuTRYrB0reDa/cnP2mNphmj5K1vpcsS5R5140r4WlCqzY/dBmM
Y9tIKU6g6VL/Z+ZDxkw7edCrcbPJ35okse/Hh7Yx2IJ/pmq/f1ZVEuxWQYOOuw4/McPcBFhY7kTF
xed/I2CavOV4MqUuZ4Io9yNrbN7BscwS4wG2whxq9xuOFaNezLApXaKENZGeEVQ8PsRwWHErNwf+
SuFr+tkXNsfmt2x2jBos5c2u2X2QbgX9K2kOT1Nh6sh5zvhWMxbSYQAiR2oFAO1LRFJpQJlRL/br
U5EXPWzgSUsu+kFjGX5C95COsuTq8HG4eWKXrZzt5mIB0T5pLs8NFzZkBQgng/z5gHaCPs2szopE
xIaAekqzawjSFX3/uuyqeIfm+7/0ont2Sy86v/xyLXRf+Wt+3yZvTle0b+/yKsPAADSEmdNlVBDF
H8DQyigzqCH1u5JjLGrvZhyYDV5op4n8mcciprqH1Z8j9bOZfw/Yt580cqmHVhSBDFEeNgGHl14w
GdLH289HfF8pC9P3Xzil6J+GyTj6eqJRDq2RwjWdqglk05umnvWegAu+NSjprMktmYcrWFKOxtW+
30wmT/i2qRd3y6cf8OVVh84QWDdkdejHjRXvP9EWZjJBIFbCTusMC6md+uRCaCkLYjD8nfyv4WfS
aMbqGXIv1eI/tycXp2fVRxDOTCQJRsf3kDI31NDDYSMlj9XCJ61PuResmZq36s2t5rn9mGy5zHrI
Xm1XyLpkv/L7W18j5XC90DPWWE7tOEHPjzit5aS+mrW2AUfWObo1PMwSKN3ZAA254Npd0KCoVvjk
d3HCzcDbUW2EmM4bLEJLU+CfeC6KXXc1Jvx9OUw1x2sIi5vGYiW7TYdGUWFpFB9zSZCzMPIfH+jz
PncufGRg3LR4iaKumc0gjAzrTCAsdAuzKV6D0lomAc2Q7Zta6KpfcC1z1YGN7bSZxQydbNENKS6X
4sQzJIjLAWdxjWWNooV+/j1EtsNW+I/76o2pMGAm0YdSX91NETmI891e6PyPt3Wq7bVHAptSUwvt
aaFPvLKsbcnaH/oiybcuANkKpK/JX4ENRna3D3R42sv/L97poknW9/5nqAddzAmXfkreQT90gija
wwAQvQvHkZI7EKgAk/0vdB5E+hrnNBcplydx+5E2FJX2r3Ed7rBGRlyA3um4bqJ3vipHF8pZvPVW
8KHUgZH44YMUfFa7Yc8R5GfNd/wER9cWtP9S8wvOfWOEHwUfokPzvfp1H24x2EK41O0JTPfjsmQ+
5ComRvrYERr3YqRgwMOHK7mUIJBvx4Opyo5Z5K6afb3ZUeIppGz4I0ZoEbnjOfFxvE7Jyr1lVYwZ
1UI5Y776v6vc8ylzZU4pHjEBaDagoxMhvpEr7RRxhbLZ8asHO8cOEeB6XlxLQ4ur+ekauRl7UbXm
HM4ta9tBuHENDr1cyP6HSiUm+Ddc+uPSPdmZ5P6M5vIchizKd5gk9FFPjVeJujXsbvsbDUcit30t
ePoBT7MXHvR0riIjmBDrr+Drcp6veIqDefFVLLyGPSwbusEay86ajNpQHMDbFIogn9VWM+QgxQ0R
Js+sEu7wjcy5BPUPa50LmgKpSlg2yi/I8zRf3Y8RyGxKW64DbiNl0NMeKEvz5jD28ITGneSEX+NT
hkxAMLkJ8A8I7IeqRrOsVy2AEpn8DtY7QzJEmHqIbeZoyA4EqGNt10XMnxFm2ugDSd8RKr8LmocK
Jm68abYX0Q5FTL4ldw7UazQqmBFCrKIAnuTt5McJBIlzEDxh6UajPBMcg5hnOUI6xzX9L1YIFtnn
k0dTwYkVrwlEXwtNh0kUrfBccxlLRc5mB3axRpqr7Go53tq1CsGhY+umOAy/4xowAaryGY5pERP5
WwBs1poar5PHG67jTP57K9GGmalyinvSvGhCuRwy8sayOZix0wJ3LYMqOw+nqqkHoQPVekeQpgBa
6k905evqNPcx8M9W0ASzqXLIckb3SX2pL5Ec1938AkveahyDJzPAvAVv/dty8IisoQxMOxrqJML9
LZONwZ+1jXvwsc64utZukTODhBJSiwRyq3Nv5S7I7T///tPjqIam58i5+xHZEiHxviAa8TTWVhiv
tFcRZe51xtgbkiIo3QHLRoY9czpAvueFHbRv5iMbxLDUJaSoYuXXkU9CQF/mzAeCJn7uTsyVwxmy
GkIuWqfx4sjAMgKto9bOfHO5jfzZDFjyrECMRane5KzaKWvMswy3urlCJP8SkEEWTbwsoeGw5/Hr
10YjGMJOZFfFjTR8+8+Lp3vCd5GXNXG1QQOWJBh3uILI7ZqDH1IT+R0/TUDjYhw+uTJt9NOskjiN
oauHV427IEh7DYej79vcP8R6gmxeHBBtzL1iq2slLrcsA1NNFQSUTiX3ajngOhDoX0zyP7ZuFpcM
LTpY0WslFUJOyukFkgKMnsR3Xb73abRee7kiM0sOOLYG48+b0ap3uSdUuvySYjrTJJeNmPsyttJj
PpnzfhkonAWozyopWWrkdAont08gCit9a0UWJ2dFhnIc3Kp85YTJk3D8xXG8g4ycSYm/1AG7/E0q
f0l5D9DHPZO34Iw1rgCH7By6ylMb4E4pMb9Ldz8aublvIsulWEfMjUSxMm9XZLnkOqeFbLD3UjO1
IiYEGg6y/xNB+bUHJAjFY0Bi2y6UU5gPqTa6wFWm+sMmKRax+ZhEYaZOTlwGb+DemzZlVeKYi9Dt
x6tCPu8+w4GjkWIoedZJcrLDeDuUKLThGo5uJW9FNAsfP2XU75yWBo/TGhy0YKIgKcmDNtwPJSeO
uKmAKmG0YiXviLEw+89fdLsQR8jZluL9jktsjo9klGfPC+ybTQSVv4Sv0pKZwexusONWzy0IWH7b
Sct5kXCqbD6yghgJ4XUrX00ufIXAXf6/DY/zQjYYKZO9uz0BjlLli0xqFsTB2QYqHCXS0pbVPq+a
PWwmEdccSstLejx1W8ECsjn4W/va1ewux6qYLCcFJ6HJ8fC+BEmgtIa7bQi4T0b7SzanOc2q4qWV
OVI11rLd2xsKxNO6JnYOKItA3ECXuf6Mm5uxxyYMRwTPISB4SHEhFVMgrBh/Jkl9l453XlM2c4Cr
dtygJU9fN6y1M30GgOzoQFrOW6uUmZjKAlnc22Uqb8xOqatjJWbZKYE2ypPMu/8+Ttdysi3kEUrz
8tzWKjG4Sd86rN6nscw8ljHqx5yZyNDtdJbtWykia/YxVYLh4XJ4L0PecZc+enBOwoITkHow7Cdm
CgmzM8QmUVNf6Rat8IMGdxlaeLn9vSVzg+fpxJLtnt24Fa0Oo0U7XZ74khMf4VwH2JndiEOMNS/3
k5GEF1aQvbSPoMPaAMSpr6l1KGRQqtegXyiZ6XIpUWxypdTervJJD7ITXFNQLjBoraEc5VKqQcDo
+S2fhFdoKIpK3jalM1rJpUAWtbctc06ezFmyBiUaI29/WMe8RJriGCCKWj3E8GRubnlVDuTOs05q
vzULyWClZ7rzrqfeayfLdRyRs6xbz4VxpvMYdDWdXYxAaY5e6xLfSEQwZZYapD+69nU7EkjLdiVU
J/+dsPn1BNMTDbZn/K2LoR6XDCChA0p5oPvqxUmQAVhQq9/1zA3bJczVsqotfzmEmwGxeCTqmse0
OjCMbxEAUH5Ue4f/JlV0y6Sul/s0FtAjpinnoiuPgrUS5AxkQYybN9YjV+Uj+ZryWngIBL/UJQa/
sYSTiSvmhoiSL90uBEIdVBxXg5sCznfFw8DtUjeIVagLDBAOXo3JxJ20zn6zGjGHmPPATQP+hqf0
BW1d+JOiMgJCgc0v7WH3yIQI9gdK/N9gV3RTt2abRZNSeE6I5fru/6kII3etHlRaklhhgLc9Rct/
wdctVKPtL9m9tehSTKVe5zuiwrUQ5Nlf4y23oi6NZLujirHSDUOEUq0Plwkv7R7sEle/V4RIQhpF
4GPzouqJg9wLzWtejsv0Ffyh0evbjU06l7x00q2lbUqfxGDpLgIyzU58kCLZOXUDAxNYsV9YTkQf
yjVZJQHz/8AZoVNLWro/vMbly44dJHrUrbtmTYKha66Puant6E+9iD1ST+sY4N8uThFkL4IvpgLK
PQ4GN9RKLBlfBs6+IZev9FIHERUJ4e4lCBmalB3ofPQXx8i06JGjS129zLQzgYdq9KtvTV1s+mng
eHKjkbtcjk5uL/7HS6cz1SxorH4XxGu9IevM3BJX74S48AKtyHwJmHN2GnB+f22ffVHh1QIV9t2q
YjUtLHCqVkRLTFctWCBmAaPWVqY/jOmAn+Rm7x6f5hrWly0S6rIbHnaWVp8wto9ge2e87Nzis9Jb
VVm/jARigS9J4o+fklIYjQ1BqMV3br4W1FYAc2vyAZINEFCxCvdsc306IBzRX328BGNHvT643hEl
Q+boWT3zUubvJ1b6sLJeqhHKwjPczuOaHdmPl1IrP2zSyMHbBN94T3pnTS+P6YmCE3nMKesbKnUz
fBVJmoPfCdJxTACa45Cf9bUiLFzaa0LKs1g4zG2pnnvWnsUKnhj/BpUwKImkSlZxxSsTob6mtkGH
hLvWlWqnvgszlQiPnBxzD3sf3njG6cmTXgitTjXK/RcFtMbH7u8edWonxv93Js+UVhSXEzP0s3kx
Vy9smwb1Xy1vdeZb4uMTOdivmbby8jG7wtXhsfoNxH82rTVcCIHEvZfv/EgJoXsVFPS0/SewHE2h
4HyKDkXBIgxVPHiXrC54QJjMcMl2/BZp495+h+sm//07TQthDEaNMtL4/bPvvhUQjEf3LaXeQpw8
BIyhnzWUMOXvQ4ZXjHnJAgU5Cv+vVxy1iKHiqHZsD5RpsfDrK9Qf9ty+DPYMBHAtQQHq2d2pqgoS
Ms6QsPFr1GLoxQHbRBpm9Ux7Aq+FcS/zuCTkry0PDLldbfatOGm+eDUFPKKtYj6W7xFlmiq+JYMM
y4HcUE480tx7Xe1towEDiBywpf6kkmph9PGzdGl1jemCAi/SBCMRnJ338MU6CyrTAgmlc4dwQFUv
s8mn5yWtGmZznJQ7HZWjLTpvTlRhEi1g1esjxNH3sqB+YsJdwyhXy2t4KwliRMuNRKPtQERsGy/f
za2/7uqP+dbjV4seAQezbW9EYN8/fjTcI0DzhG4lzlHgyU5s/5DNTskt31BAF+FE4GGTwuClx0sQ
mfbwyGCNm2p7GhC2JjFuHD5k792+EzBMfbN4uiLCuW6Tg2BN8OpuyQx/lGCqxzstgdJdAbMomtqG
xNKpNQJhq1IZT7ZIgcbYVVRLGyHeep+qM0T8Ckz0Qm2Xm13MDRqMq0ZXgNmU5P44rdDAeSzLHMzN
iVBpxCX2qP8DF+m7CeBuw3mduqEnxcXnEyQv12tW20/TGQ9BJTWYltwU3gXGC/IzXkb1fij46v81
amVo1K10jmh9VNmS1La1JuqHrX6j2lzBMhn15Npu+7sNpB4kaDGL03Bj9Oxd6S5o1VcLREnmHNXx
YG17RGB1PhxLLP46UgGTzBLlJN0q2WgXhYSnY7JnWM8PTyVAjCo38IuXt2NZojdJhHJDk3vYUAxA
rIllDELromApNLOCCe/vnLe4wQqDQJtuzvt10m21H7tsyhS+fbfOycVd+erZvqM9zVpNR7x9vH0K
+ZFaWHuIBt6Bl78viPalF+qSpmPM4+CH41bSEAfzRPpaAi8172iiYRR4Cfq47pfX7NtkHVWJ5O3m
fZs7iFSSV7CmFuZJK3Xi6d84x0X70Lpl/VTn67BycvqWTtEjfgZTc56TFt6dkOjsou0yb4fhTXV0
SyOVWPOTGa4pl34i6HFHfmL2/Ta2lN1C38IHXAjYeLfODvRScTLfJb24v6K3rHVo1HonqDlkRgXb
omcqRDUd4OqMiNeMVlkGboMf/6yLdTiPs4DRLXaxv3aB5hEpBtilX/JoZzAloSCQeb+q4XiMlfPw
HZ6Bn55D0QJ+ggacT6t8X9xT5cr7D0jvm3JBB8hwtij4ydroDfBDc+uNwhNN+FaVk8sTjQSCBH18
yCkLjyohNn6EyNroygIy5eYxnayIAd1SrzkgKjuuw3QRbsntbNgzZLEculNEEAQfXfp6Da5wI5Oo
VOGnrFhyO9940bURg6alrVMSGGH0uFKCbrtXpEnLWningPzKq5MFepmf2eWbNBdSHJszT+Vd2ELp
iLqJklZBaX/cb4QLAfw5xt/y1s9+uMk+SNljlxwGpk1zsr2KpumCSE+aqizB/tLL9SYjy8ZGjvnn
PuJPIJAlUDJBDGuCiYgRshzqIxwUAo+gUqL4/SDt66T6K3/jXXBOTH2WcopLI9w4VVi71nwjTWaz
RYgOay+qvupDn4SmjkMDv/Lz6KZ6cK7s6n+ky7X1sAD90hh0uh088MFq/YC2AUKTbphc7zWEfc7F
m/DKvIbwC91glq07FWtUI2vdcAV4AIZ1uUZfUiloOZxjcKjIdyr/M1ovJDSXkD1Ol7mEH9qgEzh7
qcuwJ+X/JrskAhxMOOOYLaaoCLbQVKWv0BOIQxl1QR06MMUiw6FbRdMWanKVG9cdqAzO0f7nrVSh
Q8ro7sj3qFCoQ8c50JIB+YM/N3NS9LBE50PprFNUhynQL6u/7FM+HftBIyLzmOVJXCYg+fA7nJ7y
ZYYECxukKCMECcAC2hoNN25b8t0x9JhChen6LUrFllPEaG0svpIVGXwRDKUcqwcfckHEpB94vdo4
w09yJQjyn8ELYRGR9N0kidgDTxyInswAjNa2123Hflc5Ul1Dct0r8wMFB4TOipIzA+XxzyLoXtRb
d4r3oeSBpLpwp38bRPdJm0DYXWkoaK4uritTlKVKN9AuPDP1OBAIJnaYS0Ot4vSsAspbTT04RHSZ
XEZw/WgcDqiW4dV+3xWVB6/kIDNiXD0njLI/SbRUa4QvLqTwfsXS65bnAS/07LLhPub7KVn+ZR0F
GVkLy36+mYx+eyGJ920Vc7pEznOtGYA5vOqc9ZihdBS/ouT86rb+6xBsQLY1frmTv60mJZWP67LG
OMvxPVdT0hbb/aHS1ZsLId1301nbk4mP08SAfAljG1Y3jB7fj6wivh9xczn7X1JjNw9/qeeIb4Qo
A4E/oR1MQzNmtaMyzQacaYOHShtnR8x3s90PsA56BiuBsec/oxEvLC9q5mOYfCOhxgsKMVqx7RPX
EF80ZmvcXmHwzfjWDbVj5YdGM0FJVdhO84vPf+9gv4TKwXEvuBcVOOljhEnU72V6AwBmpNbBLr+j
g8ntMnlxMKd46loQfCUvZKQa4I3bOYUB+G7WxUxIFsHcSrOCCZdSUcEnDvj0qPEXrfkH0oYbOuZY
yiBlASbnVXn54bnpBrQSPFAlidlIkC6sK4mv0F+cNcIIJdPEyenKoLVAuVIYHkDt+g5B0f9AKq3L
IguYPyA2vX2edfZAbeDjX2BkvC8iXm9XcVTctkmxsGSBB9YiPubvsUh7Iw5OUCz06haqBs+m6/A0
Wd7KFzqn3sEE3WPpcnpQNKwvO9xCoTCjVBLSNXalkeOI22wc978uqL/LlvlhX/GBLXbj3TfoAEVX
6EkG1g0/M8Ny/jV1lO+CubtYhmxHoUW5tsRwTcaSZ+Ym11z9o2sOP/4UhJOpW0xvnchy//mxXfrz
nn2xE1o9v0ulPb9UIYRiQEL+7ZWIRJui+TtvrPVWTZ8Glms3Ia/TnyZ5v+UPhtcEcGUF7wqbMSHf
3KG8eZnOcd+RTUZR7+MON6677TxUhfhgoBQ1OPW5FRbn/Rmebz8+kUs02zjSZDbSwTnLze9cvpJT
pgPRsP/rzUsxCgCz/mLwYFb5pdactJbfkqlXEu/5dPDBZ/1WBjZXjDRhi4YextunVzggsxzF0Wu4
D9hASRVfaM+bbyFO6/xVH/JlDOFvIHTaf5m16gUr4RvPpkENfzsVp/im/P9NAdi5UwQ1ZMaeb+Ii
0LKC5/jQdpErlUrei08NNg49eeW8+5qNFKL3n9WUT3LSgVXGXBY2MeAGdXmu5Ox4l9CoeNq7NE0p
rIN2J6mSc1e4e0/GoQeXccJ21nKGXl1XNIXJniwb9yofpxtfM4QvUK8c1u/WRB8Smn4fOkzqEy/k
EEz/8dOtD33Zoz7vutsisRLhVkZEG7xXJBn+xXJ+zOP9Vo/IXnl44DVRxIhOfkMoBVCWMADplI3T
nYMsDppOLfWU3mkQGERseA32eGums7y+CLMlUTnA8MQzS8xUJdyloKcsY57uQJJ2gJIv3GqBqIdT
5q6/PlYMGtnda63IUjeKyGwdzwuod+eoIZNwpK8+4fnDvmhpmSu+zN5bXHAnrtOa87/fxt35GeiD
J+V3ubIGFD3eBe2so2k0ZHjbZpZfVnqwdM7pjAJfwDYAScKNRtyalp8LV/kZYfAVImAFZP7DPzAw
lNH3kEHFI4V5R9OmNDN3T9St/q1QtVY+Rg9wlvZTJPB4A3QA8r9SfVB6okOolzepyTCcRjvAeeAs
SzfTRRhdppapxolyQe50dUir7RmMw8l6/ImksdoGvLEY4mJBPANQDPIjXBNl/Uoc8vJAPmjYfbcz
gaUt1tpq6I8jTmguuvQvbYfVPAsXaSLWeOyEZr1q7tqMqZ7+MX++Wemxv1ZSunyUhX0nHGf2TfzK
vM9RTK8srda3zjKqHS1nlbjNTzANH3ZAyYKbHSGwzu8B8+HgSdiVG7pMMP2E4KRqmX7Qp4AgL5Dm
Eqx/9pANRIOcmHMyC93NKonuupHepQ8Nx59XPbtCdoAeS/eKxhFavraIhxiJAI6JOmlpFj0Y/FB8
cGlaepwTmqnKkDiUbueiNyMeUXY5dfkqRwBVuyJfihJ9WkMIgy/g0zPQ7ONmLPsCfh+y2gIcgIQX
offKjkJYQxFxOMOfjWam9Edxsr5/BuNU5y8XMeygBbkE6cZPv4yJDuVjDtaSp+Ggc4HnY+OQkESD
Ne8/Wp6Kig3xWcITNtRS2ifttproxM4YcpyLSiUVOeHqg5RoJlBsCc5yvpBQFSdth3LRmhL8DKw1
MqsivKj8/x6adMkVfrRzl+1IJC/c9rWWk79OTW0sZ60A1FiGjxoOvbP29ZZDkRCgDGlxJvG/2esq
RBQAormlkfTTGZYWL7kJFfen9XO1nxjYA83nwI30zt0d3OXyf9LgtP5cUyWxfb4QuTCh7ZMDEwUc
6et+Uhcsa6GPZKojGV3pmytCg5BmnlM3RoCUS+pkkEt18uQREySdOLvvIG30QIfMr+flPLr9MmvC
lYJxIQ5yAgfRCcq38oTZwRGLFex+EuaBvQW+K/dJkB9IPCpKuWE1LFLr9ksT91rxd/HDN/XvFAA9
owOmVSst+e0xW0WiEPWgOkOzzxQ8y8+8dWFlV6wzTkWj6+99c2LpM3LBlzyHSYDy5Ubn81lxTGBa
WCsiKG1RgHLwZfisEZ9L0JbIyPsgwQ19vARuWemfqg9Hm1j2+yflbnXAuf4zRSKZZXb9SQAfYQ9Y
lZ0e61NZDyuoz9Zrfi7zKV9Sp8bGcAafHC4HGOGzEaWQ9ZYoyR8/zsCFprEudvgryWpnTCH1upRW
YgX7mz4W/WYHUW3TM2NP4977wsbAJ2G2NO7dXtCj8cNn6immYq76+fpMPq53DKLkRnt/9CAfOsle
E8vGXejraZy7UWY6yuQ90XWjif1zuhmeb7NPx2nKyROdToga9cLfmTViieNuzSzTqywNM9PN37tc
6lNJaiqbIl01dyKUs5s18ge3PcMtOupy1+QcYI4Rbah41G2onY6h0ixXsUqVIJLo1SnhLJgSpDD2
EwyXZAX2g0MwfGGaDdbAIX/Lcfw/5H+smmKoTVSdiNIR0DV+68MbA1JnIgkU8p7R1p/JYVedNdeE
Yp+Xo0LaEyNP22J8152SSqJteeBPoOp1gIeDiFHoRT7vSqJ+ALU1zPAmFwhJwespSJqwnpkIqgCv
6MFRITD0/vC2p7uhjwZlXkUKNuqZwlFfTh/xXNBDXaew6/9l1vtlz9w3Z6Ubzubp82CSNpoAgcye
dnuzq2Zc/sME7L0jvy7dbX9XUe+HINugiyo4ejI7ZJnBlfVyWy+XgM8Rw/LiP0bok9HrI+NdnXP4
08cKYMoGkgum45AO0xktRF6cWuFKal/YoFx+csBF+sgiy6kyqNAYP4Sio4QspCbubnfVub6RRYW1
m3CG3twdx4Lr+ymqS5AhfGRVGWq+xqZOxpIDTcsTk3axeYkSXJyXmugnQJX21WjYadL1qsjO3khg
b813CyHiqVpuveCfLkLFVlXU3FemmwpVOLBPSA4Didmxp9oY+mGNMHYfRE9xesHZ2TgcEQoeQXnX
ZgXuaZRqi8r8vwYEYs5zIYzN3KEvJK5cSE1N/xdDWwlxnsqMszl6EcnYanuNwTMFz5PUwkbDwzf1
CcHQfoOj8E8xbQy/HJaTTV44Mlr5CK5DwROfycpWmeGSbAGinTd45iPJ2Gyx0GGpT9E8Ijo2vTNN
all2GUThCJ8071mexDiWcPhQFIGtXyFTrzmKkKYn7bFbpqYX4uGTsYoT9l13EOLSHg1ms+J4Y/Wq
325ogQGNSP25Ds96W/0pJtJHJKzw+0u9/mrCOHqA6a3CQA7dLE6HraIS9OUvMLpABO82qwFzrj1Z
ycbFFMEDshyOWHdFbL/Th58jALiZiYH1OEFX1rIULluunkE8uh8h8KzvS6+F/ft7VE5KfhtIF34q
E1c4jMO5tzPA07jSBjFULPsBO/fwF2DZbgD61e5Bggw8PdQ1TYnPj0VuodeMgDs2MmgVt/53xN1M
yj3ogslsG8l7KbZons054PBzZKrjX5KBjviZ0+QKf4NmVUUCve4QVTdPl5i+CU43H9iXcC1MqQ7V
cE3w0i09/j9gGger3ckEOYXnlmg3HWLIdmo3zxEqA4iqBi9FEBW79DcZUk0AaJ6uA6cWQGi/yoL0
3pEOQVaDiKZVH4Pa6uAFyFRB2/OibDDs8ZtAh16IYAQkxXYfqIJ4dMtaXUeBEgMFiGxq8jNWz1um
17Hee9PKEQuEVni5nUHu5MlMST0DXAIJs47ySlnCDrdy4o/DZJiHgA+0cFhWsBLpUTxi6/+U8CEn
OALuQAqXnKCYxk4wSm/snJNsNL9lakPEF8NWnfzLO0JvRjd6BLVRMSGd6DwxY2QOyYO0YhAG4+D9
LaQmYKbySTlLc+3EWPn6JZdhFiiiXcljLpFn2UkpY5Sgjk3gzc6nRGPhux54uEeesApSf1GuTLL7
g2Eqy5a2Mx3vtfPUPWtVs4ok6dhZfJ6XLqNCT+TZD1Pk9cZ64CuoWgMEn6atlcTwdOT4V4oePpQl
ZC7/GOcGm+UWiQaLxw9jJXaudBamd3BsPOsk6qLX2jso8lhI+SrJnIiE8JjSqZhw9LPjKYbjsR7W
53viP1zjvdWAygiTwZcLjnFw62oumawTAmXXFITjSvRH0gITJyupTcqPIbFeK2xNZCX47Q6b4Bxu
KSieYYLH5azd0aRvZ8dagDWw1o4CBEB3RadPdh6yEDZUQUAZqjppJdy1urSVpIvvfnT8z3JrIV9s
wC/GwBrPbtm5kQf/U3Cao13a14OXjMAfr64pKcmT/ohmymNxWn0oHCh3iUrkIfrxEwa6BJG1+XlA
aRi3Ko6J0KghCSmEi3VZ4QXUXC1ZVLfq4xoFFujYhjbub/zmgszfhl4CafQ7aQYjIDjmr8qzv6rZ
mswliSEwASz7LxNHvQ/Ym+0z/bRisarwevuCLxO4fPjao+Aoj8N7ehWJtI32mTeVIpPUV3HGBAOb
mECSWCn2WJZ5/kQcjCJkj/hMS1rzMP5Hrr+F43eF4PC8E2G2s+jWR9WP8MffukjsidmjE93N5zgY
Uz97lvjOd7z+IqiMCVqeMBSf10TBYLm4Ok/dhh5k6lMkjqfDhNrOEdcfoYO1WENBhv4wwylPlNUn
aNkjLtfABhcEJ35WXq2ZsrB/fYQwZHGU1/gMbmPQHLo5bjZTzWni50zoY8W417QOgIfcbMzhGFls
cyTronY2e+hb6QLU+nzdVfhrylHtEofg32cI6cqOdMxT6bixmrU3haPSMYXW3GMpaRoDVVPhbAqK
oM9uyvmnD9F3JElrznhx4QZiOHy2giQyJJ8UN32mshIiUkee9LwG2V0Kr2gl8naZG4jtM7LsLMLq
xjK8e+nRf0b2gdLid5Xw4ekzIJ883YKo3ulmSjuE6AceD2Yznpx8lKnbutJ7Gnyxwq6bUqBKFfBB
HTiPNRy67b5+FcA5WGWq7GHtzzFHV3RjxA34bcQNEKwNpY2vAYoSLPfO0h6GLo4mlatuQoqApZFF
BmUySztR7tUeQowQOV+Y9rfvIKLpkPIIcbcaxqdoDD8ZhDrCp2ETmFlTJOGGTIry/mMjcOyu/r8P
rU4jUNtA4uYWA+ted3DEFEvud+kigdHkX897xb/O3SPQVxpiLcceNJCnRujmXLGZkiF4dPhZoFXH
/F0ZjSndwVaTg/m7BNufEihrDApcz4X21m45fPNiSeFqHTf/35lSf+sfJrwtPev6l4M9xYJeJ2ua
2ABB3R8Q9DktfXSbv+DM4lZ62tRC/9pOMXh5vqd4TrLC/PSBae+L5L1VGAglEweaDuOjYIePBA7R
ar8XHHsvkZH3ZPY6bMrWxe/DWyqVkWohPrDLQJ7mO99nOHPLldyNFHUaO3KlCHaasmn6nDV0SXMK
qt0MLN8v2Xm+ecbegZlZFpR1wE1rKOVFqX2PTpDgUsn2+WTETdLvWgp1dI9fpeZPUtc9F5R3duLn
fEpH2DAUALVLUB2X/SGPUu+TtLF5OVn/6oA3QfjnftBrn0SZ9me3vFc8LNCg4JchsD81T9IzjzaL
CSe8/e/CapCPFt9DMw3rEfRCnkxuQXmsRgT/kjr+NHNc9wIFGc2mgNKFmH44k8k/Re5/akmmPz73
1Jyhv7o3aRa7etadjbWcnXU9dfF5xut54dg2PDCra+ynfA/Z99rd+ywSBTszzJSh5aJAmqdKmuy5
CwgRYuBUna7bRxsd4TFDPWB7Kb03q8xBFqtOwAGyCVDnfyBj7kLk+EJor45Ft0xgtqD5aICDsoJo
7U7aOcE2bfY0kAuBenpXp0wVx4s7/BQw9xu3pqCe3yX37vGZCszoPbAcuL9a8ktAvibQqwjW/5Dg
Qfb4KN93G3C2nv8hN0sUBl3DVkss3S5M1/y+VtIf/XHqVCz2cPEOcG2phrTBr4kOGpaWT/acuPRq
wiN7tuwV5btbktvKyHz/2dXpZOiu2XfiB46knIrU8X6y6m7IC9V7N1QtfZxfxxxb4RZzibzWJomc
Gnv/h5G1F8xQsNvBiAwo1IbAwpHCnEq3Hy7eM6k1vZ/C6ktXUkbagc2KtFjC8dC08x+cpSwhLzCE
XFflgYv1bWQKHzwaY7+ekmvxTrKYTHGmxIs229cpoOjSwR6hvK82W48s/GB6/ebWi9RA3d7XRdkF
85V0i36CmawWPd1DcjH4qNRmo4gV6ImgBvR+CuqxZ1BmW6SN1sSU6zJjBTXhJM9i/hnf2XRcvZuc
dHREbJtPt4+5oQkyKVB7IFPiZtP0XO1qiv6vYNutVd6LZe4rP4/A36qp/6G5sSB5e0B8+MN8Oe19
qoNGH/CBLd3IHvpF0kAovQNWw5WRRNOWigIUFsSQ2nRpOpbbsvCk2MG+pDmrK+ZnsiI0ByhMqTg1
Rw+KYygSImMX//4B4yv6lUWSUjGg+JM6tDUyQJyjMSRJk+NEC9nGxBvbiIOrjkH8b7kIrua6Thdt
Qj11h9qv2V+iYiBAzGOKX7eEaK7uKMVpSiokqHDH+N88L8/e09L74LFKgLuNwIOY24UbenhkFWCp
hDzelRPTmb6TMRM+gR9jjr++Or9hmFGNdJmIyU3sm44lVFyN3nKcaxQV2+L1MDPszaA3bceISsEl
ho18ckxcGZ54C2mGg3AYEPYIC5EQekYy2D8x0Wb3afe9/zMPQPG4IjBj2yxF2JEbZ/xx9/zWodmo
sw6gPVfhM7/nqMUJmE1z1HRC5JatX99umapGC3CBODiWsJrEOcu4TzON1/7ZYNHrrA4bR+ogUp+w
kVDoC/VP5mZ+0HVN+9bIxT3lhMphbli1elGPth7iVq2p+6mLQcopi7MATSqMscZ2o1ZkNRUuutKH
wT3vtFf48SMfDny1rAu6siAnzwItE71IgBKRWpgYd07+oFnF0Tpb4uzKHpvJ+qEqVh6DF+ZgRGLy
FU/ccqNES5nO+8dpd8bmN1i+7dBhfgzXuaHxUtJY+brt983x2O00cID4hAV5cKbdotAQdBktNb4f
dOJssZ+rYXcPSbXlqKQUSHpQDWbI6CeXMtp6rbjLfORZ6bp4ct4CTAMMz7+LY5Cs6ropixwEhC6w
rkpvvmjQkFobepE8iO1eM+YtdIFbwwEXn/EAVykHR5jwS+DPCIaBfJ606nHLZWSvlqXpx3kLalB1
7mA6Y9NLD8KN+RxHQyHYjr9frnKgvA38iEy0XVmIBPkQIhBmAOIDdPAjmKIfiNL9VBalZBGjkqAq
nK84BCMCm+NY+eReoh/8DxFqIAoojfMUu4q4q1EYeyKkEC41wORoRI6DS4bjjunRfd5Pl0H3k2A2
DBqypfOvuhcgJ6N+8MmeyonPaYw0j6GXLGOZoRdSY1Fl6I0DZ2eaPrPvP7Ukl3i1V9HCdxBjsbG+
GVgJyK9tdsUA0roC1flXNuwJzyFJNtghDbOmB3wJwBVXvFfJ6qsZGCVM+QCyprh0nri6nFSYtSgJ
1M71sySd/77ORtSma9dOLr1KTOwqwz+aY3qVfph2cTFadrg4Gtexbch51avsmc0iL00oNPux8ocW
t9DUxMdBohMqys7TLtVkZXwl8gImJ7NJ/LSnbkmDfT/owBt/r1lpasd4ms7D20oYjPRtxk49h+7n
fiSOlLYteY9znyP43ESUtG7Q3vrM6UaGWLjHJp2PY/CYbE+vDGhKf3+EFasJxx6kSthsI2TUa8LT
SqVuYfwvqKe+KiR/lNLgU2XZ6YyBUxzLC9bKDiTdDHDNri4faxxttqZC9UfL/puWAwV2JHhN0vzb
+r+pcAmXYsvlZS3qZEDc4Bhs0N0FfBX0EE1G8QNERrbM7qDOTM4rsIuhZaLmRGNx/wDsFcE4CUeN
7y2qfOckMBz8XVKvCx7wBn2K918cQFd08QMcHUfYeETPm5clnIlBnyzvQhIX97P7UzoRZC6lr+J0
NSzZeXQl0rWqHtczDzHzurF3/n3fxXJm/15nDNmK5jnjjgRscyWL2hmz39VHnY2kZPJ/KAv0ExZ8
k8Bs9Abno0jKDGJxHTyvMz1n0IsG7XLgma/r+L76JEzIScRRnVaPexWRClK3wMIAkf7YLpesUaIh
hXFLT9lkIodZTzoqUWfiJTLXDttLjBgAwB/Tq56wmwsnumPSVR6xTKF4td/9UVLMf+O0pBxRUHkM
yl7I82Zd8FdMnbWc9EVtSSVwCV0fvN+l+J9NKXgX0UrMQQ0DgjOxgckkXjpJYYdMGX87HxmLG2fR
u0pPEZIJCvKzx12R/+0HdsZSbTJ/YTCll/n/9WP4DWnXM6BQSvEmSNJmeN7FfQQScBLc50fH8WqJ
ntcrdPk7heHVbhIG4dfhOyFaqH5HApjooAPOMSIwhwWxM/JMDA5GJXeGRdnCUCSNDRn4ULLr1T6b
Cd2kDs8iOmupOYFZIsKjra2igZCUZlWfz2eE1M/FNSPG5DOav6YF5JpZgaHzewbpLtflklbqVFwa
nL8lOzkh/MYHjPFJnIEFbZ6EQv71Th6YYqmxqwjszzKRyXb6LOu5HBdt30r/USDYxJxbZj0BTd/j
kfpEUmoD8FfORzBZbG1EuKM/3ltbPp1Wr1JwKPXZMestrylLHCfqMSDzY7ykKlisyEVML9gHdFmO
0c0HbBS+FZ4BMX2ficsx4Kbl7EDfmSNYLbpw3YE2mR5Ga0iTiwJFCjUw3t/fvJ2uN5789suNMDis
epzQl7aUVGvxFVMdXYTEg9ZC9CcshZtCJ2hmxsLqeiHJMNPorAF8mGagdTyFDO2+eA4TL8PVYwab
6L2rEu5B8b1FI65MdRH+OIt0zmOsLtSHX78DFE3bwlJouCM2he382ZrlG+yV6ZGSqz1gj4SzDuLX
0lHxEdqiRfTfHvT4/L45sOprd5wL0Yl+GN4426lwUlSoktAB4APFiJwSRUbgNUFGWe5dvEy4WpLk
HV3FA7s8LN5cZbx/svO5U3iEOOXB4TtGtbT9UL+QkwuoqiQYrkKmDo10D9ricyjzbKiEa9j698/x
BCVzxq0OqpEPgBY0OGpaaNp+O5J+I5c2+PLUl/KzFYuTZTmAf17guuRinpTK13ni2ESx21R5fpKs
+nlsorRtCog3dr451H/fACUR7Rk2xm/wHvbaOz4uK72gCaxWezO3UCpl6JAG6ycLsBX/UaHMqPAw
AW0LPt/5o6zOIxj358UL6j6btkqycUpcAoiGYGFXTT8kxjyWjBuBBeirMxOUypqJl8KIO8TEZoSY
ozaNc5u2gHjNGTwGy425b/79d5LiPb3tLixE34AyuR8dfBCLzwfFjdaoajtWwHDukPDAuLUxWwvc
CoktXJuRdklDdcVZEjn9f6gP8hIJgXpU6Jv89A7xQvY/3ndG/ofo15wOCf1GaAVlZZzYeOJExpr+
Ksm4s3zkJyygG1hthMB3a1gjUAjUwKcIW3xtZ8mvAyZKzcMebnmvu34te/o2k9Jz58wbKIAaatH+
QsB/PYV/DkF6gg92d3/LIcfxOsAlMYWErNuX/PbMNYA51JD9YEZvadHih6DEBuR088LQH4nkKH89
C1QKBuZWnj6jc/ueQsv5RAmtDKAq+SVa9mv2x+KDV1LU+xPSn4nlrRCTIt1X+31NTnfZoKoIS2c0
8irrSgoeawfEQ7wMSmYYZvknnRuz7UIhN90/PK5wnwGiZcdhpBxoa5mwvLyBVGnB8Sr+2p3ZGsII
f1a8nYxrFrckMkVMsGK6zQPN4abA/gz/SwsIjxKH33FhhODJXBLt3MLCTgUpG8piyPz91NM6TS7O
Fj+Qem5r4+nNucbeu880rnimQpbzE+DQ8k3So+DW66MFp90bNd3n5+2Psc2CxwZM1eFIKlwr+FBn
oUISmaoHj96hsSzwejqxdyInJlL+NJoz8ZyOizpdNXGYZi4dsiNxw3I/F8hgMEYe6+wvcTVE7Xz7
oCnWptq0dacDkrb4qM5Or5rq8Xne8n8SYRgrkYg3MMSaF35FXtsiLP5H8E+P4w2I1zM7pf5jfo8T
YtWfZMIM7THjmAEey3DLjJvgGlJS0MQ9eTqBTco2Ey5qfaqSsCt4L6B/Xa5fK9GrDSW+8b1kOb6n
MBpRCjz4YKYqWaYs+lG0vVVAwlLC84jBOLOBUAxEasR+DH+o8uuhZeiEnhLuG8d26zSnKzG5/cDx
uw4Gn8uJL358wofZBQXxxTvd7f5A2izrdRH3H/KSuoeJMgtb/FqFN/+ePWWLj4xoaDk2QaB7esSg
FsCoXvAcCPRmoHbz0AmxgP7R9POCh1rel2bhw3tQErWjySxaK/ZxOCPuyS4jMxEGvl+vB1Ef91fv
yP4fPuHeWy/xKhMrvEWmA9zNEtI5eaOFXgG3tnb48TNUiDo91G+lppSX+i15JV4IUo+QGLkhAa/i
Ap7U7J1smKrFStyg3pqG6H0ewwp/y5FuO0zHuhaIt81QNPl9nTul7qT5MPQkIHzcUH+vMIUMIljH
8s5jGZ1LjqbcUne5S1IPWQK43C8Lygt0SuTRnevrzHreVPXndHkuqVU0fap0g7Y6UOM0ovJRAW8l
g6j0t6XmV0qE4RfrSRB93k+2GHhuKpxepSDPDz2b2F+DmZS9qnZ2+Azl6Lkzd4vhgCSS8gIMMefF
KsHfItiA1Y7C9FxO1Kcb50/bsC+bSlCyUoYXIQ2iR4ngxyAmdINOBX1q0kcH9zAj/f/l5g6AybBu
Od6n/oB2ZSFqVl8GjvwRaOWv1alrs+0b6Bwmqx4KX7UT8xg1atWT905LOG7YdYJ6BdCzJfj3M2Xl
DMNXbncDwDHW6WXcUdcHGsje7Bz4IRRQArmd2M9QUoWr6rEFEhPsg7ZtPoVATdLgRk3OmUCoY+6e
bSgKGyXYuOw0/r1LTNKYXKIIJFYQMSE3z7FT4grDJID+ICTk7QbI3wftskRGn9qUq55z/M4FLZdo
nbAefnIe159LHFmlUw9jZm4pz25/ZUXTnc1Px900hA53wBuP7E8BY5/uaedwlqvzN0nc0jyq+XWC
Xku0T/rCigGQa4GYPXLZrN41qpcFm0AvumxDLushERrTHfcKrlRmqoNbvAA3tsQjxPoWquPZ5LrT
B6+vN9Hmsw6Rl8ieSQjd4q5wxXMprJKedIiKxbGneHgnVfzKT95AZ/UY7e3da9Oes++MJXJulZdh
BGJZZq2OMZE7D6mNnN2qNi3KvwwSQGNOl79FhI2t/N+0dCKtphgcM8yAI9m042QBmIhYVA0Yd0EZ
R4c2A+hNSqQ/LDPEWmWDmt3nJGgIO119v5HC0mnOkLxdFCYOqN72GBQV6LvzYZ9boyjNBtq9/c4e
RXDyXstp2hfN9mLudzk0xw5T2AyR3XCDc55fpaQSP2jOsetcSkeLWRlMTd2egh5njTho9DKMXMDn
l5LTPFOsAwt102pkvMo767BgBGIglbK7Lq3Rgj9cdnyLrSmXldQe32aWMDth+qJRa37WKP51lUQe
FlQbgIpt+0a104bhn7hpXQ2gHXWYN7I12+CSx/zXvo9bZvWndyWCFl7COFKKl72IywxzU58cFznW
Dh1Z+ch7Ho/i1mrh+WjVL45wLXvXPj3O1NUWBOitHnzJRDMwDlFtKqZKXRW+dBy3fapw8382b7QE
xFPigbRObBPVIlHeXxXqw9362UiupKhnwtN3PMdj4O2TJa1D7z87hShVxqK/i5GGb3RaePCUlqfY
3tCmniEjCr/DO9C+W6DBcgi6tDn4wtqyxbtXnBmuul/lDUf+VdtM/JILUMdwPSTeMZ51JbFDYee+
a777+YztOBc/wzmqOkKngvdAHuPhyJaZN1H+OpOwCQEIZdAeONF5fnHUrCIR3UJ4fA2zU9BDOiRe
74MX3HqsxfKtTlzmpGrkSab4FXJm1WZZ2oYQ1JXeIcYn5rZWp4pR7sadpTeVybxbfYiqDCu28QZE
vOktT4mbbq6CylJWl7ir8FbqGmLH40flikhLZ/ZrZBebVT0Zwzie2EYISJzGffso1wMvGVwJPrmL
72AxS+2nZq35auYxTe5HwNki9bQ19ojeoLdm7prfW0cjKsygocfKLF5eIlt9bwncwRj5QvqCi4n7
ZmRhEHyJ3n+UqJH4CVU5n68O31y1Zv70xv7udXTGES3M3EFYsiF3DWusO1HjfK9ApHmCDC1GnG7n
kvreRCRpw6paFVWC8vRwFEbzKmRpseZPFIvYSw3YR27SyImISgUf032i2zwy1/kquykhKNQ1Ql0z
eZ35+5gJv1bVwEJRo/H2jU0zHTkP5WA5V/3Pfi1i6O5prRfEeCYhydkiqDhUK+BQy62t+FOqc29d
deGRyWrGKOUuILXWI6xoL2DABipXMkdAboOVFU3c7yJcvE2lSyLe8iRnBNTwKc3G4uMITdRdwVad
HaBnPwA0RtT/ELYRim/or8/r2Bny44ir2PfVBHKYQRqn8khIGXKweT/tG+TTm00LVpdRc9I6DkkA
8MTJjkcvC/REu5k/o3hJvg55Cqmvgz8kZOmdaHCpJPqjidVBSXm0sJV3S7rLL3kuKwiyoTTCTOi+
ZtA4PQ2TaUNCocc469raGGVJSkx6zVWV/mXWVjxoQPOOLXyIzy8ACbDPMAWbt8K0BYmgEQeBnNg/
MU76fDJ5BNk3PTCEIpcI2GOvUjTpTfB45gZeXPVFT/Putusyh7SmtPk5sYcKuN1u9A52hd64gFI+
LX+p6laKRLAGhlntaHAY0D/J+lRqMUGOIjEjU9RJ5QkYqcHB274DT3jUjWb2Bs4bi1Ui2ziQsHjM
3eQdcF6+Zz4Hrj0nkHMfcF7N/mc3te4rkLcZmdRYK8BVFaix9noEFBgKHP9DZCBqdDY6dT6lyJoY
rG0UlVeu3wvLg/dpL7w1juovFp9CyOaMUXC4Lis5n/tgA2hYzskQXXMUmyhy7o+BM957iQgJbl0G
dnbrMjl9wFNCAw/OYMe1rS1obpBJA+s9WWWjwF3+4aO4a83wrOkB28I46m/FpAxRrTRsAGMAqEva
b8KV4/CI0+yDO73FhQ8IHjXeqZI8fbIylJkItlNqV5eBuyFw3NhDUt2HzbzNTti9mFInQoqQMsmI
FbUWUSRC5pqzbqPkjzWhFy0PvMA7fEImfGbdh9Pjn5iJJOy6aRydDSjGfqvrAcS9Q+WcM6KZKzpU
7KD4HQtFwFthpbQcvfbB3LhdIdzMDa0CY5sfMf6b4Qp4HUc9UYzLLUXO0vIvx0LDYf2UXMxus8vm
k3s2BCcphrVCfJWSWSfMFUqSE2Ji0oytLRV61CTR45fa4eZdTURYx4rBakmaNCv+LuphlJRZKF0/
YiALs9/ffDmUmukP86Ts99KadmQwJCbfNOmy2V4c5SlMb1JxaXnlGTVAMNeBGdrWzVlLFmXV4zhn
uR1tNCgSBL+QjSX0N408HUBa+EcdTbHfPafwfZjOM9EqkZSAg0ONSoEuhjSbc+wn5YXygJ/RKlC/
cpQHICUqcZeB162pXqE6f6c43R3Ij0B3UkGNEgEekmbDek0ZOkTJj6JtK8wQzZpmMh5hHzRpj2EH
d/wsqxNTQmg74n92ppBr+X0RDGdj4TihwdnAlLuBrCreKbePtkU7O9iJ9QB6tDVrhudh3xoBxWKC
DM2vlqxvDbNC9EGkG2YaG9SvShIVahQp0nkHHRMQMXGjOzYiXYYdX8/+L8tLRFgw8T9F72iWNTIK
/UdUXESLpoocTPLz2OtsWN3zEtjFzP511fCCZRAH0zlB8enjsKV6VDcPc6H6s2IuIaNDkV/79Pjr
lSecQkan5Pdh4qjnvdOtlOMIAmZP0q+8pGqkpb3+0XzR8YKRGwndDyCnhKZaxY41KZ8Rj7P8CAsr
uPN9XmqzcJhMq7qBak5zRnNxR9Irn5XYWzEIm/VxU7JVsMtB71kr0/5HGG49rMl3LWf7tZH6aQOg
QL9w7W4XLgMnGCxLaC+72U8iCy10i56xTpJTSciBWYfw7LCPS8CaE38oL/5O7zbgsbLemEVJN0TX
SN3sSf3ov3/gC6n96eaUkAofzptXB2e+Ziwx0p22E60Ex4drgjhyUNLyWaZA7Dn8YYba1xRFCCez
OhpYJJO2OD5Ixn4BjBWttsvxKLn0K5NIRVZyqKYSMrgwMCJCiJ+t5aoWuH3PT14MAYvMzOt0v9Hs
nz4+mvUynfnLwHmW4u0JLwjgK1EycZhF3QvWMltjy2v/aTY5f9SkcXTQfAlwHLenZ+qEha6MCDAC
jxKL9Knyk58VpdhF+GtCepeZgCbYcI438vtDgOf0BNK+Emt27/A6ffzJh81uUMQj46592CYMRkrX
P3JFIVh8EGJV4O49BEIseaIPkQSXstSwFksamuX7QvUnPDW8KOlnx+PFYCIyUdvbD7lgGXPZGO0q
EiN+vqQyA9vAqFWbai16mYv2Kj3xIQkCLeLvBDNdLRLpCSldPok2WPPwKdyQ/5cL16bhlheYl4lK
WMvfLgLF/0c3SJ3vFizY8HvJ/gJeTRsVOLpbrvODZCjAVyAfI8SF5KYL32ynOGcOB4JLce3r9xye
fXc+WxuBNNnhG7rqAHGvmyApveRnQJh4xIswyiVlkcYlf7Jy6Map7cSTJnOGRO5mlBYZ6wx2WPq/
Xpbr1f1cNmbbOFUhRZkL7upCsq9TqsfYYiTCeRvRwa2RJXI4jHvm/cPv9T5Rfv9zrW8pl1Yrcn8m
klFmDncr7omuss9gL5KOTBV4LYdyJcXIqkBAJcG83+P52NqNXcu80dHfkGZENyLbGAdeuT5UDbkQ
BdQPCVRk7NIbdfoyRhK4BxohAmCnQIJKLgEPdO7ZElZrs/9PnoJSvYViTCXExy/gsgj2gYGHFQ+0
20dpYZMvfGXu3UV8MA3BppVTBTbxE/C/saZGirovhoBbdYKRNuRdz37nIEGS5uM8fqQMmcRR/0AU
HfCiNrnhT6aIfxX+filUxE8cJb2Jd3IFQvDzkGw5epudugswTq+7oC+gkEavPwq5FgFygpQObMuV
Bq7RY/+xjQCUj0+g5sdMRfT5iPQ/H+jPbZ0ZKI092PhEYNVPmPt8AdPOl8ms7ELYirk1OV6TUVL+
C9aoQxH3SS8qTqpbQkLOeYFHg8EhYob81Tn/QR8AakA9ItzbPfy0Tm4d4qDqDbxuXzwiAkQt1dzq
fWDFPAslNUKkYAEJsKAPdFB0g0dvsZeqYZ1dyoRmj5U1qWavh1pejJ7NMU5P17eYqCiQrCGlyWo4
MLgO1uYbbvgDkxjhH3+7peSfWxtFRdzNhodGCZhJpqR2djSJ3k+oq0qTM1RDBkmCbYYd59uJQ6ge
EUVXJnJDb2WyawA7ssnLwtxe+EG2f1m2h3qG29P/StLmuy4Jl4JytWX3cvGasSJojwJouL/khjhe
sojAfQKCW991tdQGV9SsZEItX3UCYVwk4Z7SiI5cHvwqtjN3/mkMvws2e+C8YZkPrA6CgcwqFPdn
8MSWnA0VSND32vuAFsGXZ+eXaEhGAWQcZo1WcTaydnbJ2tzP4iRQw+0E+9fbSXsoZb3RP7RjsJA5
4a5Ph6q+mNH93dJnNGsIqKnjb0SySHV9YUcVeWzzjE7Q5MsVLPMcIQP/7AgbZiaLgQYXlcWvMFIi
zY77dHFjCmNpli6PRvAV9/WCyI5Hd3zWqnvguRYfSyfR1Rc3KyuisKMXcQ9LHkMCNOYm5nPAz6jV
ztaDuRWycoXdQya/T3f3pc1Rr8gAmtAiefRjPI+MphQaWLdkIdwCoeLAIeSwFp1Arhz5TIkIcjM2
z6QAYXY55JmDrR2UpZFX4mUZFLXWPbBGbIanSjib6+i7/XpQ4IgAFtZGcsSKAr5aaW/dDl3U4j8w
eUk47bdGUux+M/A=
`protect end_protected
