`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kFc5K9LvdTZe57Ta4b4w54YJ9K6E6KuiE/MB1wjL4HD6ZTzmLs1XkjmPl4LtE62Yur04bELPJlTl
JgZBPy8Keg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ifyFb0NhfgHUpJjr0mbMaFOI/NskmbnU8xR3QjvYKT9xkH3UHw1vQd9BG7/dIGUHCVmtJfIXw4gS
SUqybR+7d8FU4ja9CI90DuhGphA0AOzFxDP6/prYMyeU3eoT3CfOa5ayndqM3WofQymiXhrLHY4Q
JGk/1YYX0T/IP5SAoj4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fnxoeeqy0lIt0CRjOCSmrSjpyy5+Xt2L8J8WOsSetKdIJZIpMw93R0X47CGZEzoOfrJ/ukJ+Atf6
TLLIN+LwkbiWAJVeFY98K7tAXu0tJafNd6dwSe5zrxRnxhmaFMh8dDTOyLQ9XP+KJ5I+VcjxVFg9
xS2oldU+p02+nlor9a0xBBMtG+TfAdehZQqTF7Q/A80YVyrNpe7ZnVqJNcAdX7ZRb0WEdjyjD2Gy
wJd3uQLw3vxCy+ZTcQchKfzqk0MCrY4DMpa3svZfqhfKolUae9fnLCbWHe5YL27PZbo0aU4EebOr
Zbw+AE5R2+g/FHrgJg+bNSp1mrd3OXT6zw7wDg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EZ2vkptAJUNsb1TA7J6o5Fz+WBMu3/ERvKEQ/MvoY/XTiLTvU/9yqkm0ScjwVBb+pZsOtuDz9sH/
Md+fTWZdbolo+y8tQURBldL5ShSjSBtUmPU0gq3ZTZMuArWe+awSYMPa2pbXhF3V5tHKcKVQ0w7R
iRewWPKd8p0N0fmRI1U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f/dJA8YRX7sloRncNtKg0GyZtwkTWHqn2JPiiIpKxSpvGD4hSRO+wN3Yo0F65ZRLDYigYuzN2569
lkO68mbcLDbXprbTcJMdI4MG2FLe2f8BoRWax24BqXVxMDwE33zceFEz8hMHVSoUUuKvuL0bez89
d71tWCAada52i1FAIsCGh4VC+lZUwl92NMvM3Lj8TZEwAmgYMrlT08UswGW65ZI+u/ZzirjYTwLO
fWr0grBdpVSlClH/ggeYB7P2jtAjGtGNSvUQ0WB89C8SewKnQSw47tKSuZghALJVvd8Vqs3qJVDK
d0ZNjlufAjPKzq5P2Md0Ht1FwMy7rFXT/0ZkKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13424)
`protect data_block
aD/UZYRYhPoI6KPwKITcWqbwWIyy8i48Ge15PI/tYjHPMUKu7dPfk2/aUPxrqjN8XOyFckTH6GCA
tBh7/scN6z24ZiWHT5HaCuMySJIZ8OOndMjdCBFXKU1QH2XdJAkhnEk6wLYqyrqM6m1Aiuy2vDf/
XfO0dKTe6CUpiD6xctxVrCSbZy4SIzIgwVBvRHvPxDAguPArWCYMq1h45dTgb1w5VrvvXSEA5pa3
0ZshIVUFXhTkbsU2piJO8T7/ocV5o5bQbH36TLKm5e7sXm4/wQHu2jUF4Axb58wINMfXSqbR3PFc
m7On3mubTSc3WkwI9m0dzmPGeUue2pTeonO8Hp7OQsOjDohdOc86y9vNyoZT8jko4w6gyrtGXO8i
I0PlCCJdwQlHzGnaeGt7LlVIsjKLb2fXkiDzGnkFC6AeUaQXzzaigHFSWqjkt/2PkY5cqmAKBeIt
jtWfGC606N+a/fL8vQmxvnm5t9Bcv+MiVVmb49fxXysLazWQu9R7QrW5BIEJoE69FAf79NpwMnWg
361u1kOAZs+AO8MMmXfapiA5iarsk4bG15qoeTGmCPmhXCzkZbpPOkh1bgnG5O5f96YTdQ/2wLZv
CxHmN1d8qa9c9oI3beso5pTdYF0BF8jylRqhYdasw1hOZ6ZnA6ofQQ+UWGzdNK9IdewfjGIilmKB
O+yBvyvgYWR2R7vTZeOe/Gr0Js+Mx3CuHO4VmvbEfBCfPfLlvb+cmKsGD79rebv5ItJElz3zKWic
yE9aYCrUEDWW6fcTl1TxRBmg9ye3nE/YONDuwl5SpOTZ+PlCc4j03zWU7hiH0lSdAZ6AXsHOnYSL
OCGkRKAOuyqAynh24v8d8F+fF45cX99JqeJ0zMnG9eDCYLT9DAmnQJMhd3rklsAks/tuJYfwK2zj
3QjNWRceTEV3mSMwmP8mrnbi4UtqpwD4cmTFSKLjjfzNv9RrF3gFEZQZiL/hOh/7m4wgE23Xr7i1
GVVcROg4FWe4x0/q72Bkmouj33+u5+npCWSNuDbIvzxCeHeGDvmKC//FhJaygWckdJiAHIoLvKHN
L4KswlT9XuXtXPKQ+2WToJdwEfelXjFRPLO1Z+ORXk7VjKdSjWhVdkgDEZLDPPs5bFrYOha0zrrC
PZdK9GLrY1oUvdBXOtOXGXF/8QgJ/LFiA2RYTsuJlyBlmEtRBUBfiDxmST3Pfvf2D7ywJpCfTf1F
1cbM+yoipPP+YLzX2x92cFY4ZvrL6WsYpZ0yMSP/W8Pj1xc+YS9kMqqnZemjOfc3qs/GgAIjlqkl
j031dCRzvHWE/xHw5H5KCOkkPuXTo53HEQIV+cf7yc4D7eQzzNgTyGKa1FfJOxJVovZgADyKPLcy
Zm02lPVHZ6pCvIZmzdINlf1PaX5zgsFBFBAoNt1VSkwCaK9A1ri4BBVJlfeMvtn8aAlxpaWIRLHW
0DdCCYSeSiTuCsZIoIfPSdnc2zFovMVyDpnBKMsY1m678AM0XN0M/hykGwwjJRtpUJw9ir2/yFoy
NiBA0+XZ+6wKK0mnu2MTYVpmq4OQRp11QSs/GkH8+kht0Uq8IxJeucNjDrQUtHPLt84nUuK9gh2B
mbt+Wi6/QaKStZHqJdX4H6Xys/zXvibQylOI8tzem9RekVYemBuVHbuom3hIswwSUiZXD1H/6ssW
Jfq/JGgVtMWL/GvIV3Ttpdfc/WCPgoSQUGgZOnYW72nSWzNJS5SJ4V6AXbdYbap/0RkLJ7cIMbY5
CVqkH3iKa1d9DsjaW1jnOd0YwsTzU4Y+ESCBes1xvrWUJq+Cx3BbD/p8Uls2XJ2IBlh0E6DwrUFj
Ovva3tTwhz3KWTVj1DQjk86N7EqnWEvqIeowJK6sWCylt+aDeF7Og1U/L/pJGTy/NpdNB/rbWhP7
bP1LXPIKXFOSrudEbr4ZP4LtJiYV7CDHRs2WOiZt4JI8T/v40XuU50oHp0OWGQXlZRJYE+7LybaD
u//KatgwYJFJkyNabLzz9h6C/B5OC9xBJHDhXJUabdTrjFUH5n+Bkl1yZCsjrElx/tczefB5n5NS
Sq6YLO1uIUO3uKvS0r63A9gvfIPe8HQF+mXOFgrTREBuzw61P2YFizh+1JF4N9HozppWt3O15dTX
bO3/yBzeB4uNgsPT8swqOjXX5JAclE8fZSl4dOnwK8p48vEFm4PCtPc3Rxo/SIyrKJMexqre1GvC
aH1tOdPkkvagZY8gN/p2YSAhvKCL6qeBR4w8nog1al1c3x1iH3VgCTxcw4eqvWzqKREh76gYqady
O+p0+s1zuisrP6o9WFxVIU/dopiyWg/OZjiCah6kdNdowH5xtA3NNmcYGxewBJa+Rt5SGtKKooYP
5mudvnEola4qRhtD77f9FPTJ4hjHGhikfZa63Q3vFkmSNZDqgVbTT1UtddBn+S1QvpMKoGxrtxnu
/L9Vp6Sr11zeIFKos6jYSEMlxCLqv+ImCoQILLp0vbN50DxQuZyPFPg9wPQxQXb2OhxKqmsOYS6+
jTsLNv5hMJmTvM9DwzDFoPLlkPCFgyS6gFSbi6hUyF51AsRxjPVeLnpX8RI55ZP5TohEu8zLodUj
J84zXxJQH2VW+6FY90J0fRBt8CV1pXcGxyoL80+gB9sM/LFMpRzy6i/YzZDq5JIf6lFyzakaPTMx
gwAJA/cpuVMAYQqId0vRY7MmgaJENalWJEjn58cConIVmmRcZR51ned5BMdNsPqg0EHu3zKE7Pem
QUTuOn2fxg6O7s3+irn/w0yu5jdqIJ5V7oy828cDNRFTApq+OE/QT5PJyF9/sF/YalCJ+7SLY9H5
MdlH0VfjaYJTvyQK6cD6qpyqALOtXqMh/XzhIImwGzSGtgm64gp6CHYMtMt95JpItvEULLHItSEC
ppuLbvY+sq78uncwS5aB9dbl8/SFROu+9EMTcSY9w53G/5z98QtrCJ5reMaOLLfvUidSHeZQ7rz1
oRlhv0PiFFelbFr/C+UU4zBt53K5He0Q3VyZwg9GNI1WFzJRwiyetnsmDYjsrbOWCyK2BV/K8I7Y
NrWvqqUww6iXtAKbsKeuUSUBJiMAs02b5ORaCyhWv2a3X2rRqV/JBeO4IslZdXWPVaDRiY7FBJ1I
M39Nc9s0P8z6n9SRorl0qkZ2DPG8p73Il5jEYp5m/t2VeQ/y31qRHbSdDObRCTLwPSGXRqEgtVMa
+VV2y66iAdY3YqoS4vkemrECJUNjQuMkoWrNOZci2dLfkop5hirw7M2ZOBLppsdYLVOAkqY+qJ9K
qt63to2E08toSsznpRnitSyCFWAByQzgR/0LerUm2pQqYMtNgD0hO/ekyc+tAC/chrYJd3Vw8HyZ
vCy6U9TIlWJkOKXJ1qEfvBAkZINrhjBpSnDHCPO3MBdrfvbOhorxqhcCajt478AjA4Hh6BOTPNiU
+FXvO9/GbGq26St+0JwjIU2R8GKh5gTNbi8qJGC777PM5agWA+SaeAU4qeGI2Ace7bfhzVlIgyXZ
ZyC+CkigYgWS6/cGKkhswWCKRUVsP1uMcqZ//qk/lQGJBsM7ialNQAvvpZYnOasMJgHGm16SauIa
vEdmxKCz9fRQ0N2x+yFywIuNTtBcXnZdjKfrQ9A9qOVr6wc0nkR4PdL7QPar2jSKHS37chxUPbxr
Gp8raiNXag0d5DUgFNJ673dWB9q2aKth/wdSlRfqqU0156WAlI5kIUQdPrkDwCGfdPKFAgSGveAR
Rur6Sr1mWD+B7yhixMNVS+eIqX7bcvEjbNaxoStF3qktYlRSMFHiNDBh05DZvOR8ezPI474mL7Dw
99px7AmY7h9rQCj/Jisjp46CTKwxBkrG2xDBHTsuz0Tw3E43TPTtxddwgr4EOo+Yk3k9A1Djx8rm
7uw8ufxSPDAwFIXSjaYgpEjSWY3guzGcXziwlX6/wJxcW7DzRbYXMeWOsRWcuGPBB4Ll6HiwP8Le
W3dDDKsGQMLsgQriODSJXFfY+DixgV3/Jlan5MhnEVhtNxpq10hp9iKWLboqwZofNatQbQuXN8GY
5roxuP/Sx8+6UfQXpv84r332jhe7BULnPnu1lvB8P7CHI1hJ5CkxDCSGJfofDCFaAZPVSXuduea/
J536q3BgbjcELepy2wMP+K4NjT8gbxOrRMB3W3VsOBDycFCUuE4JXHGGu00eL/REjiBlpPJmshko
v2EerW67kqRh1A3ChcjAAnNDCG3SySVRybj4GRimg5rdeqciaXBhrhSaE0nI/Ac7vZvrwxWzEM28
mitq26y/TVI1h8FjiXOFWkCAB7Dmxwg9tQT4RSRa2F5/3KD93W/sijCUNQMaTAsImcObLtmomwsf
hUS01UHGYpXhZKKc2iIMn/Uy48RHt3AWygQ2aRAYKze4wDwAqfcmlMVmAV5mYmB5hlvszceoTFgB
Swouhluxi3jXbB62vxxJoGt3VivlOgOfJhpKNO8eozhRzqpAwDB5IcpTMrxF21CnqCDMIkogPTL1
kogJ13iYCq4Yfqxge+PE1lImomRxgMjKAl+2Qex1l+7Scjs3E9OL7VXWXeI9NAVFFTdsxltVmeqD
7xbPAibzdMWhQUS/l4LS+GCExQAwwqUthpnlyFOzF2Wam9Mp7kX0yjFqSYtxNTa7+HiIMCqgQTeg
3mvt+f8cuFnfOfoaOWYqOF0V4Fgq/M2HcP21kC6lGfnfHNWHlO8MfbD5hLjd06rf5mhp65n09qbp
VmqT/spMZ+Y/lKB5wv64sGMWonIyqGcHuKbKofP5mLpH0aemrZ3DyIm3uT/aJ/8G6rzwaNzQg6Jf
itCKVHOs3N44sYoZSf4kk+EW9n8p/oYCBkZkBQVeL0XiSWVCkfO3Otb9ABg3aiTszxQOmK69V1nj
w85I4CuXPX542HN2Lpo1xamVA+cFDHacJ1dju02eoBecIbvzazDi2gaInyCqe0Gxe9kqfjvv45ml
VYxfT/HU1+KUHcafm4VeaWZjNguQpfs3qTJMMfsNlM4Brj79+mWEY3QHxunZiXRvmMMHiq1Vn7FS
i4cCGOSx7stlAdaG2M0QUvj1wLIyGSEQuyvy9nD77fuZpi94K1onKm7f/H7DCyh0o9pQIwBFHlQa
BMdyrYTnj2LVcJBwKqMSrLMv6xuwHjr2yqvj+oOVVGIsvGQhszw9sCChPfzr/6mLXZmH1qWgggsZ
KSwOxVVjjDvAT7nPpUhSHV5wttkNZPGU8uElEkHVgKwtYyEK7fUGuLGLnMPJStlTvKlrAd4faNsL
1DTrHXxQYPCFiIVjOw43LF5cYJXKwNbISfQA3RO7tNUv8GqhKCLUvUj8bLqUDzlnn/xIwqqZTlWr
fkpIZYMz4YPUBBJCrXQnUt74RMa9GTe/86DNLvCpwMRrlfC0cBm0uXg0IZG4ITRBBqrz3QQ1R2Pw
79dvM16p67fAFqt4tbf0NuhJ3MGAL8SVAwNu5gCKxiD5Yljegn+frinah/OiwhQ84IhXOSxSYC66
PbhG24VzE2nMaPiG0GH0+TJ8DHXImyObmwjncaa7vqx7Blvn9yJU+SOUlIrsCSLd4Yyube3sqM5M
Zy5V/W7lTk51czIusMv+ychx9a+IvPYT4ejlhwucbrZTI6/INDdm17ecak1Jqb/+LX1GtymtKUsd
23K5KMTNbx4FQvvTesiH/2RLgNXL+C4qOScFpBjXIg8ODRi3aUwjoQUPJmJe6NvlgIvhRWTFJ5Fm
wgUjwrQl7HHFdut4TuTxAYoanPR3Kx9zJK7x9wQeu/saVFQ1P83ILCbUeeTYz9m4f4YK+7KaBQAw
hmtjxOphcgoR4vAaDcU7aAIIT5ZOmEwWOTaaAkPGWGb6EW8Q4xwDyYDCj2PyL856fHfyhqHUjS6t
PTuVjGJr7PfGbrfQHDxkHkvMsd9Kdhy/TCUjWATLO9Lm9kbLULdZTk0KpyIxqHFH1MZ/HUxppnX5
pOAMgNu3FOO3sioCBzxOb0SnY69oG3rF1bShuYSQlsPFKaFlPhACuXLaKKzoEw5OtAB6C5KXTQuf
AudgpAhcUidrQrSB2nOfUcGvDsyc2LzcgrMAr9r8u+6IYfyqIP8f7o7K61NXaTzFmunvWEiqgGJb
6Rs2PSe9B+dp4ySZt8jxcEI4d59YxfF05uUEyHl7TRH9ztzsfTaH8Bseb+qUYoxiY4Xr/U326UpP
/dRUd9Rc8NslIv+0prLKjOPRg6FYtyvvH4KKuv8+OdwEjjHLZBpH4WN1y8nbDJpKwM7/Wd6mYr89
sHRmtwA3HahSpk349OuZ3/TCKdPLH8lizktRMqxcj2ynROpDq82yBbHR1HYhWY4pOq1RDJmTHnfK
7kLNgUevHQUheSpZdhm3XoohXmRE62b1ct324VPIylFL0i6vAptx0iqyp0sxk6Sox6jYD12pThp9
YSC9LE499ij40JiwWvuoZRpV3iTgp4/8a2VsPiCpPIbYNGs0KdRs5Kz3blqI9wVvfJlYcG8CYIO5
bfEIgX4a3/6GBatQk3BrEDPzkQQPMUsEg3MtqIgVsuLDLwaxxUVeFPJgoKG4diC6USIeh8GyxM11
7JVOpemNeKj1ECNUUE2ZBd8LpMq9jUMKsHGjDIxbDdiTJvV/uWurGgT/M95p7oy5GbihhGhfGrJX
qzFo1AnlAVQ52mS4nYP5fJuHRk6JWo5kDZsnegqj7KG7iIbx2YVM/3IVg+QO3O3ObD4Rybwd0vfw
aWAprc14Nt6eevWCr905WeOskSMXyqjlqxEVYIPGkxxuuKHI9NfaydZGg5m5OE+CsSstu+oZWFMI
3hiv/H14dbxK/mmEijYVNYVfxYkQbiSdPn+B40jOlwDpt9ykcM/xbZhUkmainrEJCGVdoGMAbG8Q
3xBOnoqU+IUujdjSMJ06FxU1We/4kL92VD1P+kAH1KRIZhO48c2Hfb2ZBHeI/S81pZtQEs8qakVy
1YokP3MNdrZq10BpQbChVQuo+CEbuVRK9FJtmvqmBTGdmB54h04yH81OyFzhl0S7autWBiJZNpiS
QdeeqQAS9/hYz/pl3hTqK6Dd8wnliEkiZ8/8vYdBTekG0whu9AaxaewALS5eOdpNKBSAmdp3+K55
FDN/OLHSlVJFYohVLUfdUorLGZ7jooZv8I03f6nMnzOVDBacsCumhaXSQC/TC3StdESY8gxqL27u
waC5CNcZkS80c3uYmezIAOJ1fx6dmVBNRmwSgiwFJU0VpEQN/MNf1XGQWn3llXjOxnYyyret7LQd
/1iK6kD4HR6W99jkFDtpCuZDA+SuouLi8IdZNgIfBysp9O5AIrNL8ZvWsD2gjH8PoPLTKrayGhJ7
eok+6AAfo32dKky+wn5U20QXYzOFJx6iDaIfJ5bpMHVlzV9sbJ6QcFX4JJoBXXFAg7Z2rlBh6Rlx
AipUazZlmxiKKkwWgS9HRCnUwSfvJ2NxIXofenuyVZoQ3NrdDXmrPc2n6tuQASY26dfHqVvon5Xr
NNkWD7fEE8/FyTNyEJmY4q0zhWMNgi2muHgc/EKqnwFkbSbhIhccb7hUJJYsKyE1spN7nWQGWS//
qjsXsub5Jvcwt9nGDz6wyVVWiJmZZ8ZYYWo9JGbtYwqnUV0rJGnLWQ6nQ475JGm4DypnvRmKKgxD
L+HMeR1Z8xCCCvw9wSKR6g/emGsmAMPYuOu0YteOtR4+bBIuWoFUJDwLcmYAyoSQXUmLN0aGVgHX
qGBVwxNafWVeHB9DGqTVFNNBqxx61LDsMt/nfnXhJkpVYEkVTVRFyyzM+65BRy8LIqPC/ac0QMus
WGrSxJrlTaMFnRUftEd5QTtw13vVqvo4bevQTRgqX2ooNMIrqGNvia7056gPmMu1YHn/HOmIaYUu
sCnwIMWuq7qCDYhvNrtb9DuObMGM1h0w2PCY7bhCrZRqu03mn7USJpyQQFj0Wba1aziVsf/TQCjD
qHqbf+lI1Qg8YbmGettXl3NDcsXsIi6fKRZ5W0X5zZ4/6aT2489IrugPuLqg/rqWimXkaUtz4jIa
2YU3y6b0jcmNTvyijr43BNRZGj6ayyXtk9oNsz48rpwFJI1LbqfW6MiPnPZ1kS6aiRZQq6hVQjvg
GvMHIBQkR5AHWGRjWZRx+rhAQZ3paa2mvFWez56Vixty8pd3TSL15EaVbDmVdJk2Mt1EtziRcF9m
6GxD9jPkfJq1ZwpRw87sr/Cdwi3IHHtfEe5SzCOgImTFiqxQi5ENdlRkJIw8t92rC2OTGNL4hGlZ
IuALOEpuav/C6HSmOUjiVleaxxx6uCtp4C07p+MY6XABYD/gDdgU3QQN3PHxhYJBn8Z4zMsjc9vZ
qZ8NiVqcUZEQBl8lyNUye+STUpn3XlhuXlvI26pftTCd/1KQRLEpLxPBSDCyaj1m43JTnT2xG6wR
GBnSbZchV5hIlZYaoSgbTes5sbQx4xXLmJUWanTxeM2nx6SLd1/6H9CgtGAIiAKeR/1ae5JlWTxz
z5ecvvFoOllt6jI9TtcrOCIYQRl8Ir/6ZK6OzOcYJzXjlQOOS/s51vKN4QURtsMt4TkObV+wUViC
uMqgCda3SvM6njVdwiUu+5I8nktXtwwn3YmdYaKVkwoUmoU7vIHqiyi/OxzyhBWPncxt+sCl7cMA
tPuNHlf+uCk1ydno6OxAGfUAer7O328GKG7BDul7lTr3xRU5xDEpBH9DFhNWpPt8HpR487YGREOw
n4CMlwwzeaSLKb7Aqy+J57w4xCJkd3PKl8w1EcdEcgt+8e3qr+UiMUxcTBLhQ5gkAXwFmkOc4I5J
GU9ysqFmbuk1OyZgnUYU7rptgg8j2wCb9GRi6lKc+MPb9DEDeFuMpRfOfYJV8uDMclgb1ObcUnHg
fqLoPuYDHap2oJUCasLQG8rRF6c1q0p5JRTimXjH86IzJ1KZ2g4olnvKoPVKluxbwAJkrIc5gF7X
bTChzxdupaa4FTQaasUPjU7vPhuH9+l98PZeSpjYWcyo1PbosSk083OV6UyRXR9otzIiWo22/5e4
0JnxIbEZUdGfiLvsub80bYVvVDdYf+r6FGA90fhga7Tq5zM9JqOJdaQvkGPPRYf1lGC6U5TLHw05
/lVH8z5/fbuoJ5/tKgJkCfu4j+bfhXf63vcJWL56262wfK6vOefbg1EvierwiKhS7PYxdYfYRywm
tp6xKLWcMaYQMQeloQ3CWIrjJufynGKiY9DINgTpJcZdvX76AkOKqLCup6bkeiGCbnRTg+9GxNVX
D8tK1EL0ZSR4qvwG9MAj4LRs2/qSj97hT/UZ6FfxKuCfhvcj9akAaGdmH0MzTGmNMP8OCvU74AzJ
AzChr45GMlvnhYaS3pBDefw+CO4D1rNfNX/GzuigKcSNJlpO3CKDbLnXRZWk6pqk1ERY7KCZMlGp
U35sB7P6ik3pRKLmZUG5jeh0ntls6IeQfjFUlpZ8R+H0zbo8d3rjdMgs+JqA46xGgkNATOWUdnwm
T0dyr2lHCuQcLp9ffalIJwLOxjrhlNBHZKTUftSbkh3ZVeICGnJtHT2YdxSwNb8qmVLu2A1aOQYB
D/33sy8TerY+KDcKZ3dJ9LItuPf7RRK0Tghs75Zo/VqWxFvWtIfJVWEPOL1dtbZM/Ll9wcFXJAyv
0u/zyo0mKLfFH8rJULL1pmiLrj3U7jX8qneWv8wGeeVQYgVaAsMVfST8nBeDKeF+vURtU+s0i4G0
xGuMR2jVJSMAAiVxiKtUExAB2UbXg19iq/accqhX1LZHGCNJqj/WzZTtFevZyk7+HVACRqqYSIZr
+XWgD8mCYzANdHDxcdDkt+CfjDIEmicO7IcMo9D8CCZc7SmFgI0RIEfDLF7wAAUMm4d6LP4anU9C
t61m1ginfmVV07leA7KK+JnN87QXZzguMxUFZ+HFOB1DT8uaqnfrPggwmGzcDT57uKGD29JFZpa0
zWxwNAsEk2UNu14ramfpQVm2oS09OYf8wUPfH5yXDqTw6coIJCwvtKfSYQO2An0FBCAwIetAPzze
RJlmRm/E7QHw3kDWX2dl8lm4St8JN7na1imE0o8lLsTB5M6Sp18uUTjfgb10COH68j0MODKYkLJI
83fFTv5GGHfeDKQLvS3SN+z9R68BKJFrg6cZy/12nA/ElEPLL9dCYU7cX9TQ1/xhmaNZZ87as+5o
bgqeSAnsqLNC4jHaTVwpP85OZLwFETqhsPptOSxgukHY/+u8rJH1RLJCkf5GrTxpZJ25ZnSLh8AV
XgFG57yWuApsUuFt3WwDiXWBp6iLHtzRM+PVdArNXqc1ncyHvrUHG8IAH3mjYBS1tfTJS0TVvIAR
/lV86X05CBLHS8awVgw/HiQLp020vma9DDVsVJrtb7oYGztoPBMzWI7xz1QvEeH3jL1RlvIWly2a
2jj0/vKM5LSNs/hWacti4kO3AT2kfWUZ+LV084zsRTIAgpdx+ejB6PTwIxxUh4AxZAWCurGB2lYz
ZM+hqGZLLGhfWFoUnVWZxYRy640EY0qoBqWpfBdsoHw+o4JiN2/HEhaq+EtK7s2eNTN2sK/HyTMJ
FCVMX0leFWNS036k8ciH55A/hdEKRYDy+Qkdn+Lw1xH9/LGT+ERPL9EFqJ2iioc8qaV3Q8EJ1jTz
xI+vMdzZpCjsjDeZ7sgEF27N+kKZZ0WEoaC+KFhR1zVCF6w0H1h+BqVV2Y1fv6DGKlU/jjkactlq
AqylaZKpy031DwSEQWgvtPVDcqm8J5jxPNTRY0kvmVi2nlE8Mvxe8wT3/YhzMLL+nu6zac6u0zfV
KRA6YvCMxsUultY4tOCkmPwjHfwPrG2pffSlBiHxE5NubWY0NLXws2ld/e3QcZiPchzItWLW6I/n
9+AkP95WKeEGbx6dtfsBSRDZdkmRp/BCW1H9Rb1OdsTzwZnCznyk8DIMeGPwTuRuXI3QVvUJ4oaP
7haG2JdcymFDetI/h9LMNwKsDs118/cjm6gHICjjrGtUTXeeaO0Jp8mXIS1Zv1+nAUcHTKAYThrQ
ZwfOpR49dqIDbE/8gLgHTGdbaUVOszPZ1tvTJdHpWwR3hT86rj2TRYxGqu9B/9QvN7FZzqMQ8yRR
w5cO2jw9wyZnm5uEEctz1fDwHjrMwuUMBTmBAWvyclvk2Q1563sBbD3VZT9AmlY/zaFE3UsEnFxY
sDKCaUGx771g8Zj2Ci2GRyCBskNMVAKep+FjHRyrI6BlTD9Jo1Fz8XpH0K83xsX/nGsSKIO1+TEq
nu2d1dgPl7tf4EOnlvKv0/B/bQi+loAJpTk4o4Muwbfs9rtxrRwaCH/9Db2bbHxaKAFAGCuqVPd+
h0SjBJAWO/TH8eBmjbGo//Q1GuRDJ7MwgJF5xGyJTz6E0TPsvBK5bIjUbAupTWYIVlAiu1+NJhqh
3E5VniTiM/iruhDKX4JN6+Tus2hyNF6pgBr4i/J16TOk8wSWqHz8+r1nek7HjLIiewYzDcy8gDAF
XfXa8OzconOeEwCAoEyyS85XMqQqoqfNuSUo8orcg9uoK2naf9KTBnh3aFnF74cypFZB7TPNlgY1
Dn24aR1CnIT61HprhbfL6fE9rv5Qg4RY/7FIyQyCWPQeESXRqJM11M3joELeway/88ATd8kQo0TZ
AptyqZ9n8/CT7pCJSqbyzXCHKHJGV75Wz5BGAoT7RBEQ+Eag+cYkUy4Xk9mE3EZTF04M7THW7QwT
sqQbM4/qZhdYWFxdglZ6fIdsmQu4lQ32VBnKN3os8uX6FdOhK3y5Qe9yZo4URkJ7hrTCdBSgggzi
LRah/8tOzzc/xo7bVYXjFrgfMbq9v/wmCz9sIRk84wRupjAigUbZ1Dp1BsLRBkA4asgXIAemyNDj
Klw61Cf56oRJTYbJUk8ROeNZxZKGw77mdYXp8Q/pM4OsSb/mN7T4fj2Y/6NyFwsqDJt4oKo2xB/s
ZuFmMgaebJd+gYs3XQQeg+EIFhZCFbAwlDg7skV5H/D37GAnuX3NvDmwaWI1s+7qxs4NbzIyeovb
RhAJbayEu5irN13gix6MnVEbtd3HRq5I7qTAZaY2FSE4Gyd3V81V14MzcMYuYi3oXh0/1ZRS+tGo
e3PMDOQfr8XzqO7sT1ERipyPpg0TjWUVlmmFr/QOweMrEW+LFVgGpjff0/SB9gIS1k8AshariKK6
+k8uQsXxANJPavtBFEOIOysAp7qRmnB/oA2WjVHrjehz8kwvTekqL4JPe/f8QOTRV+DQMNdLU01J
by/CPBRrd2u2+alrXN0Bm41QAgV+BCz557MYmQItZZS+x7DYXsgLtchY/GqlNlu+1tVeGuDMn1fE
0+Vw+5va3chtR92OvY/8D6FnxUR1dixXYULGLEq65q3RtfT0pDUwimFq545rCQZxtMSMtjm1q4YN
k27tqXWsfJ0oudDpxVwdS5SLSq93GKegg59AFJrpyYvvaxg1drzHPSXiM5O6fyWpB0o+iSy2gNou
qRZfYupygbkom1PyDZ92tIAdL5gYewFYD+ppxuSvJDfY+VsTXXxoXtQvgOo5ye/hgA386fXwoF3A
rXjDpdPF/CK3pGsvwB9x0q358haJlkiyZdYIw5EMUso8mraOhTAonE0deRYKJIo79OyiYMdYh9aI
IJOvK2bgQGjHG6GCfy+9Ly7+FGUBI3whA8TkZvb3cjHdreOoHRYztZ5RnOCtdrqNlslS0dgsdMzf
uEhZK0wHRZZ9P98CtFVDI9U99gWFz+lOgll4i+v+OzaUJY2ioKqLyXDjMY2pgIQ+0nf/sa5UgKE/
5jdF3/C1tdRBRdr0qmtkQvMTX0cNye7xHi+nCd2gcIS07PqEcYLT0lKxFP9dIjNlyJUEVYN4sSHC
E+yij1HIaBL0zZeRTH2AibY+IyGaW1D+Zg8Fc9QkVghEpohDwj9sqrAddKUxp8cjf82A/VlCm19K
mS7VaJDNO7+6e6tEOsf/CpjoDHwDQGBJnBJR2Yj9j/hkhWa07elHRiPEY61TYTP4rgQBi36R7YaR
6Bbil0TeEhhC4qp2JHL/NSJVDoelJSJ1pAVKiJLJlMBcgOGfF3Zkn5sHGSNPJZ5hncv5m5Q92hP0
ZitRzw7kvrK2j1953Ba2oYlvB17DkHAchYY24YBTi0IZXkMu2S1taTBfgeJzIylcGCAVE9XgXztZ
ejt1o+8atn4x6+SAKz37sXe/ie2Pw7k/eB842r/NdvwDOxoZZx/6ajgpnosamp3WYl5wV1CEIVhj
iCnY/9J+nhXF4jsZewppc8BcVJrQDJgL1yFgo/Rv2aol1820e9HyYpSADnvb3y6ccvPHb4ekFhLC
lvstXjfKqrOgr51t08wZXeC+bnZyJP976SEu5WAcPo2dxj4qWTgjoxjsWWH/c6X0l4DTGRuby5jZ
lrn0ugwzMFMcZh2RcKvfWWp+cQ0AvKZkoI4PdM7Jshq3e8+qp85qIy+PjeyXyicH10Q7Gd18cO8P
epAtP7ewmTc6fZQqUw86Qe/9P27OwnEKFTfSKw3s2sywf2WNqHbKMOY84GHQxNb65Uma4NmeiSt2
71AmDuggf01vwWrK5HUFQS0UFVoToNp62OT2QB1EfAlN1zyaOR9kH6mP37N9S0cowLWwcdQgFDJd
DDa6YMa+ql2v/n8z55iYVYbasE9lFMCb/6MjezzwjgZcQQqRnYE943B2XRBCm2S16YfQKouDxtoP
e7mJw7evu47iRiueX4c0j+IU+KqBlAZhql/kyUjKo6RJKdtAtw7CXgJTr+90TGPhTym3rIjZee7P
fT+3vpatmbwjDjivkQsyLjKBRJk2x9qo598M78hqdWsnpgTr9cgVMv01GZN8h8CvECpL0kok36B7
59TbfleBKc2KiFeZYoMnN2Q5rfCQ2cRs0BfmFaOH+sM2Tpzqt3h9gQVUQqDfAq8nkIBC3kMuhNP2
Fwl7MUP1Stbqc+hmOYhgJFOu/IMzk4YiF1zuL57PWZLnoOi+q0At/KKKjobkt1+PUWMpx0EPuibx
TuWrSORYGGzuOdUdXpADvQyFoelnxeEBhySP9UXBeo6qYvBTu4ypLnOIDtdJ/FgDFbjuAWJRvkG5
IF80exPF9oZTxh85M5kFXj+HBbMYXxjxhgV7rjf2Ej0fol7XS0geUwbtLv5VZC6MwIDy6hZ/w3xG
I/ogeBAGA3Y20UT5TQbPJhe5c4Lx4vWottRiPhIY4CloBpQkPOG3Wu377mMFJ4KSMZnIrBpBRCr1
PtakAh0kSIGFsxdDes4BTv5gNJuKiawRoPI0P7Gp+Cg2VM/LbqS1Si0Wq7xpILnOm4pw1DJ+GbzF
Bcho0jjSxtOjwo+1X0CYUhbN/0DLGVhXChpVWK9/VhWF9LrzanhEE+a2n0SzYXeSKPdITagOCjUm
84KATNN4G2rfNlC+Ht/Te+8P4Rn3bG7QADWK3t2a5xdmeXYbizTqqfeUBPYgeokjU0o7ZHPp/j+6
V4fvvOaxyc06QkTpxE0Pjc5lRaSOF7KuVRRm+ILTNjiKGCLRZLH3LW1NE0WHuCnFPtolVKD/LlkS
zLoEd3zcjVxCDscvG4onrG4Z9fTEN65S/KhmC5c5+0HuUlyRVxxltXr0LqFvnk/g/q4zjzWNbi/9
XmOLKfEkX5vGF+K2SqfCvqStqh9IRuSGFkjdgI/7iSb2owXWpB50Vbe0+813UDL9Bd90GV2pR0nn
ELrayBNPOAxtaGL/YNqTZp3Byjite+AQmFjRxcKHZnyDtwijYWqcE9dLqWRjoJjrd/NYxxZJDJ1w
j3Z+H1tAVz/mgbS1nlhzDfkPyYYmw9Xx6PmEXpsXM1gWUuwaeoLvOr9H/3eauAWJdtMqka8AkmQ4
pTnr/jYp+OZAzvOkf74W6w148H1hNELiB4Q45PEtsAz+AfLKzsI8gVcQhzoT1+ItWMEaDcDpUMs8
RGP61I/tK/ez3dLpmhmUDlS3B1B62YtV8LmQ+YJrPDKm24IvTQnZEMXoOJB0gkQ7CTRQnAr2aP1M
0ua8LKPI9m2WcjRHPn9iUBFFa237UWkNZtHfZSEpJmvqNtOv+trMS242saDJ7CinWFaKXIoRbCi8
OXR42Pt1XONKr2UBMrQntNjZ9mv44FFuMF3LrDcfFWcFKZt8GWn9i/YuhtjafiufopIJbNj41Aj5
oajB2d/VOzg7cGzXofgJKrg5uvq1VrHCPV7veKFL+w3tlLIF8YSNxD+RWp7Rm3afXFmXIzz0tnnH
D56ivTTN3yMrBvYH3V5kPTzU00q7qRudw1GvT+cFzRJEpL176Yxk9Of3sXgAcaXCpPMui7wSw+vx
jCyWxtTk1wO0RjFsfD3T8expJtMTWklpe0EQPzT9HPsbexIxbQXvjsBivOuSH5OCW2J4ybDQiwe6
lVwkP3zzzQOuix0dNJdRbefnMsxo/nB6+Y4U/vo+gOPmNGmmWm4fK5bMgSMwie3rcXG+UVT36nwp
vurpG1B/2TQudCE1qJMQ8iFqEEs7YwBeSPbcFgAsLdQ/Loj/CQSSeOcL7iEP4qMAAbhD4Li1qIAI
MyG5sVNkVFXyciL5zDOVdYrTGPqygTVDny2x32Ev1vaLG02+YnL/lAUo2Voey2EgRYLo+utFY15O
3RAM97N59lG2Dj3Jx2cDavOIm+MQBmSS62E3xc+AZrpjIpFH022jfblXAXrVLRPhxsTpg0yqPj1s
gOegM6+Tse6CsWrla4IB1BlCGrQ+7F/bu7P+ZRc9RT1o5aPChA4Ioj4LV2kP/qQOMxU3PvgxxBSe
Ph2YTWuuGp7CG6W6d/Nq2w36cv1jSS7nY+rP3rgK8+cCIGsGnmelrsf5kFvfX6kDZGF2rgv23aNA
e/yrapSGEbJ602RzmsABWXmjrCeH/AAAcJanwi27SGTrfk23n+TTtNQdVLszCPJ3on5cHYZ8X8MS
L7KtVFB8hUrUsZa3cQxFR4rB9cJl1ALOXoWjSdFkg8437rUR4yckWdfyHUXaj7p6S3Jzz9wEIitS
DL+2fhSgMlLBznVyZP26tiYcJ0ThMmltWUgRy7G9Si8mz4QsuwKfr66UyimpyG4tsG6eXSlrgVko
/NoDFrtUG/ALHoBIccVKxd83PQvQLMvchsiu+oaMO0ddMyfo11T58UNKxnAswPsUQwnJQj1vI9Yc
34Yic+o7vfD0A8n8oeWRAX10aJsLvtiY8tdPvhgYRs2qjoTHcvmwAi71r4K0apWqYBRxnVV6dPTh
xE2hKJDpuqH5u4heSCmnKa2+dW5RQ0MiXorwMhLgjVrBjSpn7KKiiYGONZ6y8ToPewOU1ZU+2Ybs
u/wPzstcTHjHkMRhdKsAXyB1Qp6tgNHGLpRCQtnMi2EHLucc+707GhS/EhY0x8p6pl1STwzfmYhD
EFRk27qPCD5n9r8OcruJPmvfqVLEfkBKDBjXfYIKJWo1sqj16SsJURHgpGBS/uoonlzZoiuI991h
lIf1NBM1zxqOZF5kO0zki8v7x8nBnlfuwTsACcgY0RvuWItMho45Mbq2ldAQX5xsMuBW3k4cgonx
4UbRC40CWT2GGMc86KMnJgoW9OXfaHL4EExTjzlUvdubCTl2sAuOqWUqIebY9KEkA/DJeQTNDDqc
guFdMMCt96ORjcb1TKm6iz1sqNaI/H/2d4dES6SdxtcYH1kgE6GUVluGab6a1V39Sg5sX1g4T83+
5ewrhLnwPQpHtrHTSj56SnIoOJDkPcVryjRBIKmc9N+4VYIqt1tuUhjwDgEx+tJNfbMwfkpEIZ3L
vOvwr/IKG/Y2+3GXfOPzH/BGi1ICpPuee7S1OxiZWyPUSI3ArBzwau4r+0naUSCkDlKcHTiRdQ7I
R+eGPFtDzeFtgBrJ6lSpwVFblwWHGKLv7iro4BFnUglyZ3HmVkIpwX2wSjh9H1N1XyXaCvdLhUs0
fHn55QH8k04cariwWioIkuelVyGT63xfoGF+H4V4YSfg8w6zZtibpndi0nfyyT8VqLpwek3FDz09
FkppuJ6gMrMctBWR8ucA4ipqxYuazQNgi5kAt2h7YU5FggF96RwB8rrXP91Lfugoo3U5QMlnZCDJ
9H5vZLwKa9qwN9owtP8aA68USNCbnokLshskydc1K76g7I5AzthCxNmfcdjgUPnxGEZU0eHrd1bk
+hkwVHXGYysp3wtv0y8AnqaRJy0UKSCM1ZAIBahHZVOyQHRoKhnOivGcHCMkhI1Sjpw0NzFORPSe
HUWGRPk+cvlY8Dymd+8X5pYCo3uEqcdPdzBl6y1REmiBM4rcWF9T6hXoIQwr1y9jRVLyMU7+qWK9
wpg92cCXCdLFRLCxX1VrCzN42l45j1e97LlN/pyhLgnF4vohqaWJD93SWKG7pX0U+kWmZP45jcOo
iepr/IjIJSQBH5OLKE9pkHWMJHr8JuZsblGroP1jw+xybhpLi8KgAb8KIgxTjK5d70X+RSaSCk5y
UEb0Mk2rhH6Jh4TChWWGLGs1RXHJs0qhP8AzktAUn+MD4wMMJV1lmUwACLWP8p+8spqsKH3M6FBr
zKod2gBiO4MbxCt3SNCYvYAlH6hnYtSzqLxwTLblxM3HvIcVBZkXq1yeEV57m+Wu18F/yaENB43o
B/ezfjrTy3L31QF9XbpW4ETOAMtbHcSvjt73wdsRtAVRef2lFL1FRjyD1LLaIn0rIOmKzxo/ZhuA
2ilnXizEK0futiG5G+piBHV/J1kgWy9/QlGDyiDwQbspcu6Iuy2PGstjS2ml5iHvWFPXgDA2y2gj
RD63azI1Q/rOF9CRfNa1dv28HPXqGJ9RO2mlHHVihEMBeqJ1kv5nqQ0cb+Dw6jigNgHDpjetzlY8
NVdPrk8b0IZHyFYNyvU3i9FIkFYpuH+1dzPpT2USXu1Te+23F9kb3sp/WYiJFMjasIxcAAK+FyBZ
e8o12NsjjzBQhc5vupRafMqYHLMuiBsDZeGrmHRp65GFPXxXyeOWrhoKyMs1QZ7Xuio1x1rpdxjA
r3JPfQeJQWyi+diWSRM4JqjlCZx8EBn8lQXJAu8=
`protect end_protected
