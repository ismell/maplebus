`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kSRtqFeRldJxNwMSmZylQKOWBvPgcswwYwjcaCv++uEtxccD4VmJ9SIrpv+AN+kY1IRh0LbzzvfK
kVLdV0gL7A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ln9W15bwsrmxftclpSdCldSXJ0RM7hSOf8Kev576M9X9vVkxA94za0R/4IdNmceYoRENxtDrWruT
1UW/34cyhrTDwoh2zJHA46CoFn08s6bQ6jEQ8ODz51LlZvj7igIlswrKQNgOnMid6nf7Y+Bw9CMw
/Xy4rSckqDwXAPZXmaM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jm/xLU7uqDYJHrV0GSI6ndyHJ3oU8O8znzvl01OoyGyCtjZobPpFpxy/NuUCIgdqOHihiUhzHx5y
rgd6ZaRQl5o8x0UPp4epC3M/CasRvTp2DmjhTf8mq2wxKVsNjr+UJhUqEOBgmlXZOWnz3YWfWx57
WmvXYLveUR+8770PQbqJCeh8cln0vNbYr9bBHrB+CyTo4RRc1DcLTk59qMIUZ+wr1pIecQ65G/+u
UHo7mVxOMnpt/L7vHh8FW+Xkb89TkLkprB8eCHOpyJAuTIvMuN8TTM1ix4JbKJ/uRa/yl25Fs7y4
eFoJzKRbYqZZ1vHIiWb02ZLYuXt4ShDCbGR4tg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pMXUglZsvdvckG2gYoy06+LM/92JqvSmTr+VyEBnMo7/ATXYi6LkbsVW3XK/6G8RhHxjJdgZP76Q
r8vzm5J19MmXPZNLyEGSecU0YBzI+ZXFm5uk4/bgXWbqHKAUjoacbX5//sRZmwtzGannuiaN2uKp
lVrRo/jDL770TGnhmSA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hiLXLA14TYDfWRfBKb1k1x4sBG/sZp0xfVUc3VniU652cSjAs/1oENyUio/6or+5Ka1BhV+F6xYT
F9UEyUEn4IYzPbkUwFUt8EwkM7DquyBGOE2SIQpd4t5zrLBD6tUTlPRlbfHdTw+DyqSeRDDZNcbh
rR8E1Y6p3Jbf2zT4i/5pMAQRtz9/gVhgEioIjAPmubjIy0NNSdycqB/WykZnKJ/y7YS8LA64HQqY
hIazxWwcOxOKM5HGziWn0oQzRH4JAtjYyx+AQvUK5m4gofGqnrkU4MoM2PERQoZvCSuAH7YXCXCw
f7O2To8FnSZSNWLIrXlafuCz12c0f9RONI8KfQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18832)
`protect data_block
Rs36OAy9bUCh/vgldYhH3MraRvbG3jb0ykBiPaadl2PeegQuk10obQ2Z0IJFIddKz1BeZxEhEdCy
bIFCoPsNgBEGgyXbddF8M5r0VJRs7eaSlLClF4IbSAd7PGZJFUPHcKVULjrVT/Am45OdP42IpwQL
a7GHqpuFLBgm9BgQR8RyFMX9AbCspI8D5z1wByl54Il6oobfTDO/Uyj1lwPIe3DDOH8HE/QIuaEU
7lbtbF9qnKmv2KgTYGj7Onj7LavrFtQUgQPWwDVSUxZiSpoRCECSI5sROo1sKjV3q5uFjObwdHlj
7YB5+S0oQE2iAJRK1M3F+NfPNV969aAR/GrzRn2GyuIM5kOKiSvT8N3XidA89E25O+nULt84h3GH
W8c7n5iw9cIC22w/7UfqtkDWKc53TLIqORadTcZCft8Q9j6TirCwRBhkE7+fR8vmFTda+eZUYMRW
4I0fmjLcHUQAhubv+XC+K5duI9GuT57q+zYU1r3xuBvNWF24JWzUdDr5pQSEodjIwtANGvOcPvuq
xR5A8yVh+57VeOBdMkZBLOpzM2xSV2e3t9FFZa9/CqZRniU7URM2fEIOpMrEWQA58d5XgEBP5ocg
D/luYueG7iSVCErjN+MN5CxC0/yE2SlQFUwOBYSYRGiplMJfJYlG/RQ2/IEpof5+xud/KYKrt7gW
n7ploLh5562l+n2zVzKjiSBav/GAiGPII/eaF/4kwjcqHPTzkCEj0N3W1E7QQPBPcSkqHCwOeIu4
do+HWJlmMlT0rJm9OjIS1AKo5OST/MRhW3JSiEbtVDdg54+gf0zjo9BgXofHgXsOBokt+L7kXn0T
aytDjJPeDubUdRzTneDLWGrqJ6IZ51ouB9sMYwF1TWtkOpsbBTYb8F/iEYIrhP+fYmaAMPMsYpRF
6yAbOpFt5vnvegefUUNBDU/P74KsRdE7lBJBFtTWGQxjX0SfPL/kQWCV02OBfUdWsF0MZ2S6eQnI
Z3prlMj9uhd0opozx14a0WsasbvKMqj7h1no6JnkZDTDtTic2Sxk2YQ7yeeD9YlQPxTGc9PVMH5n
Dx1hKpwhKSjs2SqivnzUaP9SQlHGBO0td/tEp9mPQ5RZQ+5PFBZvqwU0g61EgXIh1Mv4ho/JUOHS
BV/LIXZpsQJTq/IjU4DRQfuypT9/71Je9FSs8VauRP71663NXo87bcQepTCEP3GVjvNF9gZ1pdhD
4EPgjeox1+/BuQK0EfZ5Op40Zqg39gPNXvTUjYbTgNl7AOon1yxzP0GdSr9wI7ANPFyUM35ExTrM
ZeG4aSdvRgjGG+/ulnBOjqW2o546Y3HDCW2en/4+wV5Z7zsFiTjfmb7m3wz5RHnSqjpiWdk/hCLL
StpzWaq/Jx5+0x3uMqMNhax5Qg4ip4b+WMddLgXFUIO4a6vdErr2TwLOyQaCLrxPGF3JPKyB30tx
Z5U5xb3I61INXsHKbVx8R9QeTfQo/vi7t3yJSPm5wOTZ68M+0y8pqCM0mvI5Yifk83vsYvLlTiIh
S0hvfI+bTzrB5eQwiljp4RblwvKFOeYY6yR3xxmDp2Ma5T+tOJXquYQgOcg9++ipUTwtVWssYq1+
xmfabV3Ol65xWx+o+pliEJW88V1KGfl0w+Ty0gQvGIOAG/ucTrjUcUSFaMVu8QLpgp/AL+2/O4of
CGxahaCBWNrOT9C4QJeqeZdPK2ziQ8/Qtg+nmQ9EIXdVVcSPJa7Ug7FwSuasHm9K0EQeimNO+mai
RpMHl8BlUqQsn/BohRhtWVjO0K615y+pmELlB1Zh8ujkyChhnaFma7F49T9BGH7Oe2SPcPRsJgoa
Y6iwHX6vuCzEpE3A602cC84h00gDl3gB25R++i/Z3VQWzle/JwqGcf6KAVKehD2bFTGCQqt3/YhV
KrMSfaTXYg933ji57zKi7v7ASeu9cWwgglF9eT0UJYg5A0MxjdkZ/yLRQS4LniJ6cS8j+FOKRw3u
oegfb2+7okPBR+y4x2t9g95bWbOxIm/Ciqwvmt9MKdQZ19AmzxxhrXiH1VPZjjiwMDq9SV+xga97
Q9wc4kp04CpOlbXJhd4Y6N9shA9QyyV2y+2oY+mdeIZdtTJZsME6BDQHwJAMWx0fXNAaawD1BNDD
pATKdKk1O0yLA0RoPNsyYMWCeBtdpC37u4hSATgCS6wKBk936/y8maEWJxfMHaB+0n2wMFe4X3WG
GE7BOJ02It5c2ASMhmEZ3Fi0kK2qQwSxNelI/R/kwR5i5XKVGrSUCnJF+EgJEHg0cTnh6Kv0Lsr7
FlhWRPo8JveMY9RsVowS9v9VFbiG82gYgoeSqoawk0nJgG2t8tKgLoiDMwlwxsvqvZSIoWVtco+Q
g/dbOGfLZmW/eHKuwR6WZV40pOUZCLFfF6N5S/Kt1DadGYhqlZ2ifHLcyZAnc0VlyZ40wqmtyRgl
z7eCog1w2GNqFHIssrGDCFbFE5+8baGgTINv7R75TPS9r0zKKhRDpFh+G7w/SuOrlT8Gn4lqs11s
9Oi5nvQkoNUIHdOJBvwNPxnmcagk0rbIs3HQp2q7MHZoIfUAc8eKXnpruofWOC9aSPR2TMl48LSV
CEt4egu9YxgYqdyEXyCH4yHxBt2UP+VHPj4VRkJ5pLg2JtABam067tu4JLsOCITMKksJ4tEXp0EJ
1UHL2sR5rX6VbW4xCOkkaoDabn3GdL4gMDMZ3u3PAo4+j//D9nuRTIm+hR5DotpTiviFE4SVUIZc
iiNrxW+49MkXOkyvoGlGJVdXYgkJQ1e3+osFQHAn9PEb/UBozWZCElPrptoosaAHuBWaazscNGwZ
NsavtTYFnWDPsixBnMigt5vqlz2L2DZOJoVzP/sd9tofo6s7GW2efo1xLwujVQq9pc+wmn0q1ckS
cNzOGrAydElcy2mkm5WTmGAY+foKSGZboJsDDhlPyeMccT7vEp92rA3JNRbNNYjBDj58zbwLXG7N
H8FhAMQK52DmMfEROedmYqvEFkx5mFzCkFbiTkG/mJdqa9vt/0E3vz+MI0+wFP57MDrSblKe0pdG
6ao2VQBJSWQysVhBZF3n6/DOEpLZ1u47rDhgcIbZQUhB3oniIETtssZAv/1EKqhgcTtMgnPz14+1
cGGNYbFuw80MXQGexbXAjmUV3VxOXU4UL2XopqcXKG0V3ggsqeoMWdbXFFLyLSmPrtt9zMy8H1Gr
sokd8eyjquS9RIgMTlTLmhOceUcnAnPm2avHwV8vYT7Owz87NMm/W8yOXMoFef8oPgZx6SxO1ijJ
T17C0tJRm8tWWmXlrNh43MIV6FRmmJ/DCUPXdEEkKb1kw+ujksDt0SkkkPHAEHQuVHBMOsVvkh9a
VQnYySnz4Ua0h+oN8HQUbI2CW89F3t3LG46ffU0OvBz9MBMLExmZvGlk0kIWoEatYmNmj+eyhUj2
nNwj17YxkENOE82y1I0nwNiBbLlpgTeKLeWmvmiQXP+aNo14s0zRnociQdiSmlRR+bNVcLlSV0aM
QGmXSmxhmcZQoEdb96GurZqw2Kt2GkuO9GGVFMpJV980NmNTbQXsz8mwV/m/0zRNQub33pef7U/n
BcVg8HOLgzX8t7BDDNH9uleFBmsnigSq/851+LSR9MIQnJhGV5hhU0rz1JBTuKDIThjunEaZsYuB
ADmtqwN4xE7VYtPe0H0H9aZE2l8LH19k1uljsLAi4m+v/Ta3nv0ZG+ku/yAFxZ3JWYy7OD3nwfBt
KJrvIUnQu/HWmz+VTrxKMB5ZM/PeculaVQk7cpActgQ5xru5/1IKrHOhXgP8DLBIkI+h3ZhcZ1eI
yxMn+rYkFRqvBImqcE0qIWd5i3CTc8lVYKNCk3Om2RuyOisQ+t9NQ/Ul5aFtE4f7Wo7aOueI3Dj2
BYcyI1cL06XTCFPjodCIv7BfxCRZ9A9CHbnlNHRYs7EBUSifrtZqMknUpBGkyHzX2QlKTWoCgjGP
dxndIIblvqmeQINwaUzZhyyPYso7D2tSKVWHsp1dUTRc+7UBUyxODmg7fVw9Ucl9+VEL1JHgYbwB
LlrY0I4fuL5BwHcFeuQXZi8ooWnYl8BXQiN5NoF4doqneVOdolf2meOlC+AzpVNBiOn9rrnSvIIA
faKnC5mAV0xGdMIMu4JvwyZpEtj1pjZkOhsrqzx6SwQOeJFkrv9iYYwiSSHOuPfvMsPhGMra0NQC
EIV6p53C7BF7rIciocitnUBx+myvVC8lcTvOU1jxxgSOe0jhK1R1Ib0yiCuclDWHSKvRmOW54ETg
bmIKRKgn6qAgsyIX6DRjkiSsNlWSy+HuDzbu+IJEzOPrBanVhimDnZ7UK+stqbA6u5bySYTQLqzt
fbIg474M/yUZtnV4vrmQmvHWJus/zS9ruz5pmV3cup6CsrGn6OPafFNyRw+zt0eQiOKmWcV6h7Y4
M+mYooGCj05bt0KZh+McLdP5nYsm4vYkAHtScJaHLIUF705tN8TNY4BWCsIZBToe/SeXVLT8ynny
7oL8gJeV/AbEkm0VV1YhjoRdQhHZdwcQkvocWQjRYLE2hoN/2MBziHV9E67skZWWXKTiWJ6HEmIF
3ns4GDP6r6zO7rMZI307b8R2nBu9MSQkmZFPSuUhKf7TEIUUdiRsdHaSshgjPHurGGAZSfbfT/er
zq0WXfUCtHOxUo8FNiNHJU0MchN37HOuuFiBNsPZCFXWgAWeTMYONfu9xJO5uxU+DjSnypDHGMbo
plXFIvp3t/fYWXb+gZqjz659Q19ySxj+ATJKn6fgKl8TBSg6SP8+XoVeeHQFNy8XGLxeEvoWrHku
32EJM8IXuCzY/zsob+2i5T0Fi1Trw7cauWPBgadq6GdDSlJsr5FqX15YlLUxyldXR+9GQ8BBF40f
AsLe94MEgkHfHASbPqUlmPWujwDt1GuATxtyzP5pB5uHWVnXJDu+CxABNs9JmHN14Aq3Kw4iyb02
LghhDQjKZZ54a2oCiWSJfquSxPDVuwwPKtrC0zcB1SYZfNUhnEkbRMnxJF5HJYQ9AOdl9Q7SGwuz
nV1UJ7gQtDJviPfkd2L47kZ2WTWDwmUGSMgqAAR2426k7xj/CVj1+yGskVR3sI7qM5PMH7+GFbjy
d1Sy90JjTJy6656sMj5DBu23uX1lZkIkCmEah4TIq3vjAUATV3FlP1mFosdRa7q0ODmgDwpG8YoQ
8tDLr9fq6xCvM5ao4HcZCPZW8zimv7O7ynsL92b0bR/Ig8BRBR4XSNfXRDA85PwuWfTNQVaBjDip
EKzOsNh2UgTyBiWEwaG7goMB5rbea2PxvR2TsRn17wYaDUUt9Gxpxev4sPiKWLoupVVhwDBwvw95
z47YbwK+6UE5cluW7iJ6rjD52o2A6WOqFd/ipbc+4tM8dc46Z4rtTVCg8Tejt3eoSxNlhU2auTlj
pf39YHfTV3klsHvwUTKFRm0iZH2C0KZEUgr10+SaBxFcKZ+/TKqh+F+3wfKbMT0T08mlqfdnXVmU
3C7Y2Aql1qT4pwXlq89qXStg4pT1lNL963O2O7/vLaONFpSpUkSuzUmJHEM7c85YoAsz8aMqdVN9
0Zq0w+5qFoLQE8K/rb90jwNC39ZwPn1FMQ59b7LOWpfA4pC+HeTIRVpWwhL2HjlP0T1o2Gd7f6y5
Or/mkfypD8pekT8eTo+Z9U30Kc2v7z0P4FGq9lQr1scZhk9PGOWFVtIIMupGoIXL0u+tlieP8/Fs
JIsOrA3yC0Pe8P6fcNFODP/ggk/9JLNv1AqMDGPw65iqy1JuIVexrUR4E8k3H6oVQwDhFo54JrfG
T2faz1znlDloDd4Y103iRrkFa5RSs3YjGbWJB+g+gAAj/WI8EFC/q+lJh1nejPJCTwFEnz87lPIy
a5dX9tIO0h1T5GJSCM5SQLqO+wW+oFplJ7/2SPacmOCBYL5lIoukLyU2FfdOiHJoWMR0n5NYgkaH
XOcvSoWwAaQb4Y/Du7oFv9ev3yXruWXEV1/J0bHpv9Nb10cgYdEE7eJEJ/voT7roHMoiNlggctgm
sMdKFuFPLNhuoMxBZjGuCYE15TnI5+6J7R2Q0VEzF1wiapLMwU2ok84NhIismh2pb8QlIftvz8MY
lnqW9aXC3mOn/+i/HM3QnfzU0uq5Vvq3Y0BCJzXHkLunGAf28qt1R9Xc9IlUyYub0OglE7EhSO9D
4oyg8Qb0gMlOJ8pfoS2odV9yPpiCswGC/cAjVFUNrpR4SAsIgW+HvDMWzL8Kikp4n6P0RSByRS/2
vWNPdTay7fEOBfCz7NFjSGiMRMiJPzy/IeqZlj3ho3vb5oaTSdiToEfkUjOVbzeQtFmdLeNrzejV
GBsUVngj7Fv+biQHhOHogm3tMN8dysfzVv471CciG8H8PQqxyoneNh9TaeKx4JT/Kwrg1OdcFudk
qFMpVkluAAs1pcVfszVqhaCnIt0JBuWHuLtYqqmUd4AZaUsQYNijY5JKbwIYhLKgDOB8UcqU6B9z
TBqwcYf3hQsZ+Ikw9GoCpDX6TY+yAeElr7Ih5wN9JNpleqfFMGo4hhBl1lQEO+u3U5eKlr1Q3elE
WUvVDuY/M1nD2IH8ausSYXFhA+VR9bwetx4qXpOcp+U/yg1dYzccG8PSwc5ChQhHlbuLfR8g6f4k
xtBTfoPAsh4NT3yvO/TliUieiHXrrQugqiiF3pcEV73s+E2E2aZZLDRATFHyiFZ9+Koc19Sk9knX
F3eWjuCZiC9qWyEaotwQCM7E4PAOIGwW/g8aaveOps95nVGrDUY2DZdjyhVauDBXhBrAEyPn43od
WYQA8WrL/furSWY2AdBKqmHDJiIE/oWidPoldFaqbyub2dr9pRewjFIYs7bq0tJqalA8FcMpvw6D
WT8xPCPmBSfxIW6yGE3YVKgpp3Z4iWGa9ofqzxUxuOGkUmJtddwGM9QrInXmLXAw3JbluZoPacti
D9ZJYAspdNC31cK72pvfxkwHGmXEtkqSyRRstIESif3PCq3auHjs45pEZJeSteotFU8oclhNzMD0
xqcrqZtEUtH4u9Jhu4UmeMSNgyvGhqj9E7U56a0IRB5XHPGp2kXH6pj3b4NvAaUvd9GXXCi0jHqg
L2W/8xpu+IyRWRXHotp+FzTxy3DKuwoK6Fu8SYqvd20DX6IhdxRS0k2wBLcDIXuM4S+rccu3YDEL
vcM2Kteh3k5zrn+O2CfW024XMhFd5ziZQcSR6yjd5uDZ7EGFd3ILD+RG0SztRAcbP2mkrfBZuT/F
Q8FgMiQwc2A1rDKSPQzz/ztreJmOZnDk6Su6IarIWkjAhmROd16tLwA6sNVypGtAaLfDaEWlFH3j
oOidvHcEf4Yr0VSu9FfBoEbYWSLOg1FeMPgEaEi75U9MpU4EARMYDPP+C1dgUoIa4/Pz/Rq9nBNv
Ufqe6hGpHryKXSUIk4qbiqRojSeEPonH4Y5/bx94zkLtl/90ottg37HlJLHSy6nAtaVmLFC5ZLaa
p6WB8CkGJcVW4RkjYCN9KyE1eM+OY/5Tu9roKx6PompLafAYAk0CPVJx5t34acuvQ2tlpm+FNezz
SN9haQ288CajRY46a5BMRH0lhxKAlpgnlivZBJL5Qyw+Xuw5C5Wm/hE1z57/QBNfdR8OFvwG8L7n
PeIGEltcY61U7G1BCfjpxc0569h8WEwomZOSnRgSP33BQ7al6GuW5n1++P6VPAK/v7i8mlNgmtYd
FD534X1ljg4JSGk4iHZaE70C045K+2O0V1Wg5u7ePjpseFv2l8ptWj+66/YhZx9n1qM2QRSoBLpO
ekbECg5hKI+tn2odMsONe7QEvrQTE7WHTwn2jg3gUUVGOgHgRdzme4APgRLhmt1SNUU16wvvtjcF
cfOTjMv5B3TWrd2RYkE7TlpAUqUy2RyLE/q8q2tev0Fk7VrZfasUPIG2FDJYQquWH7WfXqtENj1u
hx9hehTZ4o823C+fmwawO70sh74ruHgmZHE+qN2OVQUtJqbG2rVF1h8+tpXy6ETg0y5jkoSr5iJG
tIGnTWYDAFin9U9q9x6wVvFvGzoPcdc9XCLg2dqFv42FzhFbiRJK9NrY3BE7EgRBl3RGW/FV6b7R
ebNM7XRIHRf0vvnXIRL8RThbZJAx/RhgcNVzTW7tK29nrzeo5Vi3fUNZu/Ql7jvmWCul9HMrsQfw
cLeumQXGIRdUnLJDmaMhUSZnjXlPJk1O41ko+d+ZnZCU0otlDrDtf000E8/oNdHdj489X/yNubh3
k8WwiQFD8fVgsVRP/cfK/GTQ2V/q7LKCwtoVAJg/yFdCuD+uZT5NJnCfEJIPrFnvP3AkDA4TcTzo
N0lFHTWCVuzYQDE8suy+5zsYlGa+lx5giecov/pQo/3ew0VzQc9xmScErwbSIVt487D/6VafWROE
29EBLeR2aM1mrx986P6R+JaiVyAIlCwEhl3mltBhHcQAnD+ywilmCrL2fE88xqX3SsXbZYfmd63Y
SNvi3+gRG2/7ZpmCLox9x/n3GxI+d67cwS1FPdrSfVZv4G8ZrJXE5yGrvQotcvVV1DlqZOXj4Nq5
nFfbFhKSVDFLb8p2xy9RizqT/0h9N8W8sSNb116GTJocWwF1cCbaX6AqqDO+ik//gm7pfIeIKBz2
N0bbT2E9tBUEP5qbuDo2U6sjdBYISDrSFKckL7IrJcTLYydzC1FQXgfnzycAS6h7CTWqqiJpCehU
rtPIg+1/EH4gubWYz5j5CiAutwWePIj5BA0CS1T33jQEnHXRWricegdP1FGogOmGtbvBFGRqF4TU
XiOwnkfvJqyyf3V6/tDVCyYvoE4YJKqpYhPFl7tw91CyujI6OP3xbOxRDUgGopNYzLfLYRR0+0qm
aazsQQ0e3zhne6NzSxe4vBvCsMOdnzZbtm4gOObV4vV9iYCZUP+OS8ML5fQzWqkSq1abv3gtep0i
cZ301s5628Yz41u/w74OhIdHJnu7MAeVyj2P7up5vM06C24CMggtL+Mcur2CmjmFuEsa3mbCQUaG
F4bDG2inIcX8pDmvWoHTFjhoOtjde52pQncDY1qqOp1X0jzcoK7vuXLKzvedJUHGv86AJBTKl04B
oXToj/4aLTR9xTT4/JKsurSkd/vEVBx4il6zTTDip0Uc3CuiBG4wRXn4IpT+y8GTZpR7sCJevPgz
IesR2ZE0DjB4D8/aOEQQ3n6gXsAX7i36zoCtWRmAJMN46rPtalgoQBLOIDyajHGSMp4GKUfvF0un
XNzTiNIAGJItVPkSVn/FKQYZkSPsXwkYZI4u911aEZ8qjpp2bzs+XZD78e0fvdlyf9625XA4FQKq
6Qf6u2AaaIGixJd29xl587nE/tw3RyKBoQCxKqYBHlDawyIQf8oD8jfmBhHdhZuX+ltrUPW6aqpc
7SMiNoY7vKpF5YKBTorXWb7bVO6qUbkrCmPpj3xwMAMRuc7x+aRC1HIbDi60CsflrrmIqMcxNe/t
u1L80IBs3GoHrvExC0RKwX9xYHkD9v43RGwLYlFo5lWjWg8sR5bMhPz+Yfghu1gwWPsnmvLzeiJQ
wwhLkxcYKGvgGDi1ksVDeVlqN0kg3jDCVeLtubjKwZmclodl/A6NotWE7eWIEiEgsS8JMR0jnkXz
G/+Os3RMRRpFSs0vIsM4zSrcdUcabxlqOwiA8GPYzUOK876LtZ+vaG1+Ew/+zQMUJC9zhyasu7SV
sKpiXYQz64sUOONKehdVd4oMFM22Ifp8w9DMfSP1QmKV6FyTPBvmB7A69CyVoUVmEAxBg0SoUJIs
9tuzotqRxZSzojASj8nkRUH58rN/fudcl3dGV8z2qr9s1InXAZj/OhcJxh9QEC2hbRr3CDsKPeC0
O8PnfA2EnK2aHibF0e0cQuYIAWvoEN7U7KoNRfw7Op+W/qP5hFNqHZWwdoFMFekRn1VzSXccDuFq
6Whysn0zK4+D5eEMZuOOsqeGO7JIB+iUI0W0t1hwUXI898KSaGLtwZYVUqwrnrAE0YEOwRP/2DiM
yVpAtMpyMFWNevWUCW7D7rW30xmzz3k+zhBIFmkVWI7JKuAhFREwODaj1tghp/sRW9sHDQmnOQgs
7ZSg2aI4bBYNTkMkz8ieH6vtF3jV3xtzl56Ra1rzQL9U4dBzFyYPV8Gpf4tncLZymSM21fer/DAc
PdlL6HweShxgGldKkrs5OfF0OdpSIRSWG4yqI6TIMxeyQhyo7SfwEmDkzXHA9dkFe4F1YllqiCuL
d22pq9oXrroR+xlNamks+D6UCtKrFBjaelLZxofb72hL+9XlUeucNCkApr18kUWj3OcKl2o6uWQj
DCUhsAvgL1K1PDCknqgakcvDOvnU4cqpE8Rp+gAFOjASMnxqqWnNew4WZWQiLpV7CQVB4LYQeOKA
bVeeUh7/E23c4pqjHnzIG4d9irPMxD8IF6lPgQQUgHjmY9RcnPFx5SyAdsz6dVuki5n41LBL7nRd
R/M5Zlmlkb4dRksUAq0kBHXT1CKKK2RQKaXmVQiXgWhEqNx2HfAl/T/t7ERWgLXhTr379FNf4iMn
EAt/LvwuiCtXSSN9D07nPFAYbmXmPoZjtdfMK3xdd0DMS2nMT2YBIv20eA3KnB/kjfNrSLUy6cTG
YtuMOcjrq0JNY14Prp/GYO7SSFPB/ryJgig56N7MBefms4ZG/32B3Yy75zlXsjI15dmCpxeQfq+t
rmaqCYFKji16nSIzj6+8UKfhJXPGriwGa0l3KwptkhBpvg0UCGP5QYD5/bEDBWpeeRwSEuhxsBTt
cnhAmypvXSjbpWtv9rlOtFrLmOvU4TZTmHyF8l6bMKI+gzb/ysQuenCi6HYIU8dPIlwLkKta3hIu
psOo/+QLOVcLVyMcinuaBOULAMoAOUnkl/EhWPFFCb4Yhk14XepakFDwug9msghffWburxeZ2XjX
Eio9fPo11ia42QxPBYJWzExiMxRgBCYw2uKWDXdRjCkNu//kx/v+JRaycGd07/qwiYskVkyFgC9y
UGvivLGfNpDKxCxX2l2FpdUDmLJ20AQTD12krCar8OxOCTQ6obifgL2m1VCeJ8ZoSCPJKAsDIFE8
lm54UeUV381/68zQjjlZoU1qV4/bp3iX2uapuXi4HHRczSigaOr+Ze8k/EbX4n6+fLn0m08IV7kK
umU59UalcKQne349vqEU28c+1N0ckh9B60SVXoJXKVDXAKVFi8Z//NIRL0Td1t0Z1Q8oVUTIuLfm
vlKX3pthHRSGMmtnCDTBwUL7+HLiY6wOn5/3+QoIc9hkWmvtEcF2aiNeeLpedPavDO5ao9fGMjAc
CbmFtJVV2td4pmt6ariVhrGswLoSuB/z2p16Y0weF55yeubQSN8t5iUVplmfl6GwRiva3DvuOSue
kkyqj0soi3U7DmEs9o+lSXTFLSXuruihsSlLTSGugYDg2ZYBWEN/+LAfifa2WLbp6S5C4dKYmagt
i0VOFfdcGXN/fjcG/2HIEzqojvUxr0gUN+8ybWlT1IzK2XTHbGw5M9NHndzy5UqNRf3KsJfNMOdI
j8/AfjcEu9bXq1HJTTwPbI9dOSMCJ+U/tTBRJnhTmGEh7RZroA5DH0G9JJFzOtIaad6IUmCLQSr9
GY/WE0cZol+4sjeTCmEnkxV9af/c51s0qVG6yDWFlFQN0mO09Fy7xOOtBjZNAfKVYscacXJDJMWh
f0KBbl5LTi6tcj69ZfVjjeeykdoWzVJ+R6BbKGzzFTT5ymJ2jhmbV73s/UKZhW8urotqRZEJNyz5
8lW9aEYvwuSUmMb+Bppu/66MtJUAB7/Eyk6NSLHqtpUp5IYz8F2EnLFX8sxNN2vrB10Zb2Wyvxel
G6iCIrJRT2q8cYYhKeMpwvJAwKhMtu+gI6FJtYsN/SkfNENId1vKRkCxDdyDLQlOvTuKRUYntlmL
HnPjhHokGDesAXIyLab4x6y3AfL1Jv6tqRBMbQgmL1PoKsHeyJHPMGEO+O09e3rddlvQ1moGW1lN
87WZJbGhULz0E9GTGLhRc54cQ/N94jUOXoZ2gb7BwX2w+cMjqBmfXJtgB5/SJkSg9I/Wv4q6rkB+
WVtzVrpYCwM03nbxSxtX3lrtA3tjp1pKsqCAXBJxKLG5FzvB5UdYvuheplz2/+ubH17jMpEayhCf
Fb6Iq7BNCnehVYQJ2wOkwLzMcVJ6pdm1IUmnPX1LsDEyGYxdZccwNa6ECwlGGuQvFTwQ5u8VvNq5
tDKM5KIlvrdvuEXKdNuaIvbeB1xruRA9hYNwbLK/ZB+4LBi7IJBFr/LAVgdbzqvTVOs4lEyJKSFq
k7WWEPx7CzMZE449kXKuxKFFjs52U/yKDUQgDCP/T0yJonr3G7vyj8pKaz7bJNT7Sxzb8NVGKs41
xHR86eo9A4AuYPjx63pQCJrJALDWnpNnR/RNc7udihMofbc7Yrrbw7Keyxq41OS5XMMHc2l66Shd
+ICg9P1iErdDi0PglBzX4orh5rHZNRL7ss0/XpibBl8ewGFeZGbjZa7wofwW3MaTpyGPCfVb2qEj
d+tsgJnf5Qc3MRirf7xQXFR1Ut7/ysUnKwwY6cY2j10Qzo37imjKPdGdxkuj4I84Kk72JykbCcK4
uWRaCtebvlWsFQpYbvqEEdCFNPy57K5teweORimgXpPFNbrGc0akT8cPCQLywLH6dWlit7rntIjn
Je3UQ/ZfTmUobBwgEskHTnyvWWqrr9Do2ngWETeBA/7h3JsqfS+XVNzqfUgC/Q/sjlTUS/upx66y
ZohgWLgUby8x856kpY7mbrAdQkcgKAb7yBmM0ROoufhGp9nv8yIU3drSigFDhWuyPfXREiimQsGY
Ih4FY6VP+eP84GWiqslf0mZ4NIB0+ZHjDnyw0k+tLbxH1EGMaQpKOeB6KIQfvTAELvEfhMn+uK2d
lcUgq1OzXIE0hKkyJptX64E9GK029RoDNp5eZmzTcXGeWZbaqjoC+66Z2CdqIr0HWuCflxeD5qpy
lltFNnHTWAb4ap5YMWITmoCG+So42gg38Iqe11Be+NgyoLGnD8YdW2qU3UslPr72kk7VRPE0nVho
69fw/g4g7jtBqdeIsKCzRTZvyYMwL5XCyWU+gndTN/KAMdALRhv9xaR1hPiLGQVEqpsqqoFjNs2Y
PS/pGOxer2GIu7QxRJ6YhZU2Di7TOcJPixcHYuI/Vx7zK0wJi+hDDDjGwNyFkXcJI7+500ukZ1F3
TwUi/FadEMrLrZVX76K0pt60lqvapIGF33pQW/Zn6bQrCatxv8XjjTBYKhuKDALkRx/qlZB1zGOZ
1vUMbWtfY62IEkWtPl5hak9eV+2ZLBJo4igOPqbF1UTG0TL+rgFOlfNGmpf/LNC6iTYcrWOWaXLj
K+IzMc8E0U6ItEiX+ATp4vXJl4Z6rw4QDGI4UD6Dc2+ioa8PV8xgPFqI5Q6WmMOlPp6CQb8ob6kw
dJ7jjAdqYZ2imjwrUlZd9gBfEOHU8yCy9sWwPW3VavbsRp07CuDezEMm3k4NcsamaoFQCpE1GCBO
xHZeq9icw0RwtZUJv6n8a6rQy0ERA/zIcLxmm16U3WZ5teksXwZziwyHO+HJw4t86WY8/h7JmnB6
+FJlnkbmJzOv0ftotRrBeCU/MCpGCGeXXj3shSGXFqL/ult5pLwPGIxksJOQOla1iYpOzxe9qKhG
gayoXxpPN+s4AG/3dxNqeoq1+t0fbjc5+f7dcNSrdLxvsSWRRIp9+jnmCXUAd96dMVp7kkw4f2ti
tBXHtaF2KMhz9K4vKE8QNgwyrgFZEKz5wBnnOKiAsYTF79pOQVHTdouWSPMVBwWTyQtC4qIeC64/
vu3tTUkHB7e8z46hg7Fe45txVi1u04Qxk+ZcEgvnvHJtwklwVRBTpCXkuOZTPIiSkFhWugIGoMTJ
44UW70SaMhd3BpSDOtYcuA2j1trZ+JemIXVpIBh3h/RmOMNzsNvTNcewHNnLeYzxTr3YiVM8cxM1
INYaTM0wk1qCOaiJcYrQSMHXiv/x0rlTZrIsfXFXe4XOSmmflpBZvpPX2xj3v+HB9ooXQl2GcGCW
pIKtnLKweidPqKdi8Vque3LBt3/nakxfQo6hsWemtpw2CpPvhCChklpveI/60ZdCED4ZFjdggq6w
Pi7/6sGt4/oda40N2awj9suksVxWZomDqoSDrTS3H80TzkyHoiMkBvLZWSErInWnZHcXqofRGcX8
h/ItW5AAbXYtBvck0pddx7bgxTof4u35bCggDsCrXKpdEJPTc2Em/GER1cwmK9FlOZcdclu8vUdE
xHrtpL6MRQfW2f6tJgtrBdNe25TJG4HIC+UonCgZPNs/3D+H1uuOtoO2ySNeaTg3rHSUHqkgWFjf
7qh9LGtUTGmk3QO2W8CeiYWFnpfcCIvCAu2NEOQFJT6AEIx8nUTv2SETF7YGtukCe6KbFpAbSbOh
RvOD6uRT0hkDubEjt6Bqbk6BuDpjoZ99VySX9Hj/RBVE6xxZfuzC4hANpCqIU7fH2oseWP2Lffb4
lSy8yg6Opfkc9WeCB8KJ5dY7zg6z7/soBDxYNOf7PAMbOIe22a4mpbjvFd+dcwiMoA/dwEC+EbJT
gAuIdFHlXKUNMx2luhNs4mSXpGgBCt6SVTDNcd6NLfRVs3gsQrl/9EyqNkcVivErOXoRn8rd3Sh7
aSpj3B3GnchyA2PsaOGPueIPP1skoviNzku7kjDB8S/qxCKwJ/CpDhKKEh86tlBy5/3CxlI+8gDB
iWsPE+fPrXvJCVgPBFdwE9X7c56qxTtn8Q65Y98O7KLOtbT15qfg1BBFeus8M70LRY9EU1slKHah
MZvxDEngGF/DTShkAn02TmbsVeqQ/2T3a0argcx00ZJCbvZIW9mywI8v76L0kc8e2zhr7VSQy/o2
lF9rN3TxZuqp1zJarFRPFQVuDEmdzDZ9QoMdhWL17u3CI6iBtDA6o9ix7eL2UG+/wfFWFyVHdh4L
6IviAEPOu7J6Jrex9p6Sgv8+vm8hg1HBw7CRHmnCTJrTexmddQTJzRHeO2cK7OPNw3W98J7/ToZs
pPzIh6k/p7qDzNonEbTb2y28lzDvrfYAGuboyYhMJDUaisu3MsIj/8Z+oovQVLHfOGRlbBToBi4y
fVMjzUcsLqJ2xl20faHdtIjHacCm9DlgwdADDouxhEH2MmCpQth9l/JhnZ6CoyZoWPHIy6WZRUXO
WbiTv1VAa0ivQM0J8sJTTaRWTCmvGAr3w/Poc16gcyPnTK0JcqSgILwlOaSFG1mL1KxabmEWgn99
ZyBrpBzIjGdfHqdesmSH/PjzA/OBQDaPolRk6tlyd8zrPQ5FzbS3QRC0leyqIKUjdYyCi9P9npTl
XdeDbtdkoK+iORVo9F6Gxp52jRNlxaN4jVjWwS663qHBK5tBLggqVMc4l8U/OCswaVeA0KpVVCGG
XpoJSHXrQs+vmrYuWl2i36xFmoPcszkZ8LWAhnnB5VE07J/LBTTJujYr+95zrm4MVlySYxCuxcBo
7vTmRBahopUoP5TDk5CHJU8XJ6PYwZc8w9qEBSJvdAvTH37JeWVDAQSXAQJDVNJoD/4tr4Q1g8fn
NXjrMRdOtHHnaem+JRQbUlt4qXzpVf0IAI/mAuVWio6EsmZiaorwcMdfeNQXQGHTsFgZq5t4RRb5
uWq/wPjCKXRJr6Uf0tA5hUmS9bxsIOVJ35DQ0o0VBZGA+Eyg5X+xFkVabIO0Zp2ZJ4lIyn5Pa/5t
afeXQtqhAKe3vP9c3lOtofOyuNiYUBa4bz2fbGIKsupJaX9b1gtNP6lyKDbGCClBKT5/3SQf9qSZ
VM3xj3u16iVck7hwGZa4mfv0TIZAny+pgpMLTUIlBcaWyrwGasIcgnt0vRO70yUd1Y06CiGqeLjJ
GEKg5fqLldJhbtvW7+1PNTJdUQCQD1SJtPWxI9FAdXO6y0YyGd0xrO8FBTbG0DcfbgW0r7Q+M59E
+2LzvszXoi4+JJMKkdtZkHtmXhWJYQZWACtOv2mM3HNM93f7RFAsQO5C8ncXcNkCEk2P5DNDcmIT
PbfPWNhMnFuO4XkdNSmFF8iWDV92WEdbb3yFv1YEyvl5pTRLVzTsn4awe64hgdGWiDiIsTnoNegA
zDqP8ZjNV9KXhbqefGwp7Y0ZKcS5Th8BVaIYW0OuAGWVZdfJiBufL9bmLF9QE1tpOU+IXIZziIhJ
F1I7x3bAvJz5IsGKOJqZylYOOPo06a5MVed96hPawhKa1lnJTSVTN7mHT6G0q4/a8W1BADj+ZYpJ
kUbPY4NvTDiKLddITY2EDjvq1uolTiE7Z7/U9ekdWba2mpdxMkyF2IObkBOcYr1+JvH6Q9b7fI/u
l54xx7vyUBOj89afwXajXGO5aJUyvmYyMVk+PmD0FIkWcvGn9Jg4E4u2inEBnV0uQkXSABPUD6Fd
YfSJ7kalrdi9yZFDG4Wcv2y4UBvXnyQIuCWuCA12FTRq4ezv4HVzZEQBcLYk6BhECtagJn4lxhya
CGHTZmEU7AymWRPB7V8YMkC2y/GurWrnovIZwjquYEwjDayncVHJr8y+H2EbsJxiqAY3U0Wjxz2U
n6c+4y/iW7a6R8Tt3MCD0/+h0kfCHjCHpAC1bqgiFoeNn4hkUBZuuaJ9hKhxqiuj2xU2I5iunWSE
ktJ/gBxzydPRb/NzBDpkoC3cZFEjLNGwhKv+TujnBW7rLPXKnhroHSe2WcmZmmuAO4W3FNR+/ZGM
R7marmM+ajC/FLNW0U6iuSk6ggwetuTjmEe/AMPeaF56tGwAfFDnEnBOPvgSMoCZhSa3pHU5z1NQ
DW4/hdSiwSIp2+ekKrg4IMLoKIXE5gXD2mdVnSI/50/z0X6ALbbRZwg6yRo3nctxi90c/DnKmHkc
hX4VoVNTGXQgxa1mH4J835DTDcWdWfBrSs7D2iZWR0UDBZsURT3SHDNK5r8HVcZHBlRgpEjGln1M
DOwrqvEX2ZmtJ8CoWYq6wDYwxdFjnxz+yxKm9HpvoVv1G6+pRIq+HB4wQU8b4vwWUUZwPbT7bNCt
pHVIePTYF/tYW8Cpn4nrqzcbCU9IszGC+mtAOXzcej6ufNYWIC11Lw6SDx6lNmsYm5BdkFm9o7dC
0DIjeezVPN9/DEfGD2v5mpJP6qV7DsTI5P+cD3ul6UN3PG4qFP6xR80jm7eBuwPJWfNFhYhlFrhE
JylfRlKk8hRwgtIBJIZokt0m91un9e5hOOVxj3XQBylbILrsYZewRCZCRdBZT/TCg3J7NFdYfmrL
mu8vXp1S8gZWoT8N9hk0gKkcvXNoNmEsZylczZjv67bN1DaBbbGqjjLGbnrQ3cltr1MgVNQvIG6O
aLDqBbt4bFR7Nw1WyGUCMragvL+6KKHANzNbzU2DjeY6TD0ZIm+yV6Fw257lN18XShHRe5zwh8Uk
1MZ/H7evJouYAoEPoEHriDoS2f6LORBx7IbWWyApJol86nyfXi3x4mRKTxACShLFaasoWibky98e
LeMdoly6t6VBasvpPD05Rcj3GEnT/XbQpC2LgdsQpr4OTYBtOVc/TSdcQe17lGTP+fG5kip3Je/A
HFjmTGwNwUuY+qvhI5pnqCcJ/pQyb/1/6+mp/y7klvYMvQ620SuYCTWqOTUp5UjQPgcyW/lvj++g
IY8skOlYRNHZ+4gMpNW3lH6IxcyV+lbRp4zKnU/WnfYak14ezNy6WTP14LqJiRo/Nbs/BYvYDhaQ
7zOfv25XaIPl3nC5oLmHgVzJrDTUt2B1U5EJXg7CiBWL97dNDYAEnHkhBszSJcKhljZqChimqczc
HNpQTuaalXh1Lext/0Klc0OPK48eoS8ecN7LtksLLKoQOVF6WJKZ7luCF7PrRSVq5ilhaJEHBqz4
Y/LdxBi5VVZOaNtMHdicsnI7xSudi/Ub+oH2+vKmmju7RGXf1HH/CgtmstGUyHNTBSaXZqyDP+MS
iXZa17CaR5xx6IWOx26P6jVTIsi2MdaBtdcKx2OyZOjwKVJjgP0HracQsjK9oKSOEqeTEA2nzOcG
dXdtq22nsQJhxUOhpaQANnJn/F00kJRZ6Rj+6WA8BPdpoBD3I8QURFrv8htq0MlGRi1ejIJvdRpI
y+yQBEbZa7cSuPtLAZoI4S/ADyU4PP6MCFiwQQ/G89VhZp2JmIxZbPDW/CXx1bv+EM5r3jDItVbp
H6mUYYDJoOmMgIXFiMLqRYGB6rR1RXumzYTlFWcu4AweDlS0fGgXlNXhc6oUNT+lz7f9trMZPe1O
+/za5gPqd0aJNLlML3adE3lzbcJkGFkEBeWa25KsqNDD0zcS2hWGS8pH4OFo5zpwh91bHpQh/WbE
eMis/ebIFbu/mOFpQXUo/y9aZj7owjWcS3i3SolrSzJi2IeeW+Fi5tRPGgSqt1vbjVYEAD968kd4
Yn7UE+Lx3OP18Xn0QeEA8yRBXVeBRchWbPxsug6x4XIKv3zQpeqasFLPq71mtOw+OnWyGY6EKvww
wuitjK0z3zdffVawWybfHA34Aftr5AzX/uqeQXGV3VyhKPQ2OudH7jyipMMv6+RWaL+wKc+O7Yof
FvriCg1Gau3OazGKz+wZ25wH+rFAvT5akYATlLop2xcSlDCu+s8wXvK7YZFq52fpi5yksBmCC+Ma
QhdMndMpcA93X96C7ldRIcdzCeNYrtI3uPrT7l2ByXDA0S5JwtM0J2RXTOdzC7mkUBzvGBjzyc8C
DymX2miS9lQkFz0kZCauoMZYL/AsQUEcdt1J3dJ+gn4pcJNNXP+dmX4H0Ds0YBjIdX3/uK+6ojMu
E2Z6QOcKLMDmvayjODVSNLtFiR+GM7d2O/odoOSm0iu2k+NLCH6DKP+fHfpa7Vik2GCOO6GHwp5j
UQE6eJw87t6rTCFzDOZjA6C6UUMs7Ie3OtNZS8vRpsRjyDntzhsxYHs8l3hh4Cupx5k7w65lKcxa
68pHarydBvAaaUe8iRY5eyXcYz7zFEGw+ou1ZVU/m+1yFWP9SR7QyN8Vci29yxrWkGw4M5qbetsO
WWz/TatqADgFbsdMDRepesgteJjzca3CSTIH84OcwqhPF1grPxnnbV5ad5gWvbYYAUWi8hur2PLM
JY4NSSOeakwbQpdjpuHmeJt4pf9TDpxJRCHgCQd/eaVQJopIo18ol0OYUm5Igw97iVeqpWi99Efk
8u7Mn614n1GB9mYf4Duirr+WFe2YQyy9ehCAlHqE/NwpEo6SROGvXgovSrEjxQCNf9H/9SlMW7I1
hK+Ul9FqehtsATralwsLJSsVKRCh9p5RAFhDvR7i/efLR/ywZj7z78SDkMv/G/hST3ygentZtEon
wBORR2Gwr8nFeMeM+9edyhA9UM9WjpNYta4K4lkV0C2o69uEtOAozbrvyyk4suO3hdkgLeSVao+6
QXcUn4+oW34uCbVEprA1PByekDzZbIpujSpQYIftXRSt1I6tAk5P/BS37US0u0rOdXZH7hVZp4IJ
zh12Icxx5tcNVIuV6t5tCBivS4hqzG9G/8nTJQo17tLxKI/WhrUbz1eFXZ9WXZmEMJbVcsfU3LlA
lrBghnszDEO9vYrjdED5LbasaiYkFIOmKyk0OcwplcXPw9GV2p6TwLvH9lN3NXnOQfN557j7yKGe
AwOEgbOtdaqeRgRE6mmOUJe4oc7g4dWYbmfhVHBVAJLXRndUKXCems2jA6k0GhNEyfFJsz6W/zHi
5NgrJU0Zuh6SaVMuux6QBKE+YNfn2Uq1np3pPMu29BEVQwksromGLi9u4/Ag7v1zrH85IuorNndj
sW+SRR3kn6pLD2q5lp9vAjZUPHe6GhTimH7yEZqu+zP136MJqK+W1twVfj3EmMLDjKrap5CkEbhO
q4i+peq51LSgFD/eT/YZKp+mNZBiq5YJtOmhPv9km7S/QbgnRLV2YzTFBtguvgICgG276qWGZYqE
Lk/K5VUz55JmWuZgpHRYockc2brBTZWbwnOEjq40LaXIMbqbjfrhc0La2HKX11zKSxP5QzXfeHxd
mPkx1ltSBYJQM1WpWo25omgDDlTDgrFvtVM53AGr80ujV88NoGgb7ROx8wLKw4zgC7GkX2TG6KxC
gdmXe5oE+eZbU/M31EDcIDzYVg3eHqSAUyUMj52UlhbY9y02aJXSynVbOmv37nbOHnkIn5e2YpgZ
K7k9qF4OrZ+v8OIbm2OqSfEpWsNTVmQs1fLRQugFVuBkHwXk9cKs16zi9iDqSOD+3quPYmPkCGID
nn0ehzygyk0/eeUfO5jYrkkAPtyiDHagRWxhIQsjitRSETVft5kBU4zdnVpScqKYySGA0kIhMUAo
oKAnWlDYL3yfHqjUwj03PnRya2dcbpCYhN8ImNf3479NKUf5Q0GeyweFmAwkLs4ZUOPcOTZu1K93
pIjdhfh76oES9yjTbzGxEvi5D2CgRlWomBhNv1XpcuOMg6IZqO1YX/pixFdzv6P9vABPpw/AliTp
uJUfGLVHOAQAbK3KA1eLVDCq4B7FVRs4EOlAgo/dHXpuIeaTFFcN/tdFlUK1ntljDZHnvpmtgsnW
tw1fjdsz8v7T9IB3M0sgeeFdpivoHFl/JFUe+EMi+pwRA78wZxiRbSFvBQYDYut3OHIZvPAdso0H
uAw8KXWFZ7sO8xBnBlrSLZ+Ef/xr3UAMkhhCqGHzeae8M6wuo1tbn5Ja3tw8ZSyiDjhFObIBL/ta
P5bLD5mKsdzc8l6rQdGMRzwmJn95Qdtap07zmfpoH0wEmSbpRToZ44OVFVk6aksSNAkprHUESSvr
wFFLGBlR1PN3aEzK74AeSFxE8LRR3LUXpsspkftSKyysmhgBDkOqHPssBHd04z4yUazIcHsoj1w/
JFzPCD/lKHpd2ejOh1LvAZQ5FAMCncaMUQWldbKpfuz9Q/yBx2xNYIKiIxYoG5DYTT3l4sL8C/Y3
XWvmbhbl6r21Qy5ulsu935nFjnVBIJditL7iuA+QcD253ziiu1EWZH+Ybp5T2Ta2HEWjUHpdnLBb
2bLqSdhlEe8UFfquaLv8Rg6RjdV8Bpjo1TFEtVIoebZu8yAr+BfJMDj8zX13Tl+y7DygD6p9PTdv
riBZToMWxa9vfM+gkOc1rgKzVDP29q+ov95GP8BbODnV4dsD+nh3x647tYmSQlliCcy+o4N9SPek
UEIluGt2NkWUTuQh2blwH6YQ5lLG2sae2j5xpgS+e82y47X/1yzPhCJLn3VhUmer5h7AEeJoOKek
k+GH3w0whpKI4DfhLrxt2OS2Z3SxEcJEF9wNIL4RGmfhCQIYxZVSfkXFZqLXSj9YLBYMu/SzRQI/
e3bW6DLLaKwXA1HNnTuHnJeiVsRlTmfcPRSAHFpYVqOUb0jW1WMbj8siVTvZHXi7J8nfEjtI4muM
xF6yjxj1AP938/5idulT/5+9yt1o2ofTPVwyixciSi2p0kxLHc2X/QIkYexWJU8T15n2Z1M9LmS9
cKcW4MNd2jK651H6pic1YSypKP/KMaiHIBvtjRceiocfIuwhHcIS0TRdVFreC7+XG0eIgoXO9468
SoRTRix5hwVcAdZkyWSob187UfjT0NXq4NS3uZ69CPdudeFN8xWPTBfMkyGoNu2oc4gFP+WNyl8F
C49n0BSWLh0sL8NVDSDDlxZ1oBvP/M4aWCFCExwc67USC4oz/N1sFOEnc6RF4pf1rN6od7zbqPXD
TmyL2fk5NW2ggpQIxcQi0Jb7EWWp9YuFJs0LBVURwzTnfhzE+/R9a+R7KNnkWU6JQ/ARjwWsbWwR
1/znQbkjVnes3ykl4mlY07I00q945wuHbhgXuWRTEpiP/+tA91Wz1q6OiBtA7S0ImRkanp1DPwAo
6zBW3BCfF/N5pYDFw/wLB2uV3ifGxhBdDiDrdPZ+6KNpx2jdfN7MdrypplfcD5uuhO+FboC/hDtH
WR2RyQGe3UtZ9bNFX4WRh/IUPk16NtQ6aYMXZfcIo1Qf33srcfWaJyyblM9QbXJUAV6nU4heAVTV
4JiCYDG2CBCBGnH9aCp1aj4Gq9ehmkgD7fryFPz1ZyFUWAX1TaH3CnbXzJDiYfw9XcGbfEqy/F0u
MpvwncctxW7UklRaffxPZCc3A1wsQCLIau4gbVLLfPCqCEgWiPV3AVRYev5LG7w9m4plNwdP0ss6
ibnMrSOprZNluQVwgnPJBXm2CYLgDfe2H1eEQYv8HGtxnCTDN2R5ip/jMlqBAtE9Lid/+U9suJXB
Qyp+zr5Q+/Ue5bFOZECEU7rRR/+ut4VjEvY+OhYixHUfNMXLibkhuT5aIunrIL0sSQXnAstb9tBm
XqFlEK5NnDjNcMx/Gzo2MYOm2ieKwj5HihPqcIIPnSIkGK5D62u7EGNpaXzDf3nBbjDt0h6apMwK
o5nDZNSn6F2aE2I1YwZPoEio6GKalZxsESLgDcfO05ZljqwHf6DHMVl5LJ0aBs2FFuDEQ0spM0kB
ZFyC+nyswU9M2Kq/w+V8sIYlo70B/vIbirl70gcrTmQSCSauBbW9UshEqjBtP5xeGpQ3SThonzeP
wwpy5PwFvLO5wzOW0J18wHkaeLtzcyPhJdVwfhAFDxXDZy0iUA6JMZrWGRxkOHpEgV0FrjlI6rTD
iBV/PvLLKF5ZuNdKIwELYQwu4q19suiORPWgRG3Vm1BZoM6aOGQNWfRgi0HoXTzSfT6dfT7fwMzK
xbEbYL5hv5PGkht9p/XRXVfUUraZnOOcq/j7f2brrQoWVIFyCOsDRKJLHvESBctWKuBKhmSgMs88
3ez6jLw/3U+DHrTTrSzbP1NEJVLQwsHbphb2d2O6NvlQS0sEu3OjsAa5kz3H/QrMTKF+1WApKZ/h
RGCBoIYTb0zZAteMgNV+QkEFL+xglxL7CK0WRuO93vT7oGZNjpO4OKfvT4J4HVBokKjEddfTufhO
JVxcjHgnJLUGcQzZK6m8sifVHKjjgOts3B8UGwSqOjoMECineQcxPka5iHQ4k0FBIT8YOJVkWmsf
YjQ3+DQbAWeHQncZw/i/tQqf4W9zW2cu5+JfVoaTsQsRCHwi79eUIx+lBQZSN33KIFg5OISyaGmt
zgt7CMlstRQvoRXRfUT/rwSyyOcGXsClpbRFK04IaDTzS4DxE0OP2fr7XpbQq/cixrlzd9nO0Y59
n/q9hVQ++CiIuhIpfp0/9c7DZii2LPNmw+UQnidTp19U/+CjY0fN3Cu52JL4JW4e8u7RZwGpithz
4XCFuQrtK43imcrysVgLBPhQnYP70Vs04Je9StH07ryMOFAMQQfosRYCkVFEuo1PpWGa+wM/5ict
dzrv11zKM+hxWlr5cIPjLRs8SDelFW6lgzQaXPcNcDM7jWNadPYNaetCjgrEhkcBrusUQK9B3GNq
EytGNV3ofvYpg181jj0ZdpKAwfjoB+ZVyBD7yCWSTR+6AxrFMCy6BpVgAzdzf9Rr2m0jvkPFwka1
cOujob51VWD7H+z12AWRaDWrgygtCBTlAmbdG/uDL7YJ4lqkpsQ5GkGFMatKXloV257D2lKqz0Kd
xtk60M5OYkw5cL2DalyLMKKYVcOaXRJnAkbCULD1XfEDlLElusTGFHYyTyyoH7CjeUWjTzyB2N3N
hoDC+1szAuVPsV5JVnY8QjZwkB4TAva3duqHPBCG60VEriMKOTCn4cqy+RPkOP9KZ1nQMUSYNK/t
9EMi8OIqfC+rmgOnxAIcuNZ9fr8gRkPxmDwHBKtgQHp2OAWNVqGF6RnIJMbNHy3ex7qFEEF+DQcb
lfPzI1GDDT+3t9uods7j6grihGriClgUQJUu0mPRmMHwy4Nbqn5s+FWWGpx3SxDCj9hjLXFcTthD
sXDQV0c0vQsDNGTpgWuS7aYHkf13011BjdS9L0VabDnvuLy2DXN4IxpYcaIsYrq6Cksk4jOxLoih
Sgx0xkXMqifFiJDXXwzrEQqDG3bz6YDv86x966RVyo0IxCZcmJ8sU7MXBqOKJj+B7aroEpFUzQ4r
JtLUZwqQamAXFX1XzPjtENo1jKqoCqVYS1Q1+ycIhcCW2VCBI3xzrG2bjTDu8p2ac87apUtbCR5j
SKxLBKHuBgHuje58OxEOn7Ukr7uuW8Pg3ZnatTP48XH9Xzdf5FAVYkFlswF2CF9e0tKK1Zm1THbp
n4T4EZKr6P3o1RDnFm/toVAqy8h79VcuJZESiJZKe4cIbuTUChII1v4+ilwrUeqmfcKdsp8fMjGJ
CwLq5bbitKIPSXiMJvFb+hAtLJBuPXvyZ5S5zS1lUk8xVlUPpyjZuH7Z3gSxxGK6caFJ9koQvBhI
oLStVC5JJvuw5R0ZHEhDxC+x9VGUGvfRvV6tH2QMz0RTlCQH0cfv7yYrZhLmcqQ90BYfMA1BNoLX
5f4N8MRSO6hHZo/SmjEWXlRk4lwsEHHTO3rc+uGfqDJIc1mhBLD4zUN2DYjRxpCwU5QWfAiWS5CV
l0dsl+psa5QbXduh5IdeayEVZARrbrc//3YUoeFK7zk0B2j88m0h3s70Yh64VaycXa50rEoeb9g4
NS1nEUwZvxGOhw38HEBuKBMNew3cGgryZAeHTRXvdrghAjfzzN0HXjcIsFOPkjlqgT2er8iykMnO
DZT5YSRKvep5B0kPT7jwj4N0UHLH9IiBaqCbI9/GY84YJV9uEUIyWx/C81ncYWHIl4SVYB+TB8Zm
Q6WLaHtu2B4quq3gwrL701VARe3Bhnypm/vqUzunfhJvi4raplxmYz3osHy5dfCNCPAlmEFbT36o
yF3AMUn1VZk/rENqdkcKNxmlUyUhF06WoJtr/5RZRQUyATQoyJSjav7l7fMeEG6aCBInVKbRHte+
gSMCHyXcS6IoaNyg1WibMxsBwTp9tOJmhAZdQorXhCampHZISx1lFp5sPl193DiACzVqGUkDhJtQ
CBdU2Me3WZNNRrGYHgmbXdXLxdzx0RvSeySNXG0d0exgl4gwUurA0I83EpDmWTPXDh6OIyxEzKpj
JRsgPZEoF/1BDnTfjlfxOUUuVGG9DxA/EvlMcqyOso3BunIv2+fl+4bYnPNeBrspZnO3EWqJX34p
4PltsMsuWAuNxBDHzboHhkzsqzwwL+hfqLN0NlQjuKSuMVwiPfwiuU18R9Gjbv7j54iZ36EyNuU+
b38T4vDbACvk8vqWf+Uy2amfAVgikUcrXosR8ii2CopGhASbTeNdIx4XHIAo+2M1U0+w6YPQhjPn
Catn0DEPxE+3pQVHKDZmdzC7scLUWw==
`protect end_protected
