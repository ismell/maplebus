`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KiGptJTgfqBYZS72wh69LJC9ftH0usQfbwCqWpq6rKTKyZSFHTqV9jYUREWmB723cGIc30akrb7R
rwk5hSsJOQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oDh97TlkJefnKqv55omMQ/ZmMIg5SM6QuYpKgFYNODgbGF/5rc6rWbGwOe1hjIKPsO4/NT2klxXD
dt/hQZgrEafpc7fubpzvKuNtQF+0ilkrCJk7x82TwqQqlkD6KjaK+gGEmn3f6bTnG2oJhMHvCq4N
oHgqcLMkAtVCbl7CV20=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UfZCiEyJnA/VEE1lagPKMLZO1eFTrp5Fl/4XJFOl/8RBa04oZceVStDRlIUZIPo+k64+DsBVE/Is
RDsD2clfc3tIUHljYua9C+fiefafd0S7sxl/KDIf/ckKq6+B9ZMhQn6IVYshE4nKILXVv5gMy8Ve
CWff7IRU8Em7/9UL0d1dfiXZ3Y8j82CjbhGHczhsjD6GJZ15wF8PKEpjOkb1P350SW3C0e9smHby
E7vXpaztRvdAJmoQpW1om8fK3yzc9y0v5IXkAmckmHIquyrKkUWmpXsVFiFKHz7Bo8l/MA7tUTme
WcxrSiFOlHJJJWKv1Zi+21XopBRiPWUYLfHCeA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t7et/RrkK1Y6zv5kUSWgI+KUOfrQNKE1oxsTklop5j7rCvYvz/esR+1xd+zy2pURy+aItRfHFC12
1QexHPPIuxafV4o3ncaEzKeqXaXEcZ9fFhn12dGGYqDJIH3UU5oieiew7kPUloN9++bvo2pOWzBh
Qh1U8PoY9vRvl9BvsOA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YfY3lGfEL2wTVsCSvOs4aQEMyq5AjKxYTAmPhnUtuSw9Zfza9lSS4dUKme1tZMjup4f/4ZHcEEFf
5BDmD7MEClBNe5kobK4ccmcyDi4tOv9gXn5aulmst1MbI1xTX6AkMmg0FdCkxaA8sUIzO41p26SA
yiSDKgkccfxANLylEkrbFCz/kh87DkijKjEtWxZNYg/Uk744fJW+ABuy6iGIDL8oNdeM+Kun4ZvX
9CyHlgKbXc1IJXR/MfFXKhd+HXxrq6dA/mBxFLgexORkHopz6C0YN0o4VwiQPS3pMM62qYD/MAFi
TfU/KLPX2Tq6yP6vaF/wWpHUYnbmBrt+IxsBpw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39040)
`protect data_block
PLwkw0PPpG8za61yFvf7uHCEIsn5JyR5eXWeh8UmEpQ90SjHbQCCdxbMxVFPgRsX6dzUvY/bwUKX
73cgWIL5Nx5Bd6NLtOMmM5+HVk46iRKt6Qh2zCiDKqA1rnT+TPHP+yBHVsCmLATtxB5i1eJGidg7
Zaj3TvQz8uF0Kmr4KP4eQbBCs8UInm3ZmhMiZHW/plAVheJUGzvIBcgNzNN/b69mtzKJUU0M1LxQ
QgE1JW/Z7pEOZnqko4NvGqGdES4QRjoGHVhsBMlwWGKLzAbcgT0iWxfmVdZ7pd1gCEMtwCHT8NDM
ijkbueYX79BLUtbmLxKYwpAkeNcjTkijtr7QL3j9y9e9Rzq1CBRvQSErNz2xKDqgdcs3KWwn5NGp
CwpJglDH7bGxMD6fhywtoakENUpoe3WScMiPBa1Wd5jd5MXNCfDpVNAWZjMY6Ftj+1ootv2EkYYM
mnOpB7vr3bg54MU2nrz7uumZ43gvBDabYzXtR3SuvGv4s0gBcKCxIa0s4ifzw9s8QEsmoIfy+5rU
YvN7RNfrctwwn+PXl/zCqae0ZJhEnPTg5gAwCVf4+o3yYgUYfMR+m1Msz6uDxSSTkVRQmGV6do/V
cwldBXBF6u7RSHOkjVeIXJ9Md+GQpKP7Z5Cdy/efxUHAhBstIwfoTWw3JDhxyt2w0ZeVPQ2yguJ5
glmuPI2k7d8WmmfSHuHsOX2kC5y5ndWVQ4Wu7UoEajkp+lIK5njj2KDYMi/EWnY1Hd010539yxH4
0rERIqxhfQ12U3Eq4RUDyjDDjlJFQg+4UJYBCBWD5v2ZhcNO1O7FWFpCrKhw+4KhEhc1K7pb8p6s
8AjG0ATd1NAKkh090Xrui4AyJ10BUUDqF3y7lf1am6Ixq1aKgC9VcS3eeOhLCS93YtpsBp93IXQF
OgQR52rGHHv0hZivGASHdYpc4Ocu1yfOjDT1AIgqB7LZpdsEFwr4QlawyUsRQqqZH66me2LGfXlo
Ba2uxMzTJRxXFy1VkdikTk+u96SErOq5Rd1+u91bP2C0hp8xNnNkDaPZda1X1Bup1pdF08GdbJRc
iPucJgQDJ9xGPH2SXP8eD7v7xaYwlqZoekIdwgqdRI9EZ7bLxg2XCsOFn5YPGFmfL9rIMxesIGx9
buOfhOaTuhJdFT4ACfg12yZrn8YQGoaEQWxCrjfmqUSnQ/KCupl3jwFPEam1RrE4zwWeamVXoXi4
Wl/kGSa4usLDQL4vApePOw9urRL9VgLWs9sspqMp5psaKF2+G6+DyjsChPCgqjYy8CF6FjnV/Ycy
ROvdJE7Eo1z5h3uhEUPAFdtYYjBH07bzFBi/Mji00EMyYmtlpEIEVq+zSVBlTWVzB9XeBm+THaM1
o7mSZn4/dHZdRSy/34aQ7fj47GkELaf7fIEyp2vC8Ada+CiZcrE3pLEOSc71+B4xtXlk4h6yui9v
muYL6OTWHD/glgvcIgrqyxID63EPAc2rSsWU5oyRxXa+fOO1Au+yB406wPKo89z8bSkSPV5V0yIr
YM8JBPjmd696R+KI4rkl23gpy7kcVhVIax4HpP63vhErlnEXU+Ab/lt/omlnmfIltuPpMiGSWvjI
yrb8Z+DpSycYr+H7GBzVEmhrhTIrEl3yVDX4DHpbe12f30m9jF+c7V04y1KhuXY8YHMrBZs2G6sM
7kegM3eD3TzgftI7e1btQ9WfmQh4D36LIPMzcC9+j1tsBVwZctzCNBdHVsvBA3xJR+hdtko2kaYP
AL9wS+wNb56YAwNcIPMpewg0wQt41qnVpYxXJ6sjnCTJe2eOqseRAl5D+kG1UqXnr2GnzxQT2l39
iVr0zQCBUmiaVC6yIK77tdn9Ltwv6mYpi0tzts69Tif9X0AU9jEM66OD40LENgP8pTMLi4Xx58Tq
KiTGq0ABmWdBPfPZiJI8X4rDsrHv1b1imgIaUp8V2tJhmRabWMj7iVLlF085m8Hi+qk2LS9fkcGM
A6PKk5ui9QsXc5tZl5VJ2UGWy2uNO6e3pXxGH1f66fpz8MftNnssvStMNV/4qovaDbtacxoTohZR
ZfbDXsxReD1kDHgDuD88DaYzYQPGRY2uSnXP2qkq26ebKB4Oj4lJradT1s3EFL7AEURhzTay18lh
1a2Y4a8B9oRaJ+FeKE0zTHhFk6tdtdgOSRoT1RMho/s5nDmvWeRDS3bVXfK3tsuWXkKg8ftfauwW
HpFfWxgzV9WNsLfRS3qCFqdL4kbBTuWc9NEfUEP7o7nn16tojOBHwxV+GD4v7R+YDQvzu+TLBoK1
96xoREB2AtOruyMk3wqBjsYhq7nnXZbmZZHwA0qCyha9dB80woHzy2U1L10ynUE/Xz7FCYmlsV6G
CGLx/nQ9PrKCVeB0xyFt+epVXlKmi7Kwi4ookGZrWeoVkkvLPfrY2P3Y/sfeTeFq8E4AaBo+O8HB
+npQWD5/66JMtEvyiJuZb6kRCb2t5yfReQMf8GzHqei+q15wEDPEg2kBOeQlnUMj5yJ8FTu4tBgs
zlqzsunzjeKpjPPN6s5bqiY8LrlUEdUPpswBpXIqW7iKdTtCNnR5ZzrPafziMOT4+nM6MTE10w0q
/pPIpnZYNZZtDD/+sjWFRvWxvz7WYTk0ghcf/7vnjLXtvGNvr1f4LOMXOE2aXZYajcWA9gKyKLPY
+otHCR5Q2EbTT32dWCfUr5EA29kp8Q7Zh2WwETEyGnKI0YT532BNF3eWQAPFoXsCPEvOdiZ1ZdfW
5Tj5SyP4FPens7Z3giy4tE5C9d0CPsiv9K2pP9gDV3nOBo7m0mxArLz+r7/cY2w5BGlm/DBr4uP/
ydG+5ca50DDxsDZ8bFc4DhNkFiBlu0dEg52mmDZ4mKs461VJ5wEbOnLMQDPH/2Ar3z5FH0m3aXVf
tLQqlzvdPMFMXCh6TZKu5xN9vJxECKk9jpAeFwJ3IFRWPuOqspDafJjWCqjGxmeZqwDNka9vxo/F
ktYEeWBolZvkzSmnuivketkXdYC4KphXaMrlZsTZREIiI6S1LTYiVu+TFnYhnHRLjTWTf5Id8Lwj
6FNIu9KgUYMcBQOnhghNLsU9Tuyq8/AvgP6dbc29cZjffK/3muLG8cFRHqjNnkH0RyIUpGwecsiN
zxNY4qnzRkBwYK5aRvCL0iXBaiOVRsDdq0kOXsNNGZpVSp1yyJbz+Lo4EB9+2tcufooa2Sul+QlD
jMJmc4Ecm/FKGvXaBbIv3jSN2Izyd1PTt3zMTnaHgGnYsIt9JWUXBG+PT24zApPRysbjWcfcHQt+
hKoclalHPb11xQi6THMFIM5ix4YNJNWQIb5uO9Vc3JAOgAe2Mqw2XlUlEV9h3eKO8FuOoeix3fmY
8k3ZzKIyldAd7IWTSt+lojS2snVXEDRtcJ11FpzCS3TQuAqn4xOihfd6PbSAMd1qwA6ruG/MwxVq
ieRZBOKCp07yYUcRMSA1KMqalbQIOb3rz7lVclBBSm+T0aMgTw/9Cij/haBRtCjhOjIe8adm9iRI
IS58SPEXD7HcFoL8QLa1pIPDoX2vY4rB0JKuZfyo6kZHsNhUc0x1uy0dvQdy1GD3res+xOoLULSE
xjQXa+ggSP3xoIvapAYZC+UG6G7mO3ujuGXv3KbBQl2qo6lXklFcmwnATw1z9VyhTkNGnknCA43K
grzHNGDet8h4SQDcknEKe3u4lJbpepeQTqe7/Ho372wvvxYus8NHcRqi1TTOQDqMBYfYKJkSn9XN
OV/cG12KOqo3W6j5yCp3Jp8WdUUgOvX6kQBbFOQMqx4/jaYsC4KTF1Z9XFFWMCLiuw8s8YUWl4VA
U1XgeNjHC6lsBbUO2kYx/C46ndWH4Xm1e4iTsEXRSXpFgYbtpS0/eNPgKytm64M8rLLIH0NUYxAa
n6cJRwLM3hTprT6MYXMH4QC2aDUv3zKQIZ7F3FRHJEu1vvzVyEyBramVNqkBzlfLy+uCZLKGopNB
mqw4/0Pru9pQWDZR6H+ut1ZG+Cf2W+Rdqb/t/YRflI0ZiZy38m3C5O5ceHRO66lLtyW/er5OJ9Wx
JQKJiWvTWlIkljws72x7/T1as08g7GYZxj10Y85SnE4KjL0BjUoWSSLdcz9/ueEIO0zduhzV57ks
2CP7szD/0AZD2RuM/emQNG6kZSAkyyoh3njLm7M2Oql4u8gag4dl0Ny8Syst7h9i9wRej4+hvakg
MoMg8jqRR5hiD+H6EHvCmgAfaA1Ieu2I/L6cB14AGjpABG0qQS44SLXbw1uDRimbF+EtmFZEC/Qo
l9QALRbVOi6pg9ap1Os0gxY6Nb8ODJbQpdPEp1vqYlinHRUpE4pweJ+asEgIekKONI34sJQdw11z
ILaW61DSwgibeemf6L8nF3DAzfCbx6p+Mx0Dn/obw2X+PBAcnesZSjCPVDWi1GxjJqDn9MeMyx3Q
YnzrRUirNNHDNOD27eA19ehuBPiPgE2B4iRG4X8VBifVjZGr/Ow4dJ/mCBQFiydT/3bfYKQhiR1z
q93bo1mkU/+bYi88JR05aFbYuEhJqYwXk+rbzobdfxFODpeL/C2sWWf2r6ut+F++LCAd1dYen5lb
YhNLLXoP9dSe+AGEJLHfUYBrL0oavp2qSaIz35NGUDY3tewt/OSZwTw8ehg+l9uiuyHfxFLOkPP1
ofzzXDaur3LmJREi9SzwnbFnEheQK4stetYfk5mAbeJbe5AiStP46kbhmvGuHmPt96fj9nBwjXPW
xJxI+BCFhnEjbTg7iyEV0Hn9TdbzeIvmHUXac6WZODBANqys8Z+8YzFVvFBU1PINlV2YHltxR49u
+Cbg0lVhsTiJ+daCvpBk31GkTDbpvbD4O5/bmPy9gNCo337ajlsl3yXqQuR+a4hrEi/uB2GHKPNu
sBRYWAfXpf51Ih9DtbK/Og2gpbddhAADkAVWN1gyEY2lB57cUrNx6gq5hA8vr/GuszwnsMhTNcEY
q4ickwDOj5UitnuxK41lfAU77pgKr7dq6X61xkOhnKI+j2iqsrRimOHqfOLQ+5ZmMW5d6X5HqKhP
GJcZs1OjfUmMCbrf+n7uDBeTQYkJO/oFtiFIvvvbmk+f+kJPZAoqIDm9q87rSWnDXsK1T+JRzW+R
7N3P3XTLez2b1I5q3kvuAjwf/Vz+cvW65upALfSJN7jpc9mvhhF3P1ajq3cNR1PnyQlOIei8yXfi
ORUMNRrZDs4NPCX9BFHTcJHhmDksfVzErmy3IrJgWuIlaaf8fPXfNJSgYsjXdbGgOweq+YIxND3a
O/ZxbhTSdO7QIwSu7sXUBZZaNkijp8BMWIIrfdgmIRdRjOSxsByYEjagfw7cmyFDgiABtSa1/Mt0
toiXBHbVEBZvjrFLjE+GtUZR0KN2MSrdxBkWlBKsRdAqmxj0l1m6Xi4X83GuCxrEj3p7YUT0WuPv
7dP6Fond0KmhupuCa+nDBVfZB8Z9ged57Q6dgg9H2dRn4Ig/X/mcVKHmxg9T3KnALMPTNYy0g7qs
Hb6J+9IaHYiRVjJxnsvr+8qpRBsRdYa1hhBDT5/BZulchOxYEzG41YIUnIgT2enKESBSW4k/9Skb
Scs/C3Wj40OOJopb2+yXpjKawnlm8O39aUkzN077PKXzTPow1uDiuYF7l4Xg+HvF55G/L8FKr3yl
H7xHzHs6aBOX9F+eS7waobw6bpeuc7aMT67hfRIK+uhbaInVIv8lEaDur/f1JKPBy9rU+811YaQZ
1r/A+IbQTfcOQi2C7LOkvBr+RF3QUy5F6y8Y8jkSTOmgeJKOWP3n0vnOMhe9t48l9MFf+SOHPAzg
0R8RPS80WTISdIE1Gk415IdTE1SUmQGTDB9Wyge2YdcpAP4otTCQ9KNh8+efVUyA6EVVbEI8WMe0
C9UFjnSyzsaBbDS00id6ZSoroP50Dob4CqMWpUCmftgX1c/kBvF+Zg/jFb8kg6x4JKAoiMHvtceb
Dy2Mgm0oE51NYZ7/Kd+3wLA8w9b0ApTLjJvkSEzwkNa6JCZIf94NeHLPb6AtXRWgRUsZTnt8v8kP
mnuUqmV0pmL1lF5TFv1p4XdDW5j7g8nRyhWkUP4Oxpi385rDdq1ddu5u/0l5ApCO5xJpDh35RSzd
nLu0o19rE28iZNGR/5WLcrmXMNivGQPVBxkShNpUu2XtiSaH2A1VjGDomKXlIgwaDIYvlSUZLlaw
+ezNwyNxIkSZZFkTtPZWLVcnvUm7fKTHvExKxrf0AAfjhSS75bUIApRhlRHlRPNMPxDtNvhU9qRI
lvi/UAc1yhW+ZDylFtE5908irFbFI3E+UFj4a9guM0bwJ4zLngg55913KNHLNq5rTmrAbtq0qSRY
KcG7VcNn6tFzGewpj7w7IgAGAHk3Jz1CP1HJI7oJjqTLSXICzybojonApCfVKr42I6hNaLGw/zY2
6HON8EC6joa2meTVtMXRIyq3vBizbr8GUuJJLztIdfOnrGSYl1xHxM3cowv2IXzwOHldJICTuKHw
NPxf2ghsLswKbzu5VxraCNs8WwPJXZ84CcPWK+JBtg+paiJwLrOAEq1CphknpTkrQUa/HPL4Z6T1
3nblEpYZ//Se+rF3HNpqMsNVPrFBeuzAeAnLSpthHGOwg4DLXgp+O84SqzGNA6QxuowaWJjgBTHA
QyxFE+KOIF4GSBbzoMuyG5RGWeEGw8G86MdinQ7PRI46zZ2/5LBGT1wdRkx9GBCV5aPEv9YYPFZY
p9rusahHPJ9wuGbc3M4K0ku6oJrdk49Q3P+uJH+K7RU77J4LoxhT11CsohI4ijKUCSQufVysiaUX
byq8+5bpGDNtU55mZMNJ2tAbuemoFqrCVOvgetrPdFI96NQw8d/v5DuTwIpb0e7+TQdvifM37HFj
F7nMe3bsf1a2HBQrpRfJxZjYAH/eN9GK28yuUhafYTsLLkoZ5IMfWwQl02siIer42iEU1Bkgucj3
zCmhNrDEy2SvwE6vkJNBcZJyly23+qN+CAOEAGuHIfoXH1sVbaA2wuCoRD1n0GB4iFvTjZGAlPNw
9GiFYkUnKZUtr/IqCSwzjH4SnoYkc+RqZAyvdYd767TDluJcuHPRKmtzHhvZUD1rtckFHCZ4LzGg
RMz8LGHxKmI4fUdT/gHtEc5jV40lakZGt41jE0bwbAu31bQDmK1lkYUBTxUO/0goQ1TAH+fo2kN0
2WTb9hSQGavXmIQV1cBlOJDUELIZFoDSeBXU/iahBiEZpWdVq+ZAjcuJfBIzFCV/rQ4aYLgRCAli
nX50HkApMJYT8kIxZIgp3MtK8lkhZcKweyGpNct7Ud98imR5t0GlFw6AfX/uvfcVNcH4MmxcsD2F
K8ZsdYqBzM2Ux2BJ6BxGnOJ+okzWBG7SAltS9zlVxPbqz2Da71zSnWGqlwcdl/7NghSejVKXxmnU
Rr3rbOFRaGosflQXHwCuMDCpFFxrM8KsUOdtlLaudNI4hj5RSQjVL3/8rDFU9qWsGV/RzCvbnIDj
RLm5wqaf0lw9JIE9C4xt+nCHrFDIzex2OWAH9qyw1nmqDLoUhnQlq7aSiCLJ40074STbD5CKTkNU
+G4if/ol/LAX7lOfnnXoQuQan0ws3heILbUozc7eTbCqUyF4/ZmI9taH6wlEHZvT1HAwZHBZpx1H
wSSwgTfyrcQCvGoJVQMdXBzPq53+h78Y/4oPMukhghvKAe7OwrXLsxaDEYgi2O5n5nStLxPSalLs
OMpPgdhGM5RTcApxuLbeWP+Pnmtm86ez65wfQl9WZoVphRqsCaoo8vf6gjfJiX5bhUJQJzsmOhit
Flu81RRCWR/ZitXNsHCBCd+zXzvHY+VjW2aK6o0MXl0upPUSQ9n1YfjtecqbOanrVCtzcMMLCMpd
KtEp7WYA1UpetANp+OJIc4pVMRqljNGyTkqjB180fWy5Wz6Jvj7dzY7+qLqRVUdjmTI3OpBpABvT
QcoVRelmk4lotuNy41rFNQZDXBoXRYb2kuI/09DxdtkhOWzpJVrAjdu35NVsKdbD8ocP+QzTDEa+
UmezD7TODAy6q07tOsOf7cF3UHexCElGGNh3A8hkOElHCrDbhrGNFQrdwlJRqE4ksYOvW1c5srij
uDMoV34nVfiCnlcJeSs1cd9NLfkSMmWQ3cgzjRh0FAiU9zQrmy2aJTTgLlzE1micCESgPWjLDW5a
PSbnaX4NTaI2Lf1NV1pmHSu7GzBAiG1mAecu2ZS7+jc8UW5+ANBXniTbWUH66VwpZX96MTxee1SZ
wKW3Gbn5npOdXCfOHAlON0AtwiSUjrLYjsXnFD7/WqBp+V5CHr3B9NVUMlPFDms95Rvvmnh3YrSh
QlwyJxP0JcVPvRLbo4/Rl5S2jBj4RbSBJcp+Fy+UWDpGmFQOMVeQw5svT7ACfxE8AyKYtDbgHFoR
VRmYommKAcBuZCu2UF9FMenPS86L35WjcpKK4PTpMZARz+H4vmc63mVqZCsxUoWT7C3YBVUIPoMy
8owU7A80A6fLPw3NsWqekE+S8NYklq2dxEgwj2Usz7Yq149nALVgZ7L8Ea9SkzgWW5nKO/VC5pcX
+VvrNByBbGTFnjoU4uAh5BxhUwvgyOsidCgDRoXn5giV+5QSYzKXZoMA4HDzZeFdqpYXKDy4aNps
9hGNdg3Oo11cFZ/oPJuE7VLVIUSBtsrnWVmvsYGUhB3kVEjy2vaCsSrj2ujSZGG+Tsq6Beyq+Fr7
xnunWJtIAmMQVqzNtKH4oLLw2vZn5nOqH2ghQIrBWa9so0JgMqWKAYb0hIEUAWR6vR3pOSvPc+gq
TSYF6XQ0AbYdn5DGgzT/kXgaPoEilyWTJ3zW61HrvAgjIji9H8U8IWtFTX+M7n5mz1HP3zHkAk9m
vHx5JMeT3ArgI1QsQKjVg6Xzq1WplmEWBc6jtMrGWkOUeFuN8JGSgE8U7yHhJgoycl9LYJ8IMu9Z
EsmGw7DkafsW1BIXW07GhEF1BBnJxbgSe8IM45NEncag0wZl6DEuIAE7xm+8PM8pIcei+9+BfRIs
iLu1N8LXj0aPAOyvMk+gee18dLrv6nTRdD+t1EMtw9F165yz85fMAnLqeppDAw1vFKdos+ZaaIkz
+2Ns8Diy1c4wppb+v7YG7mMBIM8BRcNWiGnigZCwaRo/ew9RJvcmJmG2vB9v2YGgTZEzhuQPisiz
VY/3Hcg8ardcWzYzs09eyR3vr6o9goN6WHlBsHQzfHzSu+UvzvexPUpAAmzKFKociVbaT18cn8Ak
/15MNHN7iNDcg7J+CClKTLG6OcmCxbBowbwCN1/TVrL1+7PodnGKrpChnPa78AcE5KbeHw16z0Wt
JjY+jqCdG4gsOR3R+SodShdrVhDgNQO0Hfa8h7rWnDTzIFS9+ixNMBPCgfKjvmUB+oVGGe57g93s
9wNqqHIhE/gZGALJ5oz1o9NCASEEuTrIF/XyrJ0GrbkCYPe5cPieQi1np2WoCzrf8uH0Xf0bqge9
b88DdenWKNIZFcCxn6DULPf8cqefe8IKOodP1JjHUcOomnIRmsGNWJNP8PNfnrPKJ+S/vSjWlqHb
pjOEabfOauZjBpSjZ6Z1yRQ79WEgs4YaG5MV9g9xAYG3IZ3pLh3vIFsQP/GfJauxhAH847tCq7A9
IfFWrYXphbpG5jB/8ar9yS2lXL7JrBafmEdZjDN5IbDaVAPWCIwkikbXf3LJHXZpf/klaifzobEb
OeEQnHJFQhHNgkres8LMCTmUiAzQSd07yjkbM9ZYn2qTNrxTAttpFXAQqNpz/yFiY75uL+Nwev6L
widB3D+a8JrtJkrg2sdOuu8Vhj97YuELmZb0c3ycZvFvATa0Wcxj3OQLaLwD3bnsPay48I5MVp43
P7YbQzsby1hXOFHk0T1cT1phF9fX8fZQyU+8GkgsDvAtVKmSQq59F6JNnB4+2JooLgj+cBhGPhRC
atHIt6Gz+S5ZuilZ0wzgrt1x/PNGwht0L3yoXHu8N9gCgiXBJdrcwASfgOneDwTHyMUKew3sLtAj
2pIjIn8AqU6x3gx6e5PSfhZWP1d7UHpYmC7ik2J8bOuvwLuJ60cwgP769PthPPAaJkTGgxRC1tEa
SE12JnY1b8Q9UjlCdnLHrvoHYP2HCTdYUblD8a3mKSSEjH6lzlcQqckhnQACFMZ9GCjgy6q43Idv
AOH/aFocbEBHKBzXGx+s7Mhj3CAg1ywrBrDW46L2C+gx8j+GDdRyqfdkFDqeYKhinyI8p47+qFcv
kHl3Db8OXwTtQCCv6QGmZmZ9IpHWMjsw9uVHzgeMLLwI5RjftIY6y0iIWy9Qe+nZWNEJFHEYA8j4
jeEFjxmq1y33B9CmgXpNnowOoA8wqJkDNKzHaFhwscju8ZAmwb/ZF07VUDpPyuvoDiu9F//6BuQ4
zdzAtwHEca0Y8OiU3bxMKRL7JA+A2vC0FFUb+yMJ0nbmoxKY6wmI2OJt/hD5OgvWFSl5nA86pEnk
55M62eZWOTLfghSKmT1A8ND1vfdn8gZ+JhVG2NfZtIVZeII23QBMqSmAxe7nER2jpyOz6x6Eg5lN
xVC2ksflf1/9XTHjFACH5EuXd9/WjOHZqCsBW5feF8MPbDaUCccskjaMDSqZg5kU1GC42uyv/q5W
EI3CTuQRiZLhVcYpbQjju5JfYsN4KJEfGwyoInizAbj5C+snf2WQTYKejzZnEtGyJNirrVz7+Sx0
ab2PpezCPhhW32/P5FBH/DQ4RujOnAbMWjwoYUhpSpj5FCRBCkorAT8MTXwltS0KY7zt2+bn9Mer
ifPv91jPJBou//YIj/ug/Udtnl4a3nI0468dJVSMp8NqWLFWR+aASIEAlptkarAHqCz4Yt1kMxIK
WUR7L8src0g9q8fqkaVhR5VNobErsuxfqApPdCh1ffsa/+JBaKOzub3NwdNKMpPE8MYehHTbTSzd
dTZK1l8iSCpwiVvfooNsgPFBF3wgu5FEyJE5F/Qy4DNu89NeEXf+nRPvVS1bPnUzLf5hf9pauiDl
/1MrhUMGYczTcuApDinjYTAnz6BskFzCBvF5QmFbwlENWlSAO0NtAPKfw/DyeBwzP1NixM0T4ukb
EMwudX3+6qo6QGyHHvpAPHMQ2GqFmh+Riktj7PUfvRr6idPCwqYk8JqDrWEJUTfrlwGswKsrpQF/
75rByieoMZDbPXd9lJs3A+tbuqA8g14e6NGDI66pdi4dTjapCDbrvFXXXXT5ccBqvN0G7v+LfEw4
q/oNqirB1AQQKpZwd0m8iysfGY86O7UpkFi+Be1ie5yKvY9PFKcXNS47M5DUXaJVZargoodvbL0C
XPkTyc7eWpxpg/NMQZjjhvE0uuzEdg6pH478eji9tlPYD28r5JntOCxfHXgaVuFxIuY74tCGhwwo
DGn6aQMb5wLL49ydu1lok+ynUAOsdHKF4/QOkiCXfX1b5Sf6019kEJjzXHh0MqOt29DBmugZ3e5x
rUknzGPaI+tC1vN2DePhTfCgameci/CEd4Wl8YirU93/rZvTbphAZNRJO5GqMHBM8dmnIoBZqJfQ
6YwEqNt9e/uy2Y7zRHvaf7R3ORzrUw3ZRNTgW9tXqpTDT1pKpik+X2pqN2L4FWoeboF3OqHmWr9e
2K+dgSxkhNSpP9QpVh6t0G4oJXA3vVMsWkbpIyXzcl9X1TYDnFGaPXtTmLfA26z16OaIsdOeTu+0
UAfoVlx8SoIiyoiCt2Ejutwd+bUqx7EYoLKhh15bhSZ1W1vs7EpehX0DqZFSqkh50mQMMrglHz7r
sesQxuolnj+OS30axg8nILVpVwRJPdAL1TgCgLvTc7dAi5ajbpc6M1f/j0rBfNkpIfl1T5kgGZGK
MsDfgZY+HuAGN0refzBVGo7d7P8C36xowLik36vTNloBcI0+wrRyCMsFUlTyKoB8sVJMNXJerCgg
P/CNzJBIIRN1TYio59Gpwa1ZgoMtSNS1nprLSJy4jK3wL49uVRvspt09bMI2SvNumZG6aLKo4arp
Pd2DmPnWd0DcWw/Tp7q5rVE+fPnAcGndOmhuCaltS8jMC0tBwUDATqyoK6OE+ihuiweHSW5N97+2
pmrJtOAs9pQo4Oky56zsR3CHFTtez5iDA4TWZVFcgx/7LN+3bqoeig4b/Z9Px5/+6EM02goo0jlL
dEDnLwuRCV2f50vz17EZiHBImqkCI3xRdPqwehiLa59iUe7iCKvhvYwqQ+vzG/N/4thuePMT9cHs
qJaP+wFLcRVNt9eOE4P6+N8RsjjSpjob2xd+nIn/JFhzuXzLJwkFwshjhyfBrmta8Dj5AGZtinQ1
gnOxgyryYYM/scoSjXjehA5SpCyL7vTssHDTGce1/b/B5QSmlFB1svgrqXr/Do4rLe4MRM0FVU8R
v6BWihl6ajz5k+zUObt+amNaYmeYw+XL9qMkyIZ6K2xFwtfQqQSE2EeWVHGNvoswUh8rXTkryknO
wgOovPxN2nrm6MOSlUKImyFXouQWOQC5hngXLfAhJs4S9lmc6Yrq/6ugFyuPtNWpE6v5YuuFgIqt
2WOeXRB3SpY80Heslp4J3vZQP0grRLB8Kns1S9qp5BbBqxugyxVTJc1UUbAHfoT7gwIJWcaSpKFS
pit5cPMM8OYJ3ZrqMFk8XGGjegJ+xHjF7+gV2rm6FJl+Wd7369ukiqAEUAV0+9LTsMPDFhGu/2FA
YYGmTAK1xB/QskLPKqRjo0oxafqEQfp2YqOvTJILeGdSLGlTnSGHOtcBaBF5CkMKASX9H+1zsPv+
bT8Mgif6my9m19pUtLHEAMKozVq8Q/XdbCWZRN+kPpCUjWLQjBL1SiprKpW8TcLYedt7uhsj0mP3
ckqOBqR4JeOEIaj4XphAaJwJ+rLkHAZa244MnHr2REgkkTbt8XpGOU20c3CTGcBiQpIboPNKCZDF
8aqbq1vo9kmQCu7fNVrywikZd+qPSxZzoHILVrGAt50wLyrzHFMLltK4cQQon2zDlZ25SCWrsvZu
uIpd4Km5sX2Alzp1qjvnnSXsZI5kDpNt3dfRqXuLLlZFADu6VEa9GC/OOiqK4l+eclvaMdcCZfr/
fGmImVc8VSYSKJE/gPJ+E5YMfCwgNBO9qf6NgRfsXq5qZSxdHHlAS+OfuAxnFDeuW+V/XMdb45D3
Fluzha0tegP5Vw8Zutv3uJVWr6oXdpSKXUQPLk+MYmTy4b2h25q+AI7Hs0gWicU0Mw8MhhWhJ4A1
LRj3EhuHIs+UaY+qLiuqRu12XwE+MSzEf/uwNiX7l7gv1558WO42HberDmMblzMm8z/TJn/qcvDD
il5pi17fDycS/jKLsweJwEmqYUEhhi1DKBhia54Pu5XGQVMzOGyMhAfHaIPIjZDNI0vBKcSfnMOS
J17izqnUbEJZ9GqX0cNAwsUfKl/TAEkvg5Fi2ckIQ7OFw15U03bhwZAMSpkUQIgcLEEOrmM4hFgw
8Df8b1zORVAeXGApKvZDp6C6qHKo5QnYFjZ1BstEx5bWbmSs7GBdC/u5PPmx0JPXlhg9Uz33aFUT
x58yJ7K5Qp0AzLbOf+O2EJ1AtzORW4HXirCBA9d1VH7KE6TiWTGNCTdIenFbMOWAFvOxXcYvCXYZ
K9JqS8T2go9QGdWUKA7MYI7vw7UnmoW4KRv/iWNprm7AbFaW2kcy1C/fN5mVwbkbsUh3sIA6r5AW
Zr3W208IAzbkZywCLKTnF9EE4SnRcb6475B8+EI4RGSoKafa5m5K66tz3OcCZlxMw9pKorcGMLZ8
A6YNQrSVx37XaaB2ePEJe1yf0s3PWBMx2uFSbDEm/9+J3U60EGMilP9F9tw7SAlIZa7d+Ms5QkXw
tH5iSqtp9/0xiEQY/568jPSh/URg2H92tvmKYUxOrB9Gua7K75wfO1pUnLbIKxEYC047udF3WEZy
lD8iQ1vYpjtaO8hvOug324/QCqcase5D7vmtKwBzynlW4aQWzuNcgjWoViDLZ7krPmigvDf2LS3l
RIecQYzZlFc4PY2Qk7sT3AEdj90sVSxdxQfxEsKWNYIpt2WQUYcyrocoTAVTPzSApX5n6hq4UJtg
8+Pa+vWnH/In4PH46VEwjnrZoTvhAtUOXvnl4cGoXTZaKgLVz/UVre4zmarF0kFneTf4pm0sPv6Q
Lqb0S0tOCMphG3QF4M3kdeZ9IXXhG75MOvLa6Y727V4ch45y7P6JDS7ZBhCEsuGyoqwriGxY86rL
K/VUCLByyroMGjtFi+xN/TJe/ecX8UpfeG4Y4H/FfCSK52jyrDvqG8rVLEusnT11yMpYYjRYZav+
Tb1ulTgjulDDy3FCKIOeQijIaG0sBpUoC1Ps/Ps7LUHFxR6jypvq4Hzt9c1M4rJNrub5PIn/k8KO
jnbc2ajuMdVgns6N+yEe8wgkZU0OzGa2Kgb36ammm3Jbgg6PG+I7kfN4URMJeiMQ1y++m3aebkR3
QQyFifRbBp9B8P5ZhSIqSKn2B+gpLzBSsqY4OMEkYa9v8LmX6y2fEPjyv4F9FbZ6VPRtmy31Zi8Y
boNi//C3gb2Q0lLe1Fw1fGRmn/9U5iQlaWXEFApiRMVOJOR6w6OYkmFBWgjkMVKeXFlDeyaNLmvt
KcLx/WGAlPVYN98/drNvw7Ge7NhyxBAW9xuLGjcIrAawwEyJkMSsSvilU8DJB/bBzWdipV8xM6S2
y5Pq4FmZBnqzuTMzpq3bTk2Q/eO78gtohmUoy2eBKTo6FSRVF/e2kUpqeQ6rN9Nz+D4HjGqwmwcK
L0wfANmtBcIHgEVqhwUoV3nBhx91RJmIsP+3B3UCgh534Wp3rVO/xkaac5OX/eQFwRhLnFUfHLDu
NB7UUaf96LAah3PH5/jOaOu7SMNhdyL77M9wmUsOaxaqZiXZG9zTtXDPkLIASozn6fCSlma/UUG2
8ViQ1x1pocAH6FK2H3KfKmmTB57l3QKiva0ULJlVBvUxt6+b6Bvi+MmNxPc8QQpDbhZj4wXFJVxj
3SM++9bMnK8OYv4WD+eTQVvNmF8kAAx/PGMSsCrcp+L/KcIiwodidjqwkJEWBMwuoJFMEpMHkv7B
lY/DSNO6lP0gikXte1BB5xw/U8B0m79GX3hAjKMy+y3VfMhuN5Ye2V1t+lQkrUbdYFP64MwLwzCZ
EYODqO0JXM/wvSgJdC5MFsVa9w50hYfvzn0qTnhtSViuInvETZKdpM2Xqh6fE60hB0ORraSj9+yN
/9oKRcPmxC2R45PXh/niMEsjclIrFE46U4RzB8TMmNuOiRIBUdP87PA1mfUr+PaDipkZEFkYroxQ
sdbWUI0wcZx3lNAbF4oNcGb5Z3aQP7kt7JYKgbfBysmPKFg9KNO/WRr/0t/Xm6AogKLCqKgI187R
/j6PpYrukxzI2t3Vsw7NvpOc/IVJuSCxtr9yeGLw4yPVSdG0wzDnNdeITYx1wJfFRAicMojEheLj
Ht4eo3AieFgJRhVBiIba6rtWLZiFWCPph1KTHp+eBAXYq740Kx9ufDKgbT4IoZpvAZX8lCEYZp5Z
8ay3WSIZNm2m567yABtIbqPyNGQgz5NmMF8KJ9+quubK2bXjQK46peejH77PlZwl5Yv0PD87De9v
ckU1DVHiGeBnQlpz+/QXrogytfB7wfd6bDE2Ek4I1oAYJDAuHO2hE93/b31LWZOUMUXwdQczJCZM
lSX3lzkC6z9k8gizYyCVA435qgYJt52zjyKSgWLLCsW0FTJQsHXCbN90maGtYB/XLWFcO7039vBZ
2eBPjwGIGRKu2Yeazo2PITcZnl8CDWsGXyVvXoNQPnaN+RQ0ApK1OVZY2tLTsl8gPdN5d56flOcM
V81+8Ipaotx4qJST7qWpEtbNo3dqSMtzK2PA/2co147jUe2Qw01M2XA7dZXalo7814A5jSRTRVc4
MbAhZmP7ZWp/3Hjt7qHjKHNdqWMt5cpKSVzpc7gOe8+KESt8pmc/1v9FOIHA89r9pO3qxvN5irEE
dOG2WissAYi/U617ibWGxYSevCfseHYMwQvBR4VZQSPTftdokqcA3Ta5l2KfJorY2rXUL+adq0x0
Wjh14DmT3zK/Bcr3XufWYoviV7oYS/6CIjgkaGHhs2hJBOiaE4djvmMLZ6qDheBnEnT2IE6g9FoW
KgJ6VS/JCFTy63RM4w/eAWuOD0+oypWW3Vqn46W1U3I644NKTaXdIIE1sPcTbzl9AUy6JPTky7mE
7YA2hpqTN1Fl5F+t/X0gMLE0W5mRpl84vqteiYRkpqC9+soBSqzEGvqFmgf8yRJPma4taDqp5/KX
PitB/Rh1yFCNQ5uaz5uGYtA+1nVTsyz12/1V/2qk4nEHhTLLsOZM+E3GTxqWIufTG2+R9iwBjJf7
yK+bcbyNkHt5AtDGTqnhv+4fMPmwCKahgQ/cnU8HcA9PYunoBuFuNuaXqAYM3B1edToL+gDrkEMW
Xh3/4Y9oa/Q3HE6mSGvgql9a7lTowFPWgdxC+1SCrDJMN3iKafgQhH2tZVFbQTtqZZ9Zo/j1PDyT
GsDCiBvasOIuuUcRBOw6NkhM0BpaXWek2HiFl1tYl5Mf5r/WfbER3hBwuBEI8LloJjTRdbBlSRpN
4cpQdFplWkwYvK1l4PjrVw0HaPHjxfXRRxnrn/gjIdYD8GgzgnCT1qA7cd57TzbZsKmXlqHDU7av
6yULnpIYuGFopuOkshAd/CAJzbMzlnDeC38gU5VRGFR5FQLznV9LvMTJ+emhCqbEvi5xBCwG4ohW
j6d13EwwaugsePXGqC+DUeYz0iz6UWuIp2qhtQTXO2livaRsoOnYTD8zJ/qKhauQc5WWBwjgWmpr
sR1by/pvz648/i3u41WL+b4XTVdBzfYFmLx4I8D4WA2BOV9B7IZxmIYCLwOujl8zq9GXt6rHzj+a
iLgm8pjOZhbqK7vhwiRbVfCuAZ+mbgiWmYMh/RzsHRe+Int/c4OG/V9KDz44m1Dr8TpxPbjJNbBl
xPER1+ijvgLoY23jwsqy5HAhjeYWjAPGV9KvRje6VxvccOatkTIG5s0Y3kN+XqCxhHdQD7+T70VB
CTZoRwFe8WLJqiMk5WxM9J1400ANFLaTimdk/ObzNdbyGhnRs1w4xkcxmbHlDKyI5OHckDtDiVC5
AuYNfuXWv76uD7r/JqCSdS6OySVzauWZs6yrE1mQnkgUcG6pGuUcy9ONisggOhHsVpZSoLcL+AWK
JgW+XcyKHxhL5f8UIk9/hHXgrL0g9L/nYmxuNngQHv3mxmuym5Mjvlwm+e6V8bsDRLuABXHNjmh4
X6JBEDdPCPmT7ZVnloEO7I7LYoh4NPXDQpEUEjWXfTicS1iX/AuP0owGVqVIlLXbk5mSoxIBDYt2
/JcjrbCsoXyzvuaH1rDr4GtTPYqwgITDS150hinbtCwXnJBmEQa3flmTS69BDH9+UuJkHXfTvNrN
IpM/XU1ub0O4R5VNHWBk76X/piNPiDCtqaA1sRiMi+YwMxvnq2alQuvEuRXNsliRFQ1YiDS5AOD+
yEKwRwDeqMicyZiiLwA0CQC3FiCufKFJsttOaOGIPh97lWEfR6cGJTBgtzj+wFC6F5HhxUDTHBsO
6WoMEb/kQ7yBrbPQ9wkFNQG2eKs6jZuwftQ4QHmBhmwHbUsr8Adw+8UA96PW1P2hj8737T9YOSc1
bzyFXGVpTph8ln+WC+UKyE+KevUioJasiPGBQEd/Q4ZfAoPbLaFelzM7/AbLnDWcIfkfwgHAR7GE
2DKUsXjeiWQloMu0mwDUB1o/zq/jPfLRJjnG6LDUp4homWEuv16jJiszg1NmOQqucd35yoPuJWAl
4VQMfOUhiRnsFWj7METYN8Ka01uc//2R6O70dA2JArLF5YTCwOk/0wnIoj/rBvpQUTdVzuAf2Lmj
VFRVcdjHwcuohzDXy5EcCpFW/mTBbj0rTYUJZea7aNkj+Fv8jvbvEAJfOPg58jlixTSQow0JdODN
tsmh9e2qg2sfyXaYbjqsIXxkU689IqlMpo96B7NA9cvzPVDQmU0TDijA3WWh8YYHE+BXz29MU3TQ
cWMa5lnauEAEDcNtHjUj7F+oSaW5dEXqEYTqSj4eisPdXg3nOHnv8gXUXjylOqBJuOACYbXXjJ8x
80xglHFeel0W6Gmos8+utyJITLPgOVCSZYxiDIN/R0pnrrfVSxbkfoQh34LtbVFnJPSilYHcXnxA
WLslcrcXc9J9qoJydHTFWR6tmUg6Ih2Huaq627IQfo8J4ohWM96sD2mBP4LZ8U1AWy+T8tmtBph5
OkggrW5CNtEc/ouge49NeemXgcWZAGooVehuJy/Y+znLWlWgujSGEyxNdmbqrCnxt/RSAOmhxArr
IOgtMJpgcqhlBip9e2lTw+sTcT1xcSqEbXD5eQ6ZiLvOyH6Pmd3Jz7PenqKB3DF4P5eEn7QTOMpT
20+lruo2vVWvZRXi6GvpY/cKsQr0ynYQQJsO4GOWIqTt6cubC7dezxDcdx5/PWLG/sMKSgqo8lN+
/YF7qJWJ6zRFH6dUzcyiUbPaIUuG0kc4eI/cWlAEgjnOl0gNslRFOPDvIvbjm/X0dSafkdknNGHL
oaufeYYAFvpOpwNC/vZrssKw4g6aZ/f1+dKbGSLdf8/dHktKMuZeMPUxE8CBTSjAvUrloXpx5VFb
VWsofFuV/z9veco8MUkfbn6g00dvCX/Y9Fe0wBEMUicRE0Wsbd1ezYmF2fJ+XLGolXnrKMvmIrkY
htNSvGeHawix2OeBALpK6IK/rHnr4ztQTpYAiGPH/8Kpf9NIs+EDiPL362TwNVA9Ugfl5pWRarpQ
+NP8RRuznVd54evccEVkFkqkRrNRXgTtoVKmf77Df8Rj7n9sR7IosgxKs+XP4dvqHag4ZDl8Vmiv
JLZSIjpm/CqiUTjyC2yfcdme5E+jvv39AGce9KxLA0h6mu7mURgdLCH58ovRaGK05Pcj5LKQyT1O
6rjkhGzkPBQGdd4UbxPG/zsi8dgI7eQuP7Tgf5YEPsxPmcw1snZmHE/QxDRxA7QKLYgC17ke+hbU
kKIbo2X95fCAbSIAk/IhKHEJTMYc/M2rMwljFFUW1pQ0Q3PeGzKqHka2ZUGgFEArbMhMIyEeQigZ
ImH7DsgivH/MlrcSJvLKFSHE3WgtVk/WgcOJJyoFNKJ43p9Bsg/xer3M1LbwPcXSSeHyGRDk8/tc
61fYorrW8qIPmWadB3xy5DU2VCfomkNaQ0bef08OkWfDLksgfXDwMwXTZkEQxCUlEcEwuzm6yi+w
Hf437dpjB8g4ZLMGAXBhnuT8CtvVnFJsp4T1E22QgRQ/1YnHXT0ddQnV9S4/d+0E2FT3B/U/ZeBx
DtMuCb3oVX41R1CNzn8fQgOxoFFqqLBD8Eey1Knnwc+P/5mNRT9QhtPOxZ8sPHOuB48g/ImBK2Vv
GgYH2rkY0URbJLLKhdpSd7HTQ3dTJi6XYnHESbZT+GYQbNWeVwUqe+QaASpp7BYySOUSPBMCTkhA
s5dIfG4xrQccPAv2evRQrDXWj/1dm07at31Kc6fpmAoDrZbkncKTJF/nRGDx/Cs4VJJG1pYy+zR7
teFO0TKMnidfGZi89wH17na4iLYKfA/xUJZXY0LecSxdDfk5OvYYPWXfaX5vQ57WV/2PgCMTZ2ju
OXPZoncWWYuNf0XyudItF2DiIY4zwm6aogP5oj1eTTspGRwdmQ9326NztYWKt8/J9tuIP5RN8vQm
z2tlSQp5XgYvyknk0WZKWxTkTVsN7ongN/iu13AME1UV6MDWYd2J7ctXzx4mnh64TJwIMwusa8i3
mn/xDx+hZ83QPREUOGdD/DmhKFtXn8een64dorU1HNvFaf5Lfaf4lAxWEUlqxrEcvjMzdqokyp+0
Qrh93cRB0QeYuiAz+dbbQg9bFOH0V3sS7vXiJ2C1bmzkVbyO9HBFCLQVcx6Z9/dmoi7HNXE6yeK3
t1kREmiUI5FxtCvXpMAcaWIgx+zF/YbrGUnEd5VsU1aCF9O+2tHpteKmFRdfxF3qhyl3BBarrtaJ
HByOIlUzJx5OUgmxeunuAB30fT3d4/2h3tEU7sodn1LgciJpZcVOhYCrJ0rJHaGWwVxgmgRvUcYz
ZjYd2rV/3+EE0pGW9UQbhMRLwNPH0hIN/9Jl30D1C1qoiKtAVbWsSKfjs0I0Xy5v49tP6P9coFLM
O11ZbWskTJ4D9JR/dGfutc/LeSF6aOrzYClbAKvHgbiKmNeM/6QEcxZsmU8VtZVa1OMcnmqfZ9S9
g2K50qpUemvBnXnd2oyZ+6Wn8cl1uf7ve91vrYsuBMwCTdJDTXE4bEgchxr3in6wBnlpa/AUmblG
i3jP/Lm2Hu693sgIN1BGuhm8W2Yl7VkSWce52dwX9Y3/7ElwGOx1DhMGfRcnp6mO4Vwvqxeg3bQE
WdxyDaVNS6c1kvltXqgSJZKXGGW5s5Yqehj0Pru4LxmKI0ygZ5pJ/V4QjBJL4C20/gexuw/LJfDC
agvQpnUjXE9I6aLhTfEOCZqZHKltB74myWMnNj0BqKyVQX0Ptz09r2R+CTj8uJg+Md5qlfiL3Vge
LqeVbCz2qvJQPEKQKhlB+0Jb6l7pr4W7cdmzE/sJx0sW44FpoE3E8bpdYFAHpJ/Skz6jbrzGXwmR
tQSmmwNZ66RI7feN+9FL3tWp9o7/++ME+OB3ivLGD8jA9NMMw2gpTUj5+76cJU/OgyLKLvM/vCj5
g9heGF3H4ajlCReKIQ5SOPFvmdF6jTGSBiPa2ckMpdD7ltniZ5Wsejl5d2PXOYTJacYAcCyHb3kS
ak9GxLbH6ef6b3cKssfrWJ1UGgFdNqGVQUsQVPt02nR5GVf+XauG4gamplKSUWI+hWlQbQK/CMnZ
x78v3yIFi9hzVpXPUfVvI1/PxsW51862hr54B7015uV8tjt+02l6dwK4R/rEVqefd1stPyqPoiks
7Wcr01TPtsxrOcaJmH1+iZrygdrV1AzxGRXG/sas7BTOij1wkUH1eLtMkxdxH3tzSFCrNiLcUgnt
3HRE/fj3PId0hz5YVWeQC0NwLytoACmrsQE3vsGG0dFGvuFG2vCcokOOgbTeKJw71M1UB8WNCziO
Lc9MQ7hbVjyv/fQyDf7PdGzQRVyFQrD34+0arKapOwDKsVmUfIpLQLOPz7drYW58ZMhjrIBEC2XU
2/WDdIiSfpX1/OZEp02wIa6vXBKFhxMO+Vs/8ryd365zJKUzJ3lHi9Mon4ZLIjl4PJUEEe1Yi2Tr
VUV6lxIvVnqE3tXUgSDb8OmE0xT6Esr2Jh0b5/lrFZjCFSd9erf0iEEnpNzYUzVD1YcJXvuwoofV
8d75SvvgEVxbtVDJ97hsQDlvi68QCQBHbnnEaxwC1xhD1sYBRPx2Xf6Xl7We3qNz2wabewuvxwcH
B60qJf2fhAEbPmW5JtjtH644OBWCwrVrC5OCGVy6pV07GqzIDDroCIJQmvEA7yNZpvsEuSP1JarG
tHGYGzhrDuGry8ysWBUdhb09SVRL8o5WddUuNs60RXyyIxtQdNny4PRaEeJwml7ajDM1dcCXxF3w
o6fb6dji+WiM2vq1rcZc8OS5VSN7i+njQ52l1hc1t17Z2Fl9uJRpeQHS6so/vZVO8wYgMI9YcqxY
yT/T3Ruc5zKwaCGe8XJEwiSmJHrBRfOQnqs0TkKihTO+88goj+0U4bpB5zaOnpltUL06J9FQiiYp
suu0W5JaXdMnyAgRadt6EamCrCEsR5fc/IIUE0TNNRCdN9EmPpmKuQdXITxUP56uJ2ShTXYUgNpE
yB5kzU28thKrOoJXjTCSib1EdJJ9SQ4xb6bFFWSyFvn8daWK3GbYRtlBs9VE/bJ1UBkqce6mvLlu
9GOwTHa4p6Hs6OVDbVe6VNHB6ts/GvU1T8w3KziRR//NxmxkZElH4Q4aqTrPlCxHOjgaj5hCu8zl
npsmuEl43PXxESIIrn6efvxKTLGYe/vdOy8LBh68//XxrwXMQQkM/j5U/HmUVSaeLck9IqNXnP90
OakXFHcTyccqDdtl4Emxf4o+A/Jfo7WeKl0e7L746LVLJ1GT0+XTqcG1VP5FRPl62fBnnuvfHuep
UzJ2zj3PB6tEPzQN4jpeq5TP4V1pPgssOGQteYkog1+mPZSS0GA2KkFCDlpyYj5WKeI5IqGn4dQY
O/J3sEl+SNntqESsxOUgW+2QlW0VTRYeg8KFeySJ4PNQMoyN7OwTtxsXgI04m/NmQZMsQmHwqB9Z
0nClCmjlSWn+vBurZ3/6MG18MJHd8dK2bkqzFIbrOZRvPBkErvClNRfmKZCEyWxVtRhOsq9w/hPU
zM3fZax7ZEhKcvw57GDXVEAD7seSCFQHpb6usunR3dR4gfiiYF10T1FutdovO0P8q5v2dNIN2M/c
TtmXveh/z85j3DREGR6hr9TO84wBUwRV7A+Hrry/FfMzs9g7+ao40wNBgG/oHIZ4JJctfVh/UU7H
zAS8s8y5dIh/4wBEp7c5HfE3aPb4gtJvNVY+11p6BG5oabe9NzBsYcRJZYmXDeCtTehgM5OmSjL7
yGEzF7TSUR7hPjknBvD9U6dxX58z6dqdTCDC2M0ikdcBhjb/rD8r4uEqqNkWs8V5r5Mm+XY0naJF
qPQDDeIRA71vvzNCLzgrPu6RMBUx4ymS8TqxuwpNnbtdtDA/jsV2zB2uqswQMUXUS5G6AaDt3eHi
+T7L/UiR3abFRyB5BFhrrvSxPQhuzoTezExkgnuFRFt8d290OgE/isLCdDhBRZibwAbu7rtNxTmB
/XWehkXzd3Dq/OJHtsH4oSHUXQbOfhrdVaxtOO6OxtZvEDFbX2evqXGnUG3k0GB9WvkuKGdTHB5h
vFo2JnwDPDlDIKo2dZYkMTlmx3SUDkXbrhTedlkIwU1IOSQV7OuJSQ0GD0fHX0S/uVfkmdPBLx4c
83h/RihJlRA6NyqxcTqAxERALalj1w05RIXw3BoZgyQs5lXyfY592BhjXBpfqoMrZ2ZgDxaJoFaJ
vmFlnb8rd4+GnZ11tr1xfEwa+f/g3RiBwGKgF54ssKct5CA/ZMvsny4nnCfRMKZxZ9wDybUUARZ8
b/dNc3eGgvAIWVffYv/L6XtJQ4Sj5nmOubiAq+TaYifNhH5f+SysN4Gie1YzHLfkTyf4FGyUZlO1
bMhDOR66IItdluSabNXzV2mzdAgG2zQegF3KWdFilvk/BlXT2ciio3mJqnNXj+CRndflUmRvPuBK
nfQGgcnlZa+Fj+qUzqkikWlbphDCRIYBs2emd3X/CpOvRI19Xv/quVj6A09UmjQSCDxDhwGzdFJr
wltqQxHxy2y4erQpV/31jMyz8CZunPNYO9Ve3HPDrnrHAkNFMYUjUHGUkcjIZUjqnFX8ymv2YKvv
szRoJpRXFVIg3yHMVO3QJUE7jlT6rVLzGKA+0LQZbT5UtRP28rIW1GaIvvEGo1plgzn2Xe3M4nlp
er6yCe3VSUBEzk/jNWSO2/5/JXNldFpN6y6Ho31zx4SEYVyjXcqYTHqo1e8rEl5Y+roRpqc1CRBY
Vib3OOmk2YUhMUXKXFAjc8CVJpnWJP3+W+U36rfAeE+Q64gf56ldqCdqpUUIw80Gf2TJMw7qzhyC
FeX1jU+XVrzu8aaYLkSffDXK306pdoSmw1nhI4OhHg8Xlj1wtVSo/nh76SJDlENCcQkHaBuFVDG0
GXhG3IuQikP7gSHcat4D+pIyTiD5/52OdePs68wB9qyvaG3zcTCI6IjhyLfvwDTKNMbJZGAcF6Wq
r64+j/lDN/rpSoXUR6/vrbUUVu7uujnt/12r8ax9Xzlcil4yLfV+0QhEK+S7LvyxDSYShtZm0j0l
He9dhmWax5ErpgyvWnOE85h1vh7thdOPQeYd2LuoDpMc1TxVQ3wZPypNvPr6M20QpdHHIXCe+x2r
ycq19ewd9I16XNjn8xSVAXMHf5UmdNd5iyiI0jkgwP4tRNUpL6XEYb0pAdPmfnhfbl8idr5I8Cu9
fwpxWSRnbPtekLfVh4TBs+SlqXHr1QW0SxvWw3I/APp1aQ+sMc/AdwfgI6rVm0LEGuYSLPQYGgcJ
kl84SovYYFiP0Nr4tx/zCFpBv2xtYcWfEXgzKkkI9LfjuLIxBk6MnHxpkdoSIdZKDuhmKd/LPSlx
JkTqiQd0KAvpu5ivMy9Zec3MqRSZVOsSN/yhYBD6bQYGZTAwRIELppEEsp6g/i3RJVsyr+Z90e0n
pH5OdUYFtSyH07Xe5QF1qe6WiZnwwYk3xt4rcrUHVFBxw0hBvV7Avy4d9EQsW5kXlFV1dDB0C2LD
VSeA4FNBm3dcB1R1Zu5KgxbSKO8xguKyUpyhGxNH5GqfE9qcg8vSu9FHP+4RRTM02LBQqaf2QKb9
UlcgGHOy5q71tKT4a2lk+Y+0U63ASs58ZsJ74Q298FewqEKoqocyROo5qdeqh9A6HsOjYMOzU0rM
4qVcwkgsaCTvYNryJOn9Pyqb098ggcTgglGLaNhon6q+Im6ofsDeEk93V2AlyF6UKQyGrLMxQL7O
S5etyE0wOU+rFZvKqEPIr5xtNUAkS/+Ks97N/CT6tVcHsK+ubegdwKsIfsai3SI2HR+JOR+ot3bn
Os7ACYPLtu36ayVDMklnvvUS5+dNWIJsn5OIZZDXeZfnHzB31ppp6kj8lzNO8j2yo3fGtr2raxdd
q00tyCqvUn/9lYZN9mhCBtXL1YbjfSyjOJhwMkXN9qE6cUpSbx48leABT4EguA5pLzk1P1wewSH1
zk/edymFkKiqwnfB/rWDX9J1pz7UeTQQZfPt1CsKfn+GFTErpVecJJNRUv8GT/1RcSysUzM97N4j
rael7aCf2iqDHGgYjeE6xAnMlKFILRxhh4PYVcz/v5vob0O/2ue9XXUqQ2eBVdlyEtIE+QVHt5Kk
0uufdRo4HiE6ss/oIe8OTUC4VRRjPJmie/T9TWRBXtmxAuGTw8qOz5H7769IyPTdgYfOMZzK/aOg
MDsGPh/KmB3oK3S127qElIBJg/PVTDmQXhDH5spkNc9tQlVRQ3QPHr2eM87Qy9/0xCuO2z6PZW0s
flrq26xHKlD95nxZc9i1/D9xKjmY3L1NW5u4tqEwNJT6yirOvBDMR2Ti+3WNNNh8DjBeXlT1LVFS
nAELtqkbGbBuOD8kUnVhM5jGHwpNgqnUGlZYsAYPYWXoIh9QzLaq7reXziJz1V2JNoeuJ7HpULnt
ioXsLBM7AYO3brujJJ1EqbETyq+otYvpDUdK0vdsd/PQvbZEtiXWUsivsVQDA4U/DALXMkKo3sqn
m+M4nLgDSHPhTt4kQ9j5DQY1wnrKhFpglFWOBt+bGdwaKYhuArQsuaIAKSPfLuofEkXnSVOeUNNR
TUKMjZwbn1rTL9iToLwX0LEsvXgSzAkysJZ1Ol/5pY9UGowQVGOUjEYb58UcRJYfiHkrTQ3EEwzZ
/1K501CU4tVVJ3GG+826R6pWDRVvIypgEe8IUtI9cVldd9rNrqxoEV8JreTpyKqvZ0NFuogJ6VDH
SXY9mNWoGx0S/UjFQYBpebZCboNtafyCb/Qr5ftTK+Tcy/fxNOvyccnPFzRA31L1W/7j2MHtcPG6
LtS+Vj5Av4qXj8scpxnR6lVm3uNkgEO8n3MDXPmKRyfo3LIj5NQF+Ko2cqvSNiZep0/OHbIg3xok
AEk4+4Wlp3su3Uss/ANtVBd8j/ZbWpT/Hu5pSkjVtZYAh1JAdhnmtbRPRSxBAeaX0yzpeo5F8aWL
o1ZFZicUakatcBna3Wlz2yL5Wmm+Me1dQI5r0S91qJa8m3V9YsrhqHip03Io6nxmAVODPUOcfJh5
1CE3eWKfjSpnJLnxIN9YVTmUuZW0RFkvTHA0uOIJYcuoamwMe246hxT8l/k/XeZCypxwBQCbcEDD
f4vpubN3Ako1849ECoxGoGOxC7r0V4maC70+mdoXR38CJj+9vbmFVWUzi04xaGX1/l9ZbMd0HF/6
xyT3tSJTgPW9gCG1rx5OPX//rjyakIIUqI+u5WirLZxv5uFApdinxf9LgIvx+X3OxXcBYUhSNkLY
g+wqS04j+prGT5m4uOI2RDYS8qzKomN/kBX++Xxhq0F209WCv1e19cDEcJTAZomqXtqB1uzO9cI/
wLmKl12G1vc9OEO4fvgNYR6x1wRWnjMiL0jovaQ2PsU/rMmgFoQV0Ds0ffR7Kx8V/gjFHRVZVOnt
SF8Kg6H6CJdUCCt2YpB6MLNvdZZXTMTok1zmzOPnYprAHVJ4GbYVv++sfe0K11/ir3pRQrU8s9cS
tmmL303tTjBjzEZIfwT4ekvQl6hwzy5Z3+X0wFApoxuoFTWdg0AFvY2HHrVDwuKZ57etyL0A9Yg0
VW347eAUORaUJ8O4yuF7qj3MquqtxNTm9pXEs/RCQYWeX5UDRhnL5DTybdRUOc9erFz7UxdIA4bk
rC+MZrxo7XXLSRsFUfYxXaqIIuZ3rNNaIyZO9xfSZMOal7L9QTV5Dg+hU/aZXsRQq9jfmlqNBWwc
EgZilOTH9WdoIbXXkwpI3DQ4Dhqkw0KmU2oCOygtvyEOhN+eBpz72E3EhF7K03o695yzo7X4Mr24
yI56CM72i41491+Ufgu5v+tJhjC/GuXDMakG4JldxNOi6baA1EdtW3LY3nwXbNoyz5KoKx9TefHL
EFnTKnPkwG07imorcvqFf3bPP+ZCxoPuvXbvVBp4K34+sUwExIUBBCrUlInLxHSQn/urjDK3nIL8
1vsOHvOWaBKiGFyUBZw7iMxMOzU7lTUnDSMX8V/Elr2NPeEjKZ/sX4r+vSgWYPqH8QiizuQqReSt
Owu4KcfF2nNOQdusJaBkIGobkm46S5Kb2iaVkNkEMGL/8fjgV4X85Wdg7gpWDizz2Gl2l7C3cPPQ
zwxmpLSjSqJo58mMHSfipmUyfSipDL69xcv0NKg3YQhzwBiRYBecaWr/B6stV+pVr08oxIO71ihT
egiiMOllL3bg5P9UyzjGUdwkWjfydXfZxB1VMaFXv6yYWA+5I7AvRfSSQ/IkfRc4NXj1cJE/xVLA
K9L9+EmlqB81N5AHSsGNblgOCVFOVKl5A7aY04OtroTA3heOvsnQWCpOIysTAj8FrCCuIqZDd01e
iht4UtyxI1ithA+p7JbfJAKQ5p/32h3m5tdz4vH3hoakH9YMcBk4PppkhkNBtFTekQg2k+Lqh0zh
iBZvRjCtnBnVa5jEt9rfC41s5ugNnKvQxotR43dmbMYN+2zgpxI/MSkK/bTVtWUq+l6tqXRp9E5b
Uay+7veR5haDoJbMe5u+a218Mqq5Gpgfy+RWZdzG4JCE3QodIrQdhPdIoX01Tl4MA7/32XTabfNL
q8/2HacYKt85vOriUmdjAEdaelcOKx9OYQpYgweRHm/Y5d3Fa48sK8a/AYlihEzEGWHb+YQPXQR6
bqlOz3Aanpj4juwcGc+mViJwPzcy5+KB5SD9ol8lntNy2XzHKMdSGNJdNHKwjKaaj6kU2PHntlqx
UEyn69noz4iWvdWWnUT8AxH81faOB+WHjq2H+N/yxFj4/bQEBj6KiIkMBvJjr1cH207tkgemMTuH
ltha0yVEWZokmdfaL/6GttrqU1ETrr5hD3R+ikbT024sLFndWAanM91Wh7E+Bn5jc9vEjZZJGivh
0yVfdfoqx39v74Y4kTkC9k4AllBZuqVY4UzzR0PdMmJNZNRXaJFLA6uLQjXzX6xvCOMcS6i9S//E
Ja+ap/f7D9N0zwitwap9VJo8wWGu6kpqAWrdIORm8Swvla3NgudeqxGy96FU78dchO9zPTZFCC+q
gY4wEwKlbGhUHJjEd01czkbJlhMzWAFKp8UbKOEchERJdG7t3Jj6uAOyjcxjBGkDlwqa/+lPznqn
m/zpK/+qCuG+/ZHS4Y5i3+FPgiYSNCryqZlFZCDZAZnNS+hebnbRlh3kIar1oUrXGgOdtOdHjNQ0
Qr5qo0uSw4w+AS9VhEGodiMtuY3+l4DP0qeMD65FI7szTykiVsYDv0Bd5XN3Y/kb6zZp5BAoyq0K
eXm0Nebp7oDwybTazmzZpxcecIqHtrtO+tg9/3DHqYyJz4zfO32qDTJAQlwz6nqnFB2npzvIZxXx
syL0aba2OHHMu/8lNg7Thq8x3Q4qil5DR9NaJKxpF1nn5LJxVlgh28hY9W4Ckk13r76x5XMjVMbc
s49oVvs2K3Yru6ZQaIZ6cWL+J0HatdnNJcGEdn2gNsyPJ5UL2rUM+77L0+qx7O3eQ2u9LDQ3HEmy
dKXcnournUWgRCILXfE2g6/D/vdC1yR2mwkdPGzzkmbzhrqmrxTmzD5RmdD+393kTs9hRIc6G84X
8QjnXAR+c9A4XtuD4IPQCGhaMKEeLMt/7eWtol/s6N8A2E326WHiue508FfHhLZHAwpKdhkfbXXP
fJErD5DylQ5IN27XbHBfM3ZyKKWvBKpiTjcdyjT+m639/99axPp2QqTJDIt63Ay98mn4xK5YMH3a
ymxNztAPUwDsW/6qsg23VTrn+ro13mlOb9RxWIWgejupjkCVCaLGMtetVi8PfiVB6K0FDctazeLF
GADK7MrnngGMCjkvILQUNnhI7DGcoKQFw0JmwDdzrbm1A/wFsSFM2hxzC1xGO4gm7hQfVjweMqrj
QdkiuRI2y2gbQLFkwgXmHZzYMy9muingKLlpWkcf74v2vphsdmQfAttMrY5mcwRQv9+BznNZCVaT
6+y/uxMhHtFIYaS6WGiYxEN6jwdPBDeqJ2I7i5L99cKPOzvL6+HSFkD24/xX3YQfGURKZrd+fE/j
05tEdATP9dvgs/0ZzKscar/LnClz5pCYq1hZoc6+BkYYuVqKCa8ZsgLq7Dp3Cb36H22Q/mHvLyWO
rZXaF/q0NEkksBc6JpmYphHQunrQ0O5aG1ummw6z1Rbse4KxH5lQtGsEINQkuFJpn3qIX/jnHGcy
ZcpdWT0ZWnYeNYhcQ1Qet22dfLVg8ymyNnk82+RpZJZq2XB/dGXuRunuRpH32b7vri+z34ffiHUS
JAP56W3TGlCd4t6omoACWeE/NbaGlwxLn3j33191nxJ+aIo3D+2cgi7T1RXk3vrXvGhq4o6rGV3k
IMqbOT6gw9TNF7lnXcwzdmDZlFrz7rO7UeJFsW1L9tvuERb1Elfscaeb7ld5+ZPgDa2Y886lVCcu
YuxOQjcw3BPIp5Z/ccOizJiUlgnXVRx1JkmC5O7kPzNbhg2ZX8FQyFyRloTyvRJWs4O3G7e/ZxA+
SgzaQwNWAi/xbD4tok7UJDMcT3bR3jQUrUMSQBHM9wSuEwHWY2eVNQdg5mffmkeq9sc+1BmVKlbx
SgVL35sXIKDYr+D3yB8IaiQl8GSouRMC2KMUJOBslU/zcf8VnupCwtQ2qA6sK3TTRLlK+aVStfff
ogjg2pboMjvW/GWw4xfo5V1nanPn8gsMBKr6fvG/f3v/NVcJ/rQ407FmFdUUpmPEkcw1C7va2aBq
tglxYsave2nMIOrKxJSthU6kJwYB+5KoG97ErXm/f7T/nEv/yTLms7VP61ttynI+1AxLSjk1VSnS
iNclpGLYHWBR0X33HKLkDubLZPtg0+jLihMztwkHrW9SZ9+Mii6TFrfAhWQb8k6mVbn1b2PBoKoc
QiUbMo8kkS/S5aNZhPCqfONVQyNvC17sA7LvSzaYKEHbS/g3xQv0vdxeKXDG5DD+EHdWMuOVV577
4HoS/RkzZ328lOm4sHo53KO4dOd+qkF0U3nIDZiJRHkHnuDiQb6UGm1l1uBjKNM8cZJ2kZ1yKR5X
S5MrfJQgkXii2Dy3euztpt/4o7NGLs6Ng9yO5AdUn7bpp67IXRGnBtzaGouDvlpa6rtSOUEKe6RS
RmQ2N3mtwfUgZIue27L6M6r9tCeIv0pZ1BvFCFa/VeIozy/AoZ9FX4jrh9e1C+jWRwgfCDE5zXiE
r8S+b3mnll5LtKxHuvmkaSvCQNQgRj9nPrGKz5HUq4HZtpXxxDtbKastneCkRQSX0NhPaJcAzM4R
xv4d9x55DYeKjzmhLgeFnmPjImepsiCsV3IZ/oloiywoi9P9WxZ16DumYRSc+zASRN5Qr54V0Yie
va24jRYvVbaNVdGB7Qrm40o8dPDxgwpqsJmhUEzIgQahRqV0+R99gKvQtUj08FVbydrFSrvPrDgR
h9PbglSmJqYoEwp8bq8bNthbkSjdz5n+Kmz175IjRKG+yUMQXDjm6rQR1y7ZeCTkeYw/rtO07GIo
Z+wR+KdECt3kJ0x2sn4qfejnbB2Dm3O+ZTqNjV0x5ZfEdYrxhMstUYBt0fjBTy/0L/u0PgjWUtWK
u5s9okpITz8FCvZah9AxToWHvp9MHXyRCz4IGOX3o2ItZa2zLIngjgdlKbt/1ruQnpGIuf8hFc35
Tv/uA3mSCsbVpa28rWvQBEHVNKEG66D3fBR52BoM0j2ymF0NaNw6wgq1zD+9KDOQh5VYeFiGeUj4
0US4q8yHEecyhX3P4PjjixNR/qnvnFQjOKCVrs4aSck2DFUKkgxT+C2txgKyG+WN4tX8fZHFDrLq
IA7rb/rH6oo7rbuWTtLr9OWLHZk12dDL8SyhhpgAMYSDJnHgZ6y5i4ytI2VVMc9R0Vp80pify6su
jGKVJYdxaYEB3ccP6NkxvMYBwnK1NvH9ry0sadDCUDmTQNMsNku8S4x7BZIFSBugVqBHxasZzmsG
29/3k818CTmjBjmT5bgYNy0JVO+ETCs7JHGOOKmUQnuZ28IC2/jJ2MBtKIr2Bo86RG61oo6sXmDn
j7VROjRBr4AbWTGpfJe4OaOX9Z5oxKEOWaVPzii/SDmHavd9PWnXpwgkqRxXPGZ5TUB9Vz2Z6Sun
UQhdPuKCzFwXtl/Fs5/zCiJByz1Nw/H8khE96z/xXmTYK7sdcwb3PnomRtx7eDeSgWEP0JzNvN2p
0C1zRmLnl5+Fl8hygxMWV1cVCQXiUt7X47KO1w6dDCicnAnZollmQEAGoOdE0CRffAp0nv/rxIGH
WBejU4WCbuWWvWqzRuzkBdhS/DE1Uc7p5Q1FP05ZNAFz3NsTqfPVWIw38EqyNU+2SNugJKk96MAS
6FCzjIiuqv9LMmfvZ0m5GLzOrSssOwALMHENxa7tuG9g5B6ptEpnmL+I+zux2HPS9tO2XyyNMmc9
1wifec/U37ItrUyuGhw0E3vEsnpxCzm1WO1Z5A6BEZNRaZ3XtePO5Me+29kwebKjbMP4i95px7Qm
XdaiH1jEqW/jO5qb/JF/eG5vMmgyaPxbocs1hVDKbYp4nxragsvjAlXnU5V+vMwhjcDym2lQ3u18
YrhlSJOrM4FtdMfxnHkxXmW4GWx9ZZfZNyKyFB4yj+I7FEAj9B0VyciP98RjqMU/8ay87A1xtZA9
kL1TYs3NYbE8LVp9cFUAl/Ak784NdHMVVQPhb9qhxI3u17LebAcyOqhtRf+h7E6I2vjP3xTob5Qn
mGI3xkpRdgPGbYKjjlEg3wvF9iXNM5ba+XcDu06UdcOfhk6Py+G8cEkPNJ0gDpchDNAOawR0RxpP
NqN/TnRwM+Vdiru3RAUhG5ymACtp38cLC6OxtVB8dkHxBzptxZn4+J2OGCIGWGYFR+ZZztujZxgQ
Jy+vIjpOMLjmxGiZNxx2WrMhhiNiWdVNzb+vA/2KMRVoGlVovW9rdN0VBwxduqqCqrFsQXZaGqpC
8MqVzWHu3CAlU6DB/hKS3cB6SaxD0KCSimOtK5ZK01kUI/XZZLKzD/HlkihKs4UJ5cjnMIFipTGx
p5TBr0kNhjRPfIGw6dbEJUzenp41c48vifBzG/HEykxGRx0aLK/5J+0u1C0lvFwrsr2bkbfqf1Wm
8VUcSQXfLwTk4sGV0QFhC11sHIhpu90n2B7AaGPjMZndfXng83+IQfmTFzLGAphdQ8jemFrxuBT3
a8LZziVF+czl+qGtMVkRfAU0ZgPuoJA0wZCdZCVWquH/V/zgn5SXi9Y317hIAApO9ps35asV6RQ8
H86g6Pz/y1SxuycHcMpjAuT6gNUKSmeC5Dg8AKQ6eBveEdWT04lHygVi3cD7SIkBcC8XlbIXKfDR
uFnO951KpUhqor1NCti7m4MBTIlS4+oegvCua2y+NVdZXmdAydjECVN8cqFbYDDdoGTzlAupw7pD
gI0jHNGD4z/CfLKSnjNcjKuZbr8AhbWikhunSyCf+pU77FH4ANYa8dTgrEVypLXafqwhWBAVnA0G
0hO+OIzuw/WYgMhqtTDwUdQhTGMbfj05G/YpgoCdLQM+/poSSxnV/wnHfinAb/d3pdlv0pS1dWfI
UTILxKBtp9fM6EhVyGuRmjZOEHEHot4OKev049wQBW4NslXSPXrEvtfZkEd8A0FFQH0rYUgwtvIg
9OQkCGZHxRX6yoFblNxpL5dbSL4eSTQwcjJMpkS25AzNKVHeSkrm8MPpf3HqLJRkqI0PKTMyh8kD
FGBpBGyGiDzviR0goFZfqxCRo+mON6dlhf0Zavd9ZQmRTB2j0AuHQJTkLgDIU14Y2TfdXyWGkd9n
brp8q0JIjpWyMMzi/Bej+3EPTypVxobakca1GCHlFMzkomDIUJhmyJ7JzvKUHsstpaOCpxeDdFxp
n4uCcs9eCgAWL4GJmAD4GSN3KOd+wlr+ARzfqhLAuiRQTpXsnlVfGZtJSUaTYl6UXigoMRwi/M8R
hJDS7N7WruL6xRvK6UNUE4I4DLqJadNUNrwBOnB4+yiUoQjxzS6eZhQiZPbBMQzs3FFASSA2KYGM
in3uPlJLDAfLQK6IB7uU561RrqMCsQtAU/yT9keXj+UcS02WbgLAtlcVfGsuGNa6gb6vEJiLm5jM
cuLgzDi9ZSM3hq7/E06lr4A5GwpWN0yDTwWyUJXFLYi4zLYKW5akd1tugFpf6k91XSgurLeA6JTf
QHvvNdoeNGxJzyiOda9gaoTi0orXmUm1IN9/5Y02hC2PEOVB4ujGfeStIv5aknRZLtCuo8sTJZJr
KLTNZpE/OsVJJqZkeXu4+7MAkNATaPY6a+oCydxWOv9g7ieUTilNGQtH483bQTStSefZ0uFKGIhK
QsqQIoJMm+0XFx5wExyjncAYopnYzqTN7LwNVT9EQzRFpJzR6cPYb+9U6RqnEOSj4ISNjBTRFmNx
p/yuWmeARzEA6p7DuolbOAYTzF1Q8bYJr/PJpi6csTfkYRvW3SIsRjp3z0+Ip/8KDJjRJoOeZrsN
20F/PgteixJVS4qNkqvQ/5eoiTfszATnZfSREFotcr84NA8NF2OQZlSebwqQpqxBLcRWm2yyU/VY
n2A/kVQwgmjmab3zfCuPoeQVV4M9R7z7jtGyffjiAXnbpcMSeLd1CsNKQoaXZ/LQbBgatPT3PLAu
ipMKE3+phjgsx/MM0tI/XXDrJmRHNOtSHiWkAAYcymA24i4YMKEkRdeIgyo4zYjwBfB5N2lRj8/S
HrF/tT6e6oSzdA31tFpBwzzFm+WDeHfyIrgRLVc9H4Q/b8l3x+OJ0FCrvHypFtDaDj8zkJQT81Vp
cbNfOUgqhT8BQbCL6lOY9SSnWxocifb9LTu5CdQlbR3auaNb3JqLvO01V/v/Ku01V+I5KE2Wkmn+
wf69EOEzhBYssn9NUdjq3gGGkryDRzX+nYFzB7WfKI3oZKHyLT4KdTXsS1WcuTzZbcVXXal1f5fb
6SZqS+cnoXEOr2HolPT0cjDPaM4gNXoNY3C5s1uwW5O42mS/c9U6dUcFwZruHHBXdqOAZ3cPuSd0
TWXbpYt7SdXeD50ENve6CYy6tImGRL/Knn9qwLo+vMUrbLZKjsyAdXh3teODVHv58YLWRTxyRQ0H
w60Os7jihLm3aEqIDATiW7mtj5QTkXl8UtzLwrmG1trPqynEWD6JlKRdEWbY6CPfNK0io61NAki2
D7HdfEJUyA6n6BZ8BDzDpAjAmmiq9T4PDDCj4dC7DCPOWt5NsiPn7BpNFHpkF4vYILyn2d+WDfX7
6XxVRjFiHSAxRXZNVQnDT+KAeDejx+SvsO8nuSC/v9pim3i/gQLaIhDz7Xv3i7BsZxbhixwDgfl/
MXjWHbOCxL0E+HtiMkQhfr+UlccPahMWOPiASb8TJLbTlqveNjiveRZUons243tn4rScP9WalHb4
EB8O/VF8o6Ns9xhLT5GllltoX1LD3KZInnB3cL2N8sdzV8xU0Am+bf0lR1cvpICfV1/GQ7h/uvwE
Uj4HggUiBEt5UmZrT0DoywIcildhTMX0PgF+5+yBZQ9+B3fWZMra27httoWOu1tW5e/41iz9Ytwq
N2OUxPbc9tVLTnsIWJRf3t5rB9Isr/ioefjg5Kdm/kc6WkeF29mACQ+us2qiPbZZ5l5iXXXEazAt
T26K8t/7q2Zr34QrtfbaGNBmnZ/TzXUWRUEUyRm31SN4HwzI36e8B+BJntbqZSvUB0xXAP+Ks6pg
+GmVQXbuwbv+MliRLsS/cY6fxLirdfzI3DJZQLMS/vw906zcuFEO2tQ3Mzwsi//ZJp/Bf794znaV
pArLqbAk/LGUvP78FjAlxBCoiG2OMBQ5a2u8soCVwLnEQY9m62erRZD2pyPR0jHCT/ZJ/9cUOhpW
V5BAJiBFgJz7GZMhy5VpvZHh09eatFQH9Qqefq5IfvjQRYbezJQ79fZXIHA3YfGN4U3mcrkVFjP0
xzYHdJgBXGyJ/5bSDn9lf6gECEraOpTmed+u34OL66QzPvr3Fb9fRG51UJe7ykAdn61jH+7+NsVa
3sQYFbs5mzELLNHKDJNzxH1Puhg8OVS15xwUccX5wmw2SNocBGPiAllIKZgzo4kq688jXCk2eTDY
MukiomAgfl3TjqkXKY269HtacdKPC6x2VKGgDPuXUhimfqyx4kfIexLMg5TV59PKzEEM/nzxDXwf
Iz8xggJwThLm6IMAF9KqbpYaciEaZFsklD+J3iyQmLOWI6Sw33M1WEeZGmonKzF+ax8XQ+3AgXzO
O2YL1VISpIcvAQnmMVpcMpDNKQNMMp68DFpQvmB7jMyF+VWdoKXsN4hnUBHbmC13rNI+DHxx7kQB
DjGrg49ZVADwUj7NgIX2Y98AfctkyoAAv00FDBNNVDFBqieVDBt7U9t91aZyiWDokLiU4acRE2jR
FBDwCfDomFQCXG16ScBifW2YhObFmz7gRloH3Pp0/Z6yPiXXAZa7Utuoi3I7Rk/P09B7/KOn0Bb+
s2IK8GInCALJRfr2L5vNeMmsXAnORnCdy6ejSl4dVkOiWczFdLqoMDyp+H5JeW573gMZzUn8fpWn
RpM+24RrRKVcBzfEJHlvchnbCOitFR7KND4NK+BzslrOZ+Enu4j75zxD3B+A4tuQxHJZL9gOkulJ
WNv44SC3brl050qYV7ZhqFIbNeHPmp/28NgGvAvBp9wSzNoQh2ysR9CyLj+9BFUR8p1mi55x2h5g
cZSKXUrE67wo5Z4CcZLKF0rmsjXoq5656R5oyMTDaxft/1GfIce/1wIm/c7E5bevFtp1JWCyGGA8
oTAP0bEkHtVLNHY+3K7Fw7oZhdZq9lUGmEXQGiHl+bSc0ERJWOPKVgHh/lAjeDxom5UnWeARSxYa
HbOxP4P6sTAIMracfII981ng0j3P/ApBThtPygrYLDglub4u5EGwfpK037fu6rY07CnCxdAzCHMS
pevM6vzt/VB3bpbEXZHpthnlzkYqPfQMnfHb2rpCic6o5q0bm3cJag8vGIUHPk2TvN6VQI1fWqGI
7Przj4gXt/rHR9UwWPTUE77NGxkamMFf2DCifGkgZUPWX5bFfryC6AUD0qM8DDxiw5MCeYrE+Yb/
qdJr4gwh/rfEbUdDRUJlaXFIZCdaiiufrWll7RdQJP8LHF2Z9wB/Rf5CHJv9Q0UJFe0idwU0FFcn
yJaWH3vdjAS0sn9hN1UV7IBMEYqY1qQ09Qf1nBQQeCcDcMU6JHrHKIxDrOkaNRas6D2N45WJloZM
O1Db4W3RuuRMdfc34YPe7Es3rVSCCrIEVN7adYbMKccXXk+lRH19BYqC+u7oWe/NhihKbvIN9yhv
RmObVor8aYbrYHJJijjXAyJjlgGnyhVQqGl310zqjVxoMqi61VfWW9NvFrj8iq27JGFG91Ij1PDP
wQy2XffAL1aGSHcOgFkLHhmk+FkP8F0RVY3gQSxdksumhKRdIdTiUvh6Bbx9IvZRRoQkmPys+4bD
H5ZTQ0TCelaFOfpAHI7g+8tSrClZih8yun4qz5vWJGp3nI7hKcflkTF0w0LH/A7GGBUVrQrs/AqR
n7MYJeqMS1GArTOjz82BThduoFFxF1hlWjDDM+dRe8vNIvzukkpQ2pnBaqUfP1Xv/oRI56i/0k2A
5cuChAaHg9CLvfqfUkoyUjO3DeJTcDCPz6SqMQYBcQqSEZXNTlL2/QHa+UmJOODIbpXdA5pQ7Gnx
5Wxroe9QozZTfmBQEuKrda8elk68sNUGsgm9IKzyQqkiue/AjdrFs0pDfXETEJMHA+SDC0KaynLP
nrQtihUxPHDWeEgINbccZ5hDql8yEgthI/gZXBXutDolpZhUylCGOg+Tp15XpVTs7MWEepDz83qO
3yN58x5C7Njxg3l0BIevZtPsNkYFIKCRyURgLXhcuA5CJfWblax2cS/43X2q1uF67hO1hJgvEqQc
8Jr7Xi1ge0sZ1aorBAz/9ZhR/++Qt9WDYVFraTyqqUEt53j734HI8uUUoyRLQpe/wPj4JCcsDSYd
0KXphl2DEfwQO+ts3myiQ6USMa8EURFGXVKqMQDUJfWVD67HOX6roIcsMuzywqPFWZQMAIBgK5dl
o9vxmtEFi91LCwv+tY1JW9g1v940hhd/3HizxZ+G6OUw2jOByjG2oDvR+e0WlxqAEqmh3QQiWDOK
ndPTKQCjX6H+SsPQZBfakydqK97P2n73hH00sh6fdtJ8BqWQDJ0xbmCHGmwEGwlmERNK7Z+qSGuM
wz8EEPmsHLIIbcJ26531cS9N5zh9icDwgBRV+IaZ4eTj1YP7XwZHuaVcWLbl/iyGO4MmWh2BXlhJ
OYBUflJYA5a47HviFZcu6NXZd8Yo6W1t9hlFk7nWin3/B8Ycd2i9laOE8Im5/w7nlB3tPlRQ1GSB
xDjX8PGHqnTilFhezAw4uM1IdvPfFZB9TmQuzk2LK+G86QIiQ6f07DwPVEVrfRSGtoNxYutTptbe
C7biwEhoQDTH18VUYyJLlpUzVJGfm/gsj/uu0UtXF38Og7TLDwDt2C/jEbhXTzFo9PRS680ypByJ
ESnxqWriY8Sj8bFTRGWvMFD05H4+xK3BQG5GkiCEUsEDLh1lRpVzGEYGTPO2uSL22rfYc7cOebas
wKRHKQnNEX8h8Q5qJUZ9PGh9skqUdm4LhWFBekuf1PKkrlIu5VjL1raEt6YHc54owfDsyZr/dSSK
RUA6z39FUOgAyyQxedurJVHyMQA40E3gJYPbkxPw7hWCX5ux5ivVH/ZFIwIVLQIQHO9VKjEeWwFO
AwLnP8inX2YLFekHHbn58e1jedSqkRlDBXu7aIzCFc+6Rmtk7uJ168MtqklvDYY68aC+NGV8AAsx
UYzWrBI7pI8w/mVSb1PJ6QcNXY8LVcJ4zJatCWq3sQkwUHOjnslTzDbWLZhHIDikteM9W5gKP0h3
C2dIQ8xwESj85rV0yIICkqaS7NjBV8GvdVO7D4CLRKFkW/i6ajvgdYPWIulaxAI7gcpzXnLx+Gm7
al2DfW8GIap819vhB6ktHeqhX2gMjmAG6MNTi60/SI++dCJM/IoFWMDXDUewUD8a9JSvmWSyEz1C
6hs+7U3xsTXHt51LkMGrLEYZxdnOHfGIoMW1AWPMrZauYuhQV5r3THo45uUeMewP7KQ+jDv/2cOb
IK5nvVD8UHBfl015ahthWJTfs4tQvLWIgeaCed8J/DuQysSIcCse6exIAiV3asXbIYwEM233qVP1
6P5Lyk7M5KbcKuL+LiPlnRUDAfpR8RaUyXwOMPwZjwB9KlJQBEPxcXasQpcZHoAbUVgky9egOiPx
fMWGPnUX5aX9HT/RkNE8m5jSgBThlc1/HEhO368MCHcE8b60gHua5A0q2biOfTvreFet0XgGEUUL
pgtbjH3IVbxzJ4GoJgP7OYo3yHYv8e+ITeuiDQBHOSgBoaD7qy16+uCc426vSB9oJI8xSN5EHfcf
+OT313r+P18FdbMYkuyQvkFQAQ1DmmaeCvCEb+vRek8lQzs+wbx2d25axPbQUOzRvSRvKjZ3cNAR
s7mN61sggycOOJT/m8sodfaST+LfOfz2wD5X+mOySoaBaCKHbdli5aRaat8/GyNN4yj//yysEG17
1fotvZ/QEtacFCZ65h0NnCEMbrJuPrpSrmMditVr3A7TJSL1oqrK9Ke7Kp/nsyJEMylau/gkpPZu
jFKXnICl+dpUS4gfXyVE7sLDAtUcNDijKOsXxV7a68YZbRSYVxuZ2nSKLN2BZhI6Gl6MaSWpKQd/
rrIV3hwtp2tdkd0TmgA0sMiGDvZ+FZaQl8CxQd+cA+YV2bcYeDCMi0Q8Z0Y8NfJci7kmHodLD3MS
z1aipPgyBVwq8d5AlqH7hFoMCg9P+hJT5dNKIvez+LoxujzDLAJIqpliKWev5nfU24K+qrZlGIhi
+nfm/LXbQBUD95EELb36sWA+w0U7gKRG5uH/SyM+SIhVDVgN6qtOGVBsAJ+Psb5hu5CCYCfiYE5r
1hNRkRKIHKqlcb1wGk/5zFHKwmQMPXqA+1p9FHssEAT5ZI06sQZAXrN6Oyno7D8AAtKddFoEriJL
jG0N/TaUecmYSleIKi91Q5noEKS7s3Kazul53M9v1qkKNaWweYuwsts6lhpn2DSEK4xk5G4K5wN4
ikDh6UUprDq+D6nCloNV9xNcCDOHZJdrDbVUT10+tj4SqgzpeE5llh7APsz4WJlUVfr1t9LHhT0G
IwjytEP6Ojp6o38yVVMG92ssHVGeZ8jujbHbZt46r3WJXKMw045lYtNDDWpcYxQ5a029Yq+wXCL4
m45rW28sIbZu0s1PvxijE7rKosy8O/+L6fxVmMVHTveKlBjEDcnIndJ0s8fcw+EqQY9Vj9pKF1ES
pXPEEUh2Dk1AZtGWLVQ24czDsG3QIW8F1fcvmuKt5l71yZbOQypPU17kI3pOvJVd2VXu6Mcn/qpx
gZCIOa8Yq9nX22SBObfpcHmAHljcc9eG+BdPl//ti+NcmcP5boO/PDdaDX6VJoT07GBksaEgkkG2
OFnHR+Xz88cuPckSd7vcDvqizNRJbrGjpqC04XSitfiiloKKWDk9+9YHn6Q8qEqD7HHY0Np/cPXI
6JGt54omaSQqvKwIqk0W1ocpbX9js1bAox/jo1tDcrhkVyImk2B5/4wcIgTQqHeWpAOUUmoVxLg+
GE9qL4XUwc0IWfvfOWRJ5HL26mg9tX3xzqk9hO6hxCsStEd7B09zPMYhd36V9H+vvepskaTfTaF9
0nlbDa7I8FSwNclkhBfv1Ki2YBGVqOWqqFvBXKpG0pdboYcSwZlRehxMigCmZ5gDNi+nz2Zn+CRp
F9gzKanpDupNWpePY74yor4M9zctT6Bi5+ChU4E0y/KXjtglbbeLMEN+v7LvT13bmd2KF2d0rDZp
xNf3Ugec3ybDLqGH0f0hI7Q9w65+K3wK65Q5S8HM53DGnEq1rE0Q9TXmAzz8AX4A/JT5HJDJYKJc
xO2rbawCRIeOGJCjyzeomd/LYIYo4a2kwntCmIRQCA5ACmViap0nUnx6WvaG6UoyE4rqAfRTIZZQ
OJ1seqNCi+fkESOJrNcBC/Ku8kiIAmqxr6f/u+95upPgzcdxkZPtjTJT9dTWH2iGFiGCc+yA8vEy
bFPD2rJUEbTRwx0W5UMfbSEi6bMeBWys7Zg3Od8yBKkeZpu3biMf5VnVj0r1QPgugjHYXWylk3u8
imF1VotpbP9itro3rCX5a69t4xIFn+uLUYgXaw9U1fpU3u23c/WjpDjJvh0FxCbXQ23WsWzMrxC8
uuyIHgl77tTU/VGCOxwrfkxiIT9Se9KxZkuZcVErwhkZzL15/H5/CwkbIcuGTV+VzhvuDrh3pVps
9zj2/sPQcJk9XmOeWnCsSBrIzTtnyGf7xWGxNDQnAy5htlTUbzepnIamPqtMZl5Pp2aIeBMtVqMQ
4sQECRUgziETu5fgpspM4AnS9IHtWHO+Z/C9/+SS5uhpH4y9LrugYpuZ28/RDQFfUbJAsd7kFxiL
+mRhK0kvH6xtuShX3349QzTEJy01lFFLFM3qFOJYAegN5Pef9ysY+trXSjF+U/mBsMxjxHRa0yaj
s90znL1XPEXeiKYOLh1QmFAKDpNT0DQFDHcgn9yUf/9GxjMn1lcQaB8hK1JEQC3bchElRAKbsNbq
PPoPufusbVrIZAqGOaGT5OgaEwAbXVwYF5hpaiTJ8IE7a8IiaIZrjO3H7Jid6p2T5TLDKBs+fQ4a
dsfi64D7qaNOBx26r/FACrVKt7KlNGOrbEL/aYpYOFlWiVNrhJDdxBf9A16xuW17K5+88dYFebt+
KlPm3AZbItzTjbfMQ3J3+G+O+iReYrNN9JYCe8+hkyxfNHQuRNYCKovpAFLriVkjG23iJrZcj5U4
bkj9RyPEl9uS5Eug5zYGHviFi8BXQKK5I/d6GTq7ZGfsj+FS+3Em9JDozdHMmIlEcmTCtCqRiC6P
McAfhcmGJn3Qu2okpmPXlnmI9hhN0hb9p8BBW7U1WqkBapgTWToY+jBvvAfUcSzkQLJDLfTjeH+u
ifBg1W1iJn0YEXVPtoTMZhQaXZUGSR78dtvlIMAjxOv2nMZgrukgWXq/UbvWCJ3dqk7K9Z2W4xt4
GEp/RSa8rESrDjbB7rlUjBPo8wy8PuwCoZdJfhlAi4So7krR8BcnQmpu2EEZ+YXtlTVryo3JMkeS
s6anYdpm2+LPs7azI5QHxVzcGvbLKyuNd9HyoBR0Aga+dZMyUuXZYJhNpGMGWoLhsV38Ke2QUuur
Be3QxUrzT+M4FGqM6LzHaUhUW5BaaLJvCsqcmrwnxywSZUgZjzZlHS21gAAXfQ34lK3rRKo3+kf5
jSQnEbW5Yp7/mBOg7NNEhYBFQYeAqT5xo591QFBZ9P2Zj9Dixqkidpu+0JAr5HCLPAFXTWIwkm9v
YLyeQ0K4+iB5mEeBcBMIak13qy2n91gPK2x7aVYODQupswtjIwXA35TgQYkd+xjjw7gBoPIMhXqx
QrRSgl2DhHbmSNds8DTt2uE0DiZskNI3MUixnEwPMW2WBQ5XB63h7dTWcxyhpwZ8P8/Tvcy/PAXX
f0K4i4IR4b6iyJQHjbGKQ0Njgh+3EYYyq37hotcDlMqbO4rdgOd62ODpzQnXreJvjfyQnY1JilSy
6lI5+pryrPy7SK9Nee4uUtZmm6zPmDWnofPIaN9Xi0WgPcLinuwrImfqbr1xq9vjf8Vn30QUW0Ij
QJK0W5iCN+fe0xn3ZvxzH0r+d0po9pWvQVmZHFY6OuBXOlvkntRUL9hrtJk6zxO7T4a6DO3Aj1P8
PsdJBojuSAKqSW370+NId/1vMtbCYDZHrIM5VhPlunBF+1XOL4oXYNDZV1WEev488XzWom/T34VG
xMjrLE/MA4LmBEL4ASAJ0/2J9sMmjxnhTneVfvBJSyJdmL5JTutPDx4cEH9TZooCzFkCS9Uixzl5
UMHWttiXok/bltLIGavFLmm6PMhvyw/n7knxegBBQ/9z1StIrkjdStL5bZCJ9is8i8WmdYxGPSrI
gpJxYYydCecaFeOquG8KYCmwsZEB3fveQJGruGxbLPT4n5Z2mBdJzR53HVSV365UdcSA2mEhqXla
GAms+onoh01mjFHZXz2Y+qHNG0onbKko+BCFfc151/mUyKJre4MFGFc2j3zlxno1MoCpe0m7nrBo
dlPZuClHoc5POkqIjexIYgFE5nhfsXkyrVoYeFUtlZYt89r3/bOYJ19eJh/3+Nn1Kz/9DgzaCHip
tY1kBYthFRQK1k0h4MJdOe2uUNCoOcModJk9ZmXMI7i9SRWGXRWi7U2Epf+y3oirHwjo5sugpmVa
13d9C242WewN8M3+nQugpf8Hiisifm/hEGX/u7CH9ML82jnfh/PqYF4lJQ7bzIS2E+Gn+Ld2LZ6L
JyDPdiftUCvtaXVNOPSanVausvuVbncyq6j0uIi/lbptQE28fGH8HufISMU8Bzfig3fep14K+iu4
UDalOz+xbQCuTEevzohRCABZ07/Qv097Wkaamy/Zy7j24rrWaJT6tRgEuDSIbsrVMpZ256jrFhQO
NtHuFFQpzWx7ZTL1aTFsJizO4K51NXWzT3zk06xCrBcXQg3FXe4t9yTAIzHvOceqe82/CTbnNDgR
FEwO997530k2+qM1oVoI60ep+xVxBjepVsPwfa7QcejF70Pe8S1lk7byBS8Cu+XRddNyBAs54Cd3
MRArFPqCawIddEOlZ2MJKjj0MhhvCetWqdlxooiyEaq6EcMr8NegnIGUaeYSgPY6vjMyK6LONgIg
ha8pVQTk9tQPLBrOictRRllktLCl/YwyEjtS96jneXM0ayAc24waZEMFHPM/0Sm0hoI0wnyU9jpK
LgngEDShjjsgJJR0JsZ1GHeiVqf+tfppqZ3UbildjlCB08BsrePgtMjHQYURqCMBAQkXURTk2mYC
pdBpIFuEEBjh75sZyah+iIu1KgWeb2ixFFn1hgM+2BsBQDe0JzLT30f6sDCPVXOZiP1ifsjhbC84
Z70DprX1dkNo/0S/IsJmtXQ7Hbg82tn65aAMfWRhuKx4SeqPqJaCjKlTFR/8bc452cmRhML68wEi
o0NaRizJx0p7cK1lnFXIK9U8R61N3/WpPjCxWyxrHQx6RZPpFadqTIDSjROzFWOmzuVX1pzV1hDK
SSmZo5O59QbzkETXWVqNf4mVnPek5XH30AqXKqAWB9sO+kXjqcsF55kdgcs1shgNfDCT0LzuTzug
/C8eBbIh83bEguwN51XuilPuAMJi7B1c5vh7QW26AvfFM0sp9BhDfHI3+cxbHx21CXWz4beaSVgo
CftvxAByYT9D1i0sm5oXZbK+y7mwkeODn9lwYfjn8goL1qiwagqTz0v/0AXEW+F7U5LvPZZlazKF
1600BHIX+vDRRWZjAHkAZxroY34An1azxM1bGieXW0VTiSo2mpmFDXZR5YF0O68mZaXMsuCWNIIQ
TcWn5hthBAufOr+/VWc39QwxpAyw0xzTh9b3pFjsKWzgOsP2tP+EkIFkTQIh3NErNoxtz9dQFddR
yDlRFZ/yEy2ZKrJ0iZ/aWyd77zxw3RPFyIoO1aANK4k9DG3AGhcWDKERzJVOPeFiZjpPiWEg0cl4
NNjnGC+G0juyGMpK6QLAX20vtx27G9Bs4I64g0m9Jv0H4lsxTFjrhaM7GGRMEa1Du4cgn+5R9ya+
fRlbXXI6GsS0tmYBwsDEgZyA0Vk/HrIox3ux9OMFhbFZ7YGi8uL0NuQCNyvxEbaOCxDapSPfGtpc
NWXk0bGsMIVFv5r0+3FF6bEE2UjPiLeO1EO8X36arIefqOVNgHOf5LiJIZjAt9mrusqMOqCPyeAX
V2IKAdY0Mh4WDt2AUc2guBfuSmKak9cIvgKGVHMUTntF8Oabe9UxYl1KMcQD7yCJY0qE14WsqLXX
XCbnlL73Yqz5O4OGjVXFywyV9M1/gQ4cXCtHcg9RbXCyNCFn2gVIBiiBbmrLGdt+FhBDWeIvx8eI
DKG7XX4hNP/Lzj1tsHsrZUMoEeCU+B2GTRZCr20uYI/GJNmATuFFvBE+dsaW5LIGAKAQD7tRHEkm
yZcDzNHed/CKm5eYx+LXHMv2N+xrtJSCi+/HAyN4TZGzYyA8qOKuhig5YKk8qxWpjVh11NhbbGq+
2Llw4nt3A2jr/5DkJYrxvocIvTNwmE3bC2aG2023vTtdNFqc0odhKtEslJangdvQ/k9fJOQpRbvB
Tu6rXNtzupMFxoZHjGq0X+YekXY4EjnHk7gMjnTTasVeONGLsML/GDymnSoZCG52KNKBsulcJQd4
1z4sTmGkRhFOLkb+5KVIS3vjIsa3k+ns3y5PA6zcRfe+vKRaR7MpIOGXhjazhb7ZQ0Jt2sxvF0yF
itwNsWvCgTjkL77waAhEAFsUSrQu7msy0UL++T5a07UzE2gyMmRWoXLG6x4CZkZ7i2jl/5Fnpxno
aza6BdQNgujzTmi9V8tsa1rtzElBdcJdPHRRdJzdMsEf8mNs6zfbRk9S9aM1M+QqlP00IE+ZSIdU
Sd3ZhVg6bTgykUjDTQMD6rYdvmtX6snGcZgGXB4IynQfTJ7yKE6ryFcM1N/cRiOBCFycLBCLl/y9
rWB8EFY+18eRLcy4YnT+3Rg0pSYye6zI3cAjE0+1MOxck8AAdInQ2fkot8az9KGGIFitfknwJhPv
gPcNRSopWStiNt0+W/0TvaVIlQATOJooq13xdsMhRhmEJo3Do1055P04Gvbf1Q+5gDLsFTjMghi4
RSuDXylldrTBJ3tGjMAa4MIZGbQxVq1WPHCZY21kTUzQWzqg4C/nutLa6lp3YJWrrL0dMLJGkpG9
+gBwq23d2She3osLuDCHmJfPyhzlF46bptIj+Y5s5665V0ZhTtTGkIePMZymsm45c9fZegcDWjTz
mCIfjoe5p1l8Z7yygUwXYwim24Qd0bk1vvgsq0feIF8o0ZNbI5pDOgghsGcjYlq87d7gQ4Ho4Cda
vgJvHuY5gnKe86OliWbOX7WIe6eUbs+uIFFGPCufIicIgVYfwyBH9j3wImtN571rd/g6J76oREQM
swE9ALvJbqId1H4zEzpLaQVRWgGO+PMcb2q+u6NdKOn9EaONX0Vn0f5Ry+UVceQT6HRG6xePtSPl
WxQL6Egw2HG211JrnI4/EslOMTyQDqEqrmUYHNW3m02vYqSN77gnLHDjT4DxW4YbJ5gBbvSQv/zJ
J/+xwMf9TbP1FjQrwm4OWwdfPPRlIXc4N/IOOCoDA/nMr+6pAlk+r8uf/QKkWxHwqlcnQxUtQbG1
Sqtd5EGLv80pDhTPPnLqFtqHF3TsUCbgBDemUPoDouUvS6Ta4bC8YJZQl6CTIenDC9oYCcpFu0Tp
b4m3QshRotZeIqc/6ZO6lgo2V8UC5lrn2HSJtjBcoZxIPPoRtsh2iE1W+xWq3fuQA02/tKzwVIXN
wpjGgSPI4/mFXyf5XTin6wyCu5l4KGGwFMNwIWoq6bcNxYpjNDTTymse+RvDn6rEYPnzwJmTFGe2
Q4+NcuEu7alFcTEr2QuxZUbBs2WPg1e6azPmakPBK1rniQRvNWF0Du3A9LWyk3wA1AzxccNg4HeG
tuaSwJDrEHLcLm+EjruOX9PYG+cVNSYXcvGbDoMrJa8tp4Cxt3faaIgVhzCNZQbNRsg8XUqUiymL
gYuBnVxdUYYdl4bWoCMpCDoH0ce1LPiu9sokDwOCX/KnBh6Dd1aJEdySjsh+cf/gD/rDQKyZ/S1G
JFdBeO18K419j66UwBeHUMxbSF9dNXYuwIZyJqFbjJBjBAWO345S+nuMkA4t9v8HlfDaS3tdetUX
AHz7oYIzGiiLv/ZDpJWJZDUbGQSd8iIR0ZiVzrMNCuxmFcreBP4ePnximogfWXxRPXKioRltnU4R
SjeAmYXtj/7zHx2CKG4KafJ9sJPmNQtaqDZLSnzgt0p1iTKFSYG2p5a63fe6TEt2diYzrS9AJM4B
bC0wvBbYO17cYTxTjz7462bnBE+Ck4ldCvvhkGHlwaTTgEc0lAW/W958Qr3alPBts3uM/MUkHhmy
t7tTxR5OO0ZdKnL2E56isNvofjJOuKqMYAXUEgo5xhYWpPElYONjEP7n0pdBcdOJPeg/D+6ZuyjO
A2STMvmorOZcVrpscYZXyTWYpEMXWXaOPZa+EYkvRTc/3B6A2cLCmS8ZUUvE/xkviFfQxmkp9pqQ
pGbH44VqgbatGd5BYh4+7xuSHdHLYuaQFAb1AJ31BtDEKet3Gbei0fr+kBKrtBZaIAmj3xTJ3V64
0PVqG4jKwDnYaZSVNhwE/23dBkbK5UbcFICfhRs38SrVYFhIBw1p+4FuJL5SaFTkrl37qG1jppWP
EvBbMDUkfVZa6M8nUBc/Y9yP+eR5nE2VA8/SrEcdK0Fa0clL4Xo+imLtWabPWCauv9n/u4dMIbzl
IQhs9IUKU0In/ssgmF0oZJJzeiOL4BB27S0uaMakDSdR3656Bod0WIIPWoe2IqTWbziQOWf/BMEp
9u0+H9rIPaA23tW3YO5gYd05Zc9Q/0mArkpNWEhmPGJB5L04pS2bnBZQIGFkTyyYR5B9wSpbEvue
YiuzefoZomcUQ7a6G7xUctgDMCuHpDTIjdSJjwSEJfS1ScigA4275tLLo0VLZDKbdj8XUQlbz9Yt
gKb50q0j+2JAY9bhU3wc2nDBqIHFBgby/2S34Yse1SLMPKXu+OU9kBmq6YGmrrzQyrCrswtosNsc
SmlvQ9xMJWmlJmOI69t0WbKtbPrZ/YmvifMOZo7yfPKZxAMNxT/jWcOFQaUUQKCxa7yd6KYl2TGB
gR2ZpNL2kLjHjWf9vX3u0uMMVVyWOVK/UDbZ56ZZDovWAgxpwFoKraGhaWa6d89r11ci/RorXNZy
Z6AM/n0UaX21jGdHnbhsXmQ0nJ1oxHmknr0mqWFFo2yRSVomDiekWsnXY9eNqVv3W9gnT7WdiFNb
1mOQmUD6jUJkic7VhhYtP5UhAK4sVyDrw+E04pFtL8L24RUBsTyxSeL3eLcBTDIvSL5o/AVh5eNT
et6f8ZCfIxcdS6hGEIfcZ/l666oKyz/o8FWuBsxYs10cYdr8Oykef2UoR7VRR2scVxCyZjennfWl
TRWQrn/eBMGZmjfhxFUccpamOo/rWQg/0afxhj+2KXLunHZbCHngbtdxx/sI5BLUat7IZ7C0nXr8
tvxRHcWDug3EiFhpTaopr+n1ii6R7MRmjMpmt+GQhtZ4HVvbyGB4pWkvTjefdakfco+Io6+HjVJn
y2X5GQ+XOKWRpTsIrmQHNUH55S0gpNtkRu+XxaRRUG7388ZP+qQNOexdqfedflN8A+IjQVFJaj2p
kH12fg365lmafBXQU2SFwyr8gMX+Q9s6EDP2U3+o8bYAuRoaewpCKVlkJzVHYVDF2Ru6E64Jz8zk
sN+TrisgJI2GhgefRKHZmWmT7VjVfiP55SE+MH1ltwj92MNOom9u6mum3RHRiqskJFP1zln7B7NZ
uUdnzspnmoTsTaFo+hyC+toJaV5o7wmA5GFHQnTffpVEYRfUOHDvcl7Na+mqfbxbbg0CPYnoVTCP
eyvuegSCIk3ABE7cZwW+WzMM9BWC2beiRaqkTZeXBDTdmqOALLUWcLBuTX65FE1YGittCvDIprVo
1tjXwecAUALayE4NCHRbqOUuMcmexg4ne9Bv65pToYJlgXgf8yPwmatz5z/j2rSU9L5BaU0CZSh+
QODMdPootCB+YQTdVTshlkE6TzwM60Qm98E1hF9U4ZrZGYN+nIfIqYwvZ3qB3EE4/gOLLfvBm+b6
2ZdSI5cnzOdk9BqEJNNrrOwTDocu28VevRdz+/uQTcWkMJRkjN/+i36ty0xY6DEfBXDh+nm9kwmw
n+46DrfXb/pl9ni07v/aZrvyk+OeBx9rXgz6Pzei1X0/dRwLQvcS/LjV7x7MFp9TON5PHpwHUn9R
Yjtiw/8/cEGdsC0JqPKFNJotHF/UxTpUKndEUqwxGLp4YmSxuCRWO/Fhq2J+QfaRHOnScBLoM2/7
vSAkhIFfapa8rDja3rpKqbV40YSK2Ac5TiYmVAoE9r3XB+hDZP6dcp6lgyqNgM2QIwrrLCAcFphP
EgCWvFhje4+EwqsYJtME9+5eC0OrvPhiL8mDE5mdDpyHy7flB8un5YiXS8AHxPFd+/bbGWBGIkA5
KJVRLCQzwK3LCldG0Q5st2tdQuXpczgFXOm1FQPp8t2fBZT9jov2UXmGxJFfupsDYe/PeYUHrXmB
7bfxQelNI/DayCtZfSc6HfVJ+Jo6KYy0VgdYjKXwGDctE3QkhBg6+Zkvvyktf/Efp0HwWHLB/XR3
eMhVcpAq8vX9rOxvWpZzqWQZjlkqDLsnKrk8t+64g9egZrvWv63V7sU1UjGlH9vw9WG/bUMJgHJ+
kmaIBD/E0+KAhqpRKQnPAmhGpl5TDIEe4yzXBtdcLOSRJUBGdVibwk1spdqE2zkJewJQjKfAaKvb
vLnh3wggkSwLGKLyKcPbHS+s7Wa0NfbQYtXRlNQou+yI7B+6TKoOWDBAwEkerHOH/5OcieIvDXjr
ureEWhsUY/mi9BmhZvY41iL8h6o+4Id2RMvgn9VuGpjQja2VXwAZLg6HOB2FYbVnFEZL3nfQLOUX
TOJqUb68eNVau4lXtxFehXS6ZF1zg7tfJi7Rubpp0ZGxGl8+tu0vCMG3wMIK7ru98kZhmB+iCLwO
R32cowmZ7zi5+Jw4ZogUjzt8SjUzsZlM8biLOjdPdhZ6PIj1JkdfqyUnvyPggjdgL3MSPRwQ7P/Q
m8zyUq6CbliQJapJ4W0RA46f7qdU6vmRUx1vXrekwaNaXnO375M+sYKtfk7RT0ZzGwox87KJpPht
0Z26N6+BaT8BVIv/jDu9fESEWKdMjh6r377iDiMVBDqhVNR0DJnwMmBSI5cZddb+ChzRVS2PpzoX
oMy8vy27epwuQA6wYeCKn5WBXwh85fv7/Ufat6Uul0yWCreGxzKKwDzyIdpenaQccvO4Wn1iow7G
vaTHU8hC45cbMY5sjTwnuygtGqODsM+Jkq0S+/szKaOHrGuVOxQrDXPF6aswmnIzrVjmKtQ8tJIH
A0TZW+OLsP936uqRgC5c3UjHKE6I05UNcObY4hR3CXRyu/VGYdYs2t8k3MmsGH4hgJIVnf3uH/9r
jMJ2Leq7VBrpkdbA+u/JsMaxDha44MMc5DIYDFdEBuASQi+gKkcg9YXybukCt34Zq2drrbgwzZiU
BYiRj47WPcECJBPK8qoZdbnrI8T/6LRkadBjKb3kDtlG6r9CoVlwWWOaezKfcovJWNXUR2YvLtzt
EmLa2jIEt9vO5kz4oTmZvzbqeUuJvttpAPGtCqtBAtP8TvVtQnrEmx5rAA74qD4kzRaQ79dvUpNj
RdQxJ+GU2ZTv5BxAqMKT4LOZ7RszKoDC7HtAgq7DWMN9WnQc04ayi7DqoC31sK8bN3n3831rwn6U
9Ei5v74Relex9mtQMmMZruxuVpiPnkyM2xY6UHfq31piMW8m430CZFOBcHbmp614BU6WdlmR6vog
BBkTagxqCboeR292R0c/DjOFEJdJUBxgjpisHMB3/eN5z10Orax8+fx0xwCHN/rkOt//RAXO9FC5
kxhIPi4LnhM/XaGUuWNdF7SWa7a1YPcgc4bqP+KbdnCzlNsdZ6aFxQP7ZtQU07XH6Gg1QrqGSsiG
cyuOcwnvwsqFJ7OVBBNB2aiTuaoSvHuZYHoTGbNJC9uyV3oHWFlLVtQ+j+IAtESF6yNNuYnkMwuB
B0ChSXE6yFUTJ5La7D6DAH7KX1GBU0W8SNJvkC9l/9Sk4g0UAF+efjtbA1R4wcVKWqKTjVO9cUC/
yU7bLwzLervq323pbx7FJwtSH7Wbp0iqp4gUNWvwO4htnpcG2gGQs26ueer3TG7nm1rOXvRcHdu8
4tpv0V+7f+/a1ItwvD/lrJDvYAqyWyogHrdlmSE1YZ+iaZ83cK4i+kg9fkwnoMz9VZimZfoTCc8d
vE2PbYQuNn4dCKFsyYmPh6EVdn8A/ar5NWvONFLy9CnIfE77AKoct9+Sj0egDv9JErZ89N6tgiTw
B+klNXTiGOQloZ4dDd4Dd6cQB/twpkrci6EpUutEVGixJtPPXckEdviyael598V+SKkL+D2YwuNx
lH8E5N13VQ3IZIdjaCLvd0VwlD5EAmJqRRRTag48ogGi+Qfd3voDCDPZpn7jFX29FYQKRcHFsMM8
4uZtUXyl08YdroJMrXGIH0HlLTnSKY6/n2np/xc2P8tvWB0M1MVYKyU+/Q2/90He5rWQN36TkGR2
xoRSuxJkEK17oqlrIabKH0WIdijxJhCs3i8XuhXpDtYjfg8dY6pnOnzPbM2Xefxzg9socrmHkY7A
voYm7wRy7ze3f7/Xxz+p33WE8r29n6TBcHdnQNaD5AcwjTU3xYqvsxQ1xCRPSwbn/MwIfQSw5+JX
whRKeg7RFZvac64lS0zkT/lKUASbfzIwqrSSKQ4NTzYdfIzy6N/bZ71d70GElOaSOaDbGdlj1Ve/
ksz2b+d4Kgv4jvi435cVcCjEYq1Qm/P/vOW/K26coregiasYAoRdxd+VP6ItlXOXCQdFrJUcC45k
MYoUR1kmcdv9nSZh07MArCnEdxpmLytzr9cI8oV9MMmEcFhPZLk/DoGlReXkvKMr/B5Yhsq+hGxh
ZADSurxDSN3lJ82jgrIOCoeRRYXhLY2VYOy/DJHYCsnc+iNuvaboIZgatRcCo3E61oRo15NDZ+kd
N7E5Hjco/+3bk5ozJ3WagYk/nbs5iq0euczatpp9jct/fUlBiGqgaMBJzwMIvozTgDgAg/CHLpIW
BRdli4vaB8TKMsJSZyfclFxYyHwpLMjK750jsypCwXG3E3w07mexVNVhiKhNdJphoPgEfpn5Zq8i
ueBWcpCJ5ScnC+TMwDEvklTRNH6SkJexAW5v7xkW46txNJ0y9nRhkQN1LaiI6ahRmkMdOO32SSDn
H3YUal9AZlWbtW0dDGCYV48Uh+4RVGgBITImK8O0uWs6vu3Xa35mHDMInfaABlL3BmGNJJTx6A39
z6hBK2cvvG/tyW/qoIbNudCXUNmrLRhmB3r9Qfsv0wPE7Gzb1NaEXUXts9mhw/RmE+loTqERCh5o
jJdVkOxoB388o0kogeVQdL58YhSsAfTxg2Jke6izp8LY8qpuyNHDYYYJDgdMcc54+UNkPHCoB13/
S5DjoqwH8K+LYcPhhI/fy4ZGwBnbMNT/eYFohVkBJFs2/FSqhH5IX1uJrCy+UN5Hz1kiVorQvJpg
Zy39IoY8FoetVEgPtmtNASyw7i5zqjCkfXIgsa4IciwdspZ2b0lLo2jFg8mDGgo6Kz9SyRhAXV49
iXVXJGpqNsZH+a5SYT+hPRNcJ1ANRRdm9KZ29izxW3B4vpv2U5tbei4MkNsC20yvnEqb1sE8iAKH
rL5knVbo29U7zsYC5uTvltW2wed6Dq21O9/M9OUwaPbDKbsvUkPW2/mV0HHyeeGKszwDhjdWN5uX
8knBsOaBdgy4s+thJpOiAiWmVm0cKShsU71YLG5PxZ7TLTMGptH+W44UC4EH7HwPoDNBHkpCSgWn
doW4oZyvw6wtcIM1a9KnuCZ4oicqinWRZKaVLAu5PftE6WhdrWIMYo908BSQMxoYlxrAX+VfhKFg
MalNTga+Q/iLZYwEjwsHPSEBEPfUeirzn4e+/UUM2318O3yCPzJhxP7/onJAIA6CDQaC32tN+Qqb
/WnS7vLzsNfUHMFVMrxEWcdVnmsLgy92gbuEWN3w+qlbl0+9581RKhCd7ePCt98FvV38T42A+Qch
5yc9lcz3RmY87jA9OjiJ7d0ArKjNWUVRl1Z4VeS05+CeKRaAZwDHG2PUDYGo0QN9UB/ghsJqh5O8
zVKT6Hv5Bh4rqDGyfe5EzZXBeMy9ju5cc7DR4OrYGbJt//skRIh+rMeUxU1/X3oIjJG9EhVukiLf
jPqMbBs6fsZsupWxcjVNiJulYRWDm4h89ovKpWb40UspYlvRlhZE2eVyQG1Y7vrZYaEMsS3VheI8
2uHf8jkYDe+hnDI++DYNVwFp5YfTmJk1xE+Q+7fKOZzCTOj0Fvsl6w2xr29oRatj+T5hkklUnG5O
vYDdGrMI5ufnbK66Q81gAoBqLKPb4PDmpY74ZSQvmnKZ7tvTH/J+6GrR3Qew0QjeUYSpZrRPP5Lt
zjpj9yNZOzewgC3w/brzj7Px7sy8Id9z4pikTEKmU7Aj2SymPiwcfyEhxe5X1H7Bs53ArPv+9TI0
TWFn34EpFtUUr/6J/hSOqGK177yKL2inh1iN7wicIjkKZnzCVJkRABA6WqxzFg4ixbzPgEbUNIdv
/+OEbsQrK3x7LoQeir7b92huqEMlkqj3mrbwWgsFml/JFwK1QAO5HqQ0BvHPb7YgAG3OEKvsDr/S
5w5XpGL9WTO/zINWchAgtMrKsP0d20fYoohQMsVGi5242ndFD091flY5ctUwAke3oI1ZFQ==
`protect end_protected
