`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TzIiEMtvO6aATpAtL7cifRYecx7zo8XqEtOIGl2U8qAWu4EPO5yX9IJNXk72IOS1ltnUXQqR69f3
B6QpVjfnPQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DxJZUvltyEq6qJ3C722l3oEd0ejNiidFAUUWEZRjnajRyvuRKM4LnkdgMjQh2z1Z9JnU19tU0Sh1
xsX2zoJhW1PNZr3YdKS7kREU2ZaIrR2dYK7qVamHmjMmsyAYqRESuxPXEsNLBBG9bizURmqkRCSm
Yrlp1QWTnXwxQ5hvnC0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hdn4/V2pUq9izJyUhDCyZDTwujvykX/eyFQ3+UnsybE7V475vPzplMT4cOPeFuUq9BYQ4STnr277
iDaaRHFzLn5ct7Tn1XLwWw0gUj9ktqROMa1Pc64mnLuJXtw3JUM5fVEaZCR7/HZpGAtV+dHw/fAI
9Ddt6mZ5FSiEFgui0xL/koc8zo1jac4MMeBaHasqb0T5WRUws3n/yBxyACXsUpNEiEL5UNaGu5s3
S16xeAuK7SqIE4DtgxqBYYWx6eiy3Ws+k5on7TW9LFRC49uaVchs8B/AiYMXmx7Uk3R0XySa0Jla
wy3MR+rjV+p9WbTFsR0Ia+hiTyVluC6nuQ8T/A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g7/I+Zv7t15xDNb79Z5Z0LdkVeoQuvr9vwEyA9Gz7P+XXaL3mKtC9ba6fHja6T4sIcW9smQKlrpI
UIbpE6b7wC27IdfUaVenB9eSLp1oim6Ym6iOVaHIzIY7MOyUhce7HOsye7kinmZ+2UrLH/XU/swZ
CdXbYeuJcBbKnxo2e9w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OEKn+Zcnj7wYOTFSM6WyEqNWHcPmFfVh8vYwq3uT62xdINEZ8kOtiTDz/W8P+37aFQBu392Ro2Dr
Dpt22eyk8hM6CwjpHmO6+pJu8gMM/Iascx5fxY39tNbZJTPdvzF3IlurziOuz7a5UySS55OmbTSW
WhFJ+dquq0sO+XSnH0q3dR+FSboyYyg9SpGRn5PKwD75+8HK8M9Jnxd4fsxFvgoCNmXBNng0XbX3
AcX3/VkKpWTzD2/EdVc7lqcH64jbK9J5vqeE3+wIlaS7tPDigA5VeWPK1rCcOEO6FTvl/i86DYIO
i+IdRlrGcK3jiZzWJo95VidfPqrycYocISMknQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4656)
`protect data_block
WSb4NJMG6tDDjWuGtoGDDfKJTo5PrXaspzv6esWhmkP1vGrKF6CTAmC4qVCCDf4MJ4WgSwdNM5ki
fiiidiYaUn+oDj/tbwuG8QUzt3WO/HILmeEf6ObuhlsD60ijhw8ByEtRLrorvTdQpiaHbdo87k5w
y5m302HMWD2lCT0HEo12CJLE+yAyxZCYNc17s67OcbW2t0aDuzRYAiOFbo9NgUMq20qqDorQtoAc
Y5MPw9ZCgudWCB3TBZ7VvnuvX285JWC99RAnuqv1Qxl4hZpnoE5R1tykpZQTwXfukKLMFwPFxbzV
WCPeO39n3bFZa/VEX9grbmi7HEO9l3TSuA9f27YFwVZ9PxPUmA9IZjyUGgPJGDLXBagY/gWe+ngP
t6UyujhbT5TlFHxioUbwL30m3kt8XpRXDiHvu68VnHmun/zA/DwSujw/wBlQIpEMq+gjcU5bKGF6
X8WPiT85YE08r2ABY1y09QFpP3R1BTjfZfRNc3PZRC6ID5Lhw59XVACLTKFihsOG6QAIx1CCLtM0
Og3AW7i3K5C089ykfVDvcWIU7iV6+0Uk1anl5REQ4n69eelsaS3MZHo1HPnjh8fNjhLOQ0VvcLDs
hOoA4twQ0S35GTdFuyG0CKPivxEqpkWLtodYtwMT6TjTfeU23CxdLrzbZ/R+ERDpyNEEJ+9jUIZD
5HZjkLpwOVV3fHv/Pglmc+NURNEPiGj4Im01Wo/21HV7xprz3hW7ga9eaJxZmYliRm/kF1allwzt
lw1cQxVPlkoDI4MUo4iMEwjhZ5MbIFgStUOpEVyz0gRWesrQJGEWoXfww1QXo29aIxIOeTzkkigI
QM63Qq2Mm7+lcv1nTWfYP+cTV92Sl4rrAsJdaj0GUE44f0Q67mwsed9rEEqaBWxIQA8fEUY2AO9U
2ATcn13tlWv944Qd1vAyNm2/uqVofRx2d3dpvgEgIfw5aXQEx6zi3tvP3RmImDK2EL4tpLGKUevs
DCO6i+eTjB1sSf/Dtk399YZl0kaDoh0c0zqEfHlgbsiEpsBhk8AHBkXZbXY8AWrwXa+VXYarICII
GHEtdx/aHrUR/RXeHeYQp7cfOLM2eCpmWJ+2/KBJFtylwh6kzur1gGXLljDa3Td70GzRK1RjoET/
B1TMtHawAS+VAEmV/RKWjuOKVsI10oqbxEdYKFQq0SLn6c6+kZC4AevLp0n3IeHW9X+0X4ceF+Qr
StUY3BscjfRhBpVSLCPtKoYCXOApMqiwmZIxaeVZ/KWJoi50HB6aexfsUXo9ekUilC7Mw8jSVAhN
JmxA+QozVWJQhPhRt65GaMWcn/pkCK2n4tyQ5Di5Oa4t7CcwYYzEXZMIKw4D1iSo+RrcOmAArvYA
20AQyfQ7C5RsSFv4ZexQ+5pW6hPlbIkJOfn/YY3m4igIvfYBFbnE3HV0JFR/x7i5aqFw+GTTw4eM
+h1MhRZFQLDoEUoMk17F58GxJ8G1JYVI0ki8EhRGTWce/f4eLMTKdv0/JjDIUk9inxD3GeTAll7+
AMyl1iKVSIgD4moN8xwCfunj+PSULyrJkKGyohYicZS0YOJ3333chcq25BAEYPGj1JqN4xc4gjbJ
E7Mf0+BPIpRhJ3iS/Fqp+v6QDDbP4kTgSdO8wkaWOw4xJGh7V3De7lvOAUXIbxWHGUveFn8yPLMp
vEbF1tfDaumkiTvMCrc8R5rbK0IGlfzzbdUHg9ImpZRawRwtDYPfIdKXEUiEPgFBSDF7k+wvi+5l
9ofXCh19oRU6wJj0mfNPWpgXS/pKoAuAuxRuzJQN8UlWQ+i7hld4nMxMBG/xDl48gx8uArmXCKoG
lBg5WXYMzGRWc5CadnsJ6b60Zh3qRBM3xNns48gT2F/oWwhk8K+eBKSk9vyVy66fRuAzAGOscHJZ
k3b43T9ASyteJ9rsuoJAuz3vUFvrXzKyXPK0jvITDvg9/XEqIbmgePV2jCIoLJxeVxMXSWOUcAMM
IO6J4ew1E6N7ju4MI1blppHXzH8uzs0fXqFND9F0nQD1xC2wTCsC+mJ2UhPAa2H9v6/PdBYhvw1L
fE7bzwUBJoyZMfTI1X07qiD+qh10TiyZtgTQiSxi4iTs3Zo4JExuh/e94QNfekyKuKFOy3MUo6iR
2SJT63vbyC1gyVr5olRO86jWDmEYNA+xr9KhaiiuF4ZOxx0Uw/1MWkHVazA5hP2V8ENX3co/RVso
wBcc7XrcS9am7x7huaE6v9dJ7QRibQCPLOU+3YwNsvQXym/uQHA6XmSwFQ9x5GKGTL2EezfH3ykI
HIHJMxejQ7UI8ZHCsRgl73YhnfepVkCqpxkhRkcxjzglm09s7CMIK5bvWrAqdj6W6/IG0YJdV5RI
c+StMl//FZgqDkGK333NXv9nzpQHDZAEQ878tgpwTES8hNySuoaDjEfx8ju5v6tV4CA9Himhmqz3
LZPiOEcuJD1V8QeD0LrngppoLIEXMjXvnthJiTscRYLTH8zzRXMSLnJ/7byCTJ9N4rH1n+l/08Xl
hH4yTYxdyCLu3ZG1m9UarxrItaN7KRY107vsdB9bzklVcKtUgrbU2jQQI9Ls1ujaAvh/ksCeXUN0
vE1JpC/zqa3eGezBJBf4URvrXMMk478CZV0A54AMfXwyse2hl7wBEolr2I4m8QuFL16NKDMUwJvS
LJDzRrjaGYjcJu7rH+i6K3VrHH2y2SpUJEzRPgEcMA+xv0poix3ZwlyM3hyUvOYTl84YfZRI79K7
+hfyIAP0UJ8yUQEx95EKF2Qo2GBddQ8RVcpk4HvqCZRUC0pA7IyQ4cisYNcKXSARjIlR1myQA+KY
Z8i+HwrwsfO0lzrEdhmjT8s3OzNjgBmICKLYO5V/35BdaDC+ompU1GmdpF3oiOq7z7kDPUvELQ6r
1BZAV6zO8RBJbWHsEVtKdgVZNnD69drjJieN4XtInNVLu2PC1/ui3mDk9JegPDFLLq4YF+F15Y66
FFvMcqKFc+r13tTGS2PWArLt8KmVFuJ1EtlEO8fIbdaXaVYbpcwIQl8+fUBrL3rD/rhcY43cSFDe
b2NSckOcIsXAcUNJJPmCfkfVHOPNNjbENAdrf12waSSmK670lasJnY1a8hCC7WzOnVe7vOrcSOwT
HnRDjxXID7uLY2RtBrkjtzyBjibw4XuHBqwGRWxt00cta1uzi5f0Qy0rTwCDhhk7FfGAwaaISwT9
Sxu4iOlUTQ2TEZfM+fr73UV45IQowMACfzS1xtOT+2uFrynG+upDrbMPB5fTnjyYDUP9wG5CXZWN
Ec5I5gg1nE3LltKqQcpt3VCiYMjjdSPhgwKtO6Ay8d+xSHOmvNYMbEgrzrcFxl54OqKnD0CsfOo5
8i+/+DISf+o4bHfnxan2j5+L/Vr75GgGdOI32Lr972g850bfj5U58ZBXCc4R4hxQrz2HO57G8jb3
0qMN3Tu2bm/oEEKqiUxuojQtX2jUrK5utpvjBIs43wzi8pbDPxgxeQYEMQ/buPhqmvYuw+nwwFBh
p1pf+zpCjgYrshauC7o0wSVw+8pTKv4aUlNstgaiL8TbdhvAT5scs+s2JWfn5uJIHBMf2rs7LBAp
wSiEb4HRXgDY7/9EihVUgozSwiGssrNAxlh0aTwQw4NZu03zXlR6BCkzdCQ1pcCIe6z/GBn/mgJ4
ySaGW4HrUa+5mewzcnGe9wwfS8EdS8+EaL0bUOzB5QvYT8Sur9eeWjuZj1n43hSa9BZ25ySv8mUK
2DdTNCjYVdzWbde1SjB0HJDLZvnmylDN2Rzx6ZrFwJ9m7UXq3yYcfL12V+iZ68iwGl0Zw+7KuqnK
vwHK+jWIv2Jt+wizLBrk2cebRNplMCzyKinvOB2Y6wO5NpVC7FjK4H7S+iPsRQciZXf8U8/Dzkj3
RNq+pBor7AFzEkcDsHrOZQgyCNBA7kP+DCy78E5FhibSZj5iXvocNnj/FK2xHo0a4WXQF8CAOAQZ
DPeaLACjSCXTCT7z1tG7/7c5qrg9c1wvys8TOWevtOz87ZzKcYRrRjpVdgXiI+3D5phxmPP7Je/S
KbonLMGzi6rBVykfZ5u7e/viZHxokpfUrGgX2dz8kvOG99HaVvuwDptyiTLzf3FY+8K40h4gMZTS
beFqF48i6BC2JaGGJNDakx35t6s3yfEklyHJEuLdbe+UVMUFxz8bxSz81eAQ3RQF61B+FIxMyN1+
zZST2oeugh3Q+gs8yReBvkJmz2HkZonRKY43xtATdLgq7lGrKsueU2qh1WYvf87bo8ICLg9kGtyZ
tDwpUH2jAzor+tyv3I5XRGKhvRlHr64nltU5pWBFU7dbuXSBJmHRYVwg6v0qsY6aWp0MH5RNdBMW
tY5mpxplnB/cZhqqFnwt9QpjmIRo4ylZoWY0qzdlxRvEHJ88XnxcpIAbdX2tgZWqEsmW4dwVnfQK
IlXUNupNEHMBffUd3UpXBk91gNGPNymZ0SSIpvz2X37JGJBxSTEGTzCoKNgT1o8a4gpe6+Gn37UG
Fq64mD5E7ag4j9U3hSNKU+skZmtbaBr+1M3xCgaMil3ecnlde4YMVjLfEAwLwb3EdLrcshXlIgHY
cBy1TyNET0k3eLMN/81hTc2tnVDuYcOYBh6VGvJOHbAGeL5ZpGNj7orsYndlXODESTCyGZP+IKec
TBrxLxGp5KIuKzAG06k1EgfO0vP5AfOu5U0msSPV4hRycqfjgVKBRqD2Yh9S0n/KKbn85EWvbEIm
+QkYekneJHX1LKH692jOJ8Ww2RrNj11CTjjtkN+nuV5MYWodHuDNQes5RrPEVbWrI3CR4jD5lRR0
4fE2yPeb/3SWqtB9M997BrzQMAT6TRVPEhABSbdp89HcUz6VqsIguY8teF/z6121ZqCnHPycmptd
DuX90qcYDGX+pWfKMWycpeGteq7k4lg889ndD2gnh+KgoUj3Dokyn6Cf6RYceTXZovxxCu6Itr/D
lbqyoeKolkxFCslxTUbhtF3LYMF8RflTZEzMUw2eSfdQxIGGIT4zhjbM3Z3LLH9w9+6mtHiu1Ver
hfqyYUFljX3at7ZweTpaFYiAGoAN3wfHm4L3sAgrptGdhZojXaUeB4B7AJzmJl7mxzHlNXaa9fEe
lJxrcxf8VnS3rc52g8dFEDuQv4/elcXevYjPHZanAcvQAjjOHwDPlIS04xIrcmW7Jh5nG8n1kLF8
0VAUtD+psgl+EHMbNhz7C9RLtCbMBrt/+3hZT3A2Ixedds2o2jGjGVB1uaUH6x/Yaaf33FTPl4l+
r4bOd4YWv2Wn1Bw4KFvqP3np9wxhIfE9pFwHlXZM5n/YE5Rhkr6UHQwsLrX3NwV17FH3eEEpyyJ1
O55bPArqhXZ1kAYdAxBxljtUKk8LJZKuBU+RL6bwkloDa5cTDRwofRMaUrGp19rQ6/+otAgo5hH/
YFoODxqMuYWiIXHvdH150q41U/g/e5EOCMmQSnezv0jyPh7/5h3R6HiLo/+0vSJ26DBhB43niQ5p
4L3PG7yahWax1678ASiKia5DxkeeQzZMbo1WLwoKhA5ihKSMwsplkeeV9RN0qbGbvwR09pjczQTN
P78OQqEoNSTh0kfUFL9h+ljyzeI1FA3x5BGW0w0sm6oQL8jh4KPEHVqjhmMFZrx3W2ElXTwvid0c
4acTL/Ce+wwHfI12WDYeb5zYH/2tLJqVg67hUuObf6z4dKOlex3m48lIgyPWtlBQp3jGSmdwSJdP
hiwQ/tJLrTRporHhl5W0Cd5zY+Q4R3eWtHOMdMHYJE5UBzqCMAd5xbr19TX/fnAbKqSBy0U99puj
MOu3ENRx8jXc50x78BbZvnL0WgljEKKprs266I/PK+1/5VZSXcat3VAGEt+Gl4cAKnF5KqHuOW5H
hVgm+I4mrjV7YK6PXunDBFq2YObWRZHTX8hqEaAdEYLheqpQw0SAyuSCIHGZnV+PkqYSj06uVO5c
ia4lOUWYSFt40aLeZ+GO7ejhOnt7/FXSkCS2D1s7eLo8uf42GxRqc79fKQRzEajsj3ZXkeSLHY27
xOO4ZT9awc0YAZMyZHYqeSkULVfskKsPUpdgSE6Ebq6qZNpYD/ZUKD8sYrGxc8xoLG10vNNs01V8
fCZfixI1v1Db32WQLnc2YKTAAkiH+o+IFjLL4FoLUPKiEqUTpMwIOa4J/i+eUm/Z+QxNCg8sZZon
m48Tg24MSVJ+WCsSlO1u4inYDO6t6F2Ja86O7Y3OZJi8TigkzsQM
`protect end_protected
