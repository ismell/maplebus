`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UAGl33eV1kZYKmI1EkF+sL23HYyJYovI5Tt8xtrxczXuH1xXc/bv7fX3YEg0AI+mzFwJglfhCeqF
7YZIZb6RVw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GSg2hlRzoqva1ZcJLSU/keiLr7EvSxbFep6Qy9oAMkTEXBTJOmxXlOLJ5AkJ/vm10i/bC665rZEv
zBGMrGa88I6ngjoj6I/UgTwGu1T28NfpRyPOO+sYF+KQqHdbNOGpHmyshG9Wyykdsb5+ERVd/6gV
F3VJfE+4+ZLg0mar07o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ombO5+K1OeeNDLt+fcM7+k4zIqcqRFbF75DVKwx0GkUmGTTeKpJbgbwapys6S2bFyiFXzn382rcy
kzhNWPguaBweOaC5FDcAsXSObyI4aBj8NVQ1a5HHkPxnFmS9SG4nwUHDPIP+Rfmc4vSXxS4eagQ2
lQKBjhti+bQ4DYHnDkjIv10ora6jGoBG3/MeLPKa9PZvWTF5Vme/i9tSenZl9dlCDp/1EW9jGhUB
eY+rAVHQfodiuolvN/MXIvq78ZfB2cwSca9Gohb80XI8oCslPOIO+8O+sfPeAOm8Nii8qwts9giQ
YlBKwNmlHU2iCv+JFDH6Hq7qEz2I99d0Nou9GQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PbhQS3Igjtr8bvpjwV5MjRHwXvWT/MOf9aAXJ2Kgz1xsTyk1N8HAyQWBEAPnARGtnrn/Dsvo2yHR
LBp39xEOJNtb+dFsyvV1IV9yl024xYFteWNtDbS/aEiptJWoH3AJCsgu+D+x57ZPmx0r/6S89QXv
//pFa5Wa6gryCe/guBU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GbTEUk1DPMNGS54CCuFM0CVb/kcC/Wdr22uVUt43n9Gdqd+vA7U7bR+x5EcCDRn2Fy6E1kxMEMhz
HuDNxDdAUT3DimgZ6nE8kj8AbGI+vut9wt2GD4P+yyunHze+P3GSivZGjaN49dZOZXQ2iiSKDnl0
GPrjTFcyyVa2F7LukzpfDYpzjjmGLoP7BMdUkos7AsgVtLhc51aLkTQ45H130UYKg4Jjy9nJDxwQ
5wUkyz7gPbv70paH7QD3JEz/weJclOlbhknBCR20KRQfY9yRELflJtebPhgt/0iD/21/xmctMzva
dMs5CLIl348604+5N1SL3117Nf62Ud3Bi7anRA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26976)
`protect data_block
G0LRzYdaG798oBar01J0vgNEJmTee1/K4CPnT2QQ1fV1B8nM1GJW9HpJ20gyIfXknFBf9jZZlBP6
LJqBr8gETtgke6dMHDV/JIM8bsVgs61xIxErC7w2bB7nAlSZFguKqUWdM4il9vYUkXYDp5CbjEoc
0T2nt4QFqwp0cvRj0v9sH0ZQLs0kJXdgsxjxNiFiBtcaLWbnYIoreXCoUzPpyEcqKhDSerQ++Ybh
F6ThE43WVpoNqn/MQrLEosJ77WwVciTaojMyST8LRRiLR0tpGbhIkOvzYRbv9+uE+ggta8E2rfS6
Sb/oYc7alQNm+rzlqXOXq6dRfHn2NE0WC3lN4iy3fA+3CvJuHW0j4D8Jbrzyz8yJ0fYopA7Aub5N
3upKl0VxA1Hs0JwYlMWvWZY+/DozIF9y+OoFHZfrJy6jrwAOpM4k4pLQPJgIiSRZI6eOqWnEM5r6
ENSnDNgfOQLR/JKg65NNhyoye918/QEUMDWWdQokvimQKNBJju+zyaAke5Zjz92gXeSk2CRIxuHK
INjgOsvcrFs6ZmHF2EgPoEbQUK+H3z5Rtf8tKgMdXFS7qo15bYNRYqAWLOSHT3QkiUlSwugQ0zbM
xSM7wdiVtPwxjABWGGx2wTKFD2CLkTiliKvKUpwZVvsbRLAYNQj+EbT4IJKkqAd3xfM02uznIUXo
E7wSrie/H2my/BM8eflSH3HcFjel/8on6RJGHmXY6p7N8yci43TBT86t+/KG09mKlW2HL06o4GTe
xXJTRKXcVkma9HdMYyiBxCbKHHRsN4lmQnwI9dm+p1J4pPJqFziQnOd+/DHaxM5GCbzc7urZ/36T
0FehEblF1SMGOLKPMVW49s7b1G9CC8EMa/dNQYutvfmZUpkC5ZwruuBEUkcNuC4ljUAWmiLMPYKa
nlsqI/fVBicXWxWtLz6kXlmVkLSqBFEgUApqtuV2BBKMjZ9YKyjVB6sQNui4LOPSrXmAjdU9kOAX
ZY8ytzrSoYaHicCbpH5vOl8GnNz41DWRhr3PKmOMZ9Momvj/wXVTQIEbVuWfbCgKNiJBmEKmooiw
Sw1NqdeJp23Dms3E88qDKRu+WTzveHvyoEUTn2+me43Rtd2O7pkrubr7eE0mKgs4VOWyefVbGDpW
qQb4N1XrCAWFtWz9cA9MShY7k2tjYGG+u27Q2vD8/IKZhA7IwG3eSePJ+/GPWor43UKZpCplF2UL
uRl5WdUWlu+VFdY7zOK5AfRryXn+enBGD+KJrV39rbLTQgpDk6lfcP0wVR2MWiZR7Th6Hn7hzJ0k
ctNCbJz7/Qdq8b5Glkp2a+2MHaXCeqjAQev1ip5H4cWScpCTnmgAduExyzi2OCK3kTnK4I5VsnN/
9zy1jmnFKUMlQRVemuFf7dpK4Cyb1iUqxcYPp1DXtdeblooGaE4OmPmRSMH+X4OPe9jEU73315l0
OtA8k+ylRy9Mkj+dqIWOizN77Q/+vku9E66OsjEsPNUVfC/2GrU0m0i6RON2lRSq5IOQ2MoAsQou
6kPsccVtIpX1qex6giDdsPOtBoWItRZirfpTTwMRDZ+2m0q8Vv1K7z0Inh8W6vP6ApaqRSXiTWpV
rHphOvGKVEXtLZXUlp0O4se5lMI7k4/EIirnoNebPxyf4xliDrTp30XSNX/o8R73WZg+OoPo/3YU
u0aVZtfnWDOaBlw6tlkfn75rcpzsrTFF7ge41SQaKAbf3LGC2AAplVNluUG/l6SQZi5zvoMY92li
mp2DN4mW1PdhQS8q9/JDAcq8FBNIPjFHdOAhjze4SQtepGkV6VnBlTDRyFfY0V/yXgy4ESkZCNPP
I+fSxwyR7ZALIqYMdYQnz/cVZl+WOCQ2JWzQqWxscdIqwhxKfa/+KstV9ulyk0npgjPKqlszpf9a
aK5TRl2niXXTa4KYcGDKsh5b42RhRuWuIrXPhOjw1GXOmOsxENobG80iaYebuHxVbkWn8TsRLnXd
jvWuvfiOP4DWuymJ2NUHi7Rhz9vGIoGnFGsfEHfpz2lERcwOQLaGebe5Pvn14/zXhRlrtPg4xTqk
ACxP8R/6uMJ1BT6Kiry72Asg0Mgazdpd47cR+m0Y1Cang2eqTyvNBpEL9WrFkYCa0SENU23ek+tz
CTLFxUfIx9Cp8CLplab0Z3N55DahLw5Vr2Lohj0jl7PlC9L/ij5//JKZzKwwZ25AV5kTU2RLl2Gv
snCCeEIDpP8OBw4feirQTPQJPDMkipecI0blwNVmmCeG3NG0udKro7jZ73vHkZZ8KJ6+F6YMpevH
jH7y/ZQA0nt5a+fBHR83b2luKI+60YNV/AtbdkoVHtcV+DDV+99iECcwCxECw5n0GaxsnQiI7Gi+
XecV2J+5YOMdLYBdRuxQTFjeDxZSva+f3W5Au+oRhQ8H0SKVjhwmpJR+o/hZECfCBS8qi0YRQHjz
Q0cV7YrsTi3K4AxJzeZOhy/f2ACjDS16czTP6OwPu5WzJ002QTP4q6es0UT3HnOVkqm4qRXnnRzG
CV/niN/O1sYP9sEvUcWQFf8vx8aG6nAlUhfO+iNhtqoE+1P0OA6oK+TfAQmoNKelj4nY9xn0ATvo
7wy3AhknrPkea0njsjT69pvzWIHQ/90Bvw9lc+TAhaFIMiUzIonX0PLzlmVi5dll0dGIe7kwZLUI
ByOUpvSODozw3wcchv8KTq0znbRkTULNGc6YlpgqfI5zxvdU6uaGhdlrazSXWkwujo3zbcvGfr9o
rjcyR2tZ/bhfIhsBvChVpMGRRVcwCI6DVw9axLO8DDptO4u3i8m0pO7kr5/zxw7qdu+Eso1/OTBA
6zCIUUWdcw+SzN8DGyNvysJfNaqbdNcYq4fI0EJZFTMZ0XRAGXi2yq6q4UscNfSSi+AwSnPVal8q
bjm8E5/QP5icQDq0oLNRYax9IQqUhm0OYRvi3HHbQV1n/SEqPO1uO+vH2Z+Aj/BknTkyDDkNERLT
rH3+amRJmHRMvrhoaI19jooUTcFeBkAMCUivKNhJ77E1hn+DeSRM2LXWBIKzjZEKWtatVBchUG0Y
/levD0lt+hVwIafGJEk1TtlwP4/cIioQKzkp58Bf9b50GciwKBHhPZtkiloY8xpEc21d9DZH+Jgc
oTUvFIYrPThD4+yEJ+//zCU3JTxJbyrjgpTe4AFSy51CprDRGv9vSNGn+wQMQM8+T+C6vBRh52X7
41I5Lh3nREDSkHFroalI9CL4fbRPu63XtwCxr+260LqIX1l0CXKt/HmcM4FholFxD8FAd+FIXw3a
UqB33E7aQ5Orr4EypNswnrmus7F/gXuq3Kq5gj7dpwN67zwElEOanvpRFhd0qjGPfuTr1nyP3J91
TBCRe3c0Fr2O0+m16En50wR9PbzdFSnr9Ute5bw43Dmm+JPWrY+3F/gUeA7UIYFW3iDeRR56HLPu
3HiUuHduZXhw/jqpZTAXwS9ja0LryfATuDp8i7jbYDLMob9uGtskYvAsAs9KXg4SVMA0QC1dWC/d
EgK0hwluVIyVA4G9MRcPr55vQdQmGFQKpI8AUPRUoVgfLYVM7xV2CWVnOvQnJ72LS+4lPl223CgW
pci6RZTy+1yD0n/0FtN0gEaGhSCYk5j947qCUBysxLanBgn5C0RctP+CWNDZwh3Zag7w3VA1Enuy
F//85si4g+BdmiKo14I21s8fHRsJei8nEoUHNYU0O6UZJ+mNKogmsPaDphqtX22S++bmb9mg97WS
w7ACda1gXg9Cp3bNFDvELUOru8Glg2CC6pkF37vfffIgectcUsl7oxqsp1iAGBSzV4gBMWXz9hKk
ygc65UieaBetJjG8NrZ5wnqPxWHNbPnElfnk3tRa+FDdz0pJlV6IOilKEqKUdX4Xlxlg+/FsSMI/
nxf/Y9lNdDcgn7YCwCz+zUit26q2/5uQfNv/QROuL5957wEsSKzTD2VoMC9G8tqx1crjTy+tiNfm
h9aaN/ucWSjIc1XcpD/giJWqhU19CTJelcorhMpeV54rjbpOd3VDE3ABjSw3nlNkKkXaFBb6QBE5
WgTvdznV+6ZcVTmzn4nPPttF4i38YuBy272VviVF1OuS2TBBVGPGFL7tWuZCm/jdpQFQONF92MQQ
OLzPjqCwQJgAaIeheTJha/jqQNI0JWogVS0k2n0gzt8y2qVZSEnDoZFTu/Hg7r+GAcGe/wMv8uvS
CvwYEhai/0p/I9wbqux6DqKeylsuE+Qj74P/kSFZC7iGgOGB2RrfAUXFtuaaFQtqqQvRlG79Mzsz
+YF29bUR0UZXIuydod/bjyU3e0QgK3pvlBI5d5FGjsHOOfZFBto4rX4ltjs622l6uXEe2JfZs0LO
D2U8gjI4c0F4p/5+UDozchBAzdGQuHC9F/JhVUa9fqmZJj6tiVcn3z5cAw0xd4IpuMymE8goe7zZ
bTty7CIbsjYjRCXcfMXcFbVPHtt+nrDcPwT5vW+pW5C9bkXVFWYw9nust3SLdtSKVBvfR4Or0M2j
9ovWAt4AiRndS9E1pBNpkkzIXESNnr9xmMrn/WCLcrXJEIunSe+jhu9xcHKJIGq0eRlXyICpxuik
mLwC5lXo6DyMIrdjKvVI7CVYrddB1WMvITzkm0IgDgLxRFdKfur6k7kL/+QSspa7e6QyoiSyDnQj
8u5DClI8JoYo1/VNKLOf1cQ6YlJtSbsULhoIkRHeO+syPrWRuszi1scgPQ03Su3oyyeOFMAKi6kd
BhttYFL0sNh7QnHcGXemwJ2B683JQ5dEBlCYFyB8BHHy7YZ9bMQWTHwM0BJwaMdxl6erz2J3bDb8
XZQ2ovrLl+RgK+7I0HTyJIrPkzNRoibKYVH3I5dQRzCcHwBbYtXDw0Tz/S3J1Q4IxY/Yebz7myw/
H9IkK2VVdAJbIj5UxJWAA/V4Z0sVAUpIxuPWvN9zHHvbL6KAFt83gvPj6VSpxTo70Wd5ads64Hs9
8dKZ88G2a7bHQAiUn72uwtjtVi7dteWLFPh2lvTVkW0nqIWNjjt5Kyi1LHwP5frKVYxmkSg5EI3C
AwIRHbTENYmBSxHUNmTWQYV+KQLmcUDmrs4EF/jkDT+9+05taB67SecgQYRxFDaaGOmGQmMsju3e
ZsxKnVyFalS9V041De+Whb61p97NkZ6qLrVG+zN6maZf8aA5Y8QymMnmiJ0/kcbvqoUcBpJjMnmj
Dda5rLV46HrfAhCr/XGEkdEy3U00pslanpg2Z1xOE169ZLtn0+QSP1KENQVericibjCuBFu7mOhv
NvRhlR5wSIdTXJ6B90dtPEysv/anIg4IswDT0qFthsEZlIfE4IZbYDEgjnOnGDnPfH1dzh3CB+Cu
bX3QVAEJcloVJhaETqIRMAp8ILGQYWC19/zPmFdGWUQEFH3Ug4T5zT2XSooHI7FxFZDBQa6Oc+O7
PSgUNoLHdutBEXZQrJUmnIIQ0KazBaE0RK0HYtM7TdLQm85qCGHL79rD+QB9KEWe5X+3RT6qjOyo
kLKHqJFpgl35mBzFwQY/F+vzi+b0ZvGX+tn0uMDvKcDzm8QYyaUcW1pV1srbfP1zO+UA4RfGncTs
Gh6FZ1PkX0oRELkzjYto0WsDQg8olvuCPJf3Vn7ORjeocHR7PDfLXs0vtdGcOkwRw+n/ogVbvH6T
eDQRGCaUr2hMNrbF0mWdV8iDxTLnQj3ChpbbmlBypbgKbsykUetsDSe4NsmDnUruEFRcwGC5YXl+
ild74Jg8RxFDCrF+O/EepY9WnI4h7GV8ijHoAd9IWL3ujmCT7Ug9++MCAOlwl4WBAe1//s+xbwaw
aC81hWpzxnVN5as5tkX09yghGiyKMRmbn0Sg1L8sVO24aNw74yG264OsPku/bZ/5Nfl4ZeMiDsCg
45akVENkmimM+jHxwwL762+MX606e0ciKFCmx2JfHczyisN0GI+QOXl0G2RKxoDM6b99TEgfmqzW
TezUW8sKho8uNCF5YgaKIzNdXXnQINNliqHxZaRUMIxa3fnq/C7jvl2gfHmTi0kTpApczSf9zG0P
AFfV+ZLUWvxoKSy0np4strX8x/srdxoIeXOrqneMbVMdGqTpAP9BCmKCTTcdI1VaW2iI5JgR/ZsA
Dme4MZ7dfmOyGxuk6U8skErpZPKC+nK5Hbcu6jyHF48UdwGLxNsGdxT2w7mJLD4SyOzziOcEHSwq
cbMtJs25ZVX6Kt6GEICZndNIDsw1A4LciLz19jywemjHCgTILwkpTsYPQum7eVdCz1Fbd/MB6FuB
xOIeSTD8qpxwMN/aahQ5SwQ2J3qALpMLVjYDxfTcBkiX1Gea7/XeX+gj5b4c4Und7E5KKeT5nHLl
muKawiI5eklQbRI+0fzz/u3KhA0GOOI+2gIT7heVX8RUuNaNOry9WPkWfmRAoE/pEB9QBDnPqrq2
K8EZUnE4pnuuwjvKGbCmRFLXEnj6C6p1kPBxYjh+4GwBsMAsr8W1fFzPXTEADbmgXcWrWEGNXI6z
/5jrHnd3kd5Me8ALc4b5z/a+JUOrlwJwvCDCazSmCNGQb3KvnS6vIxIWSxIXKHC2rC1BxTSR/5cG
7jo6DGMeNi9SPQfhy5M4jumKqQy4TQizB0gXglUI37FVDb7SxPdQGed9SncuG0i6v0VI9OK8YKmm
o5AQx1eHnmcswaC0hC51L1EuG3iDsiA+5DuVdh1LIzsa3q2od694i4jxi55rE0plzgUC2XHIh/r9
mB1uefDRVkVDkR8s4+Pqk/Gz8SG6LEmiYDj9QyuwgFGWeASGuinivDQ0L0qndq0CU625PV8nGMce
0BGR3vEQ7z6dGs+u53t08PmxQrF/Z1WjYNQnoI1ZnUMt5Q9G6tNO2Ufl3jE0B55RsdH7UKq5oFTb
eDQVmuFTvRXs+j67epKTKOrh5dRuggZAbxGyMZuVowOO6adgMWsFOZW6DJRBmVORHDKYFf2Qestw
Rusdb37M9O3c1Sh1Y4n8UQKKLOu1slJmc2mmRPy4DPxXMkMZsYVYzc3UOUYJHygp+Cnj31hKGX8L
kicyUHTFpzC/ielN9JcoyQJ4CrgTYB1qgY59RcL/vEpTOxfSA8EK2NIzagwYvmZmaNT5JqX9NdU+
0MkdDWuzPtcfDiWPEISTS46OBnfX1pZQNStCddkQgm3/u6HndTvncpyQQ8gJqa1QOnWVCNx+XhvO
jhczzITg4GTV3f+jxK9OCjsXgMVD8sZPU9BwIHJkxdG7NNLqTJlspNHaXwxuYHM8oZbjnQ4F1ziX
bWlF2k6Ow4LUmHeNrZkl/mnNXi4q3u4KOKm7ZskwQuqGFaMfzDCJSroeNBPUJRm77MDJh6GZ+MiB
Vk4DsS9ilwOKF3FdXAThFkq72CZGN2N8oa27RyJguIeGrjZXNu0fEKtYsbINC5cn3Sl9KIyz6auc
oWr31Hq9QomVFZQrGSLL3dJob9XCag7wLmOV6p+CK8FtO5u8+XiTHOZ2F5bs7mIaHg4ntrJfC6vT
pMuSB9byUPyUCl1cnuYaBl9ZCXSbsgmUrripJ41PK9yoTnlOGn/v1foQbGgzR3mbsmhptfltvh/T
7GsosHTymV50mUxLzMb4tZFTHLloF+c9k+d4cNUjbY/qr3zpC5Gx50EJSLMZ5VC1IT/cUqu4aFvR
faVXIBeJ0ZmUVJdFFLRqmMSoG8cLsy9bI/wv/erCDFK58aVMjW8GnW98+n/W6FDTxlH5PlXr5zsY
aqFwuL9AzLBYaSAzA++n5W9JDBcPwUV17E9S9QMrAH6o8D6bVNmkGsa2yOv7UbOpN6bxOHWBOASU
xdK4uF8gG+n42uF5bzWEsLYhREjA/3UuwGDL7ibEFCfHfUdojNXUHGdhQcSdrXsN3mZuv+T2jMsp
qj+A85Bgc0B1AOAr4K/xEpj0AO1Mu0EVn17IgO72ihAQmSktngHESdWLj4kAuu6ixAMcRI6DJ4QK
AgFdxeSf3OT8mQxfX5GW+Fpk2iqP1ugucQ/7ua6QuxvCi17LuOfYa3j6ETNlM2ZLb+lVx86GTRm8
XiZ/m6gdE3df6K/jOzpQIDDr+R/F0RQJI8VjE/BBX1Q20m0jeQT5FnWk7hkfkhNDOP1uWKDkBszQ
oXXInz6kccrHkPmgGIa66hFfoJgsaRQhLhJgBUwWYX73qyy8zZ+g6HTWCOI4osVEdEQWIVDRQS7O
JwOU90sbHhsRLMDEwo/9ZYqtH4AulGqJd/LjMXbzYPfYxQu8/PjAeMqL7lskGZ6jQvVoA2sp7YdA
FfvEwnPFuufPzDZOiMpFV8ehvkZIucyoU+fw7nkKvNwRTbt3Pqk8XapioPYvE5MDe+9N5034L6PY
UQPSXD2JWvDv56zAwTR6Srf7Q6VhNSzcwHBQ/ePCSvi/Tt318uyniaD4rEEBcsxAODNgyY2PHpF3
t2OZph8kpmsGYb9y0f3juqXpbX9VEE5/pfv0pdZxapMKRkjXadBXx8mCwVE+y9ndLkbBISfLlPzX
zq4/nh+dGYti9KO5dBXVswK8D0vn5hciPPLDBG0b5xn7B19PUGHVGg6UwiqCFnuY/x/hgyO05PfW
N2WcbRigXqtbSGWzCswkja+PUX98r62m6Fu7vfwY6QQ76khCJskAQQeyYSldy1Ez0aG5gCq0KUmR
yoZ1DQ+OTjDLozcIqdgDRtEIvsOZI0w/XbX+Pxo4HuzsZMGKFiHmrUn9U76V/sHgbX+2srkCJ1E+
ngupV8GTKQONIsjUGVitBUqSGab2SpG8OCI4n+4Ttfm8BrDE1vdzyQrGJ4aE2C35JC1+c++XQB1B
25r8r2e8GRCoCGZoPjkYkv85D2yAwsZg8okdD6Q2E0GxNPTuuG+iL83RZAisDSWqMweRsbzjrf+v
H7k7ID3PKQuSmx1hoYy5rb+X7z8HW5T8le9znFHywWiB1Q02vU5lWWn4Lr2dmnS/FNHC8EB8lBUF
jZocmDVHcCklZj6tps678OdMKa5mRvPWHlkVKSP0Y/OLryzDSHTTeEPuXTXKeuv7EFMRpXw4hpoR
sMit68PMpOyzVxWfOeYEpvS5oVl3eB30RSP1xGGKZ4ek+Tnsarl6JgznGWzSdKtiYeGL6h37G8o+
8O41l9MFgWBSiqU5rWluGX5K6xGyjZ7KjDp8n1P/Cxd2PnYSwLpEsJruWsoBwo/HR2MS7GfSyE1S
f+LjTUE0yJxkQAJhikuauBvW7VNowcf74jQLBFOH1RhEZqBRYgIHLQRPLh349CBQ7MsxxgDNxJHg
Mr67Qob0ZdbsqhxNIytXPwrVojxU2bCzmYDaj/R77pAe5X29EenVbZxRB6u5ko30cfNUZxX/G8fP
JoeQRQkvUOUDDjeSTQOv04dujWi5HKK2sXxNq/IhcRcPEtgdSGQfN8GJ23S3f9BBSvucybkyg4um
k2kHE3WSmA0v45R1znkEBmIrkN6lac0ND575DnK/ZURsl/I3XY/qd/jGZ2bum/XzREq/P8haQGlv
hODtfdu8gPz4VjiqefAIeC9AEyGsZnnbFg8Tkf/RGbZKWsQYKHg7u29ugNgXhCWIUEyr4delkrOQ
N6xrNJ5JYzIR57yEJ4dEZN72FTledRig1IZAMFSqbVT47tYY6ypET/tZVUUMUj4tcsB5CCRkp0tL
sNwScHKhb9uM6MjSoMSbtRs1bi+6m5fcaoGKxwGa8rI3acnY1GjIVIagY1HGfmdkAdW0QErUSIaI
PoQqDaxJN+UdeQmsd9nUaXT2oF2nVB3nEDTx56s3EJ4dc1v2f2HEf4taKJjHneUqgrWu5HeIHV1d
EWMlGbrAdNPnoXlEmKWVb5CAtEqKYhPPNrhmZGAzgfSLaiuo8TRd3qDOgOvfaIoLaj94HHKMdUXK
dqBfd5hwM3m8lBu3JsufgGo/ZGSuQYC/IWmhxl/Ese9BABYhnZUl/Gb+StB/ovdKa0f1xm2sbJCW
/xgS2uZZUKRLhrmhOAwpYUb0CmVhloAFTvgEJ8a0vSJ5x3A4N2p304Bq+Rna8ZvfmtSBiJvn6pKc
Lz1VSk7/lKrJ8F/DGJgXbl65IP7I8AV6T81A0KruIguiJmFsIZGSCPEHqIxU9HNvV68ZATsRwAEI
6N9JaVC95vcxUrJruC8CZVoLr81hvS3gAfSAQD0++4+0ZZHO/oHk/RUtITE2KD/LbWnjhGw312zX
TLRmie30O4r1yS9NDjINvYY/b8+eH8U9L988p0LcwH0mScrxvbtnON2zIQQMB9lm9fyzibsrIlm0
mCj6+pzDHBlQGk/F468azGwIM3+oUJxPTzdQ8OrqK6BcHytquUQHZc/78QWUL8oV839dM/S4Cqfa
dFmjIkpNzTalY6NLCr4/2H03UVKR9UE7tKjaiVXSIklt2j//T3A5xiHjDqLQ6EkGN71iUhX6ON3R
KwoGO7OyB1FN8HnUbSCkpEucIQ6ccQttm4GNbXXNnI86vI9ZuePBx1Wdq7sFN2QL+1wKCNVpsyLR
6+RN+OFRRWh8xpRBanKkzWIvS6MCaCbcup+ZSrcpEWvllJ9OVDl/qgee3C4kik9c2SjlpVIUjC29
PzC8HQOIOrB4/6/EELi9px5ngBlE27TRIISQOop86nrJW5XmnPWIsMo2HdNyNMPGA0tw3mvJ+brP
gCOOjZIh2g/Qv5xrOeO61g2a8sYPS1lxDjZ4nNROnAg7+mrVIEVouqQPIF7TpR6iHn1nkMQ0D74w
JDmwb5A1lM+MPyya96fAAkuXHWwrfQp1TOwuenwQid9o59HUcK4hB/1IWSCnpheVZKzMfijmcNSD
Qaz2yyjIsDZQpmQ9IsNwNlwObcP7QIjk4AFW1N8I5PT5M1YCeGCPbS3XEsWI0zOrLqojoPzl/C8W
ugqvzJm6NJTV+QuBptjGDJS/MBhnmpjBMCj+j9MMU21UUF9syZvCx4gDsiahyYXXZQlbNj/5wOkj
yppN3sZp4ZPm54HzereHhHThTtKf3sYhJKgwpLf7Zdjjjqf26LZYiWFpf/baVmQmVP9KPfYKstjw
XKW1bbAiiioGo3KsGDhe7bmh8bQaiWIgZO/pbRDL5PPgXuv6CSaCWZwrxTDcMAU+XR8R5z8K88K5
jgqRU6khvMFmul7wpN0Lm1oqbXVikSrXIb4RFPCtY+0ZPdsti8nr24k6g9V8M/Fln3sWGRdy6Gi3
CwwkwNYlkTVA96JfFpiMOQIs90K3jvpAwcqmZoP+aScXfx4iL2v8adU/NidkY2dwwOMEUy22cBqJ
9cA12ai9muflFAbWZ4a2K/wGhGQdQ20SKhgHx9touHgpWpFHd6Yx8Wkxg0K634vwVKVlFymWxrSP
C8XGx14OW4HjmIwjEDDU8kjqKuRVoJIxDvqIVC30X1eBAakgPeBHV3UCYj1sIFsfud87GTmFgbq1
ZsN7J2WlCThIgtX0PI9U4x/uPFz6tf8vhbnn/RtuVaNHXbwsSVdYeerCRjwkRNydpPoIUPQwqGCD
eOAg3SiWwPoiWRYi4doY7rV9Er/9b2G2Pge2S6+PA1lztkL3alcuInv/hWKWeV5wfgR4fMPevMS/
k7tVtzCUT2e8VWPNvUsVem6JHf+a+loQDbi/EhH1OIfiVNWEYzUfy524htCgpeL8+FPsqEkjZw+h
i4cIcFP0F0tyzJs3JJPacJoH3faEJOVCy2IMgL/tgyLSbc703XEkpqgTAz+3EiFYKTQPLtHA4Z34
Qjsh08D4f89fkvGRuc9Rhv0nI2+Tv1dkKx/1Td47UJoQA1UvjtmikcHU1fUwKzdQ9jeW8LKcaDLN
gaFXgvQaHlVIKqYdYomwHs3kKuh6NY8byWzlonRouVvLKfPuznomq1An3rWNEJth+cNjafUxVaxV
FTo70v+lquUF0/jr1D9fG5/OSSce2w3E+YzThRUKc6diynZwio8gD/ia0BcyXlTlGK6xpRI21wpb
opQSQfs5S1iVLzc3IpsPCruWrWRLbQ9vuYpPWbzYbR05GmhbZyMJnm4u0U+iZVoOVH1GmpLj4Kv4
gjXrdB3oE13l0ix8tlJ4GO8Hhp3AZdTZ8YeajrDc48I5z38pI8Ur0q0wKET4g4JDP43cRLtghTOz
jqkRi5t39q3KmKUwUL6f6H6o+QhR1Sdw2dGzLxddr4TrQkiwDijDHWSC0vMJC/nJWoQ990tpoL84
9Y3GtReizl0W/jOWDw5L24ROt3f/q9tVfluPkr0CJUwgm1ulEv6/TcOBvbN0FYgcDwjANFwnosql
MiwT2ahwdQOIpbIYMxjDfQ+W6W2AGpeDcruzNftkclULEcRpSmulxlwh1/lKFhMTdO8hnB7zNqpe
eHnJw1HQRm1n5up83DxDitqeh8JMEMW/rjP+NIhjPKljty6jkSf7+mOqASu+BOmyzsat36LHaPQg
Z9jQ8CSCTYYiQH4cHy58f3AUjFJLMrZf9bY+55tLU8JIgF9VENP/G60XGNd/EfzyOWYyf0HCLthk
wOLQ+eldJP5xCt+BaV5x0JwGPV38kt4I0/vJjDq45681JyfuqAde6yoi4Q0xuAHrXbdauS74VPWa
URf78vw4sOMdRFoEteX1sgVMAZBP9hszmtz53eRChe5Xq5HSNAJOtVO90jin0R6MX6Sgai32EeHj
H5qbLrIc2S0gYNHxSdZK7delifPd+23QqFZMX2cIPfDlRxiW1qgH7RqeGIAjOGUhJinl9+4c/Knt
5agzGfD9e8ke359VU36QnNy++GhTOW9Ir2EL9iJEI/MvhBaOOo+B2IV9PJpJfP+54vLrT7qrmnQm
DTzZOFlX5G/TDd1fzILJlzlCU4J094ETUqvBKB+Cfp9LgXfXymjDZ9rDK1nxLWXpkAt0Iig72DHX
kyjDUq2gKJqlb1lLVD+ltNdYlHOeoZGahnB2v7W6QktcKMLUaA4q/kxZ+FNcPtKz8wBnBLKFVoQZ
CdrExTKp5dLdLhUb+p/ATLBkWnaw+yxA1dxzy1zhKSx6MvKvb5Z+MgxXOFGoOVs0sAwp/L0E9s9C
2dgwWQCeJpvXLHM2XrG5wvsxlI+7fIfHwnRFdDKwI0xUu3vCnCUlnUAMqDVJSURTiB54KL3DTimT
OgN5wCJ0cj6O2tyV2aLev04CKnJyH0Rge1roy93Jh/uJDNsjxWE4Lsw+OSyfp2nHP9QUEvXhX5Bg
zNnjEguh3iRN5DiAAebhyWm5LnuB/3d4zvGPYM1ORiIHP8OqkbgAhhhxhSp9qTB4RhCsS7LBmtSX
OidFIrmompz0M1lzBnSCsMDcWySpgUCaDw1JXBYUr0pt83hY1WWwUar58HNtD0MB/+aG1RJUR1yN
z903APoWc7U58BIQyq0oUxIMcRzWYzfvTa/YyZwd5yMYGTuPbpPkfMXgr69PMS8sCkIsczjM7Cph
xkHVZl4MtqmRzMaYd1zBve8HXxZscygBKsTL9C8geQ4q3WsWQH/PIjHVNZ7u2zG81lgK2EiOcH98
Wl3+jcmtj8x/DBVndz9eVnw/sqrnGIZCHsPDY4xClLN/Fwuk/SnW947YGpNd8mSOuP89YTu+mdKG
5dm9N78IMg7SFHapn0zg1kdQbU4F0Sbnj/c7PrP2L5zCW7NAJxbh0InQoI5q4Oelf80qJYl5mbHg
Umeuz5nw9AuRUwQ64n6QHH19866imCepWIsv9BfM1DbL4+hCrMKCwVowKbBHUm61FejcLEQ5+Gyq
Lz2dChHqCFZPB8cnpn7vQ0qIpthM8/k3WSBghEKVXOGrM7FWq3V852Zm2AABJFF+blMa+XRHiXAa
w008GylGyrCbIRtQPUgJrMTipdGp8X/sSX1Be3jCsyZIpDN/RDlvbwwPizUWLuoQ3z4ftD/TG9Nc
whq4qjhK9/8sg6xEjSe2VGbX503LJp+Gh0HLByYymQvGNuZdCCe5AnyTGaNBEFe6jg/jl/jh304i
pFemBUNHz9Ei9rCvquh7+47JXLLSxRQgqJmReabVr1+iE3BVVK9EYE37DoClNy+YU+upQRuQ13ZS
8FudRZl6vLZWj4vRAqymPCnrgg9YEkb43yZlqVwKJEosP1q6gh7lmPATxBPmiFYAJKLdvEA2P1QF
3AcnP98BrTR9pL6297K8IuF1wPSiAwnCGT0dy9BuZWeRSojsHRTudPTlFf6ZQQde6Gz0unqPQ/Tw
vW3M/dRlk3JUcZSEYHZA13Q9ZDlE380Y3sb7OIVdQIhpcKt8nvXrh1E833sTIfl3efJFIfPXZ2WI
LNA/htlef5E4qiSZQRU5geSHwBLflijOSoYdk4l23tgO/BvFVLw9v+UFNdXkUIDnhcC5v23He8O6
ypE4Wy4AZHAqddeksMYLSlrZolgkl1mbKYYzBHpz7wq5pGUf3taTkceNXKFGTLOcmNehb1PG5OlM
H5nWS7fG2jV7WGinyqVUIkveHihaggneIO1c6DkW0T7+kAa0LX4Ws4JOGnIdZNzJWt991Vcq7GfB
tlCyOKF3pPONrrvLOMJxLNI1J4oTS96X6mL02/u0juQcMEF4bMBDBflFrV4fjDKqOA1PZSJ/+GWk
w95lhoOUlR8BlR9t8M1jeJaSdJfNXjIWqzBpzLi4iJihkd6LVLUrFd7FxlDJGbfz3iVVCp4c7bcy
O3n62F7UYME3NeQwwXRIsPEI9UsPrWzQQEPln9EDj9tKDL8pwqYj2gku63cDNieOJhK7oI/3AKFj
iiNfkeKIX3zPz98A19fPP9EEEen8Wr2pCVRUx/v14RdRXipJjUGoBdFZBIMSTxgbpjSQd5o4X/+O
Mrin749UXg0JaLMuMt9AJV7quNodytBnRdDtfrnrLqPucGUH6GyZiqeOI9R+/f/6rzuw8bbxt0B0
Yt9FDucq6MoYBzFCwpu896Nmn4dfuYOrspLDxhcvWi843Javtp8rjk4WazrFxycWKkq5Xn0PAHyv
LAXB2cMWlnyY5fCaH7oLjtaldYufaSXzSw+jt0XBNnCAAMXyUnVg9zGAh8aRb63z27lCwDKYrE3g
arJ1gVmfN09CwgZynDQ43H2KwUB9KloJTxvuLAaTIAKkDAJrrM/7HMmshA01cXxEPCvksEu6h2EC
EAVc3kfwT4mHmI0Y681hZUGmqLy49SnN3aLkQ7T4Gm6X+wEtPLdPJ1AqXJVU5Z4sBmBWfF3oNfk8
pBtlt6cP9iqqghrTzEeB5t1/eGKyC7im2r+TY8p4Y48982iqXTM9YOemQtxTIAVLyC0TsKAJPG5q
iX/4U2VFPEU0uuVSBa/Z7OCEoGFU9Be2CDKcHV6dFTbXJKzwTz3wcaVYRDbQkrrvxU5NyhBbfLXA
oB+zIm7iiqZQ8Gu5dq43diMmIJrdDTj4CfH/CASPGKzX00g9709QCpszepHMw6lsYz9Yr5FFq+su
s6hv4ofNsosTRyyO087AhjUIww4m5OoZzqbryH5LHMSY5JdvosTD4/YAHdVAxwml/GqdAiraTkFc
nr7M3L4g1BCH3QbekijpxIZVeNT1cHNd7TlANLXvOUKPScPu01ofPKKT5DQaYLJm0NpBo/X3iSFs
x5pNqLpysfJIgo+EYdl9oh7QXFPRrduYrqBr76uMjp7653AMZVmTc6g9A6pwKKgT/ZZSui/S/kqu
x27kVUdZCBJbo+sRmuu3ZM5h7jfeOQ5ZIJX7rOM9BOM71czzNwJgJQcGvH3LHzoxQLlZOCI5n4+H
HFcasb1NjJ4dHS7F4pHxFln7Ukr8WyNTfb2O8LE5h3VP2G+Q1U0ReCBLOznQ/Bk7lGNC+kkub2c0
qQ61njovRQSTug7slof5MdAB3Wdrhbcu72bV9PCdQ0aLU/lCUdRL3L3dE1qfBypYeX0pby1shgaN
t71cnSHRk1uIUsa4oEZXxgWfnb0iQTCjPbHzkizSr9HvMOTE9p30T/nAGZRkS6gjrEzr2UmZG3uo
MDYCtLgaWnB91ak0pLvsx/es+BgJ2e23lTQzjQtzYGvo4f8Krc4Cc2zHXKp4iFDtZXMVzT5f8AkR
XqM3Q6LFQxoP5aWfhy4WunS5UO5ynLaHUil40EeLcn2ed3EMsROtr08FnFDNcRPuGDSKUxhBEDve
HATqLNmSf8JWPorTS9zbz0iqAX5T2+AJ5YQKh4Cnr2bxuP/6CqCszWh955Or90O24MunmpL8YhGN
Y/jJQ94wQD+pzHAluWEZFPnjHzLQh6KgtTWm3zTs9icIJBNyTnAE7Jo2qX9zD8CInNxpWGKNNbxH
IcM3734qeX4mQVnqpfHe4ze+Zl0dc4if/EmzTrQIx9VeY453maWggGp5UBfvWsYrXuM1gn2FdkXb
b4iVY91NQE7emLIZMk7En53T72UcMRqFDFRSH/TNGJvuXrU35Ygl31oHbCS84PCK8pi1BnQLvx2i
quOGiE/iFrU3mcecEkzkxtO7GXiAtPj87wZvShehjhb9AK3d/y8134/uIBqWEIOEX+Br1sDRFHlZ
nlOLs+BRcquZRzn90kl2CYP1Dl4QNYRMKOW17whWYQa+up7BTCu5bZZeYbtZRA17gSIwkYAWaN2a
kqjELoXOr5M8CYO2yQV9dGjvjQU5LdRmLuwH9ELySWAxk5gRz9ozDSGIZydmMgI1GdxQM5J+uCTO
6lNdWEksgqTetjZsQMdRhiM1q/tMhzUdBTbILb4MThFjZR15xas2fZjqNQH4KdZGLLa+18KRM2s1
u1H+D04ThwUyQL9MoCYvDHPVGOeMB5XU4xpzC1E+quxRYoH0fmRi96jOP7CDt10V29y+oHfIdxiQ
Hf+UMS4dOWfLEdrOsuZmOHHV3vnwdJ911JLu/45HU2M94A+nyjcxpLc+DvswFgaJb2r3t3PF53Xa
dqgT5TW32tzEe/2BUjlW8V9Dlmv0iGJGp2xpJeKjPzIWRq2jr0ZHzEarhRcIgR1PsQNttgn5tnEB
Yzf1OAnnAUxmEnhez8uZh8r9pPTJ1M3gTdpMzDmRR8JVy8XIfvo505iSHzdKj5kjnmx8bMFg8Xvq
k1dSK6I6Cp7PCgbvPTcJ4g474kzqdOfUqn+kModl2ouEOBvwnpAJj+BTaVd2FiEsIF0rJ8OVW/Ie
4dfF2gEDJGYuOJjy9q8VGd+KyLFj53oCf+OkfjjdW/lLTNmSNBK39XSYBPlRXizTB/fvN13El3dX
kUT4+LHR6GOn36LvQjMnEDu9+D59a/H9mUx9x8g3Yx1sI6ij7CuXr6WQleneMURWQDq0Fgj4MZXn
I/GLDveqw4q/EXaE0cuWtwARbpRGAdVq3mvcMhLG2W1W0JZzLbn88ykvDCNc3YSxOPqKwXZP4kQg
XgzsrrZ6eKb+ccUixlcSMlKAEw17/3wz6gvFWSsw/pBZXvoNsMcawdbVfFnLfQ80GHPZ6eyrq1Up
Hvwdw0Gxu05/bCba+MrPSK38Kyy1VgPQ3C1CGJYpmfJZCl6EpmK6SLBlZMbiXKi/Cfd+vgUX5Jfy
jz9j96FJ1bkvKn+P7W0ynGZP9NaQ6Hl2dNa4GTCpcR2EOHBnTq0ixgtK2RCyNarFt66QtEJrT14J
MoV3PAOXbFavNC+KNQOMwT8c7TvJIWUlHzQsHmMkPTKZXftUrhpIKVdJNioKAwjzV3jBgr7fNSjv
XIe+xO0/F4dGI5/zNInEwxbgvo4UL1tSXZ8ds0z2F9JrTjGk7Cq5gt0sbnXSYEjtIE8CUis5jhFM
iY17gSNDG4kbcBKqQwsmdAtFv1EQbdbY9nYsJNG0ZamxgSNdHnEesAd1UZ4AQ556eajm14IjMzY2
Hlo7jwaf1Yhui6bXAIQ6Nb/FA44N/aHijI4VZhYgdVr+XS3mh8upRsFD3af82e0qwrQsCZemyz4M
PySZPaYTy7RETJpLk0f25t26efwJRMgGMvIMxgIFfTbq0FsQNMR5y7iHw4sCpYqfLdBkUfJMl4H8
mY3G75XN6shH7ABiK89caTwQMkwQSFRCAbvy8xUm6O2m03zFXuMiHFDRkxyl3bYbkE3yAa0YJRxy
8OrhLE3q1htT/BjTcsqlCdTqc0vFlIAWeGfgzglGVdQcaR5j73bN3OFLVlEicmTsgpnrZCuQJQqN
+eAc4YZXNliOHzyQaAllbRT3D6Nlm4Q+e4+hjynayHnJJPxwQtaq0Wxfit9ud5/B3WCJUlhi2Hxw
WcgC1cN3r1fR/jY0rVUU6w/RmG4y1cNWqKIoHw1i8fQtAU8qzvUiSO9EB/YLyGk2N+hIxjGm2cIe
b0tYMEd5+oVXZyDbwNxkwHRziPqO2EV1SJnLUFRdoJWMbPLJAtvwAxvTLS+WM7BE3623yqd1DWlW
9nN7dyYEzqrx/t0bFanx1D1X4EprLqpaFxxiUUi1y7MBPO16b2VOdvow16hDy0wS2TcnUDpySZwY
obKJmqOMp6hE4ra12u/J/lXehrhmi1p3VyCBaxYWouCK+I1stkBeUlovKsfrsafLDkz1vANER3J0
pKauATBOrXTDtNrmKZG2NwugztbeaJPRuIzQh4P3GsXbJJHJEKfnBoQKtE+arLPHAa6d5bBvkHmb
JWCpkwKQnFzJ8SSY719AWU+EAZOxRZ1ht93z2C6Jn8mMIQyo72hdEXmU6m6gYLdxva9ETyHPTn2w
AYB5F2ZoIMQWboMaS024/ZxD2295WCSMf07OSssfeRrF84rIJbWGskA/DSiOymxEP7OdarflSy23
4wsApnMTYJ56d5kbvDh3B8vkfW0dH2++yG3/04wwSNiAJ0QKEOJ15ukEPmtFrylPodOhHXkwilH3
VRDTv+RGtrZAx7+Ta5vyjXu4X4AN2BFauxOVyOj4h9n8VEQyV8YeOC7J6Zv79kzaMp+pfywt0+Ib
5YUAlZALJF6/QJoKCM33GxEs9oayUNxseHmzi//gOlxCNeV5yuHCqHBTU51TRbGk+ncPtG/7UDRz
//fkwEU9XyyLgA2WBoDzcahRqyqIZNZNu4SZFXOAkOzts9mUNVGO9NWx0YyjyAv3slNOOupH7Y9m
f4WLxGAM2BWnqp6FH0QkZXsgRhvbvh1h+Wj+AVvhgNQ9kUeM1EAo5bUadWaC7JL3zB0qJUgD3IO2
CZJPiQ9NTEBUxNFb5VsXnx5tbaU+5TJYauuw3B6m7D6/K9xCE8A0JegpLaEGW8p8bE4tMLHhRllm
+ag3y6qK3O6Xi1mMoY7rbrOBZAhMOa2n0NW6lwf/e6nOyyLBW9r4RLsqmMjwop5Xfe65r1Oc+WGd
mOn6JEA6W5WMcIa/fLWomBBzjdGRcQo0BJ2vkYH1Cez99zR5CUxgVFajorv1e2xw2d58UrzQbspQ
rQ2hscPX4qj5pE4zxGCq7pOi/NUEvLB14VZYeBsbQ4lwEQqQegvvW9ULyy+dr2vL95790MPMwXUZ
8/kKuKY9iutRO3WAz7zXQ0qtuyUIwM22CFOjxpU7i1nNCHf6qKK3QsoGhqaP25PJhp3yvjNB4UJ9
LBJro+RhyxhISBoyQ/kdDCwEvX/8lI1C4gqZiHy4dxUSrXBiCOlM7M7hwrrs9k8E1YgVruNlHnQm
cmtokJNJ4orsuVo/pCqGRfQyokFiXVlA9hK4BT789nE2P3MRC4QN3vqCypRB61ba1O9oo5FKpdrR
w7lwXSDurRwVNbv3UA6vFwZ2X9tR+woyWP9IyYtZVflvpI3dsbA7XNAm7PQBqM5tuSueZlDi9MFl
n87QDgaEbKUV0ufYTJWB5EcrguYVfQoaI/PQF8KgXPDnOtNIbWKl10A72Y0hvlDZtUtDgH25yylc
bUOtIydudDw7FxMI2lMIWkqe3m2VJ2YT+ISj93vPNd0AeOHyYqDTBexy4NitMLjIS/97QcbE8lRw
WeKU4MPNjQzujX4Kre2MP9uYl63qX6LQNo1Xj9lxCJCPSSZCVwqnPCC8/rBUxjjZ8Y8ZcK2/oFa8
K094jEDvNayVn5ztbA42IjUmcnQvDTOxFVQVvZ55exuuaZqzJXx1oLdNJM/qxRA95ivyFjY7hMQb
8sU1+JYRh9RJ1to1dufoeVYf2al2P4sbY7PvogLbBCphERkx1vi6bkF03lcKqGlyF7m+KtBfADtL
DWjt/+0ScEKvDB+j4M95nKhopU2B00PjKybX33hqfoa/qkpIBVdCQRA9EFBdPOj772IMa9VNkS9O
Qaq6MHc2Zv6oaX0T5615h9oswdMnOEXrSMwYjakhh7WcNvszRZvgUIEo3w8NKS0Ql+KrfROanELW
v+r55KT+4q1LW8qCQQS4O4rAs0QI30cuIlfG6mcF/5Zf/NSDrwY2PAbXRNwRnyO45e7UiBdsKMPt
RCwQgkL+zoNwqtYAu6pITJ7/KR+tgI2qowb5FnUDrOGYRlkOP5BndjW8sFU4KRTY9pT/NYyh//kL
Y8dsROlAQXES7B7O/15ZAJKYXZP/WbHRSQ5ej7Ga+mervM/Ws9+4XfZpPg+KkWDF+xPI6bEQUjAH
6CopjvbSgoQ7ZCDYRNrtcYH6pro9T5HgmvLrFuE+0CFcut98BLF/q5CutbDPNFmK+/VURTIIgyxh
+tmNl76TOl0/IMEghkIRsAatmYEv0GAnJYePwY4bgzvcoaAn+1xrcDVRxAOQnFTT+328IOV4BGOh
Rb6MUxlg1bay/cTORGx3ZaqDcVEOg0R4wEC5ZOgRzeCE6FwaRsv91nPGKkdLzsOTmr5TCyalRrEU
df4TWMoMfmSkkvieOJb9DhmmO7eqrUGCXfO+I7ZdSQXIuQ5J+QzbvtS9bO+RPbq/s9LbXGjFHdYJ
tnc4KaME9sG9GYPRFEpgD9wiYhMFmtS8zyCzzWwnBNciHWf671ck8ZWEs90+jvsIpglPo8xCfyJt
X93YqJ0kmUhanxVlwW86fHRYDMOLuG/N2VMQNup/IpSNKE3bgnlXXqIpPXCSg3fJBnzCEHQ/W7H5
J2jlcAwdQny9a8TwCTLZJI+flWyHc/vlMPHoB49Mu7ndx/pkHuOHpzRsWbARLna0bCKnGVk1Yqil
avNuwycxN1kvcIROLsujyu3D2i5vY/9m0WKRHXM9qt/Azh/ycGwWbo+IrJNqpm7pNbVejuPGwTZy
DT6RCJfBqZupmrqTmYTnFPSbWqlUMB3Q0LqrTrXg63WSHi7KpLuqzGms0loghGarLIJttYdTfEDo
2622c0tDAiMyiFMEGwbxxl06EsAaARrfnuImHPKGr/gDIhneABniQULvv21Dr2NVMlM/8gF1iKpX
UTxELTbrRC9ofd4mu5dLW1+YbVLqz82wBzxFEJRXL4czV7TaeBFZZwfBFbmbVPZZYXqtVEGK8i00
Ma4vYM40AEgJL/Mgqx2tRzVkvpPrVtBK9M42yIvCOv3uQFWTWAVHtBaYKB6BEVcMPhQUWf2tJYrN
TUSJe3zA4/t5rHi59xb53q70/7XComTszKJlm4lXJBMQIbTHj/5GZVGidWC93MUok8GNxk8FYxM6
Bfopj2ZRL9M7WvQA9uXPCeeOm4mZVJHIAz9Ax3HGoBh3am4gkZ6ZZg3lL6JvRvrxLMOzpOJFENCu
4PIBHQWGqMOle+8+HtxzKYlZbCHeFbTQBkp+jNFDuz2TZYQTUpBwCYtkv+XXaN5VcuoJNJj5uHax
of6dRgqngWGkGnkyet577kV1rDB+VQmHCdA7cb2TaagZ9Oc6vRkDlnQBEuv0PMJaXsKeiLE5/C92
eZgSBvuMwvvOf7ofPdi+njuaqKM1RLuAzwI+QJHTmREopEnB3wqxhd88MSaoFsW8iVasbRoNPY0v
TbuktivkPCH9IygtG5XZ9QoWlMJKOJhuyCdKP3dVMu0iHs47gFtlxjGxVhgrq837WxH0EQGkfOEV
n4vf8Oy9y5F9fuB8ZrMXltYMZCs+ycvlkHvy3DpdX3GksyGAjrTGD7wGtdk5/PQxtzbx8G06tld1
DtpfO7oQhdtfKdTZpMxor4s4ujhI75asUxA4lCpHeEgGeJw3oqMLPuxOGMdqkGYaHP6DzQib6EFk
wPJJaq1hk4rFg+M4VAmmQ2ay/8mQaUFXp1kc8mjSMGfLuXzalZu0YnrZiz2sTZU4K+EwEYVRZrV5
eqAp5o1MTzzlocP+bpeIBz9I8H60BupGOdxArfpErv29ydPcy7ojoFpm5qSehOlv79NkonvzzJcv
C9r60rjyFCxBhEaY0Lp0bfxOgyaOEcLDFUIxLWnChiNfa38aBVSaFwn3LofSd8rZey+YrIjNTr9W
eptIENn5ifhEWGOYghxFsHYBykpIpo5lUPc/dqMylW52STLwIjMTBk9wWhQGcINKH/umq5XjApv4
8T8F2MUuzilC+davea+HwObYawVYDhmndwC4x7Zl4ec4DCAftCk0NjfkYAIfSp6Ek9IH40DV+W2j
AeG7mDq3k0JTxe9e72cHPkf34glisvurVd9GhCv99vKVnpRE7QCinV5qRGasI/j/iFPPDWK4gkW5
35f6XZ5RzAaaOAnDjhXlIQ+O6MA9soOWcMCIMRsMRi2HWHfXAdKjkDOGXKW/k5kDGcOGQxEb8/k3
CfyA0UFDbjAXzAE1iPXr4jx+s1OG4d7Uj4tALYglz3RkUP2MFA9zgxm0s5BC14UFhal1H3xoY1i/
AfvUlqFSQHV4evQ7m/+TvC2aERlbeUIv2VCpjAG/lQj1ckxj36r1y0TzDETqQVnhUhIVnYsu32bv
TdXb62nuh9sYa+onbaZSusJEdpCzaopFUXBlUhau4lut8lL02XLtFzqeNfPkUAQ+LpO6oOEZpKRn
BdFrSEI+e6v4YBwWkWAKTBCcMmDDjGBsoGUP5DYbg2DZZ9kAxM0fYYG89eIto+Urnj5h95XLlDfW
gzRkmCqUNp2wXbJGgMvsSQDX00ahmhWV+VoosE0sfd2VdjqB1pio33nn/9pURvCPSbzV2aPHx100
yLmJUt5SnW+M/sF4H8TOfDOj1nzgUqLQg1Obm3sts7N2W9QxkHQGNWGw/sIBjGFLNYbAPV5VNN9l
FVSYiQZ0FBv4/ixd/k6ulZ0Gq+7UrDLR/bGxnM+G6UoSUspKxxNWfkOiNGojdYfD2h5ok+lbz+TY
sOp8gjF7UVemVRj5RGBmQsV0841ApLRquRm1STQP3z/fJcMt7xp9FQEIv33uYcAeFhF55/nBj6I0
hVKSvomj1PDoYkJKzW9MoOqfpmIT9m7CSnQyTRUYEolrCcWVKyjiE29Km78WfA1RdPzt4MVxo080
lhQG5uOZuH49FI9AsroW0Ydj6tVAffMZg9PrbLMMm0cDBMjTHTphQW1QjSQSEJ3VJh4zN3oXrKVh
tI2qCFhI2B55QI0f8ULsEdvPCN5lA8CwFclP++1o1HkCmimf2BI0v1DJ1ppgLGjvFQ3fEL2vYTNi
Vbx61wv6CqgvCaqaC/X/14qKUryE+X90kiM7jY5eYam0DVNyyZAApfQBswzmIP+qTPd/IdOni1HG
eB33l8WpTAZB1hn+9sihzKD5GPFuF33Hr2dnkwZXy5tKjucibyYpMdEGRbGjHcGNLeuR0CcvL0Sh
hgeoV7Vk+8tyH1AP5KOxj8P3PQhHev9dhnOTlZed5ojvVxdRXHPJ3TLyr2ofJhJ8nIWJey+adeNv
chEgA5L3P83/ifzScUt4NWVSWAYUyLKOFQ1+hL+4mFivgIlIl55eSGxtA1EDDCpi8cc5uU9fyopt
hlvyodHwDe25Y/NOGAgQeWFU79noi0DLPdZWHiFTHZOskCaZtK01r/eZS3FhkqE830fnzFdO1lBl
ovJVcc/1QC1V2XnIKGKWiLghXJtUo7TPLSJqDbjwPCSiRpP/2VAk3J92/MinWifYesunbH4bt3ry
3vtNxZc+uB9CsVN+vFnnpX0Dqwh+zSEefVMgykIW3QaeaetDC94A60MIPlwIeWjLc+HwpPNIUZ4B
hu62n1ppzzyaXh3Wgr9I+CJlcyyRMFeIGOQ6K+v+rIshprNHELFwZ++rz3LjteLcQL4wlvg2q1J6
CQknPARNI6Un58zbACmeHuPfyLqKiguUIqJcgRvqL4rUXJOPZtdcZ4UZR1VGmbWlARcMGPAH5b6v
QQjsr/XmukfrN1d+D6+1TBPHcNwI17hIDIYD8zUhbcFuY2dlUK/N89jT1rsMQLFmEluViszJeUch
aKHg5UOBRe6f7RaES8jckLvykzZ/luDrxPYaD4SZBLHFPAw9Rbe3EN1y7Ip86HD0+UbxkK+RCVUH
1+TCIi9BZrUnWelFGJsaJFB5LvXTm1YXi0mlWvaktOY0A/Blg//enEpfGdbuznFSq+5lUurJu2Ad
dR7Y4ui3rOs3X/eocoA+n6kBhiMyVVWQALAEr+Uq2KEcIBmTSAJKlsX5oQ+eWQaaLCrFv5NabnF3
g1NS365AKar4pARdzOLOgfTbp+0eQqILRJdVFE4QQlSlGQbO320JlbqBkmmA4s5ccVthCbV4a7gd
6FRiyIyOFe6kdBeRvXj/MxU6s8wbUSGypu7rGl3lZ+ticJqxWN4U0AGV+S5gAdr2dpxBmKd792rF
4L+pWI1DhGWmrjk4IJqSg5Wz5YGedbUSBsYtQTV6HMla7IuZVo5yYU/HiiMyS6vbZqm8FIzP7Gl8
3zDk1/lGR+PVAHhf079qw8N3mMAFB4vacZdjMC00JQp2ZCTWi6qwl4S1yTXVsoFPHEL7mMhv8zW0
xMumyKFlm5D6q0Cwjk89V7JhR+4YUf2KIHjbiVc0dhTiBtSvae6CmhlgzQ1a4VbfURy3QmLw7/xt
gecr+2OllSQMNZyv0m9Xsyed3iVqttm3ji3imAnP6ZgJfK8j+HWtncnEYWUfqSRdWPc8EwaxAWBq
GFYliLx+4M8DmSu5AR8gKT8UnmBWowzYPl1UIOzSqsDtw/i2Z0zvUcBzr3ciYGm5NHWsPL5GiENV
bXSvQeIuX9wybRKb7s+NFZdgLODdWpCnl6WuyGzPoZcg7RlHOGd0kk1g9Pfe+rZdcViIcZYHNdHW
JxVpRPV6d+ATs/KGuEjC0/iw3+EzkLHUsrcpk3/eKG8e1LHWzOvKxK7TTSOn9JrgIqKIy+tRPnjw
1np4VKwbbYd6Od3aRwtp7lpTAnmtqkcBmKQ56Dwl+d7KDavVyUXzviQDLxv3r5f3X5BHuIXsGv12
yGFCqwQPDBz4QtrAtb2gFGKohwgmVMkOd2XvJwOIuH7VA1VK4kIY/GJYkf1sE51R7feEtj8LhlvS
J0PBlp22TVYO+4YG5yCTVAajEE4cy1oWtmuON0Bi6vkVesYCf4eTguBImKzZTd34fNTh96ntOI6Z
7wLj6ObrwzyP2nIY97s2lTuFzHjlYW3G0eMB42zE26pu8srPVayTNwCLx81sw5zmnMb1N+Gwzubt
Pv+yCAnWZGBQuhc0bL76+cyHc3soGcZBEBOVvexvHSAr35S+vzCppNIZeH03YVCidIANyAe3Bp5+
OukEfec8sodoJGoiEb9eATpF8Gyxhg4Eq8ZLJc5YTtPx2DdOeLdxkeTtNIM+2eCSi6RkkYJeb+VU
8jAGofEJ1Egz580yZAlf87adzYPwH35ptZGDDkTEAa3tfeIoFVj5Qhn0ybTWKUqp1dNlcKN6M2D/
39xIyT3S0qcBfjJE1SVEkM7YO6Q7FN5B5/YX+dVvfcRijB4Xjw5oboDV6wd76xIUzyu2gg+Xo4ha
YHEaPHeRK17HL4gY8vadE/3YIvBEn8ZDANB7wkMd/xkEQxw68L3PdP4zI6kjaI/QccOBcbg3r3HE
+1o1Y6/QzJfmZXURyKHaH5V9Fo5KdcfD2GqC+j/ECq5MOr6D2Ahldhr9TPkQ51vKgTMxowNICtaj
yk9KGx0JX0Y3zhO4vCjfYtQWCwVGsq/jwmnS3lYmqO0PwfJNE308eM8wrO28xddDnHdgtd34Qd8Q
PvD++z8WKBSZQTF8vazxd+s9xvsbUH3ApWZqE02/0Zay8m5wndrP8AGLPb0RgjUzwL3ImBqVIvs/
slW0dnamnQSgrsBPWxHv8WgHRwNLHOeiLmZ6ot//yNfbr3nxhdrQIlr4E8gGvs8B54DPr/4XKZgQ
n0P1DQ00HLGO8WGUI3bed6iguEh2zAm37Iu5tELEuXEAQvuaGFPwyrgFLvptFyL69c/2Mdl0HkAb
bxdiiFwld+B4FPc9yDJtKNRi4AXhFiIWCq8tNQ8HwFW35IytYmkVjFiXRO9utONLCWOiNfIJ4Vng
/YxrS8x1DDWNtNY8Z9cSDP9xXlx/5IZbskL5Pl8cnea/dsoBu+WYtMeH42wrtf6TeF5hWz+Qem+W
AhjJTTpbMAlCMtY9Q+/KchIyCTSJqDr3q+yx4U+5t9UoK2kczmlFkm0HKx+6baMsO5cVWk7Bnx53
Nl8lKNBNvXgh4MzPs9uoJLNz77QYS2NdeJDU+xx96A1ELSC0a4wnslrUAslDuaU9U2jbpiifxWxv
bNkQhYTdwy9DAEvv17B8AtvldktcckYg4YOnhq1PeVhAXmATuV78I/3Fo1YyO69cYwV/vCfZfx68
fb2n/vFxMdw87qWrGtC5kAFlfDZdyBapS5XR3PUrBl8eM/oC3dGJcSoWjYb1wbHet+EkQclpXZQ5
UiHlQaooHwR41T4g1jkkdgH1ARfXiCREuloTe4pE9rt+0ORTiJs4h/bWsj6u6WDvj0Z9H7vy2Vsq
WzaJ1bMkCice4mkK9jH24WWN74PmI7kN3zj/ITX4b9gIMZS3nmbedcPy8puvwQdHYN4Pee0s8kAB
trImRmRIrME3aXmt1DlRklkS6sl2TB2jXRo7Zsqm1rGk/KCW+9fx0hN44prDn67yavKpAN2elyqR
bCPvbTRSlr6pCHKTNL3vaWDgcjgbSCp9hsniaaS34RqzDfzjcEvyBpVK7OuS60tIFEPPrDWFkLX4
AHdzn9cr+d1XWOiqtHmCNqFIcdXpe7PDQCNvQfm8awQ09a1U/2LQzi6C20KwRV7m8abmirJOC9In
IOP45j6PoMothzCVgmujVjg6QNSQb+l/cyY9qFJJSpOj7NbnRlsmVgz6qAItSp9uYgwUAQkIiBbL
gBcGDQSL0MUX8d50llcSL7NCJf/lqVMuElGATJZz7U2mUOK90s1Ux0ofh6SzLhgumk6JrtxdhXGk
9sxDNcqa7dV/6zSFzU6jDLS6DqHb3vBH8/hq1GCh7JO1SduTQNfDV2DKkXbH0VUdi8w68gmMVN/n
BGtSMpAWXuGJsuluxKt0wPoZNI92jgXur7YrHekGyBla5roMBauySl5f9SWxnHl9mgX9kIKpKN3/
bCQJszEyH2rDaNLcGg1Jyqz9QpLJlVzDWenCqf4nx63Ua5INDnGudca02GOYF46OPgQcSLaEyxHO
6IvaGJ0WxSTzA1A5Ootxgo25jDR00oILKXJri7R4iaNoZ/LBzu6Xfhp0uo2W5FF3bxakG2hn23sM
NW1FGs9y4PVdEim9GYubuyO3/5+YD8MJmxwaZE7wOElsNSlrYsR/ltQgh7+qNxXfKM5QwuBCE4Cs
zAIppKEVvQIsMWoxDCpqPqeCLWucLFRUzDJDzs5F+hLNFXN+RMfNcTNMw3nSb4up6ip+ZrgXoQtz
ggpe6bKHVe23lVAFFAmpbRgLo3/kA1P26oend9KfMrrfFzniGcgOyBd6l5wnCgZi374Z8ipzE2lo
X6beX7T1CMKpAtq3FqfF5CsJb3bdEJodeaHfqQMR+KIaKt9rhzKi0HMXZTHCwlx978jOpC5rcUJL
kCEElQjxl7LKk56OuwNuy3+V/Cc45PwQ0kQtZ79UNiW9AnjS9qe+Xf+f8mCXMaq5leYfhOt3TQQU
vY35fknYOyYQl41Th5DiEJz7lGxm8chFoyM4AosJMfaDsDSLHqKsQgUxPoLA4Rw+PLjxv3mTezwV
YD6TA38Ry8xIFtN2p+FljgcOCYDdMo9gkVvsO81yi/y7VYKbeNxI/FMpNsBjs/1OLLvIuM/J8qAO
f52obg9cXrYM6idjky2v4dhk/6GxB1ARmG3mk32Te02anRC+2Xd6GPNuX4PZ3YWOSZ8QbLM58S9w
NHp5qOqjo05zeEgsmstGDroh9NJhdJ2QN1Z0g1H5bhN2tVMeLUmcwLH75hHGwPDk1LvcTXhTI9o9
QvPtlyw1WLJ08bg5XKg1cp+D0wVUwfO2byIbW1TgGxw7rGvch4+Wfd4Nb5JbUTrISmNrOXrSNTLN
vYCElSf14CNkzOvmW4U+CpimNVn7zIBz8m82/v3zXfD18e8+7b4Zr1Nhy3Bi5jLsDt5xVVzDjuFQ
JtoYu1rdeDL7UoPAS6VeRlzmcAudiY08MLoUUaIpcKWtAd/IMWBjTIEtm0cXXA6N/hIsXXB0TYDc
poJ3DfW2pK5NjYpjRT8uvx+uppZAzyndZlqAGsBe1/axsgpOlINgnOi9tN0s3y/eaCIkXTlTDhj9
HurgXLdWonD3RnccQYMPs8M9Rwe+YR9bso8VRqAjRGcL82oXVFHPTonEn1fCsEuQmu5sWn2GjGU0
uf9460+hNz8hEAme67g+du7Um6Mfs82TAdjm3oND9LsDy8tk0eyym0N1RbnXa3ZONBCb/nv+tBn6
8GLwAe1tgD5Dl8vski1zSDGR4DZWMZVck9mjo+z7TDPTxYJhlsKvt5L51DAkROQxCBrAiyScM9Ch
5sEPd4sHVDq+zNMw1GeA7IFGnhDBsjhjfDz8If7yWwJYAFxCsKcSwkOjwVGLvEmH86R1pCMdScgy
czAxfH4c+VU0WGnWwZgVkghOxVmKB8EjPhIOrd/m0m9dghlz8/Z2eIjglSakMEpOQgA4bIAzBolD
ttuq1H2Cq464hBT7p00JhaN7xA8SaPRt6nZ2plLLvIAfnnBvMAg+rTWJX/pcfbjX5S2vua6WdtX/
tWYc1DZi/5Oqg2uFwDSBB71UwbvvPDLE07zXn1/94IvGrRc+mBr36c371zduL7sJj2TJlkXE+vny
S9NjLwe5a/YSY0p5ppHTQpZv03VqO2lGtSjX2s/Q7bJQ4dMrKQskCu0aPXQNqq2rP8cPXry9BJXr
h05pkAiQV4hM2jqSCfEF2XfzV67FMtFgHBHCQa1Y9nzzCWA0ruCsjHDXNpGw/j09uLjhvCLYOvjU
LaA3NVEZ7b7E6hD0ITvbbh0MwXdZUTd2CRFqqphgx5l/BCxwg3V8oIqZ8fLEshF6+eu4tXaQ/baE
p76RPvyplEcSqRFHEo1JgfNtETbYsbYuAvUV1YU/+57QPhyNge0/yXt4QzQQRO4RhyV+qvUM+8Pq
kCz6sSdEKVcY052QfrH4y/DDdbdD1bacuv5tE1r/e74u6uPRPfFQdn/CA0uFaeWDdpNsmZKx6Ryx
1M4fiyA0piPiZekODu8FON7L3u7kI2nt3rQ01tFF6UX1spVw6UcTfk2by8HmRuAVHUOMm5xnj2d3
Znb9TNvmY/cKk23e37GZgCxYMbkph68I7V/43Eo63S8qPYpIH7bd/bab75kSP9piQaPWneksG0Qo
eYCoiZtq+a8HLRcTsEPv6p0tohCGiOJStSwbkfi3ysmJ+g/guxZZdwtvGfJvFjHXH6WU8ynrPjK2
P2V+PpQ0kPllATb4bdXqgk77ox1vSmGKtvBXgnD0ub6ujdJNrUmu2AuX/82gg6x2eLfI6lAeAQ5S
uoqhwUuD2H6/9loBeQHPxsU2e9T6IJG5/idIaQpJhnNjPTiG10xTO8Pn87x0jvuioXnMOdRD8UPb
TRkpyHl2Ri+TBU/bOFL8h4EFPw4Fda1tLEjWqHMkeDeuBvWqkRU/U9u0+1t34lypo34+CuM6tjw3
w7gMYvWjsvCPZF7+eeMPMwDdj8cEjlPAnLCOV5zoW1YrlpCxo+FXqX0sX1O1MRvU7unQvhVb/9Pv
GBKE8lcFwoZt+R9Gok7P5bYUMF1wvAHxw1aovOO7D7T6JIfq6UmR+r+GH7mmjVFIjSVPIfUMCeR9
SZpLJjYr2puyERX/uEnwh6ts8AC1/SBM/qekdsYAmJ3+yT1i7oBLmCJPN99VieHBwkCn5EO3pCmT
tkb2gZhuMwY13N8VLHrwOYAxzkv37/bh+A0Z47j2URJ/GQU7JBAMCJaWWECsIfouByjeVqa5uKbz
C4yqe7DVdCN3HcdIQLGxhnpcVnTEgDeluzGegMQ3kOUqIwmQQNDVDdxwseUWXE1eu7quKizOitsX
4sJ/TtJe40U76DFfP5EhO1HxN9W2j2cpKHZk5QS9ramZupoCl+6Di2+QrljLELwveCplf6y2rERX
MCDFtFcJDeJgR6bvh3JEhnJFWAmMJ3MhhTUa1kOGV0lzkCf/ucKyiDQCI06Ek1nMCPD9wecXHEhF
1mktTsEMuFeXoFoCAQcZKAanNY2CwifgYhYqKYNrzc0k1c+kpjiwTmo/dxtbZnpUkqnXuGSY9jJW
Ayjsg6eeU5gMHy8S/N8CXJVQ/mg8F4guKyceKf97CPVHZqwgzji1LOOOhhTisfvYjfh41l4qIXE1
3ZLCDYSTxWGTYFNpWzzRnwBkEvm6Q2gw0spXe+L5JTMgQpHYxRsAyZMAOmERnMxo4Fu37Fbe1tSX
MZYUIEPUCRJ7YzocKWdsDLoNdSJ4971K1S6duunsgni2kxwC+68c1cUp5tuiBIs1tsPgfSvfHP2W
3+NX1r9AFrVF9TblT7426xsTGthDCE6ljlzDaiJLOIlV+0tCmOcODW/K2qh9k04N54Z6h3DIJGyy
q9BdvTNbBObE2BlQ3j3MDeFahqnlDs9CxAgR2vK9sTKCeiwl9mjpVK8TgGDk5Kl6ZCS3Za5H4a0n
EMcicOYmixl5ifuF57iYTwL/RiKynBvsnWKUhVKeH8UvY301f7hp/qPjeviKnzlxxM9IycqIWAza
pcJABWQFC5RAl0q1GV/LmeZk0w9Cm+YpToZ00ujvmj1eXxJfv5RSrh4pc8Kfwb+ZVozifrXuzdYN
8vLqugEuS1nTavyEzefQyXqYuGeN4Npq7uwUg8nP7GyauKpMTiMm4tL0ADyd+Bc+7hvhJ6tIzB6A
0qmMmSy7R/USg4rdwt4eY3Grmej7TA15NRzZllUCR0OwbdZBC1i4Ti7Th6jWMKCPq0sMA9MI2MwN
vBJJXPtcIko2P1ETeFvyM/zY4L6pyUundJat+dcaj9pnjnHLQoJDX1h3moxQIM48tFKHJewxc/Tm
usygPOhEJjJ19eueugRLlfbqR0YBnPzhZFtMIOLbKtUdrztPliRkXDpxudWiDauy86QLlA2ApBDg
w5NDYGIym/6jL8z7mrEYRVL85ICA65I/gj7lWnVG66n/a2C+SKNYlwueRfrjsLQ2VfFj/KSe4qOE
WLgZp8yJXnAPoWUY3G9B51gvn1H7wP5+SDvl+8QFrfygjG4IZiDFx+f74H3N4eg7iC3mNh+ijnAz
NpvJrJqlBmx2INUqhjnoBp+n37nN4Io/Ls0lOnppQ1yWjBUUI+nhXU5/flo93aZQv+t9HtXzlLES
cm9oZr8Z+Erq/9Vy7kaEsarfADvQsaLapZOb+XQjoma7QbK2bfnAcCTInZrd1wA7owkK6QVO/5Mr
hlN4ulq1iky058A9XiEPolMD8hsrsF3WCWmOyN++IbCuvC9ansQrqzkMu9k21k5sWAjyW9BvBYEG
FuWxAGghHvwviheuq0qw+ETzKHGC6k5oGClKxnq/AfcqT/ioHzZeyeRCr8RnUzch/eIgfDiEeDNW
CPpu3heVdsbsP0l9wg1b4wU6x+9sSZ5caADOVBXhvL6Np5V5R9ptfwKIiaw+jQYpCW42nGZq49Oj
anaPxz+ip/lW37BExyPDh16dkDsDdI4SaZsW72k6V35fFl3cAW+waYcgMEjCFGywzDXuzd70VNIr
yi4lrNtm8W1HBXL/9+Cqi1vxTHUKBId6awyLGvvK3cQFRY7pSN+etXgzK7/12tittDI6WYsNegCE
hHvyN520DxxNr5vaGTAXOJS6QiYUmsCFOgUFBjg7DElwaP1OdbDatfpH5wxyhntHciHSTC1u4WMO
bbvA5tfgcycpfeGPpemUWa2qRKtn+L6g9MnDReNUTfJgv2Hc/8GlDW5qVIi+s4A4xiK7/Q+OKaiR
Jk+1Ts1S1+cpMjrbV5HMqHw16DaZf/7tvMunur6HtJtLpfLGD2nM3wKkABSXqFy9JbAkRZRBedCF
mCE+au8HvnDylxE9CbXQyAC7REn8V6JhXpsHJV0XGJg0wCKn8+V4pl2Z2ME7iRLjiCq81ZVioaYP
69B/UGHdzD9r8IjZVbbxZqU4HlHSXhk3+lk4h9MCeP1k/l/OfQJ3lH78kGGmQgWtWd12suO6Su3D
Epz2tEIrXEXC9nfGrtevmki4ZJHDMtST6bAvPKrACmzi3InHOrGxioXbHNW57JUx642JwSI2+KyX
E/wb682/4x7iLrj8TCJqJiHzyYu1LXOT7/PbNMJ/z4s79Qzy/DRjI61ApRBZRQNa6qMKvjHISa/p
UJNbxxZgFWL/uZzzU5utVqGJSzumGe3uuaXcGgbmL7WBQj+IfsH0HoNqS+QsDHeF+vlNxVw0LO7u
SeD8t8wglGayUNJZxCrO2a4zu3YK6AN6UXhw6pwYmlMTYxyRvm5VAjrONN3xEmt9bfeoUoxEDOUP
I9X8v9j95NMXYaJYYWY4wS0UjfyGsPqBCiBU28wD7Xz+0jlp/FVmEEyABqmzcxZHtsRvto/Z7ZOR
83WhaLK4vGexpoTB3UYbzpPsDs64HphL5IX/TgeVLqBP1txnNuvtsnT9/ggyTziRAKSS2NFlIt1G
m4S53KgxRVPAgbrsG4fngWO2TeiA8ejn9njIecHk8vTohDqU7PwB6g8gQ9qoMe2eZYp9c/nBNIPe
zgnICeLI0vTzQcUYAeEGmc/ccgLQlvJ8CZqBERk3Qh3P1mXg9qsYUaYqmBAfkg0fBv9tjQeajdhg
pBfbmtENRrk7CUK8FeCZaJiw+Mt0gVasXdPctkAVMVISEVTImqZYLptXADurm9FwTS7QEXNCBmyP
pnL2UURhusWMCkszv9stoYtT7NUAt+xb6fFsDwopFbaB5K6zQ+kDXy9IqIzfQSwXqeBOns3SbAik
tQdtKTN/J6gGTkwt6Ul3fVqH1gBSmqyH6KvIW7FwE6S6gAx+hqZABkv5IFIJBn80DsGolA2Y4xHO
m+szNTDam2fL/tgBKM11H8wSbxWpmujrXqRv4Rfv1JPWRXNwBqFMK5acSzV00M8LJvkRPZcop85A
MHMel5w+3jcsOhF+SqeVJytwMyi47lRFnOnrMhOoiftE1kFP+8qJvyRGB/LmCAWtwZBr/4PTxywD
05A5VI2BjjMiZkKGDjluxXB8UCJEWlHnMZcb9/EVGb9eg69Yy0x75GPdNYtbssjbknvPJzFBHhBa
LdbivrlBGzj2M9gQ+kQ2tldq7/iN4ItLokPPQxZOkIczBDsyOKeu+nAwKNUMBVWynoJkSWSm5MFG
Aj3c22HOFllM97ufoIc6b6rE6+Jh0G+kWEamhUJn48jwSlfkv5lI83jGXbCVAaqc2hCmNW2IruVC
Q5CAWmhBhZv0+HdjqNwZqQhOpgh/V3v6nHDAzvM7tppO8F/smc8DUGJbBaMUTOjS4eBc7DzcY1Zt
IPc1ZNmt5KIjoaz8QT6ZWev4+vZook+QvndXOe+VEJ+XTGOfr1XDU9+0upDyPzsCjOrnZ1fyo8+L
rG0babxTguf5TN1QwLzpZoDEs2QV5etaO7ZAYh2IO+Sn0A7VXEiIKHgSgqbTyThoFe56mNWlEQoG
u0R4SyeeJMqtC99w90KVmLM0YtKrD/2MUiI93WyELYI8QgAFm1Zf9yuOJUT5i9na3IuGzk2pksgR
79a05wupDJMuBejINtf8sRZsSqDl9CqeUosbTRlgexbblfo53l0cge2J4DzBIkbC9OuX7aVbP76x
WjgGAALXomoWuhGfGI3LjFeA3u/sMapMpoI7C9mA8E//TRKoanFllleGl/7Uqw8So/+5GM9W3D0o
96YMfeSVUxprtgDz2ClS86nDoNg+mss2wJR36TYpWaon6wbQmM1Z0tCKklUE0pRrjDfYSZ4S+KTM
Uf2GIN7D7ducrRTanO44OqHAMYdaiWmDIagCav7jhuCojXX2tITyDjMPcdV2e4eT2Wn6q20EAjnQ
UNkKJegJ/AInQn07M5/WY4FlHy6ULnK37k6j0LNBtcVwWYR+Dt0kmyHDEHlxpAq7Swr77+zHUv3q
916FKZZC6+2+NdxnM8rXu5Y/yUp7fURnWKI2kym38ZzUn+o5STIuHeudYrbGTiI/XfCXQsNYbJf8
3d6tDpELzirVfxBLgN5PPZw9QfPKmgov8rx8qmxWs6EQFDZjHPo3OUs5WweiyGZ6E4aFJmKmc2V+
805wD9CEISrs4BWfu3QTaqyhFRRhzxanZzMBCIuYWLMNKziGKlRHoDw7riiSa+Xs/KwhSdPDU45x
D+Pz/+nW2NP+3lVdLp9gEfpG8/ZYnUck+fRHcMYfrkyVOHRN345WE56/rV841T7ih+YNRvgdZfPa
vESchYjcNmJQoc5L8xooGSXu+p0Vu/KsH8Mfd0Fd3c+KzoaUAtMcfEUg159g6xeR+Mc21rl8xUKh
fTdC639JZBbq5VV2pzcZQGsHbvOGQI3lEw9M1NLlzE3Bah3WqRx0VAmmRVepa2MbBw0mYznGbiYj
GFjakDvac9XNhKrA1hvI2cg0PcEn6Z7ZSrCW+tVmjVxYoHZVf/Qd/dY9WPEC9LrcNvVUntSTM9lS
c10AIlMf/DS8nKem6HZuxSN2tu+XKrN3d4q+vkhcbvBX5GN+4xl2ClvBONlXYv9ZKYQnVTmZV66k
sgsSv4dhH7Kn6NKjOsQNhfjFwnKt2q3gk1CqXSjl+xeKrSu3GvRiDsIYj8H40MczkHy12WYjaRF5
hIxdMI8m1cmX0IoPmWWzGbCep4FWR+0d7vTwyTTtaVh/u9LNa/Itdg3YJ1XTHA/PA1aCFHD0oHPQ
k8DJ+XbFHu8uPkerqWLN4+uIy+XaK8leh5E0+WFLfAsgfFqYRfIktNBfuMkn1DgFlyJWehzHJ2mE
CIQdQEaCbQ+KgWRW7m8XVMMwRh/xC9SwtAG1CmXQymsm6+Dn5quETnTawK+9bNqs5+0qxd0GctDS
x3VCQNT3/Qdezem/yrxyklaDbnmz6XR3N6JlVSKwkuZ9/ObrTncvTWOGE3dSS1/B4E572qNFdFzx
K6TwHcuxVwv+MLW29FGoaUtCVqBLuMPFPy4Et2aOmA4isYM8SQCnI5oPsMT/tM8w64RKzrGTObuI
+pSqD7cA8UmifYEYTwnnlv3LxeQFXI0n/iO0yMlL0oltVqATfwhtJup8ACsi+zBvwY6po89CA2hk
W7KwthnX7vG04GGf28WGg2fa0yg4cZswttGPVuSnsxhSZWvx1dwZwVaQPuSnict6iJ3ngGV/Tdaz
ZbNjh/EzeMJgi1+RtMQMp9TaoH8uXlLp3KWD22H3sJz1JXaWptb7odGzgrAuScLV4qpaejzksc4A
PVWE79lS7Nt6Tfq1XjD0ovbLYJATL51IbLm9tBlFGKMp5JxcoKBkaI/LvfJIW3uUsainxhQhCM0w
1A+YCWB6aSMu5oywznKWoFYwjseXtwxfd/K2kaxuOL7IzoHL5PWkyAI7ZSTnHRUm7Ha9vTUwkbR4
EhcOzeA9qvZaT4XyJZi+ZD6oVzE+p1nzBT24hkDwN2tekvNl5F4oa8ItX+5YFeKRLe4m1hbalfvT
NvGUB39TagX+jt+dXRejkgUkQCpfaM06z4lYZozwtbDFclDA6j24QdRrD2TWCT5OHf2naePBUJN3
BHWnkmfIrL51LPQAy8pxCTFJupcMmF6SXfKFLu05BG3udYz7GzueqrreHrETrLlTTqnmxKYPGhx/
/Y9IKjbO9kBcopFTXlXqrPLr8Hwgx+tqc9nmd7mHAbXGby93Z4ELEx96mUNEdHplF5evB9m5qMKf
wkH0N2/ZFb6iqAZ4flAoszcncJ6HRAuCZwimXQqSdgK3GGtsYqezxyHEjdusc7APkX77vpIIHOYX
atWMt1wPDFZZgELqIQBPqqqs74f1KePt70EGeFcBDSZSI8q3hoG9csi99Vq3YPnc1ld01tvAoTqX
L8tZkbYrYYV97iSi/m7mtdzO6fljeQcIvQIPu/o6ajfAtbmJ6IiCy7YpE7zPkuxXEFeDBjIMym0I
H0ud/lfe9vP3PaNSEiZC
`protect end_protected
