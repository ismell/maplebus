`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CiYAnmWljK7dHHQsOvXS6S8XIz6XwCHFYinpyaUmoCpzAsKAFqBN/qZVqKCRHZX8Hqm8tc7DywZ1
ox5JUUKzHA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z9ePc5Q/axeopWzIcCyKCPUXrX4vhCC+NFGRmOLux04EqGnA/XM9qN32D1Gm5a8/VvuqBln//Jg+
CoOaX4hz48TTNVP7sPf9Iswz6zMyxIzS95DDjwKmIJUDF6tGqLdC2N0GFsVZhrFYK6wBoay/xLLi
8QdyG+52y+v4Z4n70Yc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qb4A/hbXFPzj9QjPSpEzbFfhyBouJqVf+e0j7E5Sa+lK787Uij4YrZp4/dcJEV5iyQ+J+gXciwDZ
OzcqWFn4ccNlSfXS/osTSATrtK3osZO7SW32W2w9TF6i7uRjDg2/iupgMWVF0LLfZCft0hJR04hP
mDWr2+USyLO89UbpuKDV7e2IfzZnbVBexE/L7sRTbUuQrsx3NtjkLU4cUf+PqOA/ZFSUI2el0l/9
ksLezi819FVnoA1tDLGmd8328QU22PgGWT6qZMRnDIlAVOg938oQFF/qpQeRnPKjtXubOLmvUe46
JFByAroZyXFjyMjNFy5iRY4yfj/4ukdytmhCzA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4j2biwb0C/4gt8wSc6PIUJd06XYG/m+QG0l5JFievxCaATunlHItAqHfWYu3fuPetom57QD1Z4xC
U+EjjX9xjyoQBBIoAgqSPMFz3WiyrAmtAE9zcSlDECCsnHTxG7o5FINwmVWODNt+d4FUHCvJDPLw
bRYDKhKiuUGO0y7PgKg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cPpNCCUFAqecRr6OUzt7mK0aYGDZrottoqMYdYssAH8CFVyxHvfm/n+1ujHo702nrCjtlyT3wDIZ
vx/sn6cul7isqd+Fmzz3HTUThG75F8bX1xm+tCbHEJdskGJcH95P7lKi+QBQ5DvOSZHxrXNck43J
Vl2n3dtW4bioSF/xhilDVsepTCbiyYDXGcCNr1DL6hmqUzAb+PbNy9S4h5h/oN49zcqdHKT6XEqX
yxXV9Pg02oAdWu1SCdEpN1xz1hIm8d6kzq91Cc+dGc5w4zbXpJrIElwywbTf0CF0eC36oFIRovIy
Fx0x8vUSSx57GDBJP3+61YziNrql9THWn5zsQA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21952)
`protect data_block
rvbAR8vzyr/XJAr4kEBuC2Yc25IT07JZE0jRQDfypIEQxwaIabNA+mTuonUE45UPX/hXPksDTFzd
Iz0TxvHozbfDFD+iinZWnhkZOsrE9QOYILL9yK3u9k2vDsDyX01S+j0vR17Bke+ggMVAdkzK4m+r
8jUX0TH0TH59YIAwI1FftN8vA85qIF/qNL44I/rFnlt8rm64q5sTmHs8S/mFsqQFevYLY0Tg0htj
DBi73BvJNMYpPKrfemXKMnS1Z5nkH/s2+fjlceKUXHstOdxWf0438NaojbWi5nX+deJHoZoF8APF
8get1bHaJfP/VRbgG02C35TMjUx1qslQviQeNd/vYzM98D37yRGbdgZVBISpqLsrnMEYxmCzdUXO
3S0xKvLPSJ8MmDbN2j1pUitzR1x7yTng/qUyF82nx6P52aYwK70Kij9/0f8533EXGqoxZuuDKXZb
EAjSC7sV/6wO1LDPHeLDGa/1MY/lEnCfRJdosuxKPoWEXNxVBTEYGH5+ySsH7HSQ3Inv5FWymRv4
u1izjfjbMIZUz3y9SXvp7OM2Moh2QJL53TXEUkSMWPsWYgBJ3LmFq8FfwOJ4ru0gaJ0dyw8RBGs2
lFhT00vsI2Qy/gRy5WqhPW8yQZDQdS79w76VBAfH6o8D6UfNIP8G5jqCcpFLtY8+hUG1+gM0jIwg
dGNlJJVF/PBVIZN2VC0RwTD1+JvD6pPsLrsdWgTopFVzVtxFNUvKMyJaYlYNPNy1spppiAqF0Km1
NuhaCMGy/Wlc+W3lMLN6FgPCFo1zRmVs8gZGCqIyghv9ZjJjW3Vwtv7qYPXq2Pr7HckCCzaMA1lr
RQLyKlfEcnN0U44hAZb+eqY8lsolgvaBFMg2np/mxaQIV9lC7b9iqXOMZQn/ygGWpx5bNePrIw3q
SePYJMfc66qpS7tZdW4mO6F8cgs+FvxlMfLDkWEQK7yGLXVxQKQpS2PotAGa3/IsNIEmo3TcN8RQ
Em4s2Yb3lxR+tzWIlw4ByoIevVE/E4TrxTushxySMGx5tyiOaYX4G1OsBUdeWKVuvaigY+vwENVo
g4x3p3OUw/h/GT/PSqB1/jgkWVMQJ6iLqljnxLO6ZLtFmtNCx7p0lREnaLSyV54vd9AjbEWW+WW9
aD6sShLQUrQTlDRFX8xeRTVhhps/uqeDQsstSD0r4Fs9BX2uW+Neapc2O1Rj/LL4hA9tsX3KjtcJ
M3N6tiLl4sVu7KOK2dm7MWWQ9eB0ALVH5GFk+u2IcjFBiRVLWYkM05tKbCYmDpsczHHqurklPEsh
mo6jKCTuKY0MCoCdTKw3SbZLOu16eIKL5At0b7aaaeYhElf9XukPEdhifMH6ragSA71N0Lms+9Xh
QiWLo3qxX0nX0nuQHX9hbdT1hOKC1MBUBoWkFhDvF8eXYJ+rCFXsUoheIzRU6da2+5GZh5oQ6yxy
4M4Xx5t5YASNNBML+x/2OLUIL52Y9THlBQ5aECfR++KdWv3aG4EJpMdXtol/q6Ko5+4QGGMOD9qd
xEKoADaF4MV/VxWV+MB+kuLtf24e2lz/PkOb5gcTHdyaJAm3K/ujDJ6EwErI2KjGWudAe/b1/9wt
yJ9f3MGWJ7yvBAJrqvsq0npUOKUZiwGgu8WbRuXWEwz2DvAaPT/0t/TNcglLQ8nknDutYb7ctw8O
ASa76o5UCkeubeIRE7XM7EMUcoKDOnM3pFned+QHdfsiPP2d1anQuMOTN/bUg7AICjr9iA3DuqW+
qa/uM2nfxE3vc9cvH70oOL2yS5BrUtJa8b7x72NXA5gdmefXLu0ZSsfw0RVyk2zy0w07E9LCEzkD
5iQa0h/dEvzCBF/uaCAkd8tVAWPKsdNrhSZSEM6Ss6cDdtMtMYgCb7ns+j41jRclLphlPS1n5AC2
sBagZ0MSZ+VKjY29H/qs+Af9DriR0kvfR/NKrbbGTWf4ES3E2yV+79rAwumuFo9nnfXTt2wMDyEK
WmkFTnC4ucZT+hWfny2/jWmoEtF1VAYgx1MopDBIAyJ3iIzwaQTKocSgtGdSHFAd/AUHI1CuAq4n
eHSgUNm8kzMHXjzTBkRkupV7PSTB9hns4gTXV0t4rHHXMUibtEmXmgyZ5XbnQfba/k/QgFww9U6c
4jKJoFcJbHKeDTb3wf31tpever02+ey45hXTFC3MwWYGhuqPE0+kngpu/yOqgYB+wKn2Nvfb/XYI
g8FMIZku6f3SWh7mu5WWe7+8+l2sk6ugIG4srVFmPvaEykAWz/OaXygNUQkadMg8OgRmGy+LJqiG
nUHVqmeOnaAdnOwIKOTTuwZ2yzAZvZyy2iZORCzuWNkGOgj/tVqsubvvayrEmg6ss5UgFpT8LHlE
OBIU7mFdEV0j3QJwza/JRmOMV/5XPh9uQAy2Ot6BnQT8PpawuE33o31iTyINTrc6drkJJVfr0Wpk
EIW/dTbXpCxXJJOH7T56j5vlM2rXLfk8aw8ACgAkqLP+wMCr/rUvRKorwYQT1a8IoA/lW69xZXz9
Togy4CD7uOOYtTHsMLKhG+kQ41S1bzlNqATA6kWkA2KejvDaB6ODp96e7GEer3WofjhrzZ0PUNAD
+SFXMECA88lCmvbUjbjPlq1O6Fk6VZdevj85rAJ1KYWJs4Egh/7jujIwtfNmA72kv0YcR7IXWP4y
hlhH32jbRjLIE8SG3HzZ7Y4OzlvsdsnCVcd4DVsKxzuk+gFXlUt8k9DMNCWtsGJMxeKjhhvoMty7
cd5tRJ1zY6BGm6LpxzfXcSHlB4w4g225LUjbMSV5WtypfCKi0RNOi95CknIxtMig9sh2W79lNtRe
KmX9w3UH5dplKYhkoaItTlNEAGMlhhxEC2GPWLh22zcoPOE/ejRExxVULx18zYPJPxrA2aIb9bf1
7tiMfjdDM2AjHWKyT7JAwj33L19r1e1h/pTejdNAMzWkvlykvOZpShvIVsC1nFlhrptPUui4zMwC
6ewo03L66W3rKiLmbK6Km38LGG2lXdR9tXssUADLnHgH5DPYqFGO8AFixYBEEyUvZCswvH7CIFHr
EQddYpVBrRXBSerqD6yS4lDugTStt6Fw0VGhYhijjDSeCGlTkxU+tEBxxBJQhdT5uzdQtzYAsXMv
pc7+27htM5XlwUDqcxAQlcW49on64QqobOQW5AvsrzjVoBKMcf9bf+kFfNSdW10pnwsOpZK5EykL
/kztIz5/Kv8/z1ISUsFcoIOQlU3D6vMzwUYdVdG+jHgv3oZnuDpvNiUa9+uq3CKRBLOT4O7YRtAf
1/csSgr/mXQJGI/WuVRn9+I86H4BFvGPZZm4YqEEvgvSw7TBx6TDEy9H30V4IUbg5lx5C4edoXoN
zVtnL0kDiOVK88k+GwVQHqe3qmFP87Gw4QN157GZmZHf6ApeR+iIlDCS8iEmL748NOqVswi9oP8q
tFJD58VR1gK0aYLt2GZcrF1jysfpHP87Vl1j93L2i88haTLgxnUHghvYsSO1gFfaNCwmbdCqAcxZ
KaMK+PxrSjfg2WnLqKCZ5LtEu63FreUBchSO0/6HNgthJy0SeGpUlM2JOM4X6YIVj5kW7A7cNIGd
uIqb49nRXahqpHU2GtZiKr+ObvGwpJCr1FiwtJ3z6GOV2iMpQlRT+0hLHOQ0y3ucaKnYpxDTJQye
xwFWdXrDkm4/nhqdPNM1BOcum62C3mQe5WvjeNPYEl4k+nkyTPZjxXUB0afeJgCUa8Xe1O5haBiy
AcmFo1C/JKDc0zBrsOSKkv5+VZdIwfVNK0+NrD5Ln1mwva4e2+BboXkOUKb++QkUvvU0nWDmARXN
CetByYwqQT5eTnpt9YyUujs/4pN6X7ESe+irurqqXGvY4jFQaxEQvh2zxCk6zWDzOfUDRUvcZB2x
qq0iVFyMZM43aDTq3ygsLEToFyTyO7h6Mr/0s9HtdKYB6V2vSlKamK63gGvURQAjrNETO8BTp9x0
X3VLtPpL/AkPBrB7WKD7Vw9UmmZ+cTkJ5g3Tis/zD9Z5gWfF8hxWvGoHkN2bMspFlxIXLTK8C2ff
2oIFODkHoAogDRGBBOXz2rpBFefq7vCkR8uZJSCz7UYCIxSJmOMkXXgmHZMTMlxJBs8wig3rF2/f
t4oyQcALqbdUuZHPI41kjjnC6NpK6Ja++lt57ZE2grCzHG4LN84/OPVM3JM8LVeY6e7mbmwvHoA7
FGfruGyP6PmXb+KRdjE9YpIXkbmNAdIPK5E+MpTHEJUIitUsNlwabj9wEDP18xcPkj3FGr2bpj+f
FIsUGw5vsBUGihzjkXwQwh3MukWf39z6OKJEaDVnhIe88+rhyaIk479Gg1fHG3SPUsjK/KzczVCN
WtAsDbM/ARofOwWhPZxt0kRgvViGipq3l+bMGcp+J4Q4NXAcbqM6rvnzkZuXDv53u9Qz0DbVn+rk
HEjZF3BdFDa/hVcBCp0wEIfI6ZX+IrQTcW6HnJVg92CfRqnB2V0Xo1jYtlAD12KFN3yA5EExjfyC
MW+/oo0pesqSAxre1kNRanjKOKwELg3n59sooDJOHKwLypuATtm+cTOkCJ+0bEBoDtAnSvDp49Q6
qeQWeBq9LnHW2xhw64s7iSSTO8ZVp7clkD3e2P8WTnZ2veInbADbSg6BIQpIfr39zDDza2CPaApr
QZC5T3d8qKrtYrhoOSkYCR6Hw4p2bQWYagEZtCfbBuuCp9RDDHlLtp8zQ62/e0qzDQ1jbPQ+4lX7
BTRe5IODajcF6KcHNJk0O13Xf0XENwHFRSfpFc+Bm0KjO1bvO2He2aEaJnIKiWSBwZsFcNAZ3k/g
ffLFKlIU/S4vDSXYw2MCFurL8mk28wjQbJ5PH5V66Xoo8ItxToOHfExAnjmPBvSoLittgPSWIYft
rOr3rs1IcBya1D57QLOcdNQ4vywT9BTup3Ezo20nDZIyMWyuIFJejGIeTLcqmjhVyOSUAC75f6ER
4m4yZ0rWt7HFSrUBYxzVtFhSi5qFH/nyIV3RIQJX/se468Z/0WMWsnIvP7R79iICt4/tD8NrsnGi
2ciiLTb8n4XjgKP5wV3Ice5bsS06wJeOYBKl5ImnNelVHtb6SiLHszexro8IRKtm5tScaN0DVO2D
2Z8XTGXBDr+QJUL06ypEsfLEc07I09jyXu8AON+XiOsshG3QQ0edySGv9L/K+w6YuxiC37j8gr2W
IOZA9RxCarAW1GIDmARLB9N7PZityqTgLRU/tnmeHwtWixJyup+9XKZfjHdIE4zZAurjJ4ke2L0/
I8oQUqdnH83dHOEH5kFGHuk5NcSCYABqmCABx3wXl5Zu0kWAQd6I8TA0wavKYzO4n8X4RANimC/x
RYcauI/AaTFWhv2Gi7clrjdx4xoHF6LLrB8UIZhqSLf8XSTonhpFR+JASvx/BLnA1f0SrplYyQb8
tc61i68fjGeYyVLwIgmbrknH279ahlevyYcXjIu6/4gDQe3pgxs9VlkEmoBfdDSyDOwWDFgzZALC
1a8gA4YoLrza1zhz4p+v4JNBs2DQ+YyLOK2kmuSWMHZUmVzdmpM0wyBnR/N+MD7HNhFgNY7AtAJD
Sb1Z+qUP21hfxpJ+ikaY1BYNlNHM9TqaAohSICyRa5nmpivaXMnrDagmswpDX9BMll277/BEDzGS
zF0xgndX8kBdECmrlAdL4P7FQp/vXZ/iV+ssy0AjQ4UDFbLXi2Fo0DG7fnaqyhsVONYiNfaNCBRY
GPrH7U7vGGr34b1METsPKvJSef7MCKIQmgcLvBYyUz157yJ9fmY9Y910ywyeo5f9Sc+kkR0uACq8
aI26yvf+dVwaB36UhlBTeUghwtdHqW4fOxxQaZBGiYdSGjbn9nlb47ROGWd/FW/+bHlqKt45QPRP
GQKHPY72P1rc8N0sjfI+IE3c7gatPpMRggy3kG84tQV603V5Hog7E1Ovd4of/vGMLfpm8rf8WvG4
FX2uAsT/7uCTph/vJeQOJ3+f6OKxNP5v9i0usSMi2talg3F5Cddw1KwC0ohjN8VKhyEF1dZErssG
b+SeYQ9QbbaQjygVvnslOvyQB5lS0giJStxncrs4SWh6LzE0ak+I8CPIwIj3ew2DujvpwGZNyONX
cyv3FDB7wcI3Anyxo+zTnazDLc27yKrAyYhNwt9SwvHR7vaVO9M40cGmf4hw5PPm9H+aCnEVA+/+
0Gi7aOp++nk+AXLj0CO8FMTupsca61CM3FY93e0Li7zv4xqVek1UeuJZUH/f3F60hi5uwUwnHOfN
JwrmTDQ2yDlOhDuXHSyar8uAH21exPNgAZYmNz4/K7V9fojXJ4lugIbQifMvjbEAWwZqxyNTeEc/
p4O7EoZxmtKIrK6Bc8NYRdrS2LXCweHEG/DW4wfFiqtzCREiMokff9oClS3+b2hSo5wX/yrpF2LY
1SpToEnj+/t+0bL76MVHASWfxNOBvfUh3spS06s1r6U2Lovnn/RtPsmcV5yB/s72CSC7hcoLbTbM
yYow7EcHvdr8xYIy0QtTNr0jC/B1IemV59FJBWu+naKEY3noZlU08IX+Z2abBXFSLo2OhER52QHz
jAbCA43kBPSfykyhCZJM36fZIMxViriD2uhBhH+q2/gA9nnvYCDieLg600jTNoSFXADfhkp1bB58
92xRp3surlPZmRWdYRzstmpPXLWag7Mt7AiJ9ttc88QMZQbSt2rufBhZt3nGq55mz/Hty5WCJiiO
vF5U7aaAr1OKIttOxe5B/UmNt20tNz9DG2knSBXdt1wmR5D1upwmmhND18TUnkvwmEVeTrnDvRV6
jVk8VUoV534YJKeX/HOhJc196Y8Nz7X6V5pe+VulRJE8MAcsXEXFF4QiEYxOhfOR7MY86LBgUNiq
YVHcXaTuEe2DIT79tD8K5idn3s7jsynetd6DY2mn4cnnO8xAgu5RvKvOpDbD2MsAZPVGRMDAN+Ow
SaNVsXuLTqpJr9vGF9nk6OJN2n53NoIuGNw1h8wSY60u5NPyrxVZzfIj3+40eiGjLD0j7x7785p+
21sktQJbEyXl3VUBuzJV908rWoRHr3uZEcpwzrqNOjXR+l2nqXNPA9i2t1f5oKTTSPi8Pam/8sIA
hgHHNgCf7kb0ymBULRR959Lk6rqlHlXjphlZMSn2+uCiSGMcGTTC2KfZQUPXUk1ojsxxvXCtT3Jh
apWZbc7YfP9G5GKQzJtUHMZPjs983mbBpcdZPDBjtYtdMSk6bSV90ARaNzM5Bw2MSQfM1Z2WLXGL
qkcdWae4nULvCOnlcskz9cRWZj8FQUXe4O0LTbzkQ2D2apVh1xm9KtdHbZScPrRbukASV7QjuBly
F076aZ6izjVlDGQ+5fk3/uHk+DHnEIhDmkZjYNvzHMxrqa5WFHJ6N9iQpSKgAPpOMOOuMfTxYLwo
uyfUFOX10ykNQO2npa/qB0IDt5BvQxbvAE4OxxC/s/YCUcoFhYmJe/glPGMuaAZY9gzZiuZnhUuy
ZTP9Nqm62bs/W0fK+2D9X19dp4Yl5BFL8xvXFPLBGT3yOmM6waEjqgpMPUeud2Vq3pPOSUuxhfMN
fyxbsWpPdhIEy09YHstivhT9rjUmOl3ss2MGKtdCbqey5YPFALKC/Ps7l102xWvbh9q7odl9Vx9B
oMn2XdmVNiNlIktUR70DyryRZdCQdFTtQyHLd+krAWeQ5wmdI5rYYv5PYTQoBOdWLtIsv5mbxB83
AD7RLqTli0nHqilzUOG3XtsWWCbNiMDLlABJa4LhCOLpvlkCQttodsYf5JwP0wZtOtXPFRm+us21
Ampak3LmMyD6mOYzswzHkJgoq05kDLOv26pCTY+44C8uaD/i5Ns799r9E0vbLTuvuDouEhOn72Gu
uqZAtuaj7y52dM1S0TaGpSR7DveF3a7znN7mtfGGqrrQYF6aTPRxLf038zmoH6rxsrsOTYk5qXuJ
XamBuVi66sdX5M/fINyxBX1OdhycWw57TiFD0aAFd2C3ATUUbAi61+l9nE6I62OIgivfzPWz8S1t
u8dOjiP7BwAJg8NZ4g5/Ya2vZRs5iNJWp2SSp53Wtxrakj0FiqVTL2Ol4H2XNSOyQTGcRmtOWD3k
Nx6hnb//AIirGWchtxWmc7mah7YH0d+sVhvhM6SfkoaztvD/dZ13zc7IJ5CDKFbWN2U9CONV0S6b
692iXVQ9UHKAdsss50e9m/y9e7HFXAJM+F//AICZtUfDzzZd2PTw7NhQ1oc5g7gvYWblUTjZAXm3
T3Ab2jHkITybeh/j5jhfA6pAqGEYAtHDopNB5swv5EU3+cCCm7qLyLfAM2d5ujilEQoIRxmoYyE+
7HFoaXqkvqL+9BqbKXeCJyz6Sxt7x2Q6ryq6yYmdwVUIfPcYFEk0ghGkRZvKmo8QYPTAqKLdOO5u
aJenw9rpjgIR5dhCbD3ZOwfj9qwFokbb2qy+uswWMcIGnHL98p3DwLzBQmzzLztZXcR9w2eSPqmu
kswNMDU3mzDyEGriIMKLFSXTXphx+ti6wA6Z0YQswhHc1OSm6yU+zwHtiQHAdwpvSyBPah8ui7Lf
uQlIuUJ0+u0g04VLjCUSfGCZFO/KTINvf6xDORPIztej9NMMuOmZUxOfBLuRGJCLGzJUALs1jFIS
BrKbebsoTDq0WUtPHSrW5BB3jQO4L4esmHGi+bSMI8OXKe7IlEuUSFnn8/f7ELitDW8t7quOJsAQ
++jeMyjwtp9mEDkXkP/dDdU0Z/UtCHM91D14EnIVl1ixGupXFtD+qeRmtAzBPOqubwSmAilZkfY/
Wfvihp+9fMzDG/rdEya8lBR82jr76Q0oeGKaAcmGeZPU+UgLDJV/gYFyNbJOYT2fySTaAtJgORF/
/rgGonF6n9H8+2vEIN6BhBqjcnGSjWZJVW9tYvVS7BqdhFSXLToe5BTlIgbFTaZQ98LPkYt8f8cf
FzyUy2c8Otz+VX5Zu+Rca0EjGxhjGrCQBwSasczBOsRdHzCu8GXjUaMAp6coNx08UIFK4BA5lgMb
kxkjl4VR//dsYH92c/ao39iFewqN1vjECeCEPRLp+GgU97GwIOQaTBJ+la1TcFPXJPu4spqK8Q1v
7fIpuaeCdTl6QZSkk29EWo1CGADRa6bjpe+OOU+8UC+wDMsbMHAVzZYICcAMqGGzToNQfaQF0R76
DLNYtkbPzBMqpSMd4o4gki7zGIGqvGTMrPTXhSGUsCbdNoZl+jAuw2j5RmTwHXjh3WU4tvNq+pie
GwFvI6W2yFfyuTdRc3P8DyTTBuyTc2KZSrn+Y3ActAHYD2Hry6KwiUjTH6AvsiR8U8Fmw0Tuqc3k
DxRbr7Pbjt/aSxKeUXsxtNmeLMBO9Z1YOZascuGWx/XesgksRfcVeDnK4kApsABNuDnw0LSCajSu
q8mlclxPKZmH3d5YpoOk48VyGP/touw8XddF8LmtqNF2WnAPaF/YVaS6f4OO2CScfZ6eg0xcLtu7
SKYaxmGRM17SHvUskuOouQllEB1rYlE7ZMxnVnK49fjjqiUss1UqpUPvsxXzK7FbZ9IFxuyKj4wp
G4rvR+y6TZYBMLBvuMtq+ZSWByDBZd6ZJ6pbiTU6KNiNx0TzlfANzJlKNHjkIJC9B2Fqb39R7GHp
6Mgqya2WZCbWJMnU4ush+cC0cwvNxCnYWiD+WZceCJZF3LuHlbfG6aAXnMbczh7MZLS7MkcXIutu
Neizn3ehF9Gk8kT0hFjL10eGxFiMTPFt8H8QW2zNlKitZtGaM9/2OXjsrXwZ/j7hkPA/MHwcvAAb
XOYKzE2ke+MkTVcCROJVA3sZhPn1dw3LqzjgYvt6i5PE1sFmja3xVFu84ZmV+hntgISuR2blmnYm
/Zij70925lMAcKrExFlz5Z+rdyAH77e6TF9dKOsFz92ATjXlBtaGyXGF9+mEecV4XIDJnzuLG9le
8X/IrwfTjtkJ9eHWT7EefeTR1Gcll/BQTu4xs4CZYqUfe1S6tzELsQI9D83ogrChT5krXEYvFLI5
AN/XwvPEgoJ7W1JmlSA/XYEeW8ZwG+XKreP8QY/KV5SrYxYRYVA0+iV6kUojGPVhae3AEKqI/lrN
Sjs3bw4kwriH3Z5jp6+0EFHqLoNe1dz65bEVHgEa+Ri6O/0KGb/6bMXK+jYo3s9YhHAWvI3cyzo9
i+Y0LUCOmVnveodBxZLlx3cqkCxiNglbEbk7IQ54OSouhJ92c3CrN9BT8RqRluHRzTORCfJNTW5R
tB2bTP3McwBd+pxEqf1PJvCba4ZMNgLSOh2iKTUsW8ICzlUXnX0GLoxpPucsK9X6vrThmfQxzVpu
vT+pBim1Jtf15haEO8e+eHWaaMXqI0XcDuWxPa+Djz5nUfQLTdU8lJqLIxeeCezOhsE2HcebFDuX
bihSZUez6hYuX3C2TSefWHNn7L7AEuo6ZX91z7yODr+vLgZdxNCqnJIHVTkvZ6TIH/+ccqqvUihD
ajf2hNDyfGd6zX92dz5/N4avhHoknjZbUZsoxrZT7cpUxrWqONOeHpaTlus51wbEcb23DptaoLcU
Z+h9bft1FrpSZz9m9lPgnIv0Tt/pfGhvlQDHDjKXzwJ/BkcAfD7vVZUXTJ89DrGBklaxUwk8HikF
ufp2CsR5Mk+Gz4zLJvaVWrnsu7bzETXQ76SC7Nn3oAZmlJQV8XzveJmjjVhuZO/IIPABI0fCUtqf
jp8e1cyQQ4mX9ZsM84u1TnL4eOXVkNGmwzGNfAV35yqZ2IVcU3uSmBhEC2a06nwYPT/C2aMbrE+3
ftoyppZJ2esrH8uBzJeH9H0+iSmBckxjrxdxn1ZZwyp9xn3gaREoDlwpQJYX7qZnrvwxcUt3kj/b
mvn68KGUrAsWabDNrRqTVqYe8+gtv8qr12sGmLdCIOewNYNDcv+xfB4RBlyxGJ1k2Ubdi1Z9/VdZ
7kLv3VtfBpNwO7fiYIdXtOW7/m8bjdnvzd892B9R9D+Bm2IhrentHqYWeXsGuhBPfPKGkohvRRGw
ZSr/ZEyCWTJxEBd00VCJuB4ju3Lq7TM+69rncvb3tSvRr9h7/B2olLff+PNhLAHorcLsIceSXlPD
xg5SdYCzYcoJeCSvq/1dpomWaRvgZbwGMB+OeC3o8kgYRL7UdpsqzVTN4LWrJeoeFyqWgWlwh+9j
j4Ij5DXOjE3OyVdG56ty0Xqb1hLfSKU6dGjeQKUhKFoyBGnQzCpV5mk4MvnoZmTs+8BphtBHrOVO
9CgNNWI/LRh8Or8PFZgsXEfidU4PHovqbwfC4/b+RRd/5RsNsQBPAsnkvcuwjJEoM0reb4/dS7JW
nJ0HxQXUjVI2pfMa42UkkQSk27bZqGk/+ZGbgl2jKqgT9tOHziUmJXm4ftM+OqNexUTquFY+SJnZ
Oro2pBA7mwz561XlC281oNYUZmYw1/ugiWx4knSfU2DnTsjGNfK/S1AHTYl54sPEfwWkyq+WmkST
cBBXyf6F6b97Zcyx4sggK2r8VKBWb66nOFbMOB/yEw60cWFE3UjhDCX0C28oGHTLadSOd549inQd
hfxF4RTgLqNFG6qkrYZWbVLVBYqAGZ5995nKVU8QAg1YPzMMpqk+Zzc9BQiGjkeLh+8s923a6Fvi
AxXrCHqGbTVovQQcJilDY5RNwBeaiQUYoHqFLMrEwQvXg6IqhozYhikGL2V+jEAh78Qs3iPGTHbw
eY4K9n7FF0d+PvDmMO1w3M8MvvqYLOeMBkgerwmWeP0CPzEcZ6Llyxh49m25d8C5+g9voKA3AIhI
vrMGkmpLwiDA2rcchF3kY0mPwNhuqJHs85P0aajphBAO/2B0NjB+F/O06PirwoSFnh11Do5ueuJ+
VgaCU8PMZR4kFyBqIjHIRvZdupMve3oe/ldp0ZTQ0EfQhdevIT1JNJL+MDUdeoYbJiJ26wyT7/fP
1WB/8UIzFm+C+HZnuorTxbFXay5exq+qXyJtaLo3YCjIcVYsAjBEecYKpODeqqs+GJTJd2s3y5WW
qFW/gvFZapGqT0XPePD99ciN4dfqM7hNGdaZkEFIdcrDQk+18cEjbuwyjG1PmNwQl+9eHcmnR4Qe
FORa0z9WBt/oN1TefiuxJ+susDZcZfRjN1WAwYRIDqwa+lWH9s2tH+jzPrcLATOKmjxsSPg7EXkg
SiBspFgaQoIujvz6tmkyp+ekgv4mLHb6l1vQ+AAYc5Pzx3YwHE4hs4LSVT0UHoWOLMRGeUODbgAV
uOHx5wAgftcMHfR9XMk8cs06moUwYCxnH9/dllso/uBrUyP6p6TSKPoAQ7igdU8vQYxBtZRquFD7
5pfyXEU9sHEmmPDQyEbB+us+HCT94bLjFq+Yc8hWaDRa9bUR8JHnz0fxL2pHjexK7L0Cd0SVBicG
uySis3eYAGC/xoNZ6jc3sETAzhFiIK0vPBl0o45g21mw4gEV56OzWBneS95r9vwztr30gCYnLCuN
dievFyjhXSExGFJeqsws5MlkKi+XQCvP61SMJpookU7aadlZKUqPq+fZ9qbJ1TauD09IKIaT9vIv
5ipqGaT2Ef24O3kZ+SYXJlqi4Vw7Oa0TKJIf3tME9Bz05eRwB/BxADZhEiSCYcCk7iZreuuA4dL5
m6YxXIo+z7JYYKoE7WSErNR1ArID+VHcssczjZT8UfupHYbio+zLSamHcYyi3GVT/DpYmZQaphuj
vcMqoYy8aUGm42ygZTsSQMtoO96/42g2ftDzLBbmPVkXy/8RPaMC22CcoQxLqImJcG5JbvMUHf1r
s+TeYhU8GduxreBu7RGaMk+UP79cr/KQbLP8VmJBnMgC323gR5S1Vbos66zeOlyhyHMENTW8spRk
uOUnARXHxkZ4Y/x1PJRwzMdnHFeRfxpx9gzBjMlwgTpmJ3cmp1KxUtRiHoa0/KgvYgnRkCLG7YHA
+J7z5cl48uRkG6iPaopzoKPSiDROhh5Rk+4alT6E0LWILMVf2UpsoFOtjEJxdmRw3Jy/alLku99R
/xSAT2nGzOb4AN6LiKqmTw1PshHaOXAgO1cc8iBVINr9tHi0tdiiJ6eiFkBpg3Jy9vt1336XhB6x
ItoHBoi7/ZeKTG+ooyrP2Ig9PAz4SDxHcT9kovGNRkh/XHoqRRs8qYbgwGTrAtVudHpW0cfumMCn
S6v4j7EZMmFnjzvcn6QmG1imnRmLeOutoe2SNyKQ6gomnSOfa/sYF4Sz4x+TlqJ/tytgsFV+vhiP
qGYilszR138cIUJV+JKdWPKQ8UO4qU9kmvOi6kc/o8THYsdCMFlvdkE66Dg1EUc/YePxfvKsojHx
BDVHW40JBv9T4jnUICSA41WFlc/Tkf7qm+IblF+67+RnLmhe6saq+/6teFMGcw8xy65xlhe1r/UB
PxPQUf2pvOpiNtRZahoQoT2VGUxW/SO+zTccsk7j3IWNdF7xVx5M5bkc4DFjFrldeX1jUj2aUXmQ
4luKkIz3RAINQWM8/TAVvvOykcdu3rwHDnVsi0u/k/UC9k6h/tGY/gOyPNEMwUmILSxcD3dXqIxU
inlqXD6CsKyDvk/g37a7ui7XUGJwsff86RxKXH55bquvorczCP+2p3eubXWbd78gL55uC2idSDsE
6UlRXf3lW/0rkXoumuLHnwerQmjr49pFqhUvYb8LorVeeZbGesCg3wOqnEunTRg9m77YERVnQ+YE
ya7PngtSxXqB358j8RomlaCbHcsNG/dgNypzCqoNNKoVYTFYDWG+kW8Cg3Gi83hmUsr7G3AhNvOs
VQJH2aza7/tYHcRgesgbNPVCdC77cI1QsESfNbnbJV2f3yP2hUKb6MZrjF/Lx75/9jpyr/VOTEaE
nMe1qI/wevrTDWMWW+MPMOqtP+jVkWAt3o3LVVpB2Y8gA8DeiwHaWc4VG41MaOFF83Kw+CNCkhqe
3eTZMTdT1F1uPpYmMDtHinr90QmwrdMsomrPmFpHwL36+M5kTr+o8x+tIl50mbFLIiMivRvABhE9
46tUkYSPl6bNzBiFS5YeL9NefjpyB2G/F2iglW3T4DYaoKoKPcaM2EnVVxpVK4ZEAoHsIoE4XVo6
emh9z5kKNL1REwesQn4/aeJoCEqp+rap0GUM759rDCuYKc/b0cK0n4B9nmqV7XJaAu2SPStP+VWs
eR6nXXe/zX+V49Jm9Epkrj/4zamzfhYAebObkeTF6wZK1uSMzne0z0/s73jlR0PM9AICxIo8liVJ
+rbm77I5NefE2YllLeXWqmetgyxttIkTtnT1KY921Jw8wKgefNShug+19iUjnUypC4t3pRWjue+g
WrveQS6v0zdDbLvaPMPNsrpRcuARYf8M7bvb0JG6KtaVooaD2RCAI1ti6wmALkYNEErDOIckTojV
Jj9Ji3b8fHtp2JraJmJfU4I3pWoNq7MdLE1aefCzk9jvsIN2HsTqmehaPHWQlokF5HZAlP5WD2OF
dI0JNiRZksw+6yzsCNTRd5Ju0/gJdqHc3Okwjc5t6dWMlTkCB303QtIcxLF3kC5NoHUkl5tvVHOn
zL0J6zXz0yfDXGkAIbNhq1o1Xpa+Kx9CywVi0Czo9QhnJlac74i3GtkqJBidxiBFjEn0n5UZKCaQ
rEq/sgGD+nLUtEQYyVPdnwqluRfEd4gSR5TMcum1NisCjne5QeesO0gVCc42FbcouJawNVAmKMqT
eKN2hvfZR/z1QPUx1ff3Cxkuo/vEq2F4OgSzEOM9KSv4KoSpLoioCc2gMY0KBqvvmWY2SbgLNYi4
ZHdfAFIBJIlA7eedUTU7wsbVJEDI2qzwrSnySA1tfR91VEvnK7bBqMgmYtMoAfzx5o1XlmFDq8Qy
0p+FrnqbLg/I2AMO9JVfE2k5giNA3Hlw172LJxiQfdFvMXDzahv4cSAmGcjaDQluCp9FpiYnVA+Q
gapB7zXI+CPrx6XYHMLIEMosjxorKY2HLKhGEsTVyLM2iZJCbKkU0TVymt4qmdzmOlK1bNeMD0em
0i6kDHWWbwoABlNAaAfvFfoHdPe4KL/dWwF4/Agtm69Fp/vdV7ygYj6bdPnw0JOB/tj+O4Tf+RT1
Q0ojgj5glZCA9Oj5+h/dSqNspSx2C4F+k1NeFhzWB0743nqVRMYGfzRRj/T5sA9Db8d7a8ZB725W
acJ++XkGLAawSu2aDJJxzOZPNY1unF3wqxS1eQ1iMyRnfSS4IfPQgckNp2CqWzB7BSGyjGUO1ASr
LFBlqh8pYF5d1kcTyB1WcVrrEHJsEccPPHnjMOYs51rTTtgFOCWYykyLJScVt+8NgncOF9f+iBda
zkcr1lMuolS6xzF0WacAKgKcMt+tHKvrqisPpcQsnpltDpsDiUl+H9po2V10kLkbJ/EXPUYe5IOP
88sUhJxYNIKuhLAHSZbSve9qMcHvkuMzfIlYTTuFsUsM4C0TRzyvnRdJByNB83/+3p5wnDlSk2iE
DXVWyEIE+ZSnQqULLqTDdlONUE1ve2YHiy8EeKK2AR+uNSZUARtZvToql9hqbV6uci5EgyQwkQBb
C80Re0/hPAfPOF9TLi9rKRAPH+lwjhUMbTypi1zp/MJkH/aFySwa2qZC5tGKBbxZ/KRpej+L3ymy
jUfLOXMhvVW3nnUzBVwcYlRvVTqEFxzyBs3heOhq9GKH4iNyCVRZfYxSpQPDByxy3g2v1qAHp1jU
SAJbSf0rzvwiifJxlkN8mj2DaVPHe4Sak0ZWhTZ2SiaOrW95HKYzbRxhvaoHFUcwjlt3u1bIibh0
2DqISRmy/Dicnwn7Vyz6BQ+BVTgw07hRHabQwB1KrMzfiR6fi7EVBlBVGkquUn16ReNj1Bfk0BRQ
6EBdSH7oU97G1zNGV9x8fwQwyK19VlTN6R+EGJgekHdcTJJd3JM62fRyVrlWMim7jZUqqM/RtV3a
XB1Cu3k9oco0Kl3vgxRpOuU0+6T4nno0OSfwYz5e8bFxd0BlaEphHIxI9VXShPtEWbdHgIDGWXCE
naSkmbivo7vMR6AP0DKRwQ3jYX0SLB/K7msrV4b85lecmv8/oPMpZy4fuAsFKIYbZNniuBvNBdJR
aUr/fdu/TE33UU73i4gUl6eazMDNwld3qZceXIizo833rwqf5o+oJ1yW3oH4VE0LnMKH2/sL7775
TIculyLKepr0qTRTxSys9axj1dUij7OhW5wW4JjFtGl6vCQeocnSP4WwP9wHdyWwffClfomoq54u
NrfY+Xcf8EeeK4T2ZUpDPBeAZ5EOEVn9/8mTVQxkKLU3LMO09vlcmZa/PQSOa8HlRq85kb3dxKVC
gh0gIKluEK2YA3lLhHkqXhGJjPvXqT/LVpR6WBXRCnzFmAx+oRMVYqZsZZhjMrDyoIYc6U2xZK9R
7+hGjZJ3AYDjM2osJTrvSgnwxpPqkEQR6ELNB+axW+6fCSHT6u+HEZ+INWlIECrP1MrQjixM8WxK
3tmp3AEaZkj0DoKECJr7+2+ozzoF2U0Kt8PsFJnmuFsfjh50iC1negoYGjnZ5AelCwc1k+gze8Q+
GZdGU+AwHCQZLMuctuXZ0RSY8zYCar5p5Im2Abp59s4Vyzr65xAsS0VlUlyeFVfnG3RM0DvT8kAh
rK4rLBtbcujnotqrtddlDyqgQJO5gJn8kZWbf8qUS1rDHNqNJvIlc3g5iHUO17TCtS9I8RWnEGt1
laS8TtliWqvpKYsNt/kV6uBK18Oujr8AhRI9Vdw9JifwN4qoWBV4xQff+RT4B+6CiNBUWB8ftI+C
XMrLsEQDmVOte8+8ZZv29xFpBzvMs9J14l/NScodmCdol/zynTIxerThF7gov2DBqd7YA9XjrmlZ
BSuBeRhG8KPzLhqxLLzuDcrY57SzLk5oiFi1/bIOTBMSPyvmlJwoi5PJeq3itEaT2kHX/iiFNH+I
kuhtZilQ7sE1YanjH9sz0krMBFzU+cwh50bIasSeiFG4erypeXvHPCkfQs4jIBnhIYL7Qzd7NSLk
za8jRSr2cb6y07kYSc6DqNvl2xdOzv/xwcxo3ajJ6Kd1i8jS6jjKkKL6hYNjmXHKOHWjbntZl2os
wsce9KHUtRLN5xd7k3aUj9FLKy9SC5w1nUM21ax0GFZthWTN2KwmhPyiK8rls5uWfuzRNQUkGm9e
QEKJyOGi3gI8/ZPE17bzG2tqzebnXypO27GKtR8itrZq8XsUVViWTLVsMriH95PsVByndDYz1/EM
SauP6sSo1K4Z3OEGMmGNeI+rV8Mj77wPdwApaTp40cuJPOEwwZ8EwwDk2quXzcxGBLG4QPg+egpi
hJrPpihzJX7lzu//CV2WlTGt+rCwQUui7o0Lt7Dt2sN5l5pl8d1jo4bb+rBksWkZCo5Z1ghPHyGb
wBg8Piz5+L/6fPYUmqIoVdoyasCgJMh1tX9NEwl97nPyIBGmRPa4M5rORtcPOLFOzXTmfItxX28i
oiWgVj3Ua7B49eUorvLmeTIvNJtpQ6UgRnhfHtCb39Av3Eeeo49EtAj/HD3XxO3RAuhKSMUrezGw
dYLrlB/zphG27VYI9BX6ogDMR1SwI0Q6g7g9N14yt0CcWIcmfwjg5P7oWL82f5cqN+cHK61vSuwc
x0xc03//jNGUVscvabaaOpibPW78cK82CXBa4WB1zr/5/95x96EQhFYJZmkDCIMWv0h3Q5fkdVXE
dTAmOza+SopkHRsuZwR0J4T1NLN5helAVMU8IjDQxcVrvKhTWII/YE3HltuX7SeVc6nfxPJOG/G1
/2UDIJ1A7Ltyhk/2yUtt0hRr0HfVx30a2MFCzz8EpL5jYxOtJ5u4E/8nW02HvitNM/0T56JnRxEJ
Sd8zeLDPwCslqfVLoYzoOYt0vvFB4DSd199kxpwDlyQCDZzPZs6+hQNjViwQ3fsc4JgLzLe+7t2q
ilZ/eVoTNcYRUGwttfz0uIrAZmfln+Q63Fg/x918U/KV/V0jFHxI2Z3lIVQc3A970QKsxaQ8SXWW
fOxLm+dxJ8+3T2G7eucOaUj1jKGKtRtOZkqzqs4KkrePy9oVHfAuyehytNYjdPgMdOc2bcoqswzi
x9BqP4ftrQurYzQhWQDwuSnuolJJhWZBLN01uLoY3iAG9MpQoGBqKYbZ9GJ7q9tOmu5/dpGsPhTb
xT0kNr/8ZukZ0hmlv9IKFSS0mGrmzMXzKrsgsZZ/6ZsI50QV0ql3IJCaJbFCY9j7eEP/Huqfz1j+
NowYZY7VR3nFb9ecl93ulQV0D+c/z5BvRtmzWIKmX1o3DZlbF1tHXeAEAIcRcFk8ZoobVsi/j3E/
S9P+zaqSILkQQGiAxw8ZMx2cUfcNY/BEi+Q9x4E3z0yoznJbqxWP7jwK4F3HgN0osqVwEavFmQhZ
ew96q+WRyLJ9551HepD2PGxJUYQcsa6Z+MbIBJD1liJz/mX8SC0gpGn7cAoELPKxi39x/gSTTOBF
ZztI61ozAOcH56cM7Ku1QCPbkjr1NJwy7MZBH882OnJoohm4gDtBs+bKykeUeLJVmpcb1zkn67Xi
ogBuEIm8mzJ38u64ZH7DAqbu5yvojsrPPXJkhWGyml4SKp1EGnt6f8vIp3K3tCABBbZEoiiOfhkV
2xk/Z3SekKhQjzB3rxVAa247Y1OcQ99uCrgYTWC13VBgr9AbqzByU/2LT4gPwgeYIC8ZMG1AAbea
7EHIdywl/Z+tkmPkjWMykxC6g00JT/hjBuPIUBkZglXSqy7slfvtqDl6c1pD+/X1opisFtMc/6h5
Pzb1HTacYWHN5pydtEAcqdC9uxvsGI+9Aqf5ts+WWXgtfJ81NvNqUtT2/2/Pa9O2w67CrnZ96g0g
4bRTT4D7dLKP4Kfd8TCRclfmRwYYhZ9ZbeYOy3COGfl2SQMUxg6JlfWVI1y2F6pdlUVkmNutUGlP
IlTGQ43MSNtE36UyICgOxbuwrWL61nzPBdHr3eoqrgge4ZZuSMtKnX2YZS+7GTmQckqAJi4KnSkJ
jt2cVnb8C3Br/vRAMKu+fDoGc0aPTS8FOuV03ZOSvlww1ntVzi6RBNREl/8gBXQgchTBHURODYxj
VL/WBVjYvRZ05pAtAiSan7KtSpOZK8zMWVgawxFJB0lLVtf2eTss9Prwcqjyvf2aSY7SdHNt07Km
8T81fuHr1oOQP4EiUXugIB8Ux8QqwcyQon2GBhBvF2NUgceCcwmUeXV9mzDF4iF781FH4vixJDTH
yywpLoEvASzo/s5D5LUYY8E1jvkirCSSidQGi/rQ/+/0qOI5CFLL30dYNFm6z2WPTVjdJNsQjyAn
7e61LliSRDQif3IvGHgi1g2oJVjNLIi4OCuAg4ljPTo5woEOnDTTs7ilfvxGI//YTS3Iexdi07An
Gs78v+Cn7MbJ8Omgh+TvB2RAjYiWh1O04korfO1X5x0CKxRY+y9e4dC6oChWcNxCQQ/pE3z6AoeN
I5/vQ6myl+zwrnv32qlqRMnyTzv1eMj1Ox0FwSChiDYIubnSP917VrFM9wWRXljXBksxVKFaCOp7
h7Rj2hVkm3xi11WwpO81r1tn776N7Z1lzWujkGuVlpfQSfLl7MLkk8EDnE+dp66r32SOXcQG5E4j
kqEcS6FIF8L3J3KLYVBTdTU+oack3GsjH4Fb39cKzoVoBC14k9VRyLfD5bumgfMvrXi/1NYaSc3S
LwXHGzMVJciP58Dlb2owNTerRGhiVrL4vzxvA9CwzNTPCsjpPs5KK2WUn3XXH1hk9fKYm51JwqZC
YqZB79uKYL0DKUMsFdEU15VuoMgxvEbNz18pZgbALLueiE/FIVypNC06B6c6x5oDdOYUByj38qtF
wi/SUIdKs9Ra/vI0fLmLiDpAPn1peOIqeA89LJWxaAAEVraLO81NHFHuL1jQ7Rm/WfnGaiUEOuGD
3RFdfyjKwKkbiM4Z7++cWJw/zFRiVfhWkMtbu84YOScX+94yqR1UxIYI5tTym080m31V5K+jVBGi
yePtjrGgwGITfl9tCykfpJ4tGdPfdZCSNYmSuP4xJ6GxwmWVQ0+ReQVbgoAIzfkeeYO9JhtwobAO
m+zwQZY/e9h3CixVO6Vw071TX3CVThTCODr652qbXkcz/AjX7E3t5it9nBd9RcWleFiYGNrmKSIz
0EoGw+cmNqg+WPcTEKIDo5GvHzt51tDGbbP24/oZ/Pdas88DMFqz/77AorzSk9zOGV0M9attsVyg
1jtLQsSR+GmYK2/wNMV4KWpz+5mpEFYqjuDXqk0Kg6NZ2RX0sa7Eu9lWWwFqH2sByXdSc5pdvys0
kx3BYOI/BH3V27nQIh7vGQABiZXZomoDQnhikx7ibNQbA+3jPYg2tU9X4n4KwmIo0f069K0tp17W
/RQ4ZQN3EyKThdaxQlqQV4yRmWwmzVizwLMSbVwwcT+HCk8wJ2w9XAq0MNAhhfdJE7MRmycj8zY1
lOYBM1Py7Hhbbs5M2RheDtfaFcocfDn49ZnjZy5hTyDa4A6AtoLzbPsYf1tqmCqIwqvTuawfWZLE
jfI5l/XE3sL13ooXXk6RATP5ysDkWG9y72KY1PbafJb/pEwey7Uqec0iubNJsocCy/QkavuEjjkt
YDLr7Tm2XPOT8WeUgLqwTpxftqOx6MkxZ+zCP15JBPLcsQ9HsM6BbEnbi8YnjNDB8CMlDOzdLKOv
gvxSkQRHPPkiTiXPRFPGADFuxADWYoZ0YUxP+IlXKnQVNvli5beinBfKJZ79uNNcZARuRyU0m/fh
Bz91i5MGZ4BO5xl9ZD20YgHN4gt349AzqYeeQgRiKudSluk7v88r/mav4N1kMe+nAmUKsCvsCRyt
cvuqRZMQRx7asNgrbVI4XbYNtDau/UkGGiuUZmNwo5L4elMOo0/Hnm5u5LLtEJjrSrZ9v+cfyIFV
X3NLV93qsbLLm7gTKd14aGfPtbHEDKTXtLGNYqIiSYQj/7eFw69qblGPPME5K4ygszgfr0sW1YIP
5ivB0UnNxVQqDyr3Zu9tFN/sr7AqOuJzC3u+4yYHb2CpM/vhXgSCdySBrUmA/vi0CdsmjVq6gU3l
vdkybTuDbzrk5BwB+GKmDwYatRvV545ZkDiI/EuB+Bzqdann4wohwMdKtmTgS+d7f9Ytmuch1rJ4
J3GO+RXbd/rGXKedOrIVLeJD3/KQnlZ6/QBlKX+xMLyeY6rSfs/OqMHHpSxkgoMJe7bdNBsm8NAe
7AoMslDxUOqJMydKun4GZHbODU9weoeYdFN2s5fvEs/jgO1muryGzliuj+X796txA4uazYkRmc8M
ve/cxfSgL2KTGxmp1YE6C2sEBPMzdlg8LxZxaXLtjaFP4SNJVekgbvNXpCgVb9vGTQ0h3MKL1uWO
nL8hKpKs9GuFxwZNU/7Va12hJUhJduks/1/C9/GcDxFFc4/PnVXRljMpqLIkDZm13C1kAayk9FHk
tWif/Xwa6N12xsLp2kqHZ2JpTaRIljs5cD+aRtPmE308yj3UqrGuQJ2BpmC3ieBupx5vozEzvw3o
Pi8uTD3maSvAO4sxhgO5/EZ69mMcRuN5432hYiLXskBvPrCXSRQq42Wb2HRkP2FXuIkYxwyYR66N
GK+jdPOoW3QcOFkqwc+fixdh2acJsFULXrJW1KNI+mmvmAsdBY0TCU8uVnpkzYXCK7/Zg3Ru5Rs0
5EXsTPHYYjJDByD2uV6Z5xd6CVFos+oZrU1sezZ8pofcGGoI8/+GXXb6kx+crGCSZO0S2P4bhRN7
U5Cy2+ZzLPw7+avEuHzXaDboIPFTuoqN+I1VRKRcw9qdCaqh1d7b+ZKS09IinNDoFYsmPEK0s+ct
LTW/KTuKmMY5gnyVXSTk+aD4nbYLG42d3X6HeBYcz3uijQ5v1bPCEZ4bHNRbJBv8sCwAvoR1wRAx
E9OvcrhkF+Vit8amjCuIJaeaGL0qMmJqd5cUbBuETc6HgXUrAmkY04zhXuxz0nAXyfhnTzHCXHxf
MUF5laR0GWTVy6ioFKQX4tOvAcInBprd9/r1Ts+qe9f9aQI6a5ry09XToECmDedFjcSNSvVaEtFl
Z0UaTBa3vMVo6/AK5qZFiCdDouZTQYV5EfXWlJFFmNhs05eQ6wrxj9zOjCWevLtAzC2rA0Yn56yR
HCkwTXCXRtDFMKQZzBTAGO09PwDRec2kMIkHM7dW3SXIf54uOir7gPR2KNWRgCZCnRTPSoqSV4gE
jJQtsVvK6cmFg8gDStyz6vP1tM7xYzQGJk6Ofw/Is+ROBWJ5HpFKftvpUfthUlvKGlJBsoe2Szi3
y3t4SxmSGPvLI3i7grFsPOXMvftjzX0MFUthCd3OSWX4hrN8nEewlIESbqj+sstR8JYeHib+VSPz
5QxVmIh2/gPSyR4dn/G59zWes76VC0w5puRWmAjxxj8FNVedxdawOk+N9dwoIY0cEh4U9ZuKuBo/
dX6rUScHtoNXuOl67XgU9ryrU9HZuvo5O37oxbmLQ6sAqowX6fRePiL53iaIKbR0Z2Jbbi2pOc4g
v18dZpSomtcI0d6bp+YnS578PA7VzcqP9etYmjP0Sk+C60+F3w2OvCEhW/lcKYcrIGCuLJVipWph
AkMKkmfd7N5bnBoNnytf3BvRxDD35bP1AiIQWZXyimT4918+29TH2ACwBZwNnu8xnNj9+3448qDB
S+/L6Fy+jaunoXU0CQH/6IuZG66dnRuGCHnACPMCmSUB8b7uspdJKWhLBPaBfBZm1MG3o7poqniU
/AuPldfgxTPWrvZ1ctftFYTKqvQBvDMb1houW2pktWv0GZzk+FYq35c4IKon7iRZezVymL6ipTPw
N5KGGB0RX+u1IBhrfCUM9zEBgK3JLTuE2f7coMsmO0GtoyLQZgjdM8do8SR0Kv2xbWPVtUNvTtEU
XV2/i7StZeyucP9VYVVvBZY0dgTm4mT5vHyG1qys1jdXTAZct9homQLgsHQ0+135Otguj11/t1k+
rfiWnJN//mJYb+k4Y6G+MJLvZDfjWf/+b6YZ8/aegR9nz3Zhg8ecsmUaapnfZaiPy+F3B8I8+2iC
MdjVBu9uGmKPp/07jRvFFhgQio8Ny1ePbqvBmjeN4K2wOWs5EuywTCXuNmZxd6zdiyCaPXfwV9u0
UhgZZI/LBaVDxGE+4anpLb4D9DJlwUvJt7jCxJbcnVyrPY5qIy/AxgT/VvXJWYYCNsM+hiiSJ7qg
oY4KqctBnRy0grfJiZTRDUD0UXGGyZ1f9zKzfF9SLajfjO3iR1CP0ThtCFjJ17mPpCZEtgygk/KS
7/96w2yw+EjSuI8TNeIBW0m0o1NYPQ88rP94iSnizn81IE5Afdrcys1JXMu9N/ueIa29nfSeo2pA
Gz4iq3lP7hmZ37XeL+vG9KzNZiyoOIhh4lBTWTNDTNCy4JrEOpTeKuNI0H1K/fK5D7vx/SeHgewL
cy4F3u6tbJWO0mNtvql4GpRhqSQurh858JCmkU1+ls915n59w/wJWYq2ncuZM6/gqwtWhXNV0+Lq
lUC33OGJJo/7e6gHRbz0quOnAyVpSFEqwOvvcRadMHQtyi3gmpa/2F32pdF+cfLGcPyzNn1H1z3A
pvBSf0dkA623g88oU7Xy+wEkh9v5P/YJGetsw5V/DnWADsUsDxrGtU9J+fY/CN2X9Uh7xcQ0E+Hk
l+dusVWbJPX4Ao5l3Vimi7Vsvuf+9kz0HCFOGfM9cU9JaErcFxSM+aUF6OoEXguRYBqmriRsgrjW
y8qjD0YuD0r2DErad7lnmaZZ7pIdyeGPNjhlRAaoUXUmZL/tt2GIVTSQXCNOYNGyhMC4FTr3HU86
EM7+lTjeoEHVQujwuRw07Tw87ymjnfF7Ew9PtYSpa+XmHoe1IvkglkO4KOxMpRFP1G/MjDrt2Now
ETTI/F4NqIPZpsyfBUi0kuKVCPSY6XgmuaEfbEo84hRYJZ3eUJgvCbgMt/BpHmMIbWiiPhiG2Gie
FlFH4+ZBvnjOTDN4/bADi/CI0ZqwjvC/5m5VXY7juwOH8kW2jjL5oOip/AbcaahCOrVMsea1AzBM
iAw0jI9RsxxvmDs+s5iTt5floANGKvELbg+lAXO97uylTjduWSWHfUCsekF/iSyR7IManEEiQVOS
qp7oZUdUWqd42YAFaltswRG01kKmtBDjbWdx7w4y3wdWfab1w3cV/9a5CYYJyj6NL1LtMcr7Ehf/
Ls0Z6v6Ax6QjDpeTFwXjUfD4R4e9WXFUl8ZRZCHUYRvW+kTonZLIplBTn1VJl5UQgyUwSPgqb+LK
5V3bsREOfprX7aQsT8UEdc/xXHeRFF2o/SNCgHD1oJwPndMKu3jPzoepqx+Qh1aBq14Op5j1KsQj
w6YuxShoFBurnbhihSfKMZgRWS8NgL/lty9Tun+H+JGNeoEpivwobN88KdU2kMkB2GbWDA5VxDHh
cw/nt1v4JkGJMCnqkeHY1OXYb9vfeHiJEKB75r3IQ7/BQOIg0KBK1q9hRZY70HnA8y64vQkkCIeR
lFOm3Dgvv/1ZfeywRDmYaxycEFY/z2uBPgTOEJ87i80RIO3cVkaU6g/dDTnJk0sc2Fz/rNKX4Mr7
BP0TpULNZ0rRXvxXgMHgpD1w4Fq2MzJ4/BkXGw06wcxI/j8bJGi4OUKP7/wTHXDJdFq6eO2LOAS3
TnHp2xrJwvWBJzoI9+mtvUPTaDzoNej8eROjQkHEDwIa4gOPVcXwAwEJoxLj+4V2BGH86NOCqQZ2
5RlGV3FtiIrKu78bY8Thgbs5ihPDvzl8jOJI9zUac2EZfhUaqVpUD6hiYBfdRorkoXAmUrZ2tnEj
j54yR3RLPsXI12Xr+euM5zsZTaNfuGykEALTSiNqxSaIHEnBxjX2b9pAtoUe9nhDOPLxUX5L8MlO
GwbcNqGopdxmlZWIY/gP+8x5s3PugyxW+6ZD9T1OGsfgoZfFUPxRbFlu6GPcsBE5BnG/UcIM22I8
leike4WtY1LaiPf92v4dFBD0zMlSDvwkyxkMGOeOyl9GACcaBuWDOgFzJclgHUMexjCMGi2B3TTQ
/v7xYNFjLKF38/cMJr4otTSk9Bynxu2ynkL3wDZBLBqH1pSE039wLppEGTo0WrQ5vAhyJPy/gKAx
9Ly//LHhWs4Yj3/cbYFXFF/9mC77ecnPjbK9P0p/E3LG4iQzHzmpEWighMiFLsXyXzsjdwnuW+iI
WzvXlAW2nIhvI307HJaANzgtmcKr6C5LDcFB2zX21rBy1oQjxHAUyzGjfUJjIYXvA4hcMC7at0CB
N2wkqkBKh5Qc2hnvo5c3kpcmPF9msqIvIEgYiJ25U7XxomjualGbKSE0tj42TIYAPduTsqChCVSs
AMQRwJIqPwx0djDSey7VNa8JamPu7iwV397q5fyr9jZ7wM3QfgCDbHZkZoLHVjZC61+YJDQ9v6Gx
NgQZbcA/cTyc//szo3y8SS8SqybpSDX6290KcirTp8CY00T/M2pm28wAG7GJdLJ+iVWpNVElza8E
QyNgqcASvGMI9TUQPIQfNitriyS14nmXBEKhKyCpS9O01BmKw5o/eAPcuf8ZuLIfRF1cvkoQVodK
elf6OPa3yGXSpnfTdXLqYDoK8b8Ncs4sXntaKXsjfRUU0sQ/4nmpkwRPpaiw42gKAst1ietNILkn
Eanzh/qs/0djLs5Ec1/fPen+3Bl4o6qJxAy/ajy55nYEI6Db2j6XuxQCq3NlWU3ugXK5Wyb2t4RP
u7g718mtHOaOkEOQQJ4VU1+xXRNMw3DezxvNlkMMHc1jqkMojxqhu4jDnpLZeVrPxjwrEOWTHkAQ
KaJX7KQqDBZSpKeAkdYsEGkytZbEpnxLAN00sAarFLVKZQlr7DTQ3hAvuwNduMbNQB6uCtcF1bWw
FYWeUmZhua8lQnzIStU/i+9Kj3VS3ioj5TRUK6BbGZWqASLnIzlodHYMd8jXcm0UQ2Bl4QzVWZdh
+t2DSiUYrsgP4vnNPFzzs0/keRxXLGaxi8AHqPzqUChrQTXDAMjdYwzeTSqEnekBoOhxSF/z0UyX
GqtE0F06oBA6Amu9XFsGhOkRcZty/gAhI34/IyXNh2PDjAHFqIFdPkaYZCAivhanR/wYcW6ePwUY
d0vrBQCiZqcex6OyQ2BdYr+LtGRz+N4enX0BpOFUnm9FAybj4gEEqe92c/IWsdhlgpgWz22I4Ujl
47ylJPNKnOen9i8MzK3EmPIbK886tvdJ5jZ9cCL2xbhhjreXV3pvs9zyBxZB//FgCeci0CNCeqfQ
9VghODr4nN9G6l6gMJe/hQr/zVJ7uOXOySAIUWKMfolGGf1RUpycC4AHiQ4kZVfi1qPKa2vD3Stj
/HNgvl/h5U8MYEyONwj0kbLvCc0FIk52CLAeq38tCFetMZACR2/8pEUbSM/Rja2l/ERuhHymczZs
bHNb3IzrO8j7IAvbuifZBVOgPdUc7LQpTsAgctNTSqMlEer4DTuySQG2ByJjeBW7H5sU0SM/OfN4
LqfxMx8bFXbM3jM9mVQga6DJqtOY7cX6y3n/8+YyUU/KQdc0COVkL3X4aNHtvshKR/EPatVk7YOv
bBXUcWKg2WyOZQbsPl0FpcCShgqlbtOXjin3zEMS7nFoEXSp9kevX35Pv5rLjn4Ro1a1f07Wgo2F
jf4sm/6s7GFTR27kcf///o4Lktr7Flsi5xj+VX0tVwFAFqq0NThU0gdm4wB+bExccKgMWqA5rO+a
qadDNyQVW9YGm2Gqr3Pkiwx7tUBxjmud6d0RoV1Mrmtpi7wKdYqSLdwmyjawPmIkdbdKjhxdcocK
xO6z97MvywbmLEhU0hJ2xXdtSWJHUCG+lYYw/9L7RENA2LGT+FEvmxKTqpUetn6Px7/z4NKdmCdG
k568e8p2FwL0SClfNTKhcX8v/wYPVfX0zVfdDmwotx/FQj8Qd1yeBH4BGrRILeQRDvYOGAkxTlZL
AxVg1BJn3oc9j5GQVItRLvIm6G4G7tOm6hMqsU/3VoAeO1g+EaVBXJKVj/zAhcJhK8Z9STO/ZfJx
evU4b3+k2+wQVoV5AQR2OqCHY74DxLmKvvoicuOqWXRuaJmQ7RfyYdhYQlJOJxwRTsMITJVpePb5
jXfgnZ0MpTvDLWuvL1+4sja3Dl84ZQB7Lhbv9sE30W1dbuIWFnJM5p7YTbgIxl7lB+RVq/jXAJa6
ItF2CM5Lu2zzxYedJohBnWjKntaaswpIeR/Jnjj5QEmLlH6B63AJUCD4XAzrtdtyJ8qZdI9fhap6
4Le1e1TTDBJZaGyfu6R7zpRMTZhLPX8buQLEnq3PcyXPIoQ5GytEGy204YzBT1SpNuYq9OYz6FJX
0DD/+SH/8M5IB++zp5ZqTOeaMsC2v559RYdaDll0FqgsKfaFEWWS3VTKosDKWb6IQ/Fk2XOGayea
vvCaJ+iRjXH2z/6u+bMeNQ948iqRgkyNOm/XAfPXFh6NUTR+mdy3heexirEcMhk/1VM2KDfy8Lvv
UUQ7NgNXxvvA0CQXf0C6H/bY+oBMYFa9+zryDKHIYx+/870NWkG0XEGgmK8pF14Fhj6fHjaaQjsp
rdm4rksMABU0E76vcgLI6J8UO9nk2h7+srjTvLRlHwv7L8txysBw3Tn1V58AG6ssFhvDL4QuBSuj
PvUHnS1OJmjyBFuXR3bgI/KPusKiidznfaIQIGht/tcbXbfrtq8+F+iDOXowST1jOwBQnugGza+z
YO5h3r5mAfJrkEFxUw5+kFw9r4HPXwQwE7uwbTidHGtRosWCTpcJoiSgj3Ml0NNlefnq7IjDBP5t
GBT5TX684Nw/LZ7/rn+3qdEVHnv/jWqhws0Bhar3hcnlaRxufhzKkUh17uOGTRNWemiOp1Ppq3w5
xeFDI+4SYIJ3FZAwcwcNRPsbckygbA7iMElfuEgwAnr4eZPZanWPXO1UtDuVEkja6sHZhjkJaThq
Ezs+yMoW8OMO7zJdt8/RgFXxB0V+oYF648okWYAddS89dLzq/VVkknx+6S7Bi/mTnnKKJrp1u9bR
sbK4PsgKOsnJ4HRnAYR9XQypdiIDRah9ABi/d7dkAH49yaZMBC6SBaLGcq5M7cBz9IV+B6NnaFI/
/TcjdwcwogcQOcTiVYmEfJ1H/t+Wz1GTQ3jlMCSojrD1fFBkHb9e3e6w0woGr6MUUXWJOuWTTqbU
V7uBJV/mtvwhRV83Rj/xi3Mq4KhPt96uifTzYrJVQuzpDsuNZmAZp4OjbpgRJRYxz1YLbq6rcINL
75zrhjAUyGTYlqSu2kRgU8rEDQDSN4VcCo5lQE+vLgox5M+CPqmUKsu3Uo52alet17RMp+F59EAp
CkFdBzZ0c9bdOd9HPq9mVCsem5Izy4xjTIIUNOxcZP9nWGpS6KoJzZ42r92Rec5aE+StDfu8mBt3
Gxwxy15vRnWWluglLUx+JGVNPiQpOe47M0GEO5HzvGJ/aMccZ2oLVDCyR88MTs72AM0DK8zzjRY/
ByMX4IhPlLthMkJEPm4FXhxsbaOlteCW2RrgBDoZ3tqsqwCiNCdl0ymRP41J+O4Uwevu1774sxKv
FHb9HqQGV5eL0xO8H/xhb0V2rq2vR6reYlDuCdrLSicOjwFZVgxLhN/9fpaw8aOzxxVFOpo52F0E
yVlEV09PAvStVTc06NTbHM7TKTzVStz1yuq2ECi/6MaBHXzDQ3XmzXAjmOKnntwS+OWOb+zP75Qq
hUutvnZUgqI5PO7UBT5w3ArO+8Y91UuoC9CAlP5LWj2boPWtjeYhIvVzwRSdcJtEfCUU+APajIRb
RToNOt9tWM0krgs1a7ZdB65SjvJ/XzLiXRj2b39NCCEZ6QlBMAJloydBXZkm5xkRMZTwHpHq7MFY
1rGP4q50iKtgnOMjcRBzKjk42ZGbBjsjdIa6STMoaCNitZ9GgHL4l9W/JC6mfieJnB+XZoCMUjEZ
oRrBJ4XQWTi/l5q1/sL3kT7s0QAE7+tPLL7pSCtX/IaTsegNER7ibq0COMLp0bpvoiSPSHZvroqK
cBKGupNUZXVJ6c+X+ojRo1owzgdmzwbO3UkebKr4X+O/k/F88s44KQGpQ/bTYnEZbRW/6eRVWa9V
aJPpTDu5w3BCrageEIWHWCKIhD+i/LO6FSrvPftHSjv/ohY2TrWn5Bas+A0bAex5UrJTyjvNjbRc
B5sHVRqepXGkixiqv2OLB46Kgg+wrXJlUGl0pQe/sVOV0bANd9sjvo4l3h+bbZn/8uCQzjnhLwD8
/BEe+8R46+KhnXaAbo5HHgjmxp80ZxT5RgH/DUC1P+SLZES8r64Tn+kzGsJKXteS9jtTGLPV/YnH
GHM51Da4nWqSWN9JLDBC309dbKlyHxr72QNEeOI8mSsOZ3K+OvDVUpxwzxhxTjH8zlXcmaWtuEbq
GFc/jhxEH44JBX5UaHFbvnpnpcTyjCPs8sr4DUZIgpoXsd7MRHCTvN0tOKBTtEd1lkDplU138q0L
fr6FKzf1Gg==
`protect end_protected
