`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KnygbMjgOQCqhfcawvvvOZM0kPu1gGKm6dHOIF+fHSKW6Sm6J8MhnFRV9XJQk5sK5HUeB8lTgYr/
k7iO5XNwiQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bbzT9dbI7wikdLxg+BPxGcBgnzk1MMaLfdCmi1ZHHQbblGZr9SHd+dLGX7V9yu44cjowlNmcV8eG
c93HjAr/CqG7I2IubdE40ZWEP1v7BjpzN9qqwl+FMiLo3sbuY/CUb20KIvxTbtHWNG30U+vbVzRR
Eb6rFeN2n5wrOUzoUxE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IFVfU8sDrh+QkRjdIGftK2te+VIMb4OVpyWSOlLsWXvk2BsKk9+ZLa0Dax2Y/AYrd3UWlsa7thye
dGZznyP/PHoWTDTd/iKDTLLXbB+yz4mS8KzFVJFThMkdHfmqqyRU7Ww/XDD8dycapCq7OmPsYU+Q
XPeC65aKR9GBgUNDZquWovk3judr1xU+pO75sH24qD0rz/ArCfvEo3oE0w9Sagx0PI25nQy8BkJ8
1ISp5w50Cm+BgalgBECv0EPYax5a1xy/2Z69lzPKjc2yMb9X7ruOfOcHzGHk71alYuEvZIYQjlT5
/+AnR5QVWoIKIqwScHtNK++4EE0Hc9Iv0B36bw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yaVAvYLOND+NGLsMj/M5+6ky0GlJCWlISRnVLqYx0nHFiLOrkULsQrxk0JIdxhjvRlbiHd7gn9Vs
FJWU4qQitGwBFV5mviEZK2xhw6fyTRDpdmNwG6VCMifTlm7GdGJepjbiaAMfDw0NvEwa99OTiMjS
2PyVQoMCxeN5wkRPB/U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U6P1oihChtDKa88DnN0P6Zx1Noyk8D3NRxcHXGbovk5qXBD6Eu1lYouLN0lOToZugJpYUbwLO+ZQ
wkdrFb/SjkPCwT9bahL6jiTcvd+JKk2skyBlzNi0vGWk/xMfIHI5QNUOJamEope2N/ob9AHyoROd
1qthhGG1YoouxRPxKon0WkawEzMo2zCKz+/VO/Taa4wOWTAzyfZZzsx5o9Ds4/9ebzdN7nN3hHAO
72v2APCORICIBdcXCiLqi+4eXFUEBhh1WQbcE5y71QdjRH4ygGK7sQQC0qYqEOuJAXW4dTMMCg0M
Cehkdh0Rpub+ChEcT0fO2Sa0z0K+olVVuFhYXQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25264)
`protect data_block
CeKQOQIjC9gUKifDiWoyukT/0RE0nwcgbCb7e/YWarAQg8WFg4pTS1h+wnYhelR+jr2f8tUCpbca
oajFoxKM5gOiQw9F1WhtBPcJpF5+PJOyn+DJS+r6DA+FNFDEDCBFYbQxmHeHwuhoQRMXNyu1E5s4
KMoX/mgAC7W3W1hkYECHCkvvVXufNj0LdoPFFDrluK0IbXzE7icZ46u6VkY92BErnWo2L11jSgs8
O56h/fd/CMiNuFnxpQuhycLH2cZ1b1/OckBUwx7z7GJUgJaff+Hj7mwM5eZZqTg4S0+UIFMdrBad
o0ryWA1RKL+RjaeJSbRL6n3AEgPlgPsxwN5ffwdMqVDl1g3+lbmdz3kLpK5vG7SaO4rIPeMphVUJ
AY86ITxWstZqniJcPqd1oCVjkVvgIosH1kh+JM3uaAtcTF1Q1kYMGm13lJR3lgVoXb2dv13eKdMZ
K4of0kp9WNUt5RobBnstFXD/3IUn4cUb35F/+XBtaBFMd42+F26NrxFFyrgHlhGN16JaJNGh8YvK
fmf/YBzIEbonH8cSl97mmxDR1mTP64KkYIQVAC4iqXuSCVYB3qa6KegQ+nEDhqzJqBDM7N05A6VL
MFM9vYqbYbwwWHNsPWzxUW1kNxpqhfQl5PjuYEkLzpuNTxbfb/8Jwa/tHPjNogE0F3KPoNUe/mji
i/dFEtFKM9VNeSndT/3KjFHBvfUl1FElhdwUInqn4Pj6mzyAvJNF6ON6YbRwlW5HuuCHgBgkrBy3
4TH49bFJd6l/a7XoRvTvDoU8Ts6hx0pnO0FPFcq1WmxmOZ1lNmuQ9XL1cqwcCKeEBJoNOpZC2nZ1
e7kkUBpcr5NLb+q4Z+9nA7SoHpSdwmtlNxHnxRfLf1YGEmMyT1mt+50fflCUeoI5VLSr99uf3sUS
mkDnbygZsbZtB8lzwhmncdAywAu+yGN4gm1FrMWSFccWSqFtRw9M7PzwNnPx8qH4x0SGF7XxqGsG
Bs0GjT3qd3O9BdADTVsHW6gLQeFLnIzlgH1H5BpiWlPIAZVvCbmhp9+bLfZfBN0HH6hnFHq2hpi5
tscuvvezcwBrKkhp9uLDCja+n6wQdzmSoTB3gHDGjIjZwy/GBz99HJ+DR53fzf1qQLRTH+skGb0u
+6GVV2j0apKb+hYmJfzmNnHn1IPk+68MCIpurAk2+r3cRhrPvbeGCLJOe/Y9ss6+7bV13wkRZitG
VvMNjaxOToTFCDmIEH3yLvR1ntfedh9Fe5p4frFHLkSYETpqae/XzXzJ+Ep+7QAFFY1y5/HiHMhf
Zr3V+aLM5AuaLzYBrtZ52shJFIRBJmxx11FjdJBfGHavGe2lH21Hj8WzwMIGeRjsqWhiI9c4//RC
VbrqIgpnJwzpffqS8z4WOhs4+HbAu/IGtCD6u+l17pF7F3AlHK58huJLxs9k7pzfRGJmp47ogOWd
ohf4Vsj8AYZVkshxNmpiVnpMogvRRcw4OCR+p9KPYdsR/zXI4I8S0s+uU7u3eOpj9KM+PsxD/O6i
TbrG+YV/YZBIhgRzz/n5Z5Wy59C7L3aOLK6GMDBRbEzbukqqq6cgroAxeGk1Ne+RHJGmnRct8C6S
CEyTOfpbmNLcSVkYCG5uOd6a31vPD1xzzRDlwxuQtlfNa+iZ2Lg5vTD4eL24wWn1qiDpOqupeb8A
GPQwYq7QlgS+yhYN1bx0tE19RXIdFN9r7q/JuH51zJ7H4XAxxu/D8SisTFX/kZbRGc3X1Em3CVfZ
AokETQW0QVvft9XM5fSor+4v18u+Cs6jRi+adxfkws6MD9Nr+KpzRUXHLI5VqDwPXyEs6foZz0EH
AB43hdOoNDYgA8aKzNjwqbtjwo0dH46TYfLYqb4kdK7DisSwF3Q9DNxPS4lmbvls4Uro+QJXjAX0
b+yGea6oUelqaKg/1vFt86WOEkbvypfFWM2kMk6n5o9S13rz3nai9TKUKSJIhzS60VOkVLmPAvod
joefHYc2dcz578q8VO5GlNbTIbbSYRCs3toMJ+3Pdjx4K3NxZt1F3HsEf2jtyaiuy+jwxItZU+R1
DDLLXbaVktcexrqiqFnOKINxCxWedXSjmnJHJfWzh+2PBV1kbDLLlyDhadYE58QO0eFmbd3fUlRR
pbpiTFrKZmie+8C0lcPmTcnIeCCnUc0JzKleFJ9hOX2Z0qU8FfCcFdG1kYIWKhvlZwM7oNkS1Khz
0Z3IIuHqIt9CnYjKUqNUOz3J8Saue1bIF5Uu0GnAh1UDj2U7ZRvg/nYz65vgYR6D/sCD2C1+VfaY
7Noy8IKz6GT0+NhzC5UzLI891UD5VpM1J2qBL+D6iqOzYfw8gD4t4xWwsu4BB7Mh6NBSXFyZQhLd
1+Mza0gD6W6dgTwEU4kBzaIkd+q5lU0kKzwPlsrBKxkM4spuf0ceYagxfHSyO2OifNxT4tKzseco
QJLLl8Xm6rYA0TMrnVzriFr6g5AOiFgXkEGbqKehnf5ulFP3uadOQOdmt4k0ugfScalD/+tO8WHa
AxgLTqoTjFyhj/TvZRx8VG1Sf+v24rRLP3omSOvX2089JxUn/E0d67iI3ETuJeDaBeQtndFYbOUk
l8hxjnqqnIsnINerOSdIr4ElGiW+mBBT4nIo/K23Zv2wqTU6sSQ9+UnPdGb4DpfY3edZszthEFCM
Xe8iNeAi1ztJNV/apubCyL9ewkQjHXdspuoOp/0chN5Z0ikILyN+e8AHHxdHulCefWl6KPRvuam/
OvMwB5F5ZB+/HAZFqhElk3Lf6qHYJwRoErH+pd4+NolmsU6ksxGeflKibLJMXGM7sL7GbtuUKXY9
b7d5ZYxLK3wGNuhJWltAA6iQ93GlZYoADzMchlLZe5woGHWLiuLgG0PQ8fQNfMLgtKQFGLuVxmV+
JbyZdWrlfSRfOlpl5/e+JlB155uGkeVBt8T/z/Lc8So9ea5zEkJS+L9Q690yRos5JRBHDxjzdu3e
sJlGHLBHQP68NgqKr7nIdvhdNk0EH1yUaxayjke9hZjhNztXHJrr3uG0U/axSmC3keJu9zoRsxEx
5dFjjr1nACkSZyHO9L1s20FOtKzTHWnOlJ3BHgWvhIJCxBxgxj6mA5aIjwjQaP8pr0gXPGiD0pan
HYTPKz61cXswdvVqran9mxrR6jzzzP45lf5p3BozDPO4Som0oaNPta83tUN4xN2W+BboHPSsBJ1n
5yoK+Rffr8e8PKHL9LvGv/HAhgBXpgvNIkfhO8/l7ldyrOamusSLJerFDQchn/mKMDF9y6Wd5Eka
H0ypLMAKAeAHatKYOy/iYshJtrdT1OoOaYuKs+psByXJb+4jReKdVp/dgxHr5xIZl350cgoDcsC9
3kSEiay16Zb49bSDhaT01CqGCmTMjYCT8Nh8Dvo5opUq5l8kr2Z/2skFpP5Bg6hVTJyQaRtDOoMf
Wys9KT5HXXRKr42a9IXUe75azHhHgTBagx5YWv9aKrjGJ9cBFXypnhtz50S58HyXv7zLwbtmjjpK
3KdSYK+CI6vPEwFk9SYJSvK0lxkDYDUjfHQbm2ujZp6+4JH7hlN2V4h+4yDxzwyl/c+Bm3mOp7fK
fTu8fJvHR9LW/DcXLOk4OWmvpXL+xkYJitwewVnQEJW268LAb62Py6ycWJnvPhxRolm/+5r0shPF
8ahcPPss/IxlFQzqioTDTv/GH2VAHVT3QJP5JzBPRxxzGbdOaJXit+RJCo6VRH4426QzF0xfpJiQ
feiVdfq8JUIpb7dnP1j46+7rkDdV5aMeaKQ2th4cOUjCOAU3LsudbWiBgJpsVYqlwomrVRJW10vP
+O1DTdU4qKUN070oP+E+15ALPSGN1BzpXmZ3PfmrM3buP9lndKO62WkgwuUMlZixBAnQcfC8bYit
7SL0bb6qtzT+PM15o8bEWmw4v06z6ZfB86TP9zF7KcULFhcRI5pFLKHylYYp2h9oaNoaTPogDdti
H2VLrZirlTMpadg6ApJmWJU1bN3nvuQti/tS7hYTZ/GXvLOQSFnN7frfKmnGfoWuhi2pQy3cIZ8e
GRem88XoN2RgV+nIkg41ycd58VAa0JX9ApssH41PRdX8i4SRDi/06iANRO7/+SC1V4ND7tw8c4xS
sqF+HGtu6JNVFsLQeAtN6LXLiWa1dXUKpowRkc9Z7WFMaaxQsksFM5HJ6MUspYxA7zy/XKtVxCCh
kYh5nMPfY9DuNQpbYr7ylRI20ce9zd9FZ1Gchp8h2AmG/mGkmHM2k5y2VOkFjSBSLmFuQjMnruhz
uayxj5kZpGGCyMaVtzcACb3affWEvaFEXXK98JIG9QHJdavqgJuOFvyvVRN1BajCBzwUc7pD3Jeu
gHNZzNPlSQlp3jhKUZ44HLj5sK/4sdx7fjk4R19ZsNyhP9AULR0JFVJCQUpq5Nfk+Pi+yJJ6W9of
9wXIaC4HuRNuOtftJkYYj+a1pDTRiJOstpnyzityBR/2lbH3NV1Hek/Bx2NSpqSumIFbmjWiLnFQ
8H5J+23onoWSqxoIieWgwds+h6AZKPyciEiafGCEUlrAU2AzghwRkEek5g6BoVpFt82Rc/9HFr59
s1sos0d/M10X8iDfdA8EElz5FxkRyjtUAt/brYbdUSZtlkWzilnj/M4xaIpN6Xh9GAitsB7Ap95j
bahkTFpNORBuD0Kk+LUH1r/Ok5CWlRp/lQ/ntHe2s/XDOxA4FhGMuKJLy5KRV+15eA+5B450TOar
c/JIjPM21cZGmAs+dYA5yZ2D1VlU8hBfjuj/MHgzXMHyVJpkoT564VnSMLClh93QRLvR9V7YHmGK
Jpz0PZtPN6JmCw2dSolmFfk99/qHLX1Sxsg98fQjJX0lQwlKokbrKrDVzQ9bFlBr+HeWnDBOKAg3
FSCgTz30Iqd1VqX3if7dSB17YqpGwckgACBmz+ifiFMSZxLBIPDfqu8LLKCduqTQF6qLnLlWxvnJ
Uv046nJxSnHdRzx0MUzzoCR2COYr5M+AfcoRUyaPwFTwyn5ZjEjhn7O5BXPXqXJ9Zqx0xgs8qSkB
XYighHmc85gVDWYxnqS2vcOnFWSz7EfuIrxieSO4VN5CG4C7son12TKPXYAEe2ASP/zle9UM1T+8
OTl+oZqWMLYDMCfrhIuNd/DaBlEK36Ddt+8Agf+vvhZqoDSal3otoGIeM+818yJxMyP10yojcpGJ
mZlt5uSJL6N4IhhckXwbS9u4rVi6KxNM6wT1KJZXxKtzW90bYlYdgJzcJY0ZqgjP5AA9lXhdqShd
ZrUpXkOGo1+M16fLikaWmhDWA3trCQLQgzw8D4Cvlq78nxTuAc+kNI9O/lOVVMrfZ7yi5blA+5Ci
3IAxjxAHWfm/uw0wzUYyYzsBKyY1PJBWj8WSZJMJXZhRMkluGxSjKgZGi9Bn4bd24wj0Fe4eMEVO
OzseIvQkMhzi4FMf/CZ2Nz4lvt6r9cJGMEXmEaa1/xx/nqE7Tb0E2mwa2ArOSkVdYZQGzSSnPfsr
91oRPVpb5LSB5B0i/jh8Fdb6qOVu8mKkdGuPQ6JAnDcmbTDS2+CltyRsh61fdi55Vi1b1vSmIwYY
hzQlcNEKPhUxRYalcyEAqtkSvV3h2fKhXOaLRcVDH2l6PIIiaElDj1lZc15hIv5WFcfFyLb/U5Mz
xUD0jyyhb5xB8/9xpUZGMHELeC2rgra0L54vnX9f1YbU5EoM/nk6R3zb8L7EzHvamKZqKd0+uibc
c6/+mKT907sr+XN2Wy+bzY8+1m4u7ftQgs8RAt4Bd9LJUCLIgMnrRMbcXwn19K/DrbyPOtaYKPrN
4PfanwcqEu/KKhMHQ0jAlHkcdEDZo/V3Sbl6pXvIhVNXZeFWtkEGjabtHxdyQs+toRECeFX01/JI
Hg8nDiWNtSuSGB4dh5lMY4Gngm0IX1aQuBh+tgONa8HraeYv4NubEn4/GN2RSg+97D4ztZW0yOoM
ZidRgPOKsmbS2a5epDmlUyTLrb5KeScE9Xa+aRl4QUp8YUpYKxHqOLYBOaM+38g/X10QQ+PpkRX1
1XYLZ22OkNBINnRnTgde0EZ0VhgDTA0pKeQ250YW6itIgCrXDDrH58LvUhl1nB1U9CBwoC+TCL/b
OXKSJb7TkX3bhyO2W1GMl5qh9eyLhVXb5h2FpwKvgJQaKWGbNbPTm/lPbBBs2GNDQ56+2NfpEn0N
Fwnhq/ohoenrR7YG8Oph8Oz66GVjibsK4/GNx9phd31LJJX7+gI2RnYsiWFB+uJrI/Qxe/q/fhhF
2Rr03+HLRdnjfLtq9F1+//kDQ/hOQQ8Yjh4rXq9QlCM4j6lU0EGjhF27ClQOkmJkzsen3xeHcifw
a4Ol86ChAbIgum9P5+fOE2LZN3SZXB2kYygZ77A0dNhFXhxOEuz6hDKkmPac0eB/tWTMnYJQ4qZc
zn6y4Q5BOiBblhP3tURN8vsxdW7C+pzzsjQi/vOYPuT/Jgwat2WK455W7r3FACCCm+uL0UMRMuFU
aPP/t51AH3WulgqEjuj532PywxOH5MVyIhW8N4Iv9PZKIMUP15O/sLLmRxRd3+J2pcr9pTTGc4PD
5C+4tkt+AJOdySwnaA+6k6diZLC7WZ3BCCfWizSfBmuII1Gm5ku4SeV6aWWv/H4dCMYg+awxFme9
OasN+XoigeSdbpy9Mb6PNcSDALIdDF0KFRvNp8EsPNb0VazhHdffJnVsUyw+VV25kRUrxeE7OC7S
YjiFyRH4FHU6OuUS8bDJYRxuGUDcj1uyVNf4k5w5J4RoyI1aSY78EqOZ0ItK+UND7Uwltm0PkLgR
wg+IqzqN8dXfyQz/WG03OQjDsOrDB3My0GXp2zPblJAL/eRj8OzhQ6Pp22CZnYdMWYfIMFaL/AIL
6T6p0xj77MTooRgeXPUmIWeE1RWKjAe8VrGV+qtx2rd1hSb3j+g4GSHC3+HY+RCMQUzN3HO59uA8
SXIXn9sZCT2fuciCdrpWjEr4HZLBP2T3OWwmt8v5r0bqDtffojGrqviMcBOl2omHnyWLHVpogcts
oS3rVUk+SNA3TX6eJ+NCtI5sJclLkgyjC573T0MA6yhlWbR+NB/feiK4/xgES8DwIMyWsusxz4Kq
hkdyTwabdjvVmRYgeXiILh32ZJd07BZ90NFV9L3hfmNRWFBlPqPe8avDl6KW/I8EiL7WRnBf1DM1
BZ5ETIDA4IX3Y2z1Qm5cwN8oQlMFt2u1Rl/VXgIyy/JJVdGUtuCc3mYJm58ZGkHdRf8xb1z6PO7l
gAkAI/wSb7icSfW3U/i3mWHPlj8UuUBNe6BSmnzuIqg/R80RoBCiVdoEOl70ETayqcyXscjFwHEh
+nR5Y7l/KL7ZLdGDVI2cLCvrjrwO+sz+h5GzcIWbuvAnje/Y7IJNm/6X1MhaAJSDer3EUe1q7Nj0
Wasw6btjT48WJc2QRnVZ4usJfkTVQ4wzB5tdMAJ6tqbjH7ZxnRrLHaSDU1Kpw55Fo5MUaNJTTqdq
kaiU6m6tycQQOYfYtbfux/HdsaaYiIopxgoNMPqMgL2PB9n2xMYeSzdY1G0kS9/VJhhFETI3A3M2
Jbj1ZcWWwF6cfT8EzUUelQLkvp3EQftJKi349Lp5cCMMwNGMorTfihcSYM9mTIMgSRtQUJbxBT44
iheXKCNuaVOOK4v0Vh3DZ+A5r2w1aahumavsOYvvkmgr8YRO7bI1ue0tv6fPRNSWA9BO2QQDTypQ
4cgnTy82+/FFXW2plr9z0u2R31V5La8eS3VRU12b/UibFQFHnvLC01eXyzq7dLKrpLb8JHhROOyB
lV9MTbSTM5nFZBIRtiiipoU1bS5MNnDdaFmAuSX+Az14SE/bW6GEB+S6v7DZ15y08gsQv2ZFS/gg
ToLDSLwHSg/Gr8ILNTRT3EW4rRgmtCnoT5HU/3r7LkE8s7Sj8/Cgi+n7JYVf4VZRlzCvesHb2nDg
PTJg3+PddMV1RuMI6gkTEV0SDzUpFFTkV28+8Wm6cvvI37dlIIsSMfvI6EuUrRDXgHyxqAjyJdJ7
gtTJgTMmO5b+5xhabdqpkOkSoNwHqXNSvQD2H68xVv+pAH1k9YCswzu9JDeIuiDjDznRrwveSw8q
q8wxmyLY77phlF4PAf3i83T533hX4zOUk0dTnpisW3gu1xsaNcmYOS+2vPJSmpXo8Vcz8ZT8dRyO
pUnwQItdGr+cddYeQIPjenKCRzRpFAOIDrwu9wMnS36asZT0cw6P9Yo6F9t7KQjZw2TQ92OEfzOw
bv2vQY0DMKty+4URNhXK1DS7xziam/9lUe1Lmz5hFrpzzBgOh1zG6wuAgZ7dbhcp5CRNP19Nzj6s
pIkqBUXpfMvM054BErgzcYtfF/KQIvLH3Z+IhEo3d3kDGcfisYbH91Xi0VYMQnFHYr7jCmY0rQTq
GUGtVbnLidkccPBeHz9MeCqD7lMLFURHclDFvFysqa3fEW5tcu794mvORN3hxxd7gk1sB1D1h4lc
P/aFlNScotdqSbEv84yfTJh3eOxYp+JlCxG5NsuPhM3f2q6fiqGte3D9ZSi0k/PZrvdpqrUVnEB8
H8PLjZbxXSraCXUNsjwzs7HEAK6gc2sLWU8a+jwi3yhPuwVciH7UCjp2z1ZUOiYCD5/e8S2cTWyA
gxUc3JJ4iPbfsscrUMC2mP1Hdg13psHkMeTe8GHTOq4wOVmq63y4IhK8LzhsVDocjbwAMwPVr51X
cEunxeu+aC18gI8bU1NdK33ziy4DCko+qDn7TXk8/OU56AJgF5AhyHlk1xL6KyFLUszePBalHwDO
QLyLoYp8fOyQaASHv7CauudnZutl2lZSuMNi1DStkmK05JC2lEs7gTV0snEsjqWHCjNxzo5rSGjG
Mn+b/eKvNFIBiEnE8gJ22rM6HzkCnZyFGVt5I/swH29dnbcdh4OE96UJGUSFIC3USyNlN1d+4mgs
rHrqNJGsFzL5HiaJ/oIWXYfHAnsym/enoTeLkefZhPs2r80WiDwmzSBInysReYjD5/lPThVrmG8E
3Bo+soyEWz7JMPLSoMBwvp1JtF+3pI+RFBmcCxTT1JYCiEd0QXqPvNAF7fT+NP1HL3+HqtHj9Pyv
ZEFe8JeJ/ZAvcwWNtDViYQhFD6aF6Wb3ck8L8iPxUdEtSqNciOHX8cskZo1tGYdeqK3g914w0Rfy
u2asCufzbHoGK3IEPk/B5OjRFDsEwpx5eSQqlfTFA7ySFl8y/48WhYmGwWihBzIJgj0DwqHyTdWH
g7HO3YHXGtlnB+KmpCHQGotnqIMB9Q62EfsGCuo15gdCFFSqNOtsShOp4tkoBxTtmtaoDe9K8yac
0U3IArzeQobRj9a8AYfVHIZU1k8OG0h5ZK90+cPsTZsl3pwieu4b0Wq2hiO0ZLsY0eIEiR6BH5FB
UMyYOR5MG2nO+s3OlJpep3V8rfBqCjGlYv9LNI70mAiBi1gXfId1e4ieGM4vXbfl8D/o3JW5RNmo
NCnnJ4zhd5HvqLI5XFdnuAWsOEAb3LuXMoGDF/kBCZPPS4HpKi0S22uExioaHmazVMcaWzYWVLbu
gxNVo2Q6o144aKHw1kakXYoYG63EqRAY8DfgCcrtfhghWAFC9BXDKDEinNrZbLqym4z69PWDH3JU
0mbN7ccc/nPugCr/NSY+HAUIoXIbGwBZdAbtNngPcq5DwxvUXCGAhM+3Kf7agFvBDSrirk77Jbh2
6UIKB4Ofor+L8ZKlTq042buPCO8HM099knByb5SJINgqJFuf9aYSkqr91mqQpdMlX9GGxgR7SdGA
9UEwEztF5PHhM7rhPogaIlm34+6O14R8gHe3PNGZoLvSrwA58xmWhn3/fvr/Cpnu8+4Q1heEnS7Z
O9IegDcHmvpyHHQt04XzEdIOOfY8BYocLzFkII3di9Jl2dyBwFXaz4EIdzgibhFqCplDyq+hI/z4
IQCvgggy7zPKzuVmrgBDKWsxJ2CKUKyUcYeqoSmOWMSuV69E43N2AZHIwcITdr0sa6olLJjqyc5M
BYDi6gCUndPKaAi02XZec9jPd8HMfULick5nnkYDmz5ckRJgI6Z/FHjx5EL3p9YfS9F11bU3T0Vm
NBmPZXXxYpzzBQYG1k/IsvNOiinrjwChm1UJPFtagk/fDZ0xhqAkPLxOeoopI+ZOJ8bz5pntBXpO
Z6TzwoC/duYOCNbyLob4FNgqgFS5K0As9goe67QrsQFEByso93J5iJfWzCr4EO6PuLOHLrG9WO2I
thHMRGz2cOZGnKNZVUyCVk+LWaO9s1oryug7NUVNcXs3BaLVc1Z4J4NWzNzncrPRxZ4ASCwKk3Rq
M+LXLgPRi6NS/H+d5t5rYQq3tlzXKfC+/Sc1hyeqms6K+JEPWjR8jV2VMl/4ycq/4a8g0oxds1MF
KYDENqwVXCluYgb6su+DcoMLTW/5hm7tZ7rgVZzlg48/0shoHUxE74vxSx/Ms34Hj5x4V8NciYtu
EuWyawiNGz2fYUaG9MHgIGWaC21mwOskRoHjlaRW0YhpK8eyiF3guoNsDmkcz/BwxIlb/rZsQLY7
T47madRzJrSYBsYTZhZcVOrbVdVb3I/PMGvFT1xgqCQSM3S0bPSRHYkzEQyxyXqLPEsWtOYAvf84
d9bcsUcvCaarEDDJ4PcQkTXoC9tQ50dqQGghmpRrIjKpunW4hAFTRwMkHAjXcFgG6Yegtbo0g4p3
QmSlkLpiK2OTMwpTxdBfDF9syMeXV/UpL1cN11QjQ9zU+FEpQt1YJ8tIa+S3pLzdOPpwTrUkUbUq
8Ixj71mIEPcUNIvJ5ww3m9a6NGXqvlMLwMwGIBqO4ddMDP4ozCRyWw/es+2e/irUttnEK4Q63HpF
ElQt0xpf6NwAFNFqUPdcHNSHJeCH0KWIMGC5dPZCFQYtbNjYvSkJuVN+r84OVwxXa8ct62YcAQzS
CmMVgPQipdZlUrxX35SSdbhSqL9TJF/+9lRuyv/RFPle0rs2g6XYsvXT8Ho4HufL+GydgB5ggAEC
eDzPq+wPhAGLtdL4iho6uSaXOPK0sMmPlCxym1Cuqo9sQsrKysOCq2ymullcSu6szs0/MRyYF9Mf
5LkUh0QkthnjJsbT12xQefYWwjYvjCjhm9fahQB5ig8QtDc6OA9oBFjSzbPlydZA9A4uvMrb+/sR
fMXzEfWbeTlGTL+wjwvSILm6Gd56qr7oFiKCAr4VMRY99iEwDSPg011k4NWZewMf9YS5gSF7fdfP
bWKkpdceY5UrbTT05HiF5ZCxQcZrXZo6GBVRbS+5oyz91ST6jH6yjbtBsUEUDGlrBhOV5NGuTvQI
PGEX4VP/YP6V7TKEzxmHttACklpTzRkrHhInBLVdilR9fXnkNHEp3sMwsiViMir3DYf92ktejval
FINCSfe6p8AaVz3leSgrl6nxa5uJKe5HQK565aoyamtIMf6iFrFsHCgdvyh2wd3ktWEw2SAEx90G
IJI7dnoVrgxzW1OgiVFc8mFek3DXdK523l+kmo2gl9UGQQRoLH1mW69TX9Pn2/GrL0z47126/JWt
xooUTJc8l1wpg/44fqhdAxKDED1PjVxOATgQ0a2w860ryhcl9P0xGerX9LaeZ8wcm5o1aoP9WBO2
hU6CY5zaqsTF+L82pnNaE3AbXECkK5UHWTE6nvB30whgMW/k09NHNfWFafU6VKESuUVFm1TvHott
a1V4WanvFVvWVN3Wi/dJ5dN6BtRrt+tiBhucATiDtXp/t10t6pTODaSCTg8KjUmy1caaL6EePgPN
wQTLhaSVh/xgKIu1KQ2DRftFGkzN0+bR9Axoaj7mhFI5uOFLaZXThZGF9jm31PRbk1Q0ARHYnXxZ
982apwu1/AcjQxjOV8qhPjibhvT1ZdvxkxcF1Vr8aCjcr8WjxjIUH+m8ycqRn0UWpyNfUkrATByU
0NEMxDHvPMLKYcaVQqXzHGGFXLnPY2yfvvbchGXB1A0HS7de1aTQE/cmgb42NKsamnFfzdtC6u2T
DDRB22Bvq5eefOIbrQMPlxPr8CfOY6Df2cZlavqXyAj6kh9uGvJvIi2+NSywK1R6o6VH8X4uIjow
LZJJ5Fa05sJQ4U10LEQb9BaA5elqvjGObMnjzXWPfOT5iHc6q2nxjDZnrAqzGyrIJGvA2yfL1/tv
Vsd1LHgY3tDo5O6rcwBC+H7udSPGWCjr3OXcCG1yk2V8XtxysS4wpyvChJcE3DU9XIs6dg+L8kwb
Xge8/XwlHz4999MVierOFLy5v0JeWUb2BBPXOo+694V3mC11eG7LZmQBWxyvsMH+io2jZr7tbmXv
B4X38KQwxribbFe0x/tz+JLsaRZvI8w9nOHvqqXLPGFPqd9E9K+wtF3Nwn0ddC7eFb/c/9iQvsUW
9bZXBMb6b974wb27sMO8FTYk7+kNj4O23JUaBhzgGeeOG8qi4MvN6nEvfKs5rRSeShYqkXpirqIm
pSCaSj+CBNSwMd1SKeLP5EUu04Lxoq8LVCLvb7f0HMqClG/vMxDyRVTcv2jBWAPFAgsNAzJQj2iJ
N8uJK403VkfhVKWskYJp6kOU04TtRz5QP+xOIwkUH/J5dAp8rAXNdW16AKFgPG/1POZVXmr4GZPM
fKb2AZ/1PeK3KTGDxP94Oj+hijxHIzG+IatahsXmVFgJriDcA2CYlH3bP+PHgZ4qHdyroB6nOu7k
S0MDvwplhFyiXnKTUTKWmNNhm/BoW4qLVVYv+7aRj5o8XY2s16nMYXJCfHVRUzNHJ6IkkADDhG/l
mV8frELIKJgizW2bFoPz45Kdv5A1E5z+FhCnOMy9kOPowi1mFKgJ9gMRPpotDlIvWWbeEIzChvAj
pHdDF+A0upCWnJDmYgDI6btkexwz/TyHwhTMvXuAGxiegYte+pFsUpHIodt3pIB1x0q8zzfB7rTN
P35AsmnSVHBAo0N7IsD39/kzdJmtQv4h0zj9rH3VCsmcfJoZMRPOqcRauidOWx0Mp4mzMNl9HmEN
Lg9yTanrvxnCNJ9qi19nLboGY+NTtqWkEN893q04RigEiNz9n5orF++mNVL+n52yASF5BNB9Clxa
jN8cjl8nXPbdzXp+wbY3fe9v3xZQ69FN7i8GQk/CfUETWkMqlwpiCPr8PGYpQ5KYiTmV4sA40Yhs
Lf4iLhnOvyQW+VK5Eyy4HlLfpbhgONbtB6fdGW6ZQAe5n9sQ+3U1HtFIkPEFA6jzDnGkx0kEDpX0
pSvaTWCWtX46XdQRhfv21L8Ag/15u5YlgCGgQAIiDH79F/Te/jRodS7adg9zJJ3Ifmb+dXrIgU+S
ggNtHNGDvDuObZPdJaFzX2gxWbrYgrXmC9ilj/lMF+i2zV8InH75Zqw2QPjLDn2QUxfbbJlFzu8u
pFSyadRTXDDy/Mx00lodG+Lgx+gZlUD7tC5B89mpUwr9feoQWHQN/UTAaxOjm9lCmx496+XLVgJm
MlUKKpv0jvZcTYqdPOPwAX9I5t3PdS6sk/Qck4RxWw7dz3Bom5qfw7CShDf4stYbPKLePAKnK76+
wQV5qHhjTXeDxXp/PvvE4vbpPRNDMbTmCJ4ef+FsbYXSqoH6F1LZa/234+FYH02O3lECx2xgtLta
lL35YMmeCdtJm4Op5mx9DPqECY/T/SjeYsduJ+/oEGQLMcn/kcYEFZASpRcmbsc4B1PJQq9ZBVSZ
6Blkhgxi1VKNaNLpuEO2NMmwy4t3G6aAGC+RUxprJx8hWjzVcFrH87X0/cpWa6UEKe9mfZSrxBOQ
JWPEpe2r5139jgmG7qf+3I/8RfX/GL0R7YBsh65N3WSyREJLjYOKmc6Gr3csy8kiGdTXMEVeqQ0+
2+uZQzS90uqq7a5qCEnIIau8Mo0uZViuz0/4glWGI/yQtvtY8ZwY8+xvGERpD7p9CuSv5ieFmGX3
F/zBtHoR6OvyideTPW/WpriNEuuxfD/0SnnBO2mr29XZUbXMXaCOPxo282x7DtSe72bt20Tb0aJ+
bhpbhpUNZQov1UkSvS6v0l6URQCdJPa5AhUymaBsA6bt6cKAErASJK/W7XbAexybA8v5yBrKbMtk
Gzp75YjD34Oh96UgU7SSCbQix7lPwyS6Frm40Qj3AGE8ITBTOo+8SR9WfF18bZhinvWTKikMfZFq
4QHuGKTTHZehXjpKb5f2duqILTCnMyr+V8g8Xxob1zuVZTfZCplQbmQgJ8OeysEnnI1bmk6sp/HA
6PO5G8RyTp1k8BAN/mSDlGgc0oZV9jM1RuZR9wzSFrhDe1r8Dv/urkXM09VuB4OuhC9jtclOfgky
SRCY0urDMLHHroUV8Yy+BCcBmiWFfNVvQAwAl6PgRv7yhUD//R4xxm/mTF60tWxhL4GwTgD3cS+6
01TDJtTSDcR3kPsXrXIyGOeMf+cL6+WYsduZK64Gpk1VzSJUkQHItlT97pstZsSYrBPevQWny3Xa
taJSE8R0B/uHGT3rlYgWY6ROI99Gp+hwMt+U7kizdDseRwGoYOJ1WK0skYGhDJm0m/dD0s/PP8jJ
WJ9EQ4YwHr2qulgJb2GovUs/6a5W4LMphPGxZdc83hYPilnZxunlQL1FgKAIQ5Uljco0QRJzS3R8
m3wQo/mWLAZoZUUPPNatX9alwf5akumXjzQ12qGcpusuk/1UW2wY+gcNE+SecA1Cdq4pbiAckJLI
sdL2WcQ16H22eRFyY8udJ2cD4rHTPmZ/G36KFJD6T+Dv0gTmZnPu1WWdsl/TN++yIoS1hRQG/XXR
/xHjmMdszl+MMgqlwo36Njr/+mHn94yvafZKK74S9La65heBgnYb382Yum4hDudFuXdJHTYjwir0
6jquNBBN46f0Bh+h9TfRrRCafPKDE9Eg6lkBCatFnaTBiDDQZTb4IANzPC4uLEHtzlKCTXJcWPwQ
LrhAOE+btxiSCP48kLDm2EaVzjmWc+t0qZhJmueNT8iixE9Ck2QufCkKgJUDfg5q5XJzW8qhLZhh
LDBzzA1OCh1PgVdx6sCrO4lcEDBjzrXZn5w7wYjtTTFBfQ/9ovNp66Boa6towVqBncmElwvtMUXC
Z7b8QVn6y90BI9Q+lbs+jd/aJ3KCG7qFcwlGtu2An68r8vuHosjUFN5OVvmVP1xiOOcgFKJ000J4
CyVoJltba1NdRWCGSzWpxhY/7HQiKkY/Ir+0+KPxgHUvOcg7qNP5Ym2mrG4kdUwMgNgDSK6U4QfK
2e5QbE2EXZZjKzPXE0BK7jIX8vW8SsNvGsBSpy/G66Z9acI6tptrpmkKS0ltQh6zv7GrKHnQMhOk
GbIahiDKOYh/slf9+R9pJ6E42/F2/O7ahSbMIMbaO5C+jcm5cAsifQ1nhmosynBhp5sgcq4ztBoF
vD+djIuzC3QIPp3IRiDQs4h1mh7YaQZ3scrtgGg8i1WiIBWXfbmMR9BoXlvUZEruMB7qxO25ixgU
VCy5pcYgB1MztSFsAyBsgZjEVho3tS1/sNmnOb84ZAjxlsvpBvMpCaxTOWkvtC112ZdwoxNFqjWR
+g7Wt6faHEExm2smI+oWdrPShwoCRjVtP4K+NrZPABlSTmz12oiOg+iWatwUTS9EGOIepIhDopw6
Ef3vMHC54EmjkFAlEC3UctAMudGgyqRinhOPooLNOJhg477+YB1Eem/BVs/Qmm5+WeT+o4+jVxOi
VeUJz8arIWfy3m9KIo3gzBu7MRcJsmnB+px01u2poHWcJci9kEFFK/gqrwktbuiYK9HRg948jWNy
u+vjz5XcsbR5f96EipxXO9DWTrExN5SP8qZn7za/HtZJZf+vOOo3z0OIY4haRhCDNYFkhfd773qp
FcfMtXwMlJPaLzi7DdVTuf68mEafJheyrBgsfCZNkMBxfcTnXucXFqaigR9nz7fxDTC6NO41bIbQ
549UedaiM5UTKvjPbDIYp3w8rxc8zTTzur4N2r5fg69eapeGTQ9A05JYa7qpaP7Jh5r1yoaJ/7fg
oPtp0KcFdq6+iiKf5xDO225JYbhG7f5U/V8UGgm/koZ4BiohZcqJVCwXDcXAYmvU1p0BEiyhn1Xr
IPlu3oos/OPA+MNvIzQajuzqa2QA17y9A3cvEIXUALhD+PJXz7ebU23MtokjNkvXz6CdtAgBImQH
+LwsWpr/ZODlSKA7UCncVaZy4JD3LHMeBkheHMDas1BIAOHSOJwu9dIxC8uPcuGy0QnI6Ec8Wk98
suchuLn+0ljRwoE8xYMSuzNgZkX2ZLKcNy6R03fjzSGOGReA8+vQgCYbR6QWJr0lm3ighADUJyg3
4DYLSo/roKW1PN6GNAwhwZHA7qspFv4aTjC2UiaLHsUsveWWYFDOK+cl2UvJVUI3SbcnljJHo0Ul
zhC46Ud8B1X51xRafjXmjKSsU7watOYz2Bcq29o1uRVaXNNB1oHrsMwy3W/bVXUhaj7jHVf1gc6g
yMUcG9/3AH7vEa9HII8Ym7xDInqu4T7WtmNqHOibGrYl7IlsvsnIMLwPlsjuPMnJQsV7nOj75NAl
8fbCy2RNo3VIrPAQBVedb+AhSNVduwrdU0FHEAI09rDs38FHhPwYxdjRJNnzMPOINJAjYfY1c7h+
vUwa34RJn/ZTChqlEj+fVYFRZs98leptWF8vgHHAKI+Zka8mS6SoyX5gTxXdaZWPEbWp6dBpJDFe
GhlGJFBAh7SdCnQu/O2MQfGG3jBOf6OoDYI2KXUisTEilcHgWRD0B+nMV6FWq4SVRMR3sK0Q8KE4
oZZWfMq+bW5xJrOiAzramYqw1N/iaGmZvVvVFnqND0kS9F7UeVyo3AkYQkN1IXM4j0G34Co+XsNB
pQl8xybYR1xqONB8vZpXp9CVFVklkSW8grd3ldsrN7jVcSPgvGOHvggBXWMKEWbrUDIPdpi2IIDV
SlqR/tGWK7P7T/iZwnVrw1W53i4isikY66BkJ+VmShk6zmaUSUdCdOTBLaF8qTG+U0FdyJdojIDH
1nRjGKkiJ0CIey81T8vBYTmFXSnWHd1fAUoq5a9Vh0opqRQUg6daSR9u/ncZfbHqhJdKijgdMDNF
5Gw0MYkIyy3gzQbQYLNKCG0RU6q3HiIjM82uqR1fa0H4+sgAdrWZQxmsBQN5X3lB1tvaO6KFG71U
OA1cBE5uWwpvOWKtNwqLrc6gngB4W1JSsDSh+0yiudJZCeRFTV2nBg59yWaMoKV3itmLri/+gT3p
LkAkNfmDxHC20Q7tYYu3WhLLn9sU+bAoSHTU+lXjtAu/Udb3YYu5rRMVR8eHtsgMcMdS+YrHqczR
mqLIGo+jL+dK7dQ5vcf8IdNio0ajnDoQBFIQB29BYNXdhOc86N7jGAM1zsgUjVkXEpuZh+rlHSgp
Pq4Mc3XNJHA8xNez3kqYeNXxnbLMDl7ldqAHEyvTp0vJYQ/rdbQSCVPHSZTLd7ZhbfoSEDVrvdy+
e1lyVUffEOz5Gd2mSSHsrS9GkvHb2BBLIl6yZtG2usa0UV7eVNiZiFfX8mWcPHn7BFkB6O7A+HQJ
oaIuJSZugML9PCSzo7Ug8SuEql0no/UNFopfJJeLw4LAzcj/S3gbx0wabAfPbNnN9poHph5S/RXv
0esa7axCDXb+732DkUStizAkNTC9gfFBHVg5zK4cIP92jrjiG7XHggELn61gay2ld0sL8JMcAIfH
eSTxF4wq4vkqyVOmjwtVqJi24VQCiHQoQM/xVABHrJWG5ZsQYP+gJrj6hxR0kwktUICeUaJotIVK
oxmC12uz/FpDTRrSveRP1i4pd2NUfJs65YAUx5Gwx+gqEEErWz2UO94GYDUrXgzfINvsWd1Gh9sf
a7xi2U+H25DnYVkv5V77/TvvW9JPrf6T1Y0RAQGjRFkWjIM4eO0uhKe+11O/ssDDGh6Y1fcRTQ0Y
LCkixvaEao5qgjofLduWwFm8IvOMi6KSBrid8tT34gKeBVxx7bqSb5rCSBhH3BrmbxfIn2ZE//Mw
DqkFJe6G3K9zNZapZ8Lg9YjxdQLHpEnuMQbh5sNuRZmcZbUKDv7XhxHeRMGRQePHrC1r5QmCgIxp
zZXOAjE0CgyM6K0SHCWsvOOTIqDD28sCUjl26R4RzmWg+BLyVf5xPntnSfxJqCVmTrPFqlRyNHRR
UlGhh8Rj/XwRconBGzbVLP5ddMmJdmbdIUqbrDtUUXwY46M3mN5Kl5VPyfGNf22VY5J6cixLW8xZ
HKwy4wJyxJd5Mk/dcO+8uSZQ7Ndqt6HGwTAatIYGrpRfolpryc8wev6FyfCcfvYPEWiCG7pr2SfF
MWpJzfDCYVVjbxnXpoK5kyiyZowg0TRhjkGyhC1yOODAhRVqlgzdUgbWQ1yzyvCi4JubzugApGgv
iO3e2swykQ8Id4xfxM+KWmxtGlyi+c4fSd/Em/AgqEHyx6N4yjOlSVPS+Ca8JpFB6QOn/ojHAXif
rlM8s2+JFi3P0dbaZUKCKZXWpV9xpQQefXcsUB/GiA1khG4KgDALZK5kkxjh4fu6LGMyD8IXwc8k
JzXYGXg99C7/iTadGaXUdlLRkHqfRSJvqSey8qqMM8g74M3BhO4Q6eFhzY4Zb3iWkvOcy31fEHs1
iOLxzimaS67oz6efCTpULa6KzjZQzNbaj0Wa/9yU0E1lTXYoafObGPzpKbRCXGR8cJ25FVEx/jge
M8DFuFC0StUvhC5uIAywdVeH7gyKpAYjZsHIO+S6L2CCPPzEPmxBY6lKLG1s6bC/DfUl31ckce6c
kUN5DibxMQzkvtSXST9RUQLR3OEx5MfneP4RSo3z/JhjiLt1ZViXu1ejPiZgZSzDqoZN9CKG4ADA
4nWv0IT3X/4ss9MR7L0igvsgakFn/ksdsBLK1pMfnBH/NjVzTC0n69JTnt2acN382eW+EhiWuXLM
H+bunaNSTf5bavE9u6fHpZZY2L3Bhf+SR2pov5g6iK7MF416MMDLl04os359w5Kz6BT34aGXhWlH
cQqSq+O3pYv6VhuJkCaGwpkO4hWtuxbexUGFUGKxFn+Y5JDVc9ATzPmE/1NinS942N0KOeaG2WyZ
EFzjgOchWgpPGNBfrKuQcoeE4t4pcYa5n+8a/gac0tT1kqbnlM+dMgSNVzncOtHWV+wKg9kikREL
9btCpYkhHCuDF52ES4tbi+T0g/r3PrDH7wO4dIIbXL6TyWza26HvI/Zst2dAdocd14poCGNjbPS3
U8hlAGdWCZeF05Cgy0Kc9dDEFIPGhsawZxJgfCj30RlRPZkou/n9ajyG1H8/OxGTGCOVRTEB9hlT
TE159FrT8tMpndfw1TWQCN/jSxEuBBZGtis/dsGeRazcKa5teugjNM0vQz5FkD++kfwi5QsaEsC8
tK9St72p6k1EK1IQT1YmYvqKj0y9k6Mvn6QlvvVwlBeaDXiVy2TJ++CYKCf24aLuLG2uRIA+IWO5
TB0adCGY3udu5Q9/cNnQRA+RBB7ps5b3X0KK4t5pJ+onep0qFpSuOBhmeCx/Ad1ptwL9KNkcGwX7
9qZKIpxIw0okp64I/90jYN0cidW8uyZMurkiq+KaeZcMtLf1Bwo+J62wLoukN4fd3qSDoMiEJcuJ
AUU+K8RrumJwXMm5O5G2fFA90FIz9WEthhkxIXeNxdm4nX+tgouKZEoWznltRD458W8WnYzH/W/5
wPPqL73cUYWRv1NFqe1oMZW1NdNqxWBq66TwyiEH6ig879MSFX82xl9VyzNxsCUfZ64TIbJBDAJv
UhwIRSTss/osU1sBNutCqp6u3BXmaUPoxqY13XFu1OTKGAcII0FqJiwOeG0tm3gaq7S/e2uPhqcM
J1a6kdyxrTD0UkmJ9Duh7auPSE+GkfkkAHZkuqJGct3LW8i4lgscy4hA3f7szyTA5o1IbpvwhBtk
2dtd0UBixnesHBBlssUoMrN0RrMwKkkmQGDdCllS6beJMrifVJILaB1o6I6eLUqh9oGyAN0UKvvV
gqD96mYsk7NhzG/tEuei6pwva7YIN/eh5IYNrCdb9aJM3OFUn3UwALCtRrxk7/Yd/ujU16Mx6hMG
+B3HzNqupf8ahEivtWv1UsBDShOwU2rkZXo5trtfCn2SQ6oANIWoyHMB+6HKylFfWUJNKGWnA3qE
9pG6zfm46cKBD7S+PUXKy0z0y8LnO62gRiLz6UH027qyfut7z1kYk1VjQ9RBQk/4EpOUPap4511m
YuqQuoxD+YxgjxyqG1+7HP8pfC3/AjUHEclHH8tYEqpcM3qSjdbp0iYUwhPJrBiNn2djJZ/qCUKk
X3Pt3L+PUako0mlTnuRrBMqfUn42HdqIdLXVeDvL0I8zgRB0i39jTPjMnARH6H6rhnLk5vgC4PBu
DIg/sMyVLmNAh8vibCIJeMg8hlr9uYvSprRVpeDKTKGp/CF7NB9uIkfSbf+XzfJzVcDdISX4em5/
oUdPkoJieZv9HODz5AgeUW96CXgiv6W4/JxZ2hJQprZhdUmcypzuHrfLEkZ2xNBMSvHkC0/AclcW
s7oLjkuRiaiGGKp9qwuXxuw1/feacxxpkPgdSV49q53B2ayNUNfRqSMrgwJaezeip58fv8R26550
t9rQhI18L8HGbsecNjR8vhfkg8ZZvglBu4TsAr4uZNyWSZwG/JRD7PLvVi5XD97ZybHjm9cV2M/3
05KbEbrtSYsTT1HOfJjp5d3FV/5JkGz+f4gHzilrSGVAiE+CRkXNRQAASRqgG4U305w3DU7ZUcGS
ur6s3Ch5yujrkwha5kcUoC4WJN7ImDeEP92kumijEnw6sgfo75jcQj1BzNPbupTUz3vlEf8PBmhn
SzUitikKL505gAPdRmeq0LJkBZU0xdUHgPfskfus1VH2RxRgVKLrmAbYz8oDUqqc8X3eshZdt8VB
w0d89t6uBcno7b2L6oOQuWB+iw1cN04wL10wLaD8ZLmJa8LRfAoBGiJlC/k90kMZ9Hi8lvCrTAUL
0Hb7i28vXNi73PglkSuwfQaE09UVoagDFnHzXFlIN6KyRuDDbuQzZnNb6gwZG0SqSvmQQU4HF73B
i74R9rG76KuLGjqxaDtOwASYZwZwDSSdYA1G3mrK9teKBK2invN2eXyf7eNdwSB7gJnJtughD4n6
QtXe4fpKZLsL1BgOth9fxpK5q299sHRHIwPnp17uJV/GpePDIaVK6y4WTnZkbXEtE6BzM3FVWcKg
FYW9IOkK0S+umZOIK43QsHdMWfD8yGgL/xcrMxNQJkGy56eG6IEsDfvqgneuplh80BgmCLDsjDl9
vK8MRek+uLk1UsY04CEEWBznRZdbOxBEEjYvb5jiOaPfbiq2StUkT3HNa6bHoij8EfuR765Ki7Qe
z97LXznP2sxkNLutnTXhi+vTMOywFMYh91h898nIvCgj+VIXU1hT88logWnDxu0Gp70RmWzT27kv
cayajUUyVI0jRBQEQWkx0It6Ivo65vBzK7KttWi/HiWOGzWwJJi3ZmxOGqXkHVcgyecEY/f6+CAb
BaCvmqCFyO+FWGdks0X3P/oCFgn87A4BkuvDbUYJt4J0Qi8pMfvE77AH87Q/kwBuVoBWtXEe+BWo
k0IILKYiVUJI5coUQKwfJSE0ZL1uW2UX2ONkq+nr0b7NWGtGtqt/2D4nsfJ2kmyBANvbFVNd8aHI
p2tK9QzFUA0s/+gsFzDjx0Bg9p6aVxwaAzrWuxlHeaKjDMfm9GOCOaCQKPbXff+a32gWNAcrPUTL
6qysEDwFK7qvAILM835NufEquXxDVwo2pciylFcSaRSPmuFhSKwli738OA8E2iQBptCgtbg2SdlO
ksbxYB+neewB9CyELQajeRyc85O8UmW4c5NjI4mEgXfqh3l5a94W+XboYWwsfHgNUNfbqPXNNmHW
OsJ3huNPrAQVvWm7MaCLgKQXIrTYiZvFuZnkGgzOMn4rOCp2ruBsOUoaS3nGCk8AmloDVt1ro+UE
y8z1Q5UDbfWOMrFbzf58ZJc6eSDZ3h1K73K5D2Q+XuHhkTyLX9eSrovYxiwy/hlSuL22r4nt82yy
RKZGH0PTrmXJdJuytuPnjrE/GSyL2/M4tM7Ed+/p8BUfJKltao2BsGrx3fcBnFH9ig1qEk6r8idb
8llKEqFEIcGnJ1ufJHOmCfsChqObNDHSWH3wnWVy1ewRg/8OuSpMe8A0DEfviHm8hBg0W6t0HLFS
y9wjDYoiFb0p+RGpRhaTzDF8pKO5evidegPec9l9jSPftdTpVrJ3FyghjUUeYKe7E7FYI0RnfONO
CgFXO3KDiPzAn+dNrLPUJmJRom+jwt5tFCCxxdt5epNkVFg7xh/plnAaWfZPH9FWogNQkzjG9evX
y1PoDXviTpMAZb6icfsWSnC0f6hRVJ6VGg31kMMZ8wo3NrMuzyLhFZJfh72tAYLRvFBMItFHiFzb
AhDpT0txVpNIBWq3pK09w+mMLDA/QztLHwZ8ACuHvjKHGKQrgJM2Tl7ptqTe0q2N2vHENVZaCsCU
mT2XChASbmkVf9xv9qDhRB2e6LTScf3vL0Tkz/mg+pQp0CXsXbugeAgm8/3mQHIuHfR4kdxDj9Q7
ybtLdxwbe88atHXScYcA2iRaTo9KTSDUl/QrhdS6HNTSKUnyKQIW1j7UMihSpFMeoqmXgrvgB7rF
Q7OrwR1HUUHDEeyn3NQPidGOQCp8crrMJrsvm9curCYjhCDcZI0o+J/tHY2iLDg/82hSgQMG4w1F
rK4AWGTOlmakuNwy8L50BlQ2Ja64nwQycQ2xLHEEBV2Xex7/iLNYfQdWXqfHcQruuYojEndIKM3q
0LX3MKaFItestP6IWLrvGA8x6PlhVvINUKkFEktYVS72DttqbbVaBOylCyfsukZHK0lEjvzTITfs
gqF/HaP2a88ph1CLsR08ZH/7TFdaRg+CLsKtJ9ngYFtzhEYdZVixWgC2DYxRjF6evNJIiqAxlL9D
apJk3w8Ya6AScpL7vzVdYouahu0uByMsRvnIg+sfneia0kbRI2v+nOc5qeyfO8gIJ4oelN5jRzFm
xqEsfN0AYzB+Ns6jNRuxd054B7xMiDjTmI8PbXPkbSOMm2OIHidb5eQP95XT9vdcwz69K4uoqyPC
EjxOYGRDOm59s5lvHZhXktWw0wHWjWZ1OL52vlPt7H2/bVRh5zqDjDcxH8sRUKAkORvsCScSJtfj
67OVYHZR3cuwvndUt24IYC4Zz4rKD7Xv0F/M5Eszgc8ySaxOYSSdQeL3Ut+zeNex4kaWriC/gcFz
XyB1/uE27s6B4pUGYf74+lLPwUzUcojO1KXN0gUVb4HLj8f43DiJYQK0kxpPIMX+BGecBYIR+OMU
fYf25GfjKdvkOFvz49jfcF7QO/Z0AvEC1uhoJuAT8j0lO12uFEedp5KnzF8vpODUAeKjMhSiBUGC
0G/QOgC8p87x8zkLqEyY5eLEmM4AiKrftK1LPOlvmKG+DEPMEYbohh/DqJeoXMr9xGNf/fete3kE
w6XmPzZ/fhlE+djBanQu+DNUn026n/fIh7o3pU1bnz9WNF/Jgi1/LZBz46H78lvDizNZkllbY+vE
AxoqbAuml2ZkVkkj/oK8wnW6NMsunOZjedfZHnRV63vEgCUttTt6oeDJOTuPD6QFxzmSMCQ7Zeqa
q/fSehLQsUtzc7IhmHjUCixAnN2oc+hXkiVavuoWFUHBe4CvIfdRDJOPW1/ajUzJHjL2pTD7QNoK
mzSksOzhNT4Bn0UJccTHpblHHyNlkq/1MTXTHr/ujoDq3pFlE3j8UHCUt9ablaQ3k/dWH/I80k46
zSUSbsG6H4pUX2WJC3aWsLSNGy3vKpq161YJmoNinRxiUalQceW/rRIOTzseiL/9B/r8erGZFWKW
Fb9I3Er5/zfpitxaJVAOOTX0BUYdpQUfK3lw0BDC1Nup0RcWQPwQ4c1zCDLsfDsAswVfaNBtlDi4
n/Xv30N0wYR6MapZde763QyvvQxJX/HGvlHbNXZBtkkvxM8qlqXSO9cN5pfxkDl0F0IMJ6jqvWvJ
h0BCcDZcZj9iUVd8tBgXen4IlinlJqOIUFRjNr+WXxvhaz/UdZgNjfB6B3qxOxvNXibZ7QYwV4bl
bXmmflcs6f3O/sgjMgoqH6j5Px5MXb8hgB1w7oU7ypmLhgoPA8cjF95TnTUGvCEscNVmkGZHGG27
Ib/5Zi5fDxcUb557brm+x2znHMB/Ch3IWr5+L8UbWqT54DJZf6GZfmqQqr8sHH5KJHI/hkrOoO3T
Pi1ih+LTsllmzazfuKzbF9ksE9wK0zpUUJZEFskmQTD4o9VDuySqXsdYoPYOIfYbm6eqSYB/SRTZ
XujyzlZFrpu1k9G0/B8cps1VMneA8DIErUxX/ba7+rXUU6sNMUFA6I7tLwkAIjNAdbi1VnD3NNZe
KIclb3Za//GbDx0CSRMUd7+yzenrJ0+x0lSDS1zoU18ohTzX/NHdQWQ7t83TwFjFARriv8w9DNBF
7GbKFTQL6bgpBVaSkOjfUX9Y/z0zzuMmQq5SnXkgBWzn980yM+ySDBVrI3jUPa/oJbk0dbrSIgcW
jk8cFgSLes7mYY4nazP+BPeOQGEA60Yg8caO2FFZonPRKG9HKF/XmBIfQ56aKBhEwf5hywwTHxmZ
bUNJbqPmmZk46MdDoVgH2xDqY58aDhbYn1nN8BfSajXZzeTykeYDi2gbJ/dp0ht2fMtkpfDFIY2V
6QqPVrrdJBfhE1L4bCyGi8CbFyLHLcKpyHPenfGfW9kmWvbrmLJYHsOrfwsUUUDyhmL8BJJzwyqn
sH6m1b1mWQpEsjjy2L7FWQZNtqB5LorHZ7lfl1p4J5e0/ekoN1hg/a2JvLOljiWadGHMZZuqxGHT
/uWg3zhETA9bd7RBaieuHnUCQqzNpTGR92V8hnO/UeZJKuFwQi+UwhQyLcp1t3vAbazudfARSF8L
z7BTYHhpdpL+v70GFDX9NcvEGSaqax4dsqNDlrvUDxEBzIU5ZMw49H1KywK6Fwp8INjydIndByNS
ZYnygj+tJiXsbbwvRUuumFqV0qbVjjf9N6FMv2FiIn61tJ5qP81gPJW9d2U2KTeHwdA030dCUHTM
a0oCiA7nKMksk0UNydumv9Jwp+UHU8QXrOeY3uQlcyk5378nTnOYSoyBYjdanu/wl+2g928LLYci
ePhpuQ2FJ+rum5qLlsXo9b9uzuAD9aUND4xAbCuygyY4PFAIU7sTqe8Sv6RD7VxKSSuUsSgWkpxf
Uki+Qe1l2Z+9go/3fyGJjBhkSmZOuC3RvMrcc4WllYzqcH8TzyBOpe7Z9kX5Cvu/ugFfcOTti1lb
RC/nln/gYjedurK+tFek793trAKwMQMiJDDvzl4ifsQgn/xidXqHmvBignxwHlvT3QllaYupAJ88
2xF0UVgRz68je2ZlG1lFsjMbGhi1liqa9qsObDK9FzOXD29drafJ07LQHEzi6RfY5JC9fYS4scW8
T4fgJXHvwpqqcUgKRH4SYC1kDX9Pl1kdPsyfpbPCYaqu2SPDNcT+KXFEsRQTBtK7H11pU+snbWep
C0DK5XJAYG1Ye83jXR6pVDZZ9h+7LCkgr/6FnbGz/sI1+ZN2tOnPNPWcae1Vu+CmvqL0tBoPjuhY
QrpYkSIP2MhRqrahOCegZx1B8q43RXsGtN9hy1PhHAHh6AXlW0M3QS/2iC6U/kdFeYXbXgIoYvlD
bEiH8ErgwvhgoPIwjNzJOoIVGMf8chW7PSjiqTibBTXazmPm9Q53G+3sodYo6pbG07yXZrGaUoVL
uDkBd3n6bw+Tr2yJ8pAgkRo2ap5y4GT54JkPwcwdUELVt94RI/lzuaPLjGSMHlzbaCgjCKSDvwzl
vPol3YjG2ef6S6gAXfF6mAhY6VUc7eBV+KzlrEQVaCyH5PzYMDN2je+GWzlxGXyOTuXVzV2r7RLd
4Q4kgzY9gSn+cicil692Z7cGtJA2KDpWQlyw3//6nadf8wygyKNGyFJsb44OqOPBHtEO0Pa/oEUM
SBUA3VeFTGgWg6ikU8IKHHfih/MxFAJHXaiC28qSgIK0LAnUWwOj4Ubv6U2spbD4nACQzy6dkim3
SKTCYHe3QBpyGbcAoYuvT99g3xiq5ZZfsJG+mbNTgV+UVceLNOJ6btp8CNEiKBKA/Bh27xmfTYK8
/4pyIMGfu5HOAyk1NZ9HPKE6g0BLttAg/G/WWJqKo8Tfc2+NPG1GWLXRAs/lLlnCjZRHL43ddA0R
NfdYK9h4B/Bpgg2FeyxvcE/dbEfqM/hExSty+OPmzEIsVA8MFZ3MtcrEQmGSMUMoToPd3Mlb/ALQ
OJDwT6BM7kYS8OPB8xIp5MS0pIjdQM/KRbzmCgWMHnUJNkwakKS7WiMsI6Gs2ljD6MAilzzStmht
Tw5KvDtB8CD3VYd+9zBjwHslYNbw1WqLClf0ZesO8gN0b3GCw5lo6dZ8HDY2NgAHXJHuKfmm07fR
CKAQrdJ/o5L4vYp6EPvdRwHgfyDErhy8TjYUJCPhBrVUpduyxId0LnPBJNFFXwGLPUGV+ExQeJoP
e8VnDJe3LntsN0yHRfNBuQvbqDSvBsUFBcp51BiZdXdfqq6gdrwPx+8fewQCkp7N+7VYFy2zcJSY
v3J1wpa2ExiSEWO/mTsHsDyTp2G4LW3+lgwqDDHpfwiP2qvL9IG/qI+NQrI6+GSE3kak4JaJe+GD
OUCL4pjLzW2MEbqz/3ZLhjVcWrkdVqwywAvkCd2zhOm+TNTgY6GXaDfFnN0DLv7LAUyZfw2ThMCs
Y5AlFkwxAJ/LgRmk9bQycazxI47QhDzXcPhw0L0GfS6VfxcVB3LCXHwEHdjmCY/PsxGp5AD1fs+b
wBxsduQzFA2CmSgsBfv+nVDRyZyEdA1PIN2oNkbD4bECykL7M580q0z5giD3FRuycsAHeMkZdrVp
Wn9l0zZWng5kVLQvYKyLmwbDLLHylScSK6Z9EGaJZt7n6e36v11s3i5kNABRDq0Yjjnl+pOrJbGQ
EPg1N1SALwAu9MGBjZ0xUQVaXqH72yUDepDmwLPfFRu3C7UhM6KwuQVZP6w3cE4dexDTAlYTkMoO
YBEDZsSOPwdlh0inePpvLw3qodRk2iUPAflOHs6EqI2KczwxabDPBsgHPIiPrAKc3Qh+vmeI7lrA
4ZWUGyEhIn6Tq3gLuh2FIsfIyKuWJ3eP8MBvyb5wYhKjzninfrUc6SfhI5/PAhuydeJdKEOfgjdP
yDAQ790fyUh3Yh8qnrxZS8kwaZ/2FfDJQHjQz9/REh/D+wqLxOli0km725jxV/B+5Ah8QCR3uk0m
WTHDzMz+H53YlB27C7oZt9hcF1luDbagbqk24R7x359gP0Qgi/KVhHRJ9mNrDzFgdbzlkZ2IUZ8J
ucDXQC8ym561eEGq2xTplby8sHDPgbg+5aLdDardN7qj/4AB9ROzNihwhFffSMqjnHgl5hFXblNb
YzWktM0lA6KgWglbWlgw36pZZuohFaEv+lQOFm2cPXpiqppAyE0cj/9st7e/oYeaoQAj5aLOW5GL
N7H2dHY850WSV+aZ2qydskDU7yxepEh4JMxnsFGieGCWAzmoYyvZ6HHUb0g8/Yx9mRnvynf/KWLX
guX0zWaejBLAKQigRX6EJqPVpLSYHfPdgesjOIgbDrrQnd/yvh1DOqNp4TikSIBqVkPoCpOyhzhq
tvr+XDuJcHCTQc+PPr1DImp5SqT5FSuoVTZPGm3Y5p4bO4QqVuXfeK41yfCISNi3q2oUth8ou2yS
c76hoGTDd5hKrp2XPn8i3tvmymt27S/sSFom1Sc+EHnbCsU1bcxL1IFHQUH1e7CLMQ7UPR7y7aBP
gcRtb6DpHX4F1aID9Rje8Imjw9AxXRadeC2O5VNjfdQlEZipx2/5ThT1sShbyePWrKe5UOBI0STz
5b3iH/RkeUabR09qNxA5P4eMnNq8osPylPAxjdT633HOyYnihZqmJadjNsWcQ4+Lj24YbcV7mno7
dbUGvvWS2vByC6Jp5nboX6UJ6ij7E9DY6fnwt7EZcnyLQ0N/vSRb9jPIGpdSbYKvSzERtR0/sgHd
0+Tj+VkMS4RpeKavFPdyxFVH5akDl/Y3yJVyyqHbUUjQLMEyH3ikZcJUefQlY1qPPzOVV1BnG5Xs
8MUi1ohZazXRs20/sdOscbz7tms1cmktWfhxldCQ0DpC84mTbFWjK9aQX+wETDL/rdN9t/kFgHzF
aFJZhpBYsfCPwP/eTckxT+A62hq8FYTsf4h96qbqI0Buv/SToFBXUeoSUgaWCzDhKUah/62l1JW8
zBbe3VuvLEzAEUI5LkfHnA8c/ksP6ob2cnxCrT/fk62vTV9neZm4GHzaDg+tDx7G6SaDEAZjLYA8
+XnIbGLcNvylLBnXk7AvNUISn4KDd8tn3uk0hmuRBGKbz/qWApoCSoGlcVgCR4+Etf5qDGc0QgkU
jKb65hLJ6JY5r8RIge5nKeYlvC2jjUiFC7lkADf8kdkKThg9wRGZhcxyL4kUTiHsEubR56IoEOGH
uTzgfxCeMtvd6DmtfOCVCdKy0+R/csm+XexNT/+QuiFOwp3MvsIPgl+W0rbwxMUTNlccFDtAdTLq
vmgTIQzEOdRWxT337d7d70jkeyK71+4Y+eBR3lcbrE3WLK80+QrnH4p//I8cPt7ifZ92QoL1qz81
b/AQJhMDqAUDb7tOPkofAIzT9tqI3RqP7mR6+jul/bt7JVJjhTuaW11LtrfSVuQ3qyKgVp6lrZto
XXP3j4Afie9l17cSY1L005OokIsPOI6TfScLgx9E5xMBwrQe3bcXWsHasqLXgBfkO9NlmPJsnspw
pHhOXiP+dT30+/ZXdloH1cVlgGC4Z0iIICkpyKhBkyrEU9gDUy+XarffDy80Jb6UtERWJmfCLxo1
E83jjc+e7EOfzJSac0u2+q9a5xVgfKD0SLMXxTUIe5zJrJ9G5yBEpg+yNYdUzuaE7c4Lxzxx2wZV
v9dHKD0w3IMBFQjQKoCn0oOnQJy1i4bMf2fy6jdZOYCgAKoK7d6CaMUwngp+78lXvaWVoYKBM6Ol
r6WGjoEf+2hH3zIWSWNkskgefZT9NbA6TGVI0UBHNxoy7MnmPwhk0FwWnU1rDlejfNLZzzJpuHdh
5gjiQwPsYF/KXyBycv24bqGlKchTl1o9Q/UjULrLsab5rP7Eewifyc17+MLXb146s8y9DkzA/aNf
YEaOa3t1dC8YNcK0DTbNVZbd3MMbhqQ4DY/5jMjkhBmC2L4ghC9aTAIXYt3My0kGUd0eaUy3Dt4v
L90jcMFNjZC5x7JAhI4Ka3igVpAk4YnL9i2pPJQxQ76jVyQluVSiMI65R/t9H8OuQHc8jL/8gDBH
AAVBHiG5gQmyP9EVGvAvJPqx1cjSXhZ0l6zLOHk0Ekvy1UCpaCTebRn4esz8ELJJOwgnnpaxWxd8
qghPXxtj/ZHENDu98xvm+VfTQvxcPhKDLpC2kz+mKRX7eVGgslf/Hr5lg6Cc0heQtcnkcXSgSp9c
Bx4IdHdWNM2LrAnsxYVn3PAF8PBh5MTthbM76dwyt8u7jte0FP9pjFKzjaP0b46GbL8JLXoYH7qF
QJ3K1eCutP6i3C255b7++Pp7o3MX85/NM0Zozci77w83wVRrB4bEQ9bKuarryg9B0dGkAih8jGmV
+qrAwVNSGAyCPz/w7oL3ktNUL9r0Qvqq7PqvbXt4O6OrmaSUvDd1jxNwHN2rTUTBbocAsifUGoDR
foWkHEuEmKUB+NJZElxxcr28YY3MRI3nOm/gGbzKdDo0QrTdimPw1ICOsiTcJeu7HQzYCTDUm7K9
o46t7RHVLBPEYPDvPaeyhtMIFfPKKdLROxLBgorknrCRpXCrvsTtt1YJXYUbZQAFv/xHmY7MeLK7
QU5mw8ItqZFQ5G9VZwjzyTsOnagX5OEU4g+PMqVTBp2HUEIu9QNY7fCOZTryTOm9OKGyYy/odMFq
OXphHvnxyLdw7Y6gFf8XbiV/3FoiBOs4ETXDc6QQ5PDlNjePIBEV0JJERbWTy7Y0qROToQsTkCWu
2UYi7zEYDYI/JliBqPg71ssSRgj+hxV96YRcEQ1mMylLXIBBsuadWWwmK/LHnyrZxh1PqR3x5x2I
eh9Aat6qQ6UNrPo7QveaWGY4ICM1o/2vKrgBVX2vM8e1DT8gPk5zCDhm8VDC/Q9IsnB7eTl3qXm3
RhOYIyB5py/c5AqP0aotArKu8bcUxufTj9GIOsiw6gBES4cbzzkg92aAiElc1XnGqdRJg7TcQrd5
9cnjo2IzxPpLJzutx2riAULdSUU1qWo3LH50Biy+bQLU4i9CEe/wf0/Q8W2kzTmuDS9n4MKT6Ti1
DcgEX/5g0bsAa0977+kPxn0O10Pc6U/HoJx8el9q1s4gwwAjBtXFzN94GAlNgVAy6nJ1+5RZXxoL
hAigZCH8790qFLafG/crwdx/uMr4oGtv0chmYNXjZbxmFKfp4MuWj2hzVGInmVUZgdR+7f9ybUOA
21ywNguiym2HvabQiRvqm7RGorDNssb0KopxsYPB9ZIie5sWmoMSJKn1JaHTSLpFl0F2oFc7gHTy
zjlJeevWDD9MzgvENu3fRIIbG3rfAWgKq0ppa6qmtISgG8IivuVClUp6OebXzEHNuTH2C+QhjfTU
ZOR3b+EBjGtwlJXxgty5lnvkCI1eIp2cH6bT34Of+/Fe9k4zBsZITyXDo1Qt2O6cbp15jIRh+PFf
J7udQoMakkZ9D19Zvy3bUnSO+D6EUNE/daK4NeklNREwd/BcncQoO1hHPxhKnXK5Su/Z3eu9bkz9
tZJr5SRhtSlpjpAoDUNPTYd6zTzSWne2Yljt1zNIeKo3E/eLPnICBMpgKhLIlpbLagV0fZwpYhyT
eaHN1p2y86dr0L04+yObCHpTcwFHAIlOnWRJjxXHR2ybRbHkLNs7rrWAs5qFD5DSU0GkRyCTtx0j
r7FS8X5bSVEcZneblSCC3q9GWKKNoUFiP/dUXJiqfS+SvSU5inEKqeRLWNcwsptLQKStcFzIx45H
mYCNzcXwbHKTyVyC5Xo1vjDV/kEUZO3CDYLHGSG9gk3zRb+AOQk8ONc/sagunBtimeL/nqGFEe2V
sGFDhArj1Cgl+uNMQQ8HWT2f+xkEqrmA0pvo0lMAb/q6VknERub7nWdf+7UkUWoAl3uaJ76aP88h
RsDD+02ucq8nXjpiEvYmBNd2uPE2NX4Z0zqaYdP2gVSimqRvo2dRcwTrgBmiHtFzyKWSXERZ9z6M
8J/+N+Kbdq8RtJ2zFMPHR2UjGmN0hQi2hjOp7ggOUSJXghDXKSjGAybpOLoqUcoKbAQKTXDeNB1t
6GTeHasBEGuKatE1CBXkgCYOSyUmJ1EhN0i95Z9wE4/tAvf3g5AKShJXnr7+/L6kLkeIs/CRfHMv
4sJUO2z4jpGbKuIjG1QzNamsND9Hwx7nHOqPDwLewVty761Pi1wxapUT4WdSrb+jOpSFOmSYWY8S
Tiuz4yr9yKhA6RR/vUQRMXCYi+fTqiJjVvz+OPFaRsjPQJ5ohzd158mo22jSnp3pNRDU6uJ/YYNv
9y1fc8W4PcrD5LVCWaYPQwxf3u5bzOUoqjM4P4zRqna9oWqJHqHBjuw5rjdejqLejBuRy1c2jW7u
sjRP0xw7av26BLFQpSYQWsiL6HDZR3X+guYDS72yDQQ1ytqYDfDrQdXTtVueQ65G9QJLH+A2ZuXx
D7mdZIq2YahihD3d8ap0ge3xWy3M5iQg/iHDd7kVKLnlH8Crq0o9GjHFC79F6kH6QEEMpWVu62Qa
KrWWuS4InrPoPW85GCzLVpeE0g8lIaMub1IBXXQIESx5gbSH1PmxPZgeUqI9ZzfV68QMfcRP/fgY
w/39qM5qQL1BVruv7ufOGJ83L1yZuRf+Ow9f9BkPENEaOsB8g0qmwNUlL/5bQhGGRj2zqQocBE1j
ZKPbhB6EzXdQ6wlcvbKOjVHuELhHgLDp75DqRQaYPotlMPoFFTCbeiRPN1SXgZzRkOvLc9K5N6eN
Yrp+kevV9RVxuRh+r7H102GSuzlvBewlG1jwKfSy91GVbQmrK3/KXWCO2fnzAKHSGRED0+qwccq3
5prUAeQti2m9TADEPm809llK0qMP/TL0aXfAlMFLqB4amojEzWMxezCSY0NRn1FAA3tT0KL58gN8
TLnw/K+nA6MAzLtSio4gDrWig0xHfRkewS3f8hQxjVCZL2etVgJ00Bw7nGeu62b/J6liBHKg3ftB
VESbhFrwclVjI9gvr7iZ6UxD6LJFPlyBHZOtcwp3i0E48lBIv1VLY6kpGoMWZvehtajse1eEzmy/
ykJKFb9jx1LtR0gxYMcG8F6WEb1pnH+y6LdM5tJ+bQRW9dLqKUVRmDknF8wB+AqyJCRtggi5fUnd
7i/N5nYHKKzHdLWEbYdss0RViHXckhWwQTFATdhWFboJcglPE4GIUWWqLgG8Jywog70joJeZV/Mb
j9K03fG5ILP/900mlh7400UUs4EcqAvqK74JH2mV0Iz/03ZqtpSHvRdZDckj/zcuWt0x9apHlqk7
xeHuAWd6D7eKqF1fHDYV/9FGdyvsMWGfwyLVSJ/boYnYSj+FAo4xRvBKs4tBYTcwsDvt/fzpv7Ls
glCWoeCguevfs0w8Xg5ImlbQyHqVCSO88KdBLc3IM+kgmHwsN6s0D/jVeyWrXYchBq8JvvNJ/rCe
oouvC6MWjKSyAwE9ifVJTaE3sUDl9Rzw5CJIWclX6uPzy/JBC8mY//udBeNNWLnb1y89tY05KKo2
L4qKSoL2Ob3aLGbQIZLZLkyxQvzSNZFt5WDBsTXIE8oLE1v0VHMq33TcjTW0U/eQFie1g6U47p6C
IDh44L4epKLnaWNcRmsaeJHfb8RO6sX8+tNviPoUUbZkRkGirdCFPfAEPNiHQ4j2N+vQwiBdBzzT
S2izI4gn8DgdRRVbN2OkEASs9Nxu3QOjhYTh0i/k8jq7rqFTpWtEuLkNUuhn4sLnTgfkke9Bg8IX
Kccp7kAIPIhYGWygJHQtkvPn//QsXbzJqq+eNtD7cffautMySYjc7s05c6d95whqig0/UfW9i8CS
I1PpWOEU3e4CjlYPsUIhxZnv6+fP21ahGKAryOByqUwLxGmoz631jZMErOcOwlxBcWbeanQybsOU
iZpuwt5orYvnWAc284dkZli3SuRYT7/5GY6n6UG9akY4FNlaRM9VDpYMq16QKRg5nb3pONv0nP+P
59YhxJ9vry1D3cw1f3clotvroeY5O7CXFLOyGU6/13xDzCfqdlNNjQ/iX2dYfyWE8YNMUslHr9r2
dRH/rh8G6/RGxWfJ2DHS1Fpge95rQuIGHqfxRDq433OuKGASzdLZuNy75n80vJ1eUiXm7reByJgi
cr97cNoSop/+EYiiOy+mRPoXoSaVWj1N6KLxAUGZTmdT841bK+vYgc4zPQww1W4VT0UH5RODmpIz
QtHdAEoW8zmtWo3XAN1BF9cRNkVOyjOJT90GIn6qUvhe7WTQM5O4PxwLG3a9gdo6AH5/wiAXPsXT
DmJUPkpmjDegBifDrOoQkFDj/CDWBrYdHLS2HyPPmWMv5KLfxiArBXfItEa1QKUJENDLx8vFIdf/
UJQks0l7EcD+AbueCvZ6oWaDorrczgVIgiwA1fRCXmmohNoO4Wm49IIWhWf1UUNvFRHUfCpjaTQ4
/g7qiut+ZR4naN6IE5IQRS6CyMXMsVrdZ82sbUnQro6BRGbZFk3vSN6lL/s46635PdgwE/DYKSHP
6ehKkPG73HHBVd+LMC7R3QmAOmvheCSGWUdWRTVBxFTtaCK6tNolG6jNxUOsfObSWPxtZUq4G4xj
Ov90gzcq/chM5e366g==
`protect end_protected
