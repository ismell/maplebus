`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SUXCb2jBIUqUBHVlN0KPH+td3p2TKZFkfevOFlKZ2ylGNwbKusPtMhbEawoW9JJ0K9Eiyz+toT/p
7BwBjMnW9Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BcT09+p9KTltwYQFP+cWp6ldOVhCR3aeYMfocuXkweVU4J1pKGI3DEKzmhz5NU7r9XQc7lkMMb1t
Hn0hTUFQVI5e0mSUtCkS8sen0DLuGCCmCtzblkhAK+/QVoPp0mrt4JcZLjmR7n45JcA8hZDVsKvB
WRTNHU2saP5hajEOils=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DOrZ3ipc0lp5XyWYVtHWdLeAzigiDawQXTBrb7sjhbm9nv/ZmWoHNirIqbodPnMJ6e/tWquICHfZ
W3RYlxL2QzrlClDCNMIzCVaFqVdGVVVxQ1CJOALPvGG3dltR/Rb24nT0npXJAs7ffleb1kqf32I1
XtNO7gKq7nKKW3YZ6qAzjjtnOcaX20zeVWRBOC6SKJtT29FQVwapEUEsFeZyaRCXwgyJAlnsyi4A
weN/uNGaosxTeyUi3CfGTgwoX48cmI1bJWYaPt5q+UkLp7oRJ5grLNaPafzQniTGGFClqQxSMwzl
bG3UJHLqkTWALL2O7W/uhHiwpXdhUDcqNOh4Ng==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xjlzt8Vc0gLNoLfvlgzWUtUEK2+RCkp9337xEPMzz1K9oxxwYuLXr6wg6IfA2Zr4kxHLpN/FnvAb
H3kZfyvE3gmi+BXT89f3QWXABVeRQliOMv+mmBn/OLrjSceJoBB2E1BgixJyqMFMZlST4UnoaLxf
n+GhuQ7Pz1izATR45j4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DQKDJqOXItRBwnrst9GQlPLjJsR1Xdplvzd8+wGTvl7oPLUIf8+bosi017W3UEjnil2tJiF5Bc4Q
SHMlS6sr4EvjpFVXDCxap52Ze7PXfGkdq5RFJg22dsmozjQzAIBN0eoo7J6WNMFT4ezK/5ILZbhD
s1ASzUJUaIw66Y5bcGrVM5w6STHYbmYPwjr7fDTbppkcamsE3fx6eFcDB0P5vkoeZ/3Hc4vWG/WB
RE0JJuXLcoE4TM6Yxvt6flzNyus/j/ixSZyA1wdjP/QnLoxGE+wrRsbdw28w2/VpBJmOHR5yGx7e
/IC+kPGNoygynH4b5EhwgTJjZjQZJvKmfH1ifQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26736)
`protect data_block
i91Ajb1vzx8Hv7uEUoeJjrdn0kzmcJB8ecMMfO+iUabeludcx5u05pPnKylq3Nw9D8hrIS5YSfIM
DHH21+Tld1ZgtGsxliDpU2pVLhsgElz9FUjnDKqt3vxr7i4fCGULgBJUmGskS8h5VqHg6VzshtR9
heBPTlj94l3jFviNru1sz91Rvw6lrtZg2AqvbL6cFRMZFE7YTtu6qo49MjSACyqkNwT6ioPkDwr/
3j52Y4i8QzC57kxmTzb0rFR70BMvbgAq2UgxWjdIs/55anRuTwdpJOm6qCZLRQZsCm/0gxHePBx5
fpaE0jHoppDDBZhzZrkgr/OGNXDqtIRveNVqaKe8b/7nhILYewzqCQoHPoLSKuXgVS+pWac9Xh4W
78rwdk+Yzrj0oaBs0pdTyeiDKfsHcwpF9CVs3DeLSW/1Bgk2LKpkOvjgOGGu9rlZiRICg1R7/LqV
vlMXyIXCE/CDEHvDBcFtCB4KmHlxP+ABiAZWejGUkcos+uYIH8CKHxZbsGEAQ+Cfl37TSKXi+2G6
GykpixGN39MIMqDh5BAROo3aOfuIxpRh5kqIXErg2gThNS/nF1eNh3XmgJ/qJuvW73m4QwzGXJ5G
Pauvo7w9HzyLDR6r/E9ZInJHennTFPInfNDI5hKHhk1PeL4eMxcugOlxUz2OhEGwev1mZP8DoxyE
vErn+UIAJnAUxpfZ/gGBFU312ZtwpzEwv0/xRTzXlV57VtFsHJ3xeYJ1tid662zaXbLdplc5emzE
NDDCKT5crzm4jaow3z2s9GoUwibieab2m2d0UeZjNfYiBZrG9hR3zzi3Gjzpf1jahi21L8DCTCxv
Di9loom1XSumIhZu4fJMQVQT2lhagBbYY3RtOQ60jGP7LB3uWbhqvpbd0JzTOfSbv1bhFZr9rBLz
oOKNrYTjQJ017IlwfPfuJdhQmukqOzPH6Bz/v2LvgtpTrx9q4DyDqXLsEM5Lmu8fHDgysAQvr5S0
rXNE4Pgji8J3QqCZXhMXnuBETQ66dIffrqLJUhTE6ZJc3WaKEKTK+kTIGvjjV1I5G0arT92GV9aT
veP+LmDERP3py4h8Hbfh54rfr2UnDF3f92OOR5hQEw48q5hLe4ye1c1qxv2sEZtslxROz41G/jeR
ioghYzuBrCtS7XmWRBWkIdQEUaoOqrVr1aYZbQLPJGSt7xfPUua8wMXF6udumbQ7tv1BonsiPdza
axgbe98I3j+XgU2tV9DtugtnpxFLkTujJQRWNn41uQ9v2Xf8Ex5UZ040ZgONhZmWRvkS74ms13n4
nrKekO0XdAL+ImrWO7XUjLsDLQ/sz6lxt65Xi0weXiKNw6rj2ldSdqyYQsmlsYuMs/32iXo9p7Wj
F1QRJOVO+JvIFa9xt/vQBjedjuwjQWkKaBV0ZI2+BeWRbs2Kkxr5YK81m063Fbu74g4/czzht8uK
8gMCiWikUVY4FAt7orxTGoVOFsa39b1uIENDkUXx3GmZwLyOlIDAilRSXPWIIdy0pTRUFdYGoP2f
/mSwWpOFHeD1x8kePO8mlohHViPRm4DZYGvy5Yb5o6w5Wsc78LLn43PjuqmRYJ2FdMYHG0j17wyH
84jQA+LShsiuEWRZwxpGL/WxvqLThNMoGToso+I37nBbFVQDgGUU7YDrXQhoxXmBA4kVqGMhYSRS
nLM7roQLus8ljViuxQWmoAWyDLyTlw47SboC96Z+fGMuZNGE2xN7vzuC4SkJkEO6FcG+nL5gB3zC
PTzgbniSXuvb6GxygIA2K6eCZ/bFQEZ6yB8DQg5B0sQ0noKHNunQiyHwI0f1nhTNL5veNU3uH9KN
3lFNwSKIZ/5nC80260orqgMSyY9LzA5DrG/fD1bxKX2rcg4nukkb2+IlV5aztaLkXLg33KVL8q0y
0X+0FO/BFKLXv1ljWM1t+MXUl/wT3ST1ae245IwKLwskDuEDDBZjIzoeAmWmxsm41SGuPHg8VOHd
LIwUoIJPoyRFEei2yJqr4sqyO68l2Pi481VtmzVYzRbnwv4qvD3trUlFMPY/N+lqOmGbsqkjpi6b
x0/0WgojMe/XpxOAX8LMkwlDGydy7bIEaUHiKe6DSb5aDAxqhYA3KjFI8cDqKhEX8MG1GNLVYqlf
ewuVa3UDJIgr72BdYo3dpt0eMguQau+X2aXhbiEhd1jayl1By5sHxj97Nrnu0QvytFgQHC+HRIYo
58pR/LuQ5Vp4jqzVthxqcVFK4twi+Zn6Hw1/Wgc5+2QWTdSmOcSOM0vZ6sL8V6BNmxyyKip1SW/Z
Np2SRd/WBEhGU08weIH9PSApOTWheOSX1jQ3NF2ojkHE+nvjv+2yUZFuGW1TEQ6NzqIfvnED/HZ3
XLKktbNP2BHc+5uzZOmI8hbFzTqSjUHcCoHO3jcflRMrVEZeJm0WiAYKVLynv4EP24a7IFcioMEa
BV1Lc5CA5Q9fo7tQe+bJpZK0R2Vra/oiitquyG3Ee4O6AbR7mjwoD7ttc4/VUvpJr+rxZ+VvC8Ap
s8p5yPwYEisbHMMWg/yWXXuunBXN1piCJGEP+2L4v1IW/csFz9v2cAHgVbFIe6kOrF9Jye6j/Kcf
6hdiTugJDytDbhdCQDm5JJkmRU6runoLcWBp4oGoMN8rsmmVxhlpk75g51PvHSbMvKsU3a73KMXx
vA6ZS58FZdDD0+65o9vb2r5aqaAjFhlgqCg0/Ch6k8rw9kMt2LLO5DbAVBdoLIiVEt6BwNkCjm5Q
rEZyFjZC5B+Ms3+g5GSlopuOob8z54UrdRWMGyouF8G56xazH5XdJjG9dDmegd/92ejMsuC/gzVO
QLJya8GSptv/ZLG/6jzCK/bsOgdQ1kHrIq2bLWZSGXIul8IfX6POqmspyNlT1F82lJlDJqEf7csn
IqLGKdHK4b0RldXd4+LH51u6CoBa2GABlCtrpvcloZKfqLhUUJrU1AC7uM2tmawHMTS6HcvW6q8t
IHgoOQsKVGdsuUUlebv4VO/tj5efiamzlZWnCCOKPsOgNUXG/ywZQp84yZJBk7mboCB8u9jzuvvT
RAIWFjEMQvgRMhK0N9zkSLjFBIkUHuWLV9ofW1CEGjkFamy0ZP5+/3KoiWJux0jXCsVuxNIV114e
Rd8QyV1Eb57GejasC5/4+frKc3HXIlh6ALYsr12CVsyc3WXmTw4Rh5TOro/8ZtWySIeGT3qoKSKT
ddqXReOe1zO2Y4Bxs2ht6+/2WOIvSLXe6G1AHfK7eMXEcGH8oJ4PD3SZTqcDsKoJ4yAp8FiI4RN9
VggAa+Ii4onxsddULrINr4Euc1vShQ4U0jqu9YoflpPiBsQTlepuZRrKp6dv4ynIWzjIQ0SO1WlB
riJ2C7+QVOBNZ78qRDeLZkWaCH1p6p+9WJq7tZLygEmlXcTdwepZIw5bPmPTPGjlO7sX39gZlmlb
tG/zTb358iQUNRdu5p+hMw7nfsL4hOlgHmGQNbDEJ5KMLz3lkEN2sBxBSr2hK1ra4cCqqF9zp0jQ
tvtdfMd0GGCqXiRKPsi9Pe9wtUhP5WbAzNLkrovKDxJOSXJ8jSLsC7c2PnwwVPU3F9NnpbNloXfR
M7+4GNZOEsRoV/v03pjTiVXkISiWBGJQs2IcKcwaKw1XiAQX9H+X7i6ElusmW3wclayBmnJsFOG9
2wMJEFeaWuOifBR+ui2UV6k8oheAo6nB1LPLD6D0STzYk/hIB9p+4cn2M9MIS0enauYbEGN+FgWX
eBWOGrmnEVXd3MZj5qZiFF+m1EM+ztKo4eYguzIP+uyfSS0QWYgzkDjPdfNcEY94R61WUKKyzyrE
Q0JVdsbfE+NuyKOm5Ggv+toV2IOIyzJR+Y0fC3uH14ETrEUjb1XovOeRWWTvqTJYgxjDeUPCLlA7
N8xI/8JBRzprclk2uSuhx7Z9F3ZeeGS+vjs5yoHK9/0OV+w941nKHL2YJ141+XDxj07D27KtbTRA
i6hgnlry+GkL06hBkeenweIfRxZW08jBixXg6NaQ/ftDNC7ZB8IvAlFB8382YKgirHqQzeDjdkl2
XwX/rdIfVovmORc54mAdImlb+P5v3ucjRt3x4LyfiEdW5zqOHY76WUt7t4IB22CEd6OC/TI7ABbB
VL7SU3GRvV8QN0MIpXdxVYDoS3Y0aRovHLsonErca1pBR0ZyAFQJD7pYNVb8eMl5rKzeMu2M4Zim
GKLDSNp51wE5MrljDRU68GYAynL5bL80GYabH/WP7/v7MqpVncefqwnlbN9sDBzKP/+BE1R1Jzml
f1QflOQJBWmR1w2M9tUFThgbMo/U3gTo9FqUKpG4uOIOGUzSgGJ0PTLE0+UAAuCzvk3T/IAIjuKV
DHhTqC6+yTvsHhfEfbz75SdhZovTlpwOobzE/URLkW1vkr1a9BjFcLJhibUUaFW2Pq0cx6S1/ILz
2GxT/Nw85qHcjTE3o2uDNL/GGnnIfVtCK+9nWBA0KJ1ookyWovwOzUI08wDIJRQJe3dc8L92PUnv
kNVdcD/KptYckmFWyVPkR+C6h5KMOAQEqzW98oxbtYk6sVGo7hML5ZBrC5V1H9pgx3acPt4YaizK
zxgjpoTL/taV5rOlzf3ZEFNee+Vr7L1MElZQ53zon15eXGa8sgX8DGTm0r5nQPzw62EEHFKvIr6Q
w5psmSTk8TA1gz+l71OIC0A0ZgaPHBnV2b1L1ldB8j2N3Dxtw/GONEhfU3T1f8d82VKKMJ2zxxFW
E/flOEI9rcD0RZWoFnDYmrgRe8FfVbTp2UMO7yhASr9J9OQDbC2oAtaJsWA0vDS3psXqlIu7XCeH
MVXCSE4xbZjgP/YnX0h89k7N9S2ie46Wt2Ou+oVI/jqhsXrFpdjC31pgYsWXcOMhNd9TyCYVM3nN
6MQ2f8auLfrJ3G5kuSeSL8lotBltF7M3AdXnsg2I+SJ0iPxThN+EibssxvI8fC24cNhkBL3mnOqe
cafYAsUW9lnQqUztVBfTurm5rDB0cx4/JRAuwSXEwwlFtI0s8yh4bCdc4+JJUalG8KKrH4tlInvv
w121V6+0iXLsMQ/q1hNIvdJ1xA0yod/n1W/KLo6UsGQsPa+0RZ6v0tklYwbi+pgks+sc910PF8er
ZocbIAN5o1havgNx0aeZ72c2TXas8ekrK6jtNVBepwz42KxSBN5K+pcAwr9ob/nuDZ37eX8MKJxM
eLTDjZIEfCrCJNjFxeqUc4i7JJXiZJ3kB2zB2CDG7B1sBJmmqJ4g3P1qM2oSmMGwZ6LTuZcaSmIT
Lgzi8fsjBxT/tFOnX/9AB6PJcrTHdDQpaHVjW/Y+ARJ3bwxG5VwkkY6PrZoQzyqU6NY5QVpit42U
Kwdci84ZVbVZmtQB6IGeC5nCe+yF8YGX2g/9nivGT2K/FF5flBYnW72zN10cxiMdVu5RGnulJJDU
VC1L07suwBMaMzhiQi9jYBkO9UnF5k5uxMGUeaIIoComdw/tpmBKLvuqKYoWG2/r2nGn63Ysp2qA
1b3VN8GZUyc7j/NbdVDU20Q7sScwXZhICN5hsKZi075hJ8b7n/MerPEFJmcyI8X7Q6KwWD0wGxRq
jcM5mVI4aGka+LPwt4W5ZQbMJ7FzQukPtPuTrLn8WLgcg6y3Aj4A5m9YVjsm0KzLYFX/LNgPeywf
LOk6E2xPV/jwluqQiphU4wyoFcVk62XDHCfbcHSNLMNcI/6+9CBehhwSUP82f+UjSBnjm13e267P
QGBr8x1xEAZbDJ8LW9ZnjaPxE0IEvPTpX3EHHYQPDwoiEOf4dKl4MdtcEZ0EaVMObuxpuVSg2++a
bwBK0VnfaPB1g7HjIEA0fWQsi4ysxV71kNH+b8Tl1VvTxep6QynmaVE4oTlJ3BWYq2b6hSMrshCu
xEzolYVZTb2TvxrkYYtH2lCpTroTgXIU4calCrggQ7jLxIJmGcf8xwMO3xPe61kO1XhNCSx3m9+o
vEHeBgiHjkIJeu6f33SwrlOW8WtHeIATLZaq9a8OEPL8bG+6PDXXmYZd1bp5Ly/CnTbJ8HjaRFCF
yPuQ3AyJaFcXm/5VCPFNbWe9uqrwKHd1wHnPnM90YV3bgxB902ZwpqNv/ko5TPYrPJKoCjD/Ln5/
XIebL9ttnmTXB/ctbk8y/F1kVELJBKNrcozxjhy2bpiX7McKsfrrXmiCFkKN8PFwIRWkbnd5Irhe
9E7lYFuZcocKiGGvIduHigkfQ82gO9qNnHWEsGDdbGRziXhJCZrtNzrM7WLajMuOT5mzQqb97Q2e
mUnDRz/Bq371mYn2N4ru4PYtVhYbBOVUbS/I+Xj3uYM0m5HI6yOKHPUqjytdbk2yQUxFUnh3FOiF
6qwAOLXPQCR2VeK7C+/I/E24+irf1cTMIxMWKR9YT5ppiC4JvG21fHfvIu6e2dCXzQmAYweD8rZD
587gHZaY2VcGxFVin6P5oHuGyXIt1xTovK4QYYdrgiCpUTzkpNmr5UrV+wylTo2nbdFEut/8jnlY
4nH6akbWVAAEokG21paC3wfpuK8QoBkHz4NcpQZB+I1ZDwAJWoC89JtnDgKK7mCPImujPHJ5lGma
qAqHMZKqW7jFVwPkeNk5M29JUq0M630tz9mwRURNrJS0QmWWv0st4nbaqMLCDWqu2ngHuEJXsf6O
ckJiBVnAACdJli+UC8j10sN2gkwl6puU0tUFyYjHgdg72HSxT/eby4uqWf8aPPklFrPfIq3J1O9J
k60JwSeAGyyiz+g339OnuT4pTd/HJmFbV9NBbPNxCMQlNhaqXSYyy+uXC6WfBoo0cy7f0X8/y1Fh
OMggylljJhDnvllc7z5T91qp27pulX/7LFNBWygmprHMnhkpN7DnciPy3m5HVd8gkakvv3tF1Wer
M7gt94VrCiFY5VtjY2nUmfasj5+sxM4VvOWWCCoWqI8mLVbNUPwbnfcm72T3ctpCD+WzmlUC20pv
Y+5NjrvkPyCwmcG1rHL15W7gfwfbJ9weuHGJhCQkSofHIKDoANAFhaXD2pq35vQtPtq5xMlrDsHa
u1C/251WckjRnKafEG/D/W4R2KNpTEISOGZy1+J5ZWGVNX53+rQpo8UAbzczRmcZKGk4hEghxDKA
S5Jm1OR5+0W8s86QsRkdoXiE3kQjh3wkwaV0lPnLedv6XmXYYS0cflQE2RjsQXTwCqe7mJKQF6iW
SdlBE4roblfCDyQLZkLGZmPMIO6d+rt1JM0IBRoU0/GUCdl79b3UtLMuvgwvGSGuQnb7YBGf7yWn
Hs6Iv3h+aS9jIuTMRx96fuH2WyhCyYKBvV1DCNYK9g6umKk0hhyyVNthDs3ZiK5+wu6SiV0YLlpI
mi5DVH3d8/ozB5oQpa1hiikHY5WS+yXz2nGuC18g8Y1Oykw+bGB4bp2sIHVdwl5ThucI3U2PPFuT
6kdEmUdxvquxS4zQA3FFg63wS5+12eSlIRb4qYVPVAvD1d7nKrN2xOKyJP7JEayC9FeAeg9pRnYt
Z4vELfW+5Ru18v9yM4hriQoPnU067cNSAr8kiipmlqTTTULUhUnvaa/WtvKFIzvavalTnkdcIcwg
h4gfD4N1Lt0yDfX1xHBqwB5n9TC7DV/miKg8byz7+tlxwnTItH0hTgotKTMy4v0i/X3/xgz6FkLB
HdtY4HrD/Xud3zLfphtqEGXNmM4C24Po7WYYonnBQfRbtCv1e0L+FLKsYpOpHfc15rTKFyZW1gSt
FGGtEhKo39aG8vC5yjkTYFnXuShdDCveyOaKCETnxdMky76Gb6ZhZ15LHGgsD38F2V0ysSikOBRD
nd0IsArwKcz4WtE2c6MVNb0a/Yaxo6m1ufsYLNBts3kBJwcpl0NXmzZk1ltAJbrhXZJ/+93A2k3q
ALdfSI/v2brSB9Z/7emvR+l7cppsLk82n9+DZ1QhC/fZB76+iGaV4mJ8ycxdElOKLtPUZMxj+w7w
CcbkAsLoBAiQ1OtUseoIvwuITf/4x+Q4EJmW3EZybWUveSnAbmP5kdac6V6yPUuDIjVX2auH96ki
8Y5MwPX2AlbieGdbLdF0g0Y7O1WFNHL8RtexMkXrtq7Oxcm/VNleKvApcqkTsP9AKbTDqjlRa+Rz
C0fcDGIUe3z+vWj8t6AVjA5yNI22Jh4eIse/g6pDrT5cQ1wGNZ1XYf2l1mVDmvfKCB32anHLEfyo
aHsE/0oi7JaAQJU9FcRUJfxSymJj6HwRexJE2NxFI7C3DVc1DMeFQ3JVtY3QEv5u0Id3HUV71Lvr
2lib3bUPi8H97GyLRJh38YZAnNG8U3whVB5GWiamkD8nKRQiAFxSqljKgs/GeJ2ENRdd4qZdSTdr
xDMSGIMKVSvLD/pD/dFx3Apn+nxWDzodPaSD4XDsqoFLKD9XJS7YjeclLN+bUHkrHHKhZ8KnPyKM
mhWYnQDI3YA2RUG0gcth+aTCYydDECxSzRvu0mvxtF4rVTE8qrrcNXhpt5eBSWcr7NbJ6LQz9KdW
0BTWkdlRrzFcmFwG01RkXW4j/7D6aedBKUJOK5cwOgU1hOoNXk4zORjM68lY+w+TML5kXtoRwrEj
AL7wqVClycUi2VHvVcX9i17+Qp+Q9e3/HaieMB0DTKfmX+EAi1PipTgmnSG1WM7Soqv+Tc42PfWs
F2hok8GSYUyQbbZ8Gg6UodxI1X9OxRkwno1FXHxvla6dJzZywHMZganOHkcBgCSf5JuabVsgcwwh
DubDqanLm0txQ1kEKqS9zK81foru8TaQz6bnkXOo+AiThwgozKjmRSIeNsKB82xa07LyBP93ZaCO
oEAtbEX0ULYBGDzD8jiXRZy0xj1R6dHYiNQj3Uz0cgK5H7vGExQu4yuTluTdciTMtt+XysPhCSUw
4VkcfbQnbuxPr99XE3GHlSJNxDJYVMAMap8w0WYkH5VyiO4waigo4GPakAf3hiCxwjdtolvauRjy
3zpqa75fPhmD8DH+0sx/kNBiWZvic7xOVuMFxe+Gns/vL/Q1B+LvHSd91ZMKvlDL8TC0T5nq/RM2
arcVcy1KTDhN4EppzNYZHy5WOLQyazZNKD1SQKw0apzUShce6+yzsjj67ukk1EospCweWV4459r7
lbHbwbvF05ik5s0dQeJsVcRCSl1rtGxSNhMQs8EF+HnteKAxyWeeum3KfGKlaU3+YUqg7rvexxhc
C7JShgMjDWtfyIxiymL/xmi944c2bbSUut3GoKX2BicP0CqyTbxTVuTPLQL8JFv8VwZuQaIRRoSc
Y2DFAKoWWorcXUC/V9APWgh8aEoLPg2zCX7oejxxKemTrAqn50bgc/3Ph81OYCxoTw/dYpGWOmwU
es1WMyTKKfZMMxHCVSrMU2N+ib9mb7c/rEwL+EBJDy1Jcz9qqzUhFfKZrAI67VWPu96MQiI9tyr2
FFrhCsxLDyJFH/QSrAchcHcd7eDTqpN4yiAEtIaNOgWBi80lv70dVDLexrftX8rJ5+qhU6FhIm+/
eDZJme9nurjTpzU728JXGB/L9NN4hELjQCcRDky8eXVBWfGd2FzOio84KOjV5esAQCEQZatNLZ1v
xNP+kWQmRzHQVyWZ3wPDD6uAmClxSLzTlkrCpPukc0L8KV+88taAWtdn+lcd8MDJmVAtkAeNwH6f
I7lO04rdj8nSylJFZNeJU5G6K4w80bAZhF48rOkqTjzx64iVxWc/eSWxOWZ/cyAv8unyCO7/UvL4
9t0VJXB1R0SIDOpjn5J+R2I6gsvOAi71x9cOaHk9d9MNm3Jz+vJJ7cosO3EMc3DTv3jHrBaCDpeg
kSNHcTrOPC1o/zqKXjylAyTaWKDcOQBvoFtSlzcV2fWa2y3bGFghk315sFLpIxjJxBmS8CSf4yKj
0gE5Hl7JwiYcoefNINyknoYTIcf07i/fvfjoTRbKGbJ7dioJXhX97/D2fw7TPKGvE4pm7sBuHxYX
jsQGKCwmJs13S5rYrz7Jeju04EeRCMRSbl1t4QuE4ma18sI52QLZsqon07+ThRThHjNDOjxpkJfS
5HySuZf/GzPCgprjCPFpX23+PRUDknLqH5R6s+izzkvbaNt7EoImz1p4pBLmGKvxHF5tQzua9u2S
nITlKTSt0QY3WlluMiZksMyGdh2XNnI+/DjT2PqqDaWAAUVVGrFW2gghjXgzC8qWr8fh1/5lE/wl
qj/2uM5LEYm28a8mcUjmiR+z01iNMLEZd0tIj1SXBf1fVO5woRn2YAQRCVWn+MRmBdUz9EZiXDbB
8NbPkfoP0v4+vGTSHZkw4SguzOLIpFOKDPy4lKJNo8tiwow2cTGYFR3uaaZRONZbIfQEjsw92O6c
kqTjOGwhhXrjtzjN2fjZzGr3H5j8lMo3bO74WoTCutj15Th60NoRiHZM5baRoeZJTaDL+OZodS4q
PrAr3hyDjQOk8cNocCfJJfq/bUqZlpyOx5xDuhDQt8gys9QPwEmz+UwsWhz6LbQ05n038i+ha+LE
SIVqQrnulTmfBrjE/tLCgerB6tcmG7aSV0rCnExuJ22xVSjpJxuYBRVdIV0vacdibbDkRdckpB9V
zZWgdTG6a3nDo3w5GmbeYq1YdcCfUBQ8bJJHG2fYOXVOEacbrfvcxrJdjDMqWXHz5zKbVFbwU5IN
b8s67ChT+9xn3cntthP82v8IaJ89k0D/1Z7VJTdRXJ/fNBfGHmK4GSbn7CvjdTFae7FHpCnnkQB8
FVx9HCtO5gyDDVi4SviiyCkzaQxflFxIj7ajDTlh0WTZGyA2QQfPn6XJMKLs3cX7QWBSB4QqwDi4
Pm069m9EPSry5uC/TMi6bzl5xfTyibFTjelYw2mDXCvWhU6PcT3wvPDu23IeuHJ2eZx4fWDbq+KN
rCImYvNFd++E47i0L0SHemrxV+KfIfx6sIwoAz7ohVo2dIb573X7G7MEj/v3N19DICME0AIAIQDC
9PP7rB8P+pW97NIF4EbSHhjl8b94kND1N70VwkWzmKlt5IljIZx8CY6NUwWAWVww+mKze9KwFN4h
6sPpDRiiAEUuD9TErtvmQGqga2vcU6E5JOL2E+t0y/26xc+hMwCi5q9TC+D2bdxlVNcjminGxN5A
xei78lcBe+559OTFKoR6uO6Uxb6ObWq704/y+kN9htXqiKO+EItVU+vsGVRffmeHQJdjzrDYFU2w
GjbO1Kb9HdT1TMfPPLb8H9DB+5Cg+T5aKvDN6xKDz50vdX5PejiSUw3sx5QvH+Zvi4+yfl7feO1X
16ItQYOf3Q0Gyqiv6sou7hc6FS2DCjJPZ7EsAxDpeAavDqjVwmQ2zJw2CgkqEiDTOCOeumyGa49I
pwwwjSOit7rS44v9mx04yh2BIbWAta42MVwtPVEmK4ZqvKlQTXYnc17zVDa6oWBR79Ju+JvXe42z
+qhvKmYjdBh2SsC4oveGPoHvld4MnUau55AOe12K9oU/EO07snjjPFTQQL5QklwgdfQpLxfgrgIN
7pfO493TdOa1JruoIeeyQF3h2whOfYwHAlZ8M+VKSbakbJGcjDzqMhNjGE7u5BD+cSw+1iKU+her
1YYjWMzFwadkftIm74YodBn5/R8M02SezmIZGZ+tAO2aDbJQMDVvFLYOcyemqoy9+YuXby4lYgIr
2fki6+I7qmQiWbFfN2oO1OJK62vTKqcBrKYXPvoznFDGwX8on8bu5liJZS5CenTPoyOLJmslCTXR
c0iIXSg20ViMhhYn0NaVoa93yEGpNpwlS1mTNyYnevvPBmzflREUTW0lVCOg7jZzP8ojWpc8wqZK
WVWeG16VR3G+LXU8nT7f+i1lH+S0FGAIw0E4TIY+ivFinMlYiLwUrDC0KOiX0oy09Whl6KL6/Puu
ajBcL4DkzxJSvxYNTettHQzw+pKarbgywMKwp9gjZEpj/qvgj2YN8zERdTu7SZWK8T4vrCguDWpe
9HI1G26Qbcboket/bvBfUjnAtPbY1v7Hl0hLjcUkRz5Ezq88jyKvY/8tPUz5D2GhCvy2xdcHIHmv
bTWhblZP5e7wX9JHSKung0RE4Tv8+xIQJtTB++Df2/ySkz8NnLacmnJluBl1A6TjkknHIDa6Mgn0
6yaxsSVvPTbJfqL85YbvyYJd6XZLSPrm04wsJL2VIYwUQAnwzqALhCWatMCajk5swrsMHrZcNM+5
5lwR3il706OApQ+T/1NLq6BQwnFDsKkn43SuFICR1xhDccM7atl41sxzrgrZ13VU+Idx6PHK2QJz
I16UF8Q/yi7QkeD6fm7kVujsL+2KWpfUqpgicvoYvKU0u5HUAQcBRGgFCxoEZYStir8WR4Ki3jhR
sn6G2tCR3tkL9D6BYWp8Kh9fcJiCLQg9zVZPlblBBvc3vfRRPtokqUwEh7MyI0R0oJu/ZWvMx9Lf
N0MO+sx98ekKa65p0cALO9KwoaYZrGssdSN5dhjGkCxI/ikjdgrOLTeWS1cTiCx+Vk0y0AEeVCwW
fvRTgCEn03S7DGdiP7/fyqA4ldvRfrY0k1IEY+JK/WQx2E0BLpnoMTrEO7ZdwjNmtw9/1Nafgxd+
LEi6sgTqNDaFIrzGLTrJaOsy5QvreMcKob6ogkjL/m/BcRFD/3MqlDZ6zuSrOShebz6he2BdpCcR
RDRHohSBpqkUrU6j1IG31a49A7IOQCqriURAFWVdDXQL/DoEyIId+vkV1Zrz61370Du6w9OhVMfF
sP2iO7E17IEOYep6NAOfxP7wc6chphR4SoZLcUmDUpPrRHarbK2PMjUjiM8X+BjuwU4fB0qyrxDW
V4Gdd6I8JbEx9WF0iqlMo131Ir2r2pdu+fDzJOmtjJkHwYLVYrkngHuBB02cSnXCvzvAe1QWbebU
VrheC2EIr72GF7JZVQ8OF1i+srygFKwmhg/nVrL9/f8LL1UBeUY1oDxVV0mHoiot0R+Up9u7z10O
SiI9XGzKu3pdI6QmbWP1xz68YacTjQ30VaSbIzDI3YCFswkSXYQg09XgJPySWjgxnTDw4jmcpWND
TRez+5z7H+SHTqM2Xp+bmchXMU7C9FEk4N/x+tykg87IG3TP83UN3nim6SKW0waPvk4yLXENE04B
kaa41fd0yvTTziI6qyQgvr6gZ6GpaB1WCC16799gX9EBkXKT0u1UPff3ejL0plRpb7BAc/RIwCCi
h/PrBdjiMy7VjpnE0kDQu1RIRHEvJT9ZxSWOVdVmovbqC74GtanF0jVosKuBnYo/JGst6Y7JANei
TuP/rh5dxRrg/mDNgoBkg30ckhK9OVFQllb3re0gRwz/f8FdMNdGlKmH2URGos5VnBZiTenkeGse
uP9RCmQ7ary9kCXEFIn12ADkmSopSe2XEhyBw92K4BcRbZZGkmxveBX+WyJhg5Z8FZ6bhx3G/nCU
HkqWCrCY3yvuT1P6E31k+atyRvyh6cnJ8yJdq5U5mHh+u24sv7WxzK2URm4CXOk3lV6GPi0RZUqe
oBnrXQumeu/mo3KrCOgvAHxzM6NlQwYtB7x9cdtF8IRO3VzLO1AUI18ZlHiYyy9j2cL23ZbyabWt
72S/wgbOiR5kULkaHqOEp5T293u4m0kf2XkO9HST8v/GwkK24xyGphYfJfAAbm3zNl4qJN2ojRk8
+RPcmyoZ1UwmrVk59Omib5VZJ0hbItVQOl/kZ3ejY0zP2Egrfu0Lk8DcvogFCwm5xSGNCkxQuWgn
EB15SvuF3BrAyKkhBKzv2KFv9sUiypUObyJPIKm05l8rxpnkg3kHlU7zf7MnQCMVWyzPK63eK9kt
Ft3itHE5rmCHGlBi4ki4CiS/X4sXr0abI2f+bv5LwNZ5aHGTnFy+gvSGh+/BEhDEAGodFfV4fU8t
Drrlzu6K1kt8fdMHc+MDCEoxXW9LptZgR59L18hzDHkvkGLdRQEUT4Yk785gn/TQTzcK9T/hhQlw
WRu4WqoHSPuNT2NfD4vuyxbOHe40/QsVBl4Nsy7rF86/pNS64fN5E5oPXCq7/VUqFzcVgjJMr8zZ
EHHx9/D3t7yYRstY7iEXSOD+DaGGIErORQrvPgBkqgCy35luy6rje1Ggtqx73x34I0hX2AJ5YKSi
g1CiIJFMhdhQzu+FqUa4zs+HUgitjdEdAv00nj9O3FJEjtA/l3azgU4br4Fw+lB8j3Yrz+nHH4Yj
CJ1IQhnopDyFMZzJXdFxb8IPDvYQ9WYpI95KzAXR0tnMyXWTxVxIIpnfwAHoEuBL1+DiKNP1qFTP
+Ca1/aCR7HztOJJVphsFv9r1NX0CgR0PapiZPyrHppMuYasGo80EGY/uJE5PjGqKJ2mfXQiv+29c
wZ88v/Q3UdthjGBdJ3izQ3T5Pgnre3OFtUzUObEMwf6MDSmumHkezuY5/CMafFZ7/WKLNHoxviqq
oXikptu+Zuxl0J/fSG9V9u9oEnx0muJYzYFGpWXkdZJhD1jKL3jL98VDQRvJtUPffzcI2TkmL9kJ
z8aIB0II0sHo3pAHbZqSR/5O5RJp2IaQVFqU54W8pnFxC8owq9KvInse9dNbyPP0suBp9b7dPMux
jIIjWsvXpNP8zHwuTm0QhngaTo1OFGnLcN8PqiBJ9iZnmVEXr7zafj4+4JhtLAwXDCORrj9g6MuG
xNf6ettDbWK6+k+pMdfo7XNTa7NV7REzt47wwYUZL8FNoTR4r/yjp++eO2AkMHcnyo7Z4SzV2pTY
0jkZnD13MrOTLrN9onO/TV5uPTjwkjaJF38r8E/RcI4BKPu8Q6Rvz9XW2TIV1JnDYBVsZZnOtWTX
h1TbspVwB7FMz1n1uouFBVzKM3IG7P2Cfd1wV6zt8w4TKRSNHTGQ6qEKDnLSWtAmclN4ZUxZPQnb
qxkFTHKC5A3As/5Xw/rTDS//RAql8AUMe2kTGh4aNbs2nSg47TIZ+55X1DBD/FPZsb2HixRYtwpr
3lOfYTMF1VV/j/FbclUzNcGnv53ttj5dISGnWMFDor5/GH5fG6kV4BHdVutXtABrv6zlvvJHA2NB
zJnV/Cw2TkFM9KKm3yRiEEzAk8O3lnwesPDMnOaL2mjNXE3oA+EnZ5a9PVaOzU7i5G32mbRO/fal
6hz7MZPESyEDelWoRcY/AucwyNg325G7eam1fVrxUEsjwczxDy91/ZoqlZV853E/xF0R1bYmj7y9
usrO/K11mAngdXc7sTl6uxXezPcgyVEnLJUkP9ybTB3jf4WLRwc4kxWYFxq2+3B6oZ9NocmF+0qq
h8583ZhJ78hUWJ/Og+/MmxxETst0dXOxAL6QHFvEMuJORN8rqYfVCNZGWgz2VK5XrPqtRX3xT/ba
H0X1v8kFBuu1Tl2t6zcuDOoZsIZPPLhbscBgHD7bp28gF5EpRiPe6XOpc/dgfBhCbn3QZyHTeuBK
3jb0KujM8eikCydYFMNOFKGywRAPMkAb5sC64saM6NLsSPMvdgdCUjdkQl8pQhMvxwaW6In6+lNN
n0iF3lxXyHs7igO0uqpiw4mWmScH9iyYkHg8Q3OIk4qPqZCgQTk2G80+lVsKViB7RHjuJ2eJRuPr
bcknYxja8UQKdydmChkw8VYKr+sSbTntaEIbdVXmKosm/MZA+kgfYl8QFSvrNVnIpwXBCvN7ip7m
MC0/jki1lECuWwEcYxNpk4DE52de+tbH4Fj38RazNK/fWgso8EM+aasFnTuADdoIm4XNWtw1u03w
jUNksk2LqRnUI3jVkwAsf74RZKUL+2fAx4LUvXUeT1Zr2LeNEcxDwBXGHooMg11ma5HmINlNgsWE
m0WCpQqDBA8aZN7wG5qh2bwn7QQtzCsL129ulVLF+ZpQKbQj+7v2s+XvTTurp/on7WKQzRi+Taf9
D+x/bqDHK87rdd+2XaGqTepTLFlQwWjC3Zb5atgE5nUlOAXVrRYRzuIb7sdgv34ydEtfOMHZODAy
hGMrj/xl2B7Z26070CXotbLwLZ2S1L3PW6+72UZ0rOp3BqwJXVzu16jDpG7GXi5xgeNS6SUPE57f
EVEW36LnUOoiWwVMrxIRH6EaI2qc0LOGbwqkqb5rllVwm4/v6LuE5nhcmoEz9rFyJwB5+kJpxl1U
J59jGCBdIzMEidMDoENiIkBw6o+oFJwm/TivGF3XNQg5uk+Fd4DtVQMZX+AnXY0Fx7f9krncpE1B
Nv1YDg/I6jgC1lF+iH6wEEEEOjCow+cIqZl9pYsgvco++SLZNXItSY1zIY6MxywO22LBRELdtLsg
SoXRKVWkZDS+XbFxxQxUqqqPFifhN6EVZKB5CDN2maOH13S7X9nUpEn+kKhAfRDWGZv2wTyJ2K1k
aeLxKmWaDFbSOW6MsvqumzKYaPjTiE7be3n1Y0AgbS4aWfXG8LOhbvhSF7UVJD/2gGDaxOwBCyio
PjxPKGFfUh7uIG3TuQdwPwJygoYdqjDMcUkPxYiNDIEd/X2UCac3cUdDezd2Wkl3LVg2jqx7Wtdt
fK/tZoT4BNG0TZhhitFFBC3Rcpa1ZCkdPCHFazVzka9aqITvKQ5o1U16e0QP2vL+WGzqyQ33Ohnj
op47MvAp1UwxYwOW5CsgAoOwMEsqKiK3OT4lLZRPk+4l/A/10YHsAmuc7EIyDew/JTMZtt1JCO4Z
xjv99VmDQPq6Pfyoh0iJ6hwjDJCJcRi4hTYrMyNoHAtGi8UTS0BlhGXDOkB6E7bgeKMKcB6+11EG
FZHvB15iuUuHSAlMCmIjak6lhQe9c0UAqhc9Th252ltzSAlkLyk1aF8Y5vv9peAAa59YteW8RNbQ
b1E/N0TxNh5/lQEM30XrZ8QcFXy2EAizHWPhZfEA4G6JqPzUOh8qCQAOsVMRavP/6hLP62Dnlczt
Tt30DQUFTugWjQicoWzE6fM5fmNkkfmiAZ0PKeyZo2RrxFaFJm+oVG4nEikDvPDw8MT1PKLS9KVZ
tJdudH9itmVBrE/fmOsbSTtKGut797rcD6z0dQWSbAs/vJPVkuBW6I6bhViOTFbrbDCewsdUIu3l
xwMS2gfQUB9Tta2vj7kTlbA7scK4R5BtvtA8HlQRKcUT1f2paMa/6meqwpAqY0oSxXSU71PCLRjo
7S7A+gAjHYL1m2jyjJmUzsMssboylsr6/+LFi/FamsJ8UKGJBb/psWW1w59p6Q1+T/Einx9PEsmg
ucAF1P2o1zU8vGVVmjAGUG2f2070DfafNw7WC772xf1o5bU2jQ7i27an5g8/o43pAam4OqHupTzu
ghXgyeGI4cs2mF3gm+kx002GyIizy7TjCFXhm6tph6XRU7Tz9Oxebfs7zRWEng1QreTlo1vniO6o
nuQHs3aq5KWw9BzxErvavE9yGZ1IsQqxiapaZWkMLSGNIXd3nScJIGWLZQZ3VRTYDmVu2+wk4L9k
Y8MVx3c4xc4mAEefO9lCZ9H8DF8rSE7jJTTF8/Kx2EumomL4KTPqPkTOdDNFOkD+4pyne9kLmJvv
ibdv+aIMoK7j+aWFxj2z8ipm5GrZwbbIitlvz1WzoadfNm1zo0/SGww/s0ZZgsJPPDT/xLuUsBzc
HAOWcETQSh031vu9rGY0/0YtFhlAJDaK7dz3/2ZGfR4bQrfdUmhyoX3DBvqejXtdrWId5fvzauhF
Y27LZQfk1Ds1sH2hMo0C0GKSJUufC7GIab+w84mbiqtMSuwB0fVa/UaRAHw1MwpiO7oIJQM8eBP/
bpIyFIfEO3iG6I6xN036HhwYiLZn+o/HSe6V3WR68xlspMFLe09/2GxroD9D7s8vWJH0Z0HFH3s4
rh5vzbxCREokBovCeh6Ukpoli0egThPgADezoMDAPQ9WAgTRs/YysCJHunncrchwpevk4Ygbe7xv
5jWtnY/k28XLfdn8Rio/8Pi3ucz/gNjZmuBHv9Tzrsn2m36l3Z0963KGsGCxCrn3YgrhsZ6u9e78
ieC3ZB/Ls1jjsdCeacacqOosvIH4co89rO4ulWX75ngCPBpxdaLfXg99Wisy85V9Cz3GgzMit0FK
2ONAGk4DqTjKkd+uKyOAES0SsRgGxV0VgZKci3w70Wnkpfkxg4w9LOUvOEGGEHCgovtlxY+vXNYj
xj6QVUc4BrkgaoE0iSAgidFcNBH0yA1ek1Sv2aa4LQVhvS2n/FTbqR3p4qMfsasxNXgFeHJcrVYZ
kjcDlV9viR5rm5YW3n+BoPZozLUF9iESbhUD1gdjjYvwBMgEoEsfg2lMcpfcD3R8ha0qEMEAMzTZ
wOK5dgR+c4Lj0WFDFETOBmaaF+gu49vekeSFktkbSJ7aalfnBq00SwBejGaVkZ7dJ0rAyAiXmVoX
0JuMr8FqJnPxDfnnre9B2LU56k0ZANN/7V2ZwU1MlM17o5jwT7cAwLjH19dmYQXNqrqijfkLhmsC
8TIthnX43IX6PZdBdV5HO+tUY9+TynZ0NuvFGMrh5dI90lDKqrwGwau6rWxdFQSeTw+BKNissJQw
1dUW3CUwbNpC6aofqGDmpioHUscppLepBsk2GGXj9ihQApM1/W14bJnR9QqkfdOYih9tfqgMmB8+
7PwCQMzC45cPINYnsKMQvW7cPOkl7tJu+VHnL6jbfE8ZUUeq9MAfTgVfz1Iv7pSBwK418EC8PP0G
Znqk/jkGenZAi2zIhI2tfuaRimWHQZ5q+GO6swKnSQKaOdV+s52dBAigaBckmT6NQFO0EspS9Utx
ASJMtBhZlnPquo8NPyOiSZd+de2Xf0EIrVw2pKx/okQJ/jj/TEfQu8GcGcujokFVFrQokVxszynk
KKD5YF8gp6fJG80BUBcbbJWWKY7QpBoAtifPKMnHSKqrNirULsaXR1CG5VzqJhz1M12oT6HTAbUG
XD8Xn2w9Mo02oT/ys1MmEe5vf6KqpKg2Gk2mFYg9/HWSjvcFezhmTl0ZDN0RigvUDtdhQOgWoMHa
2ZKmRzjatlw10n+zFbIfhIT0tfMjJb8MwmZECa9PGGKqECewAKvU6BeRN8mQv1WLiRqDggOmRj04
M840+kZSQk7ZjGVhJAmkxcURzxsuSKrfrhU1p8Xkll0XyvLaHijS4pSuO2Ip7e/o28pfF1N5lA3n
fqmvg3k8gLddGfY61Da1cqWS0NjzUuxNVPb8qsAO2rt7l/qqfX6CWSS8SPL1lGPFJIXelxGtMgJr
MEKnIFhy/ZxFdFFloff2PKeqGdfsXUWgkRDlphOokMcE9IkghFDRTO72SwdQITS4dHY8gw4MdIee
OfsEQFwBR4yzmcoW/ume3qs2M64QdHJ6oonRwj1Y4q82bCF9QqXuL6+2tNb1o41GStgqUrCp9bay
M1Ufgr+MNOkF04E/wTirGS5MZY9ctIpcpn50kxYlDxGZbwskIvFRC8mRpjPRjdLCzIWI0z6WYvPs
Oqw+s3KE8AUFd5V8c1+NNKnSrLDKjg8Iv4CodkYprM8gf/a7SkkUAP0/vrVtJd9X/ITD6dJq7nFM
DSj3u82+a+4KeXQzdnFPr0xqTw16nWzpTPt/0TQix0Js33527eCaOTySdYiV8vZ6egEVCYtxXB/N
qlnWso89x2mEgz1IGZgLxh23aWRUXtwTfoDth0Ctw3pIeHdBv2Vbe1Vn2EkDY4i60iJ1O8r0AVkW
LOhxqh1WVHBKWdRKQXfFu7T1SHgAf3VFPJxjcOI43BxOqFafkvTcKQE3PvVzu7Y4riLOpmxZs+OQ
DHojRkWhmcArkgcx1AwcCC4vBQJ+9vlckHiT8iQU2XghGf1CRPtQ54xihVSq1autFWWlu6MDC6oO
6fQPPity4/IbSWuG5fcVdZqP4zuiiAso68Ys6Dy1y2jYFT4dFjMwVtjfp+fiCHX0fIPOE45ca7v6
rrYw9zpbuvA5ZpUarShXzxJW2ZLn6kUW/2qfLglZAWiySc+GURdnKKckM73hrEXvhVkh22RcLdf2
0WqLwL/lhMXPwEDq7NnoqT6fWFBnXnpGivykiYxG/u5S8d7jG9xPKqC7n1G0rWBvxyLLJDGjGY5d
NAAz2yhisxz9ko/BKYkDmhe4Y2CaAGYJPIA6EbJMu254qahLVwAVRQ4+NRBteeQexzDFfUeEsMtQ
KO9Vg23O+D7SC8bJz0+aFVX5fgkEU1oC3psFt6G/yaLeKQ6pypGIF3rEIzA1AQZalIUVT78SuUCk
nPQt3TV7DzYHhLTUE1H7GgjT+yZp4bQNUkIOYqW+RVHEgXR1GFiLowf7c8Jkp4BtNarc9uYfp1iH
D00hU6J9QTMpX/Bix6sJwbZHg/Mn/rpdmiUIt0vgcgj/oseO2IXCkQTGO7qRnjPIXNbKLatymHpS
MfeRCGekry1k7Wyu2mBtQhOeCYiiOx3ypyZwyPewbx2t3BBhPEKVuwJwby++Z0j3l6Uh4/JaK4uK
Y/bTs1Qtj0k6pDLYGp8Hk4xgk2JN9KqTnu2DLvBwcYTyW7IAA6akxq2/8z3Q5uQt4e27F3rTWarL
rxqgo/Il10GbrBHOZYK2Q+zKiCxkNC4rtzjrQtvBSD01k0mWmiBw5mTd7Jxtj2lz70zb8IPrleRD
YWhASXmhBmsvpNgFwav1PzK+rtHbffhQLNcv4LPISuFbN4Xf4fKO8kV4WRCtqdHbutI5WtDJgHyx
YW4qmYX5pzxSpcLCOynKfVdDSwOeEg8L/LmAnlvE3jPS1cQpdA6xV8Tq+oGqHYBpYbMx9lKevbYq
te0MDUL/gYnMiwy9t1YIKSgAj78eFlXrOEGPIHw/xDNZL8uk2cUgt66sba6ST7sd90ueCxX3TgwM
PlFwzQwuZWaQp4JWefo+Hbxh90XGKUwHFqh9z7FKnMYKzeQzZWzQPS670eSiMgLrFaJM9tilQYax
yFGUH7vBKusjaYVeMadhDJ9O7u7NU6Db4/lmiMIXTn9L0aLbQz6HAKtS7QpKDIVwxaVCUNTx7jQy
IhGdQeFRYbR23iNJBZPOWyIyqjYwkP/Ujx644SVdwJ3xfoHYgLjwhzXg6Jv08G1uoAJZ16SJx75j
kVkqfBuD7EzCrGXo7jreU6thikkThW2oSsnHr/pm1VMrHoV7UvyrEOqts5HWMj0aKb66XqYDQIFV
acahuJAVj4ZG3cFa5WU9HX3XOd4SceMFqa7/VjGDLY0+IGcGMCCen4hHJKKhNSjrjv80mCtZhLSD
SfLjVD1b3FWz6yWaIUnzcyEL9Ud3e4uJ58RRWRnckZirYnRSyYmNo4msgezUAW25aoW5arn/hx1/
AIG27Lh4QcTdSDoh6VMewPoCghd8XcmM4f6Wbh40FMg1QU+bVALqpul1gO1PW7k064HSYXoujHH7
dp8ZoTknA1n3q1+LMBDYk7JPV71HY2N6VcBjWcSjbjNyjRJCFAyq5KZMTAHlmI/KDj074Cw02Eab
QKO84owx+5ad7W98oiMy40JsvZW/a+kRjYbd+HbDCLMz0dKQkR41PobRkcJJ4L85I+bcFU/FSuDn
fyEHB+WLR05gMqUyQ4AwDFMLK859lRKFgzCT44FOM97FwW6TvGBQs4zJb4Vgg1wbKnv4r9ulv33x
DXCgha2Tn2XnCGtjoAqvAydkbYtaatbvewPNdzFIhAu3XIh3u2HheRu3KvQlKlLRTyLTOvgeUBgp
Eb4xqbx9HNDdgN7vCS/QSF0UDLYsGKlDQfAnGEW6oVXFNeTYVZiIQY50K/FX46gGNbHVcgMUeLow
e8Y1IzvS5PRPApbPFEpdPqCytjrmI1DhPoD+V+wHG2BunY2YwlrtgOStP7Vef2xAgwINMAaoADDW
egCHSurantOWFOB4DAfR68ma8GrQz/GukwpZN4h6QUVMpK9XtDJaoWAPC+kk4SyTEHLIUBPS09tk
8h4Qo0I1/Z/hBedpQvhM1keNsaRrvmXA6cBP+5qi1EE7C48NqUEtZyodaVePZKeM5vh0dbEbCPI8
1LuvLSGDsSyYjD74q2li73EopFH0So2Ehu01dXHnEwtDZPrAYTCjgpuwYz9ViCtCRY+HEB/PJfj0
66DNb/Z0hg8CyYLGQV9v076YVctXI2TttKfO/qDK3rCQJGSJ3kE0RAybVH6fBvXMKeEdijdCM3cg
3OOwLUYwv3stFX3ASD2d8RZNpLb/yaxeMvOB6D/ZLzpBh256Nzg5YpJTiLs9/g2u7OllOtzDoAAp
MqDKNI4UdWj4NiQFrY3Nt5M8vKImNqnb3lvn6kRK8tLZkXRAkDgiks49ajWT6APGi/5o3zW7KDF1
WZESTC4q/2jaGdAUzl1+STT+IRGp2GN+jDLJ+UnS+MwIiXJUslaRsvdYrUC5ZQEf5xTjK/cL041+
eJ8nWlQK/qbssUa8UkXM5rLS4AsiDH1i2YfZwzzUpbK0FKC+vV/7TuXV9EJD/qOntLKATm05nZyw
XPH+noZNqRhEtBn7tB7tnF6cUw0mBfqyu9s4MtoTiPMwosuQKX/x7qelzimamqaxl5qGhkQI3lvS
GLjCQhOeO02AHIzqrEJuO9YYmjSM7mwqfaJh0QhHv21qloq4ximmBCgZAgcYDVjg+Ruit49a8NuQ
bkpnQdfTYVkl+xc+XX4nnQgo1tfDvGEiwCuVUrIA5ReBZND0J4VLwovuSQe2G2JuvZ9hhnbgfLO4
9FPPKoHaHUAO/eRIsS5yRI36C8X5av1CAtakURYevzlktmzK2AjhZi/lb2SLcaNZ3XWGB0WFGF0r
cUyYNxTHmIaOk3kPNxPFrOnu2uvduuzt4K+3FZ6DRSEVCIJmaKFqKQy3sx4zT6iOw425U1CaGynk
qRGLT7LpvyYGbfvwXTDQYsBP15SAwwnG4zx3km0gNLlumscXxmUN9jDVqShwK5Ar+v7iFDJg68o4
iR4mN9G8OASywtLaXhCrkttQpxf/Q7XyF6aH0joUR+/RmC3NoPuQQ+y3/UvxQOPxo468fN0l3zKT
F86PTTVceyz5jUl1AKkKJXZl8mhEZhLEeY6EThPzXHd2Fb4tMM9xunpEc0eSNhEwWcTFO18xyRRz
vH1gL9B0Ktps3yeNEkDFOOVBBLLXmDPk6mKTEOdN/MTNFzAoeQLWgtU5VP7CO34Kda5MJENoqMzl
PP7itLraQ9OHtHnPNIcBeie3ZOF6JRToEzLgwz7+UDWxTUAdk8T8f5wKjMI+eS03bpasTnWb8r9n
rqzAZDoLFJaGTTPiyGXIq+geb02GO6aFj/kmfQPy69732wz5pqJsf7ih0V9ESPUefZJAXVBohkdB
dg+lfjHaugPBECdpoOQxtvEt295fIfvjAg4RYR7lESsWUXcaScYjcLCDS2BUBPCT4y/A1BDaRbyC
hSj3HZ/Xe5vxLJqtHXkpTvrStzqjKdxQgdkFZH5XrXFTC/e9esb5AjWqeid4UmGVJRVAFrZoAoKm
8lxB/BFm2mN7aUzXOlpKQtSXWzZHyprn4uxqAjMjeu/BjfJka4HJVp+aKeoei4PFz0dLdTRVJMKv
Tm1uGlWJLbObtJxProzY+2Tsc7HO1NZkXDWGbcvtB7p2CovnInoivuTD1tNmUksHD3SSfBjqTa88
xMrdGVXbzi965VbIsaOjtAjNVq66vJlf2iTsE8YKoxxunDoZjV/wOPvcQbNLqNLwYbeSiWfuLqcZ
wLxaOKiqZLNLUA+E78xbt5PJSxzgKbVOWj9NJLs2i7q522Z23MgzHOcJGMAEr74Bfj5BaD7bRm9e
Mc982NhpsksSDwe3lBWYkERsrYgis+49Rh2dls9l3ejuxsvHd2DkLlwAmBE8zDCPuEnNOUCujA9y
m7YFpKFm+Tz68Km26QX0yIISYyM57GhIAER8RXdN/UAqXkqyybx6Tuv6GV2O1SLPC/hmGRi3au/9
kaP21q9kg63Oi8QpXgUQ5rmN36R81xblyVsT7HmdwMiU+9Sld6W/jol7vDx82Ykj59JwAKeOZVrN
VZcLWjOasX8M/B9xpfCFHx/7wml+zrXjl8/afWlnpouPfrKBVIu2sqKWq3SCiQu4apr+gVjQX7n0
Be42THu92vDtwxuQgI9qMF8h2N6EeEbX6sV9X0vF3uOmQk/2BPZGSl7GLkl8VjWugDAHq8Po6oWP
i2Vd2V9IpOxbZMP+s97eO0JFLK6mDHR9y+b+SKGicMH6Z+EvJT90cBC+qFstfo7Jrt93JZVxQ1Hq
mTTuDEZQ2ECmIqqOVuG1hb2XPOJM4XcRyJY5EaIvURb6TtJvzU0XMOQberstFyhgCKGFb4SegJuR
q4NQjQX0A2W63QLwIZ0Nlg7BJwzcNxU2/XH5MPSzSlSEGmS3cY0uuxER1ONHUavHy4WpsXUBoR39
r56BHU9d/LqPK2OzrZ6+fkqbQhgbBsK/5rr5UxK5zKxw1P+Cft7kYE1n2xwCtsX7wbCYfB3Xl9gt
PbkmjVqO/LvgQ8XjaoNB/TKBEZOT/+naxEUxZEW8FcBalCvAqyKvO2PcrvJBULouRpXP4Sknuozn
OkXa1e1lel4RxqnRZg8ecNqDnzDOwsptXgjDx0M1eE+JBcwxAzmH73rYhmQResKWyt08rj6XaDxN
BEU85CWXCFHUZQVD+w/BTsQZlU8Ubp4gnZflZqkC2nHZBFVWx37nTAqrJPbf7lAFRiIFoDQPn47R
dUIA7LLYVWk2rjl+EnuwsL+R1ED0PZEAknzC1AnvfwbEepBDkyRU5tgZ1ghwKFpec+KMZvxtLY1o
c9BpD2ao0lZzaMzCJy15I2FuUn/i1rQ7iV4vZWkNuSGbtuO5T1QU3xSMSfU9EMpFpwkezaKL/5F9
IFeaaASAq9A/xUz7Rc0QbesSQK2bAh34B6sc1b/IXe+Q6gkyYEwMuifevJDrqIwz58ljlVokBp69
LK7zF4RI4NjZzqiHfQl3gigFsYMhvFdcVmYKVOkmLtNwTA/d5zHvz7HH7vETBC3H1yh82gy2cMEj
x6K4XPwQxHGnCj8PN5qpPaOTPjvWOJ00jCRF96WCtISEpF+i6bCnMvZQe5ftVTksO40Oj/nnuNBf
eoN5tqzrGkeUctLBeUPKRBJDH3iKLOzLlPQsrnH7Nvw5xMr4mMURVgwfAeiuDDeY4zNd1rc0qhVE
yF7TdozrCRh/IeWhhr1t1qJoc7TEtgF7sJS4h50n0Y6+qLIQs0GWiBYkycfSQCqjijfP7P4HLfZM
jqY8ZD0+oqpyT2y1IjQbgVX7Wj2/c70Nsc/Dx/pAXjy/ORhBdxSydqUQMY/RuSk+c2lRmd2oz/Gt
7+MAP3ZeL8NSCeMSj1xwVCGhwz0+jy1N5jfTuNp709KQTV6VK2eM4bnLV/OrMg/R7vesH4P5A93p
NjbZVbSCCuahqSJaRN1SLBXV22LFjSDxGun/67yiFSY/EdqnRmKynd4iqCYZ64kPAIEVItCxJAZE
dox6YFvLywXA/SX7OpIrm2LEvG5h68ArAFq7r5gkdmKOIqGIsWMfs8TsqJQT5olySTBvau6ufWl4
3pOCXwxVTcnvRBx2TyumULEmuTJB8BCUPmIMul/npD8T+Kmv60exiwLXwmR5Hafr0sx1+rv0Y17D
3APVCreHf9Pw/v36HNLH0tfRfB6lX2MpbnX8Gvclm1izon/StjpRQkpMvwxAejAybt2Jv4RPRao0
hdU0N11BUl+N0NPRSwZtMqSeYx3tbCrDYblAzF/8Vfq6FowEUKp3uqt9KO7mbZYDmYPYXW4fxouO
no2qoKHLwGUP92tBHF9jyOXtuMEO4QeUDONo2yhaxrLU7x5xnHKVyioffp/wUJ5Luv3Uwx8+d/Xi
oX9ux7xAgfHRjVudBS7DsIMB35jORAtKGAydC2yrtn3Cbj4PDH9wGQKb6imHoljEvHf65mDepDqL
Kux/nW5bt+/qYFuW6jLWR8kRZN2ODgkCmu+nWt19dwmNQhQ8esp2ZY4eQAYJ9c5wxfYzKFXhtx1z
vAs17OSPWRMM11qdJZ0CVfH99qoyXMzBPLq1Po4/2f46PnABdWmYLGbkF9b3CuHdFd5AYD3tmUZE
49jHuZFI2gBaFgWck2jDdxg/Egk2OfaS1vkENBcGBPZXCI4JjZaYODJM+0YelwT/dME65veywWfU
Ji4j0QA6eapkvLzfdF3ms98Ns2BoKR2DotyOVFk6ErskCzw65vDY+013IKh9e9kUILW+8JLciB5u
vE38Th84EZ2yszVouPrS0LB2ylfd+6Y1UWL+CtnNK5dkXpDnkaeuC7Bggpwg/WP3YcJNQdj+xHqx
y5dqHF8dwzXY8YBl+78agUDLziLa3+aJrcDtOmkFFthuswzyMHzKR8MIvcn7wARAUocrkdaG1uxy
h9ZlahPhAR7rQXs0Iq29h38Tlzj5AqFYDwdEbgxC/jgVaXRSpFV/LqWLR7KDeic/H3zjiVspklFB
ssvju5HbkR1MR5nrhXOa7ZKgAE5WOVc112NscolQP6fSkocSyenzBECo70mD4w2BcUudxnS2V73A
9ImpLGHuhxuponyVDaz/fQTsAEIvo3VVBDfxYUjm6cL8kEcP2wydJpGKGziLCbnZj4oepbTgii/S
EY2/iUYOZuvThKi+cE74J+bEWmNAjZJsoax6azLCByB2GFU//QXMqlsQzmwVQHgH7HkR4FpcGd4a
Vbd7DZUDUZZS1pg/kBb8QCQmlfb0QBFO4mYJqOmuql4Klo+5umqxjEg0qvqBedG31NsG4XFXra5e
fTltwGetlbXBGO5vyT//zI0Wd89AIyHhpqfp028fmaVFp5CcJ623NdwBQ/EEr16GW4arfKUXniPG
JTvNOwBvJ5N6YTRjbJNqqYJ1/gRor7OVy6zSLC8/a90raBtcPFlcqkjzlmD7Nl7tQxSgVj82vZ9D
TN2aEhMMqbAWwvF+Cw+q8WUN6rCHgkzJTtKWifmHpbXNYohanhLBznYKzYBvngeOM6MCuhtXiYyl
J4K34IRqpfoWKQ4GwuW0WT0Y3UpiWmSBTOXasI7G0FT8Fp2F+AQ3ZSXtZLwSzLray+Aix1ZKSThE
OLr9sNJUBE8V9EOUpsE74WTzzEqwcQPJYaXClbsS6q8J3s7xZPqAI5rpD0w834pMSNv2LOjrK6EX
Wls/ni3vu0jtnP6NOhxIJX2FzgfwgHNc4Fb/AHtSsuuu1D4y6GBKQ4ZraEOA1FpGzwXD1wnQuYEH
VcNKop7RvDZosp3XSuR+0vLRSpjhC2TQKGNHbXycKe3cyb3mdPHOjtOwYKwCw2kUNH795+8NGcXo
0S2vgb6kAzNJuD6wuAYovDSeXVmBxa/ouYnSjfSJpgyDSp5JGxSYQOOpWtYTIPk2s+86jOJobGic
FDHJ4z7chCiFMpbsPOkFtbeUQBz4EbuFppNGhGyDsnYceJ88Ca+auAqm+D70vAUVUFOC8cuCcCXW
g9kAJcsfJvijDgMHqkMg/hf2wemGqPDjrDcdmWWptLyT+NC4/D2sPV7z93/UEQyTCO7+j1OaouML
2DlKebGoT3L6ybSx8q9whVrcZdkN3u+0cInA5h4I1nq24/i9wsrpUyCrEk3q3mC1xQwG/65v3z4H
F+LOF7QRL5XiRChDV6i/RJzkIp1T6TTTi5sHQwgyuuLVwLow291i85PxIe7MIO3kIJ4Li/lhIk0Y
ydnxDv5nKa8i/ENRFAzvGlrukXp2gkO6AonNsU6E+ybDzTXQ70s5zwi6unqdc3Lh9qiYPhQiCGY0
mMK6hfCc1ThGVi4fOyPj8rc4by5CXAtgCR/5eaYQxlWpl4nhbcVfitBjV6FDB0X4fK8ulf7Hul2t
+EcrI8masp8CVbXVdUZdkEfvJQn3Obg89qHZFdesqQUSm4uZ8eWHG4qxBd4U7DSzIrKu9PqUv2jR
GR2nTquYD/rjoD2JwrqmXn/30kL6kXmc8d/GJEryjYVBRryx9IWzZP2FShsE9c0OF7T1qcp8jeBx
TKUm+tPF8bUpt5d3awH3bjp6JXrx4a4KSOPzLwDLeZhh3AwhMQoL6jOPQovouCjHG0D9cgKhXkL4
fBLHjUlf+9HmpDMkEhmJ9+HIBGEnpRPMSC58CaicxoKhekmt/MqFWXkw4GJ1MqudfI2EYh45iysZ
z2GMDRc2UdI5sKw8p2pO1QlJ2h/JXoAW7uq3R/vJD+mXdaAhBNy54OaHBkZrTXuOUsta2VsY1uh+
N96CBxTdO4e3jwuYHS7zyg9gTukYCKtgrpEyAzustSQUKLvlwQw5JmuwT/TvtFC7dLRsnCZPm2X6
dfLPVZzQ3nzlyLhFI6W6MsWmqe8yAXFgU5cfRmN6rdVznxlyBHudM2zGuZQCPEXz9fsSK+G87ibR
t7uQ3Vd0vAauRnyVtq61839NfJaFFBi3el9e1he1IkaO9yVtjruRAda18ZAX6WJdpUf7mYALD+Nd
ueJo2AX8KXpSn0JxXHIcQOH8ajW078FeL8LUc04v91MbWeTNP5fAjQ97E4XbvI0H+EDdNsJEcnFo
XD3n7UGvLnU1H2Ms7NhEyuNheHst3MisJOeX3qKtqhmlgNuUGnDRjG1V5OAYq9bgTfqBYMQYT8e+
LRTQS40UAorKseCZL4/uvyLFgZAhtnmhNDObetSWUeGN6ZN2XeoJvTqo9I8aDkjsqK3UMMHsKo50
s3fgEL4pbE21dhoF4MvUsVakH7f1RRkRxeexqGOcjCZi1/uggvyPPJJI6zfpqmvJykADjqjIAvK3
uWKROSgC4uYVligqKIiwUuoNzhVGrcuhafbF8Rp60wl6f6PnkROtuI7o14yoklxXSqLPZhwjdGgt
7YokQIrJbNK4Nae5RgWrq6wlCGlCu8YqccUspVXFrJHOfaoVtLPpx6FaA3P1BHteTEUe5SqY1QhT
aX/KVVKeWpJ7kSPv8spYMRWlkBMH6QUvH8HTLsls4b9YURz8Zlku5/2qkSilj5hH2W6oADPOERKU
mtwi50rSldUNdsnopE+AgpnOCs4nHblEuDDWsvSdfYDQrfzWn9vtOCbk3bGEDhEyGlzSvInpIifi
HQXL2hHLvtXEPZ1vnVcNZp5kmM+/z+15uI1TOYplvR8M6Bx1hDeB85JYQKVM36M8kC+VmYJmjl6X
d2IKtyqX14ZEcMo2Z14aQFO3fIUryFYfkW+Q6pVck7cxuDH9DwdjbWjrW32XB7XVJDpR5+R5iLiI
E42eXNmSvcoIuQPdLtsS9MMT+34mYHIvwNb7sc5lzWnoGb+Ms72mhCwIZxJsZ716LgyJobwwHYzN
ceBZWCJIi/cMwifMIvqdmdc9t1PTXE0m3CR+SkcQ53RFkbQhWHUdzcPntmuQPVkdumTX+FQ17CFn
cAIC9+F5hBl8WLiRpqP25Lo94BSJmEssJb3fbufdu8XquYaGLEYvcM2RSKWj3LIZBZgdkdeaCLdo
HjjRkNB2icqINx3OLwHmhvEeEuv4uLWmdHdzoR+w/kmlaIQZ6DNwDMyMA9UOgwqIEyNRpCqeoxLn
96G7Q3TF15MAeaQq1QESvQl2I5rsDQ7sMavBEZV+KL3vfl8Axjk/WFRkutMTz7VK74OhydV06XnO
iX3U105NiqI/S7PyorOSk4vtDIWxGDM8Cs4qcu76f4z5mXQ/RvJtsxN8q84FZXANEV1pRlGePPSC
we+d5rdXvgzNVkzyoe9evQFUaKwiYVUuc9GBtjtpMiQVQ3DRISNQmj6yPglikHVQpOvn+B0jaV4G
laTx8ighNr8/Fo+yX4gysTy8bTCitsOoV3ANFGNG9EpfVaKAweuxwVq28TbKyXRBFQ4RitVwe9Ie
mq2DyW5ApJYX8PNa2sjk4BF8RwPA/JOMVLfsMtENvsh3Q4/jcNHje9fyDZW6zg16Vwu6El18BAiG
9jZipYc8NV+i2G5qCPJuTKxhl3+yXNXWnucbztk9vBbSd/TT3nr8O7DcXsR362Ll4eAaWqSZT3Kl
RoujaO/cR76hZjVAF7TgpGWSG+hHg8/HVI0DZY9yGNo9Ed1oo+t6b4el1/X4ocjS1VsPYV7y5YBS
h2FM8y7Haid1i5z7MvjsgkqNunoeGQ6c8uGPF7OpRQPVwlMAgtCssfPx1kUQKInPEXl7JPmGebpI
Medy9rH+UGfh2mdWpqK9Nt0gfzfIWnAfXRaPcoFy1N+erc0rhmjNT4JOfUk5i8qHQaFv8gPMGDqm
vw0u5RTEGWfIA92v3kDHC7H0gDB5H+X2cOM4WNLiq+lX6s5RKyk3CHRsGkTK7F5q8PdrBe1dfWWt
gIkYs5tJufrL7duVoUJW9/7IYtfnpth8eKWMCTxRif1njOquPsgQtjbAYV5lYUbd5SR5CTZ4Ro7A
+StEIqMZbbDKuAy252JavzuZbgZjEZ1ixBghJjfDWGhxmW7xMkSqbXJCTeQ3JEfGf0hQkC8Ua5vj
wDt6x11rckRDxAqcQxDCM7aY8NrVX/5tQawKc24xYmaP/v+naD2UxkGsGfcbonY+zdWr107LWXR2
aQ2s66PhCGK0Dj7O3tOD/RBCqxfZm6CrIAvqAeN3YmY2VDZZ9zZwAF4yFAF2kS81dqJEFr75luKy
IrdRwTGKcRZMVOjedFgK0aJOjKfnBr0+68L4fi6LwpHI6c0MOX4NfA3YMXHkspzU6j2r9+pS+Fzp
XG5rZhXkniX+tjhVWxryqC8eARvtSfsEYoXutubdbBSRASnzEBGp4YPDyV3nIQPunAdMH1GbuZun
fTirVPHbUxZX5LjpvBZhcGs9MrJ2LXVpnwl/ny4guei+MKaDaA7TLIF9J2FSKY1NMYw+fgoaCOW7
dg2k7RbznZBIbqHfAwS0o5zHANj6LaJN9ilL9Reo0RWcXBw844j8of/Vl+C/PQg0wku8uY3uzUya
98qXwt6iOTOLnDzaUZ5Sv7dyQkPmnyfbTTVpWfliiDxSwWSSPfrxyXmc8xLw1rw9aS6ejwsY3OgI
sB0LzuRh3szWnfSs7naKaSty6YPIlqsn4eagMMRZR9q6ZmhZnuySda7/HeOTeWvEw4jgZOcqBD2N
u3COPvcQEEwkK7ym4z7Rw+2GJPr9G4vm/OBr8rbW6ebOkCF1ezDmRnqeC5H/x6yqaZ1wHEhcwFQo
Q8cg56qOtwwCjppzqJlJ7wIV1WApJZ5i0erU0VwXbRGzg+Kg1aXbJsEajV4ozEStKFhPwfYnVZ9H
FKfr2XYiR/q/oO/wmTznf0uPCsLCaEuoLM5jDwtUv921bx6Nd7ipjkNCy5Fq256XrPACK6PkbIOS
xeUrXDUjbU2UraFDcV2XtbFLYKot+7OdwbRiSZJzmlXwQugYvdXgrtjeAakNIPQrm4TPDtp59goA
yfexi2Mf0Ga3nfXaSHSt8gOclzcQGDHiOh8GyFKaIq2rPaiULUtVOWvnA3ct8E/XAePo/jAjXFLZ
43gLL3fAIQ0jB717Sr3Du+JufIRA2J0XgeVbOnb2p10UQ+2dqoggrMlxFXaIJcR08n+hcf9onSA6
c1UAiroDQvC3W6itdmaw87C8ASBIJLNgaJn6BhuG6zmAvuzBz/2Ec0QMRrgjof0a9u2UqyY4PnkB
fID0aesun4n40v8qKKEi24utzosTLA7ARD7vDUxH4rtYzEXHFXKVbJjPUndC4D5P8j3S2CvQNkv9
ivR5WuIiQxreyK8rdLmcZcMkOwicXMhlLReeG+hjuGG8G2JLfL5PVawCWWKQORUwOfU1DG1tPkOo
ECpRlAMbfOdY3E1YzWQlKo2w3XkUVxbzdkbiT5fQoZjP8b32qpcSQkebJD4CPQfDbyecrzcqBs6r
eQ+qfjpyurDJ6XafyXWeY4hZbcLMEO18FLk1js0ZRifNo+LsC+VJfCx8UJDODfPfrCuuYlE/Ach3
NXbGrqCFrXRZRos3QwwJZWozc4tu5XR7nR8bwmxRp7zVdwr+ftgEmfpCz5qp+sm9GYehvXpbzxxJ
FRIRk4tF8D1UULopyraS9bugi0MYaBOMCqGhXRuL3Pt2rfM0o3HFpM0o8jwIAA6WtRBOHWEEBRNW
y+q8UG1WgTkJ7/y+s6s3s0kzkPfr5Dhjuhjw/lDIJgUWULmcaf0/VYtIcIOaYC8aUqm9+exytqoi
HLasfwJ97KL2ha7kUebPZIp46MO2Tl1cuSOS0fZiGf3rvPETjsAhSSMEK87OgDiPDODDdcV+U+Qc
MMMUBX2fzsEUp+M1lR4T9RqXKtLv2l+VO8JmiA5bCspb/ZuMFQ8OsuXG7R81BhVTi99NAzBMGfb5
8XlKZbIVfeUJHN13g0Q0gA6h83M+BLdV3f9qq+HewzC1sfpOGu4w/8ssg0poaAQpsRtjIGI++vou
lMk82mMuszbVIxXIP+VzMOhYQHwHkGYbugQd1beqVfR24UFFfe1pvHpkmBE7xn/AtF1eQUrVJR6i
VKnV7ZETrrxSDTpMuB2r7MNiGNH8h1yowQ2L4k2Gm6+3voUQxXEwLEiqM+aZhd+ENF/o6XXXz07J
LGmRxuXqUghEYg0x3YcmmkHbhSZEjgJS8W1+Mglv2FErQOt0yx7ztSTcBr2zMo54pLCPXZJI1rwu
35A9Rvfqj+s6+NtemcADETDMcM7GC/a0TziLUaIix2NBs95918w3vhZCIqtcQBZL1FR8b+skxqlv
BmsK87qEWVEPgPIbtw/UrG3xURgfvjugesAcXISqH3J9/esdrbgJv9/KD4eEAT4jEV9XM9LIo73J
U9C5BffiYrK9Eshn3BpbEcTEHwWwZi0ABgehV3DSzEdH7y5CVgFKUlyiShWlFZksPZ5COQ8xA9od
fU6TMc6gY9X00hRlOUGMmN2yXzrnkLasGiPc2+/Kymp3Ob4i927C7917n29dqlI4v4VITG5F+jBl
jbcW81TxYaOIsEO42S0inYfdZx1s9bjMYDVyzICYM8gi7m1EfjCb9bMCjkWleOiosKVnyJglB1LV
0iiL9hc2bTvbc61+i9oARK1CpT4BCFL3PqKNKgSYB3VzmG2NMEsxKoZ44GkK6vDhl7g31PcNnzGX
GjRJ0p+CBjLttynhA7s0YZuVMOvBbYtbwwWAStnx6tXVlG8RTs8wmaMSofssNtFsgVmcAU2vOF5b
O6xpjURUAnDoUGlooF0L7D77bod9scbp+s1OAI7dQeiaE68sBbI0t31hdkAKVZabDG9/eWzRlZb7
nKZoxUPGY7j+cW7v2qODJibJhdeB8W5VYrZcRW7C+7mb3f73C+n02FbJOhDBg/9+XT8AecXPWfjM
NbEZ1GBNQ7qgxhSkLTNYlFDxSb73Ee1gptmkzvD0FognvkKanvqSA2b5ZBuwcDxAw1H0uSsMSq+4
7GJm6r58ddN3nu0cM9t9JrheLLcFio1Lf1YMdkGnKAmf+9lAlriTRiYHR6HWmnRbceWfsAWpz/Ts
nzdMC2XvTbjdCMerHJkUrmW7IeOiCAuijwrhY8vqXR3MojAxSr6FrcPUpHyHooygpMapbb1/tSDP
+wQwUoI3dN/EFjGDidzqauCwf5LNTb0Him9itqbM3p1C6RYOMLc373lfOlpx/Oig2W54aXOnb6H+
jcNPKu3/UnZLn5ac+J6/sJN9nnA3kMnYRdsJHDC/azsuLbYkjDwmPLOLJQseTzUT7b3yH/KMYhbS
rmP7tbLgBtKQXYX71ztqKQYu402jHeWi+gwFiUMp1DFVmZPPgkZNQspZqK4OCE13xcf67avAcA+Y
onNglZvpXac+mDnqFTAm6ruQFhiIzdoGJGRXaHNZQ3L6S00hJe4/NpS2FvtKavTR3mq1yygtU7se
XmEjPPhcyRcDw4Nh8JSSykl0WVObwNLLg5IDhBkMBlz5WqMzWv0up42x4g6xgUIqxN/fxbLjoSkS
f4krw44AyQbppUeCKDW1bYr2hdqX6kgq9FL24Jfa6yP+BG6i5L/TK3x3GWTmQYXeP2bHRVRrQOfe
VZmANpvMSlxqQNUqaQPxqPbBu+/yIuFagUbiKGJnC3db5bKSkxgaojBA3F2ebJpV+7tKBM7nyai+
4jqXyIuVhVhBDCtSpRKCCvFkfhxIJADzS5ihJQF1aP23AvyS97yN4qSH8rhMpwlUnrvOwx04xjEK
OsCVLtR/XjnBDis9q6BdAjANz87UJU1unMq4UA7bqarfo/9kf/N6k+5KY/psVkwf+A8+GUJRPED5
KkAVCkk1qvshXnTZ6yAW+JwNJ+XAanOwV0MKHxuY4n+zUlktdv2qQopv5f1C1EyZg/DuCrcRTopN
oOyGhizy4VZiwAm9PZScAdZYtfa/yAZIBUujXOt4rAo1qEVrrKWlyR8isNuclec70P5I/vJs00Ts
1mUMwGJ7qNpudB6PIRAOavdUGi6GZtPfHyIt0XbWs+mOpvfzEEoqb6nfv7zvEQbn89xr3ct5kLEf
AEBVO/TYLW9QfEbp9PG20uKYfQVHKmX+8T7wghnn3FXoMfBIm2e/Dvup6i3VSpH/mA85B5VG0/Cu
muZsBe0mxcUXpV9ycghZIrUgMsK7HUCHiuv5XBeUsSCcaI/blcGGDzbS1Z4LRr0l1ta3U+vpyMBU
1dVV9xZu7ymo+LKIm7Q0bIFzYkGxWthDfbRryzmRre54bHXxG2gM6CKBN/QE+1IKNtvVw9HyWtec
U3UumZTlGLpJ86yfRoBRnlOxd0RHBZ/gHaSWJGO5AcELr0SrxdJdRG+4qm86A34WeduWpoB4QMMr
uYPph1feAi/qzcToO0kzHMfSUCyhdFaPX7nsAU6ZzeUV9Gq1hdYRLOIKeFm+ET+Gm7yHWdPrwIFr
kwA5QhWLXKpSw9wQwLZ0iM6OK9RB6YIUNa9U0yJZzrXuXjGXeeU9WhTh794iCpOYclYhh5JxicZY
RUPytd8+lek83slT+KNrAyjDBZpEt2of/jv6OCe/u+9lpgAJNvTg4dRzDvtXdmxFMsjJpBeTHKGp
Tf+qZh0r2aUwYkZxBsH2rXJhkf1Fs60Lawl14N/rBTGJmjPysnJqZKsVL4fB6Nz9msRp20Cwh/+X
l/U85E9h1pY752vqWfThCs5XpCxm+L80OwZDqoSDCW8PcTbjDT+GbajzbCLl64quVhdoaZdHCAbQ
R7xV3ApuHbs7nxGpMJnKvTj+5MRyng0EIU+w4i8xY6Y9oWZXCMwFHFcKB5VTOpGfh5IJpNJPBstT
4kD/SMmpbben8bwwUAfXEqf317//2Ru/XP9nMwjaLTwSQgNp4wvOdyv09+89CCxJD0zrI+T23qVy
rT1dPkbMx51erJ3RlyNlE84DZ2IFsDgSpvJEAPxUnWoANg9J4WkFyuN86aJJ/SnSFpbB/huc4JqU
ORnr/mG7b67n364RIpIIy6BAF0QgD+hCwAwefRT9hUvhFO83b2h4amhl7yH7nGT0K4q9pcoxUpps
zw44nZMj9WeAz8WZrUvsqVaRj6WIFj3xO5kBnl2Xk6euZ03gXCCSYaiTJWxLeMB+6+mXjtyLL8AU
c3iaV4/bjZ6oUbATaijCe+vyI9lCeXIKuuNsoU1aHQuO824uXy/EQOO2rd+xW3pDgAYGINw77be5
gBqgb7G0DANBomWhQ3MoJFudhmbsjKEPWptzEF6qxifwudvxil/UpUNeklEcrBNmsySQuDH1g1nk
EJkNKFS2/Ev6wBHR7pWgwq+GIboUpDibtFpS6DlGgh/76nq784TzzRN81Kk4eoy+m16PJM6bUB+x
UI6U6bbdBxNaWgFo69Lz7S7R0oUk79AlmvlLLYh7P9yTPTSm5GAJOntV/LaB3YzIdbXn8/C4BLra
G2emUsIiNRGZzhC6qo2nuUsNF9qKO4BOEZ9AkxA8jatl/oF0+35yAWlZmk1MpNoGLcy2aY4R0rL6
qyAt3DlhE8ladOS3cQBw6od4z1SgZnCiZ0RJrkyFBPlzECMfTtpI12dKsNVKk+ghzTkPelApktBz
S7Z38ouqWDyfvo9oT0qmJr4gag1hNyzAHrCam1aL/nFNn59zhHrvGLSfcyeNSe2B9jCbQzF9Wn1t
BmEN
`protect end_protected
