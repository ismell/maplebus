`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fpLVXmHUjNZYaHG83u/TeuNWOSz6lkSIauGdrAhwbr2dJ4fecXpc3GWO6skA5m0g/ifDpYiKnHkb
M7uwMlgcLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R0HmhDgUaVKY/vnP0VYPBqVPAM4D7HubyCyc4cq3IQ+82/x6FCXxTxqgUIWi+cADNskY6Zd/LJPo
OGERgXEaWxaECtcR5nNM6juCSUKoatv2fXui86uocluAEwiE8keRK3MDn8hF9JYgDVaZ08gAp/5r
TUVejTgQZlASVg0V0s8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qh+P4zwUHmB92dq9eyV3fQsewyiB1qCB4MaD7V1y4PukTjMaNMLi6fRZrxWIkjqhqCLoe5ixShrD
eIJzP7w34ulNXkSJ9wCaG9ggcLwpVxWmy3JOLpCPjDskIUrd2ouCHC6vIB/FOZ/GigeYgSoSZJ+E
8acTDiRJwjtcNfGBE6bgomgU0qwWvo9TsCj8r0Kg0oZlVSbGUdubrBRi9qATpdwBptMQRHunT+Sn
IvTqy+nqSfgEkIjplJn9eSjmcFVljeTQNCkCaB/m54FO/iM/+QeVnLKG4WSJvgWE8oX8E94jA191
vyE0MvHC1JFxVZEVoh3oyCIv1QfE3AvkBuvOYA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tOkpeUSanlCu73mPmCZkdlzsKrAItQbA1AemEJgZrVD3/awbVG6J26coX1nn7AirzzA3ILmnCgCh
+CXSCMsthBO0sNdDfx4gVT6Cs11W+eO9OqDBT0L4EqaPK/QzRXXcinFsg92GoZeOsidLiSZmMkqv
cb0G8Knjjy6Yd/agz5g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CBq8V9tNozEnv8P1RwyL4lVr6+OFNwoVinywVPoMQfcGqDFlBStuWb9KLW/u4FpUVQ41F+qTggqR
cug9ubtRJecS6G2I7+XLQemrvIzPNesE65y4XHMzRWJ6MXFjaqkdTouPWbwnna8ejO7jy2DHgItA
GkHtb2MtbnSgwiDe31AAPaKy1Q2s8Yv1+7HQK0jTCeT31cjBRXGflhaZ7EAr5K/WoQgYaVmoZ5vQ
+hcC/AvuuLkyC+iJj6QECrT3YfIa1hQwNeSbJhpHuNy9qNTYJNBET6Pz9cTf4eJnk2VdEif9vtD1
XACp1SfcHr2k3CvR7IE/R6ZBtgIewr7ITq5Zig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52624)
`protect data_block
oOtHYrKEhLvCrRvtxdI4rjJWPavgBfRmbNcCW0XIiCpQaAQHxDjbz9UB5Shi+bPo3Rp9uQ87cbET
11WDYPSBCAXFNEMUn4Qei+m51v4GkZ8OMiCtU7vLZDuCM5e7TOm29Gz7zOWpchL3brwDp3EMxfM/
xrQpktHxohc9PjgdN5lw3WQKg1SD0GbRtTpkAJd7fy5urTpfq8zhCr6QNDUOx7lcLH/aWSapQGaF
SnaT2whE3dswr4ruqP9a6aaBXG0OJjLoy7zgZ1xeemPzHhfmvCwBw8I7k3vg1oDm12oywhwRRg7E
2b46PIloTnpycV335F9zRFOXi8Ze12Mn/DfW8dhJs6aMWMbO0CnFmkjHHgOTr4V4ZdSZECSr2bmB
JDljCSqDYbIHAgd0CobpJN0f03nPdmT1Hf8EI22VL+6Q5eacegRCoPHessfD5hPTiJoPZFgn0ecL
PJrhzNyqXYHNCjA6bPiFfTORBIhUwiyTCAzxT8I1ltiVImAJBg84i4LdQSbQhvbPbhDll5khwKId
kLem1PKLWp1SXOwaIG4n1PVunekWsmSbAmZVGH9ChdyDhSPwl7XIeskFs34yLvTb07shgYchC10/
IInyJn03CgsXWWVkhdw85X4o0UGBLZHyJDp3w689GSjB4rlpPostI7pehGbIPfasfHxNYDgNhhTR
U0WnEpsj6hHAd59bFmp4UIu7sFTaf5aE0+rAbpOuwAvfUcq6DSFPE+daTwgMI/HwRghA+NVSx/DF
58JTiqCqHqZwS9649xxzUsV4/ikgNMfiJ3QQU/8vpJwfwYQ7JMgYMMR11dhSGaczCmrtC6UPDTT+
gmvsVfdwr4igx5C1e7T5fqk30gzOtcmov6UnjFC0swlk4WBB9fF+/vjY6UwAnoLO40bJm9a8Jtx7
Uw5RpSr0TMFQ2bRD7RFc2GtukQDyxNEKUGdeVLQUdD9iD0TXJNcJBN481Ta7ee6GrXFTpYxaG82o
kC3AX39MtVxgrP4+viZnWLWw72gmSTPEg6LYKt/7nDC2Ltrp8nOXTO9jeOyoog+A7DE2E6sIvARc
glhBApVMbTH3L76mO8UHs70ZwQ9hWSLlSvUjncmjUYthBz25e5I3eB5lTFY+zS8fEUwYx/iwba3X
CJbiEeCUzB0I2HiP6yjOuG0uZUNK/PuLaHy0rOpNbGuJLHTHIyDH/J/ZZpFVG98IifGycF0TpF4B
ZSazOVPT0wKQag2dMQzf7XBwUltrVr2v+uY7riJ5HMPm96rXP/JFbgQ5vyLLOO9lpwkytxV1IRCN
BncxjNeq/aPHzoz4QFH4LOUiWijQ0F1jFD91i3OJWKNRyZ/uFxFCHhZfbN4x7DDoI25SEUIG7Upc
YjZ9m+4Sd0wM8AcM2SZIGc0KczNZRtZUd1neXH1dmILOo0oUk/Cz6/pTzqZWgoL68OzKGVaoyhoz
dpCaO59YBBNE4O0gOj2eOFLePXSz+OC/vqzGXuDQlrBMv7h5wlDCnVcnv4mmsu25rSc5bgfAKPL1
v/wiSUpEnPxC+S4qJRYbQWPHqkHeODiZf60j2Oy0nflGmbEp/USfkJP8Jc9fNpFdUmz3a9pKqVJZ
e4DIlpR7bGn9xYmNPckA3YPY7nfQZrTNi0V6LHsqlpI9AGYegMkj1jwIjgJsc9r7pyx4ey9U77ZU
SM17zQjiV2wTxTc9KbaP9QX95/sIWGssfMn7pLK1FFBBz2f5EhyuYcb8OgNwtz9ZNUHVwSONd/hi
7P235wBhsaDcrevHZYNXDaOkGEDGfjtkpcAQbQJOSikQQmN3nW0+VgOnwD28UKVT0TV5sPVNzGOD
axmLWVc+XOV9BgBzcAhAjHLRpijCXp94d0mIRKPeAnD5De/6qPvDmLoTFIVNFNyhSvj8+gsCsvJO
6dhrGZUwCrLzc9pf/x+4fuK1L7XhRvxLebzUdTxcspD3lbl9I3hxw31t7M04ErghMieoV3BOHCTp
qD8fEb5SwSoBm9MciwGFRhLQnIYKwqWd/GtHNlV4oVTjfR2CnPKZZGmOCVOFOx0xY6LdZXIkSPjr
v3vvNwEXo3oQsGa+szg7QyUmCjsEzugnSV6y7mFNNdMEeP4RKwJO+dmH/0J8yYXFO2name8YVupF
7/NMUBJaw5m6V7mUOrLSOchODJ2vHdpbz0AFxHjglNWdVoOzerAIjLH5tyuhZR2es3vzGOI1y7q2
CZndROVMURcFQ8ZYuMqWliTZyeYRQwHsLp3s0wbOsPkDr3psRlJt9aizMk0RqUZ3CY2ii2Nw4Ze1
G0nX3BfW09+oAh1PW+Mw6RfcZARXch/dy9AarI9Cvkj+AVefcnlX7Ns0aZ3vk2/AAqzZXWy/o+zy
VKBvkOYo61yz451hUlv37KNybDhbLtgRVE8c25GNsw5xIlx6oBYem2mswisy55lkMuLKnRSk7vvU
bc6xK+5s4SHeweEHcwu/O4ngGqfvj6/pLcm7mSqsgjJExlHLE7c3EW1NLjzW1yZPUjmw4oz5haLF
BZhYIphIeI+Ox2FH1WX9tjBztTWxwBnp5f7my6RvWiB7ZfBGRRP+5DmyeS4e2vG1jYHfon0GEAxn
mnwQ1ObxuzJNMzpuEe5Zsok5Dnv/XlsYlH0bA8Irwr3hu2XIymqVNB2WyG8XWiaAvrmlVBb/ncDX
DOqQVOmzIm8vq0RslndCpvr4SBkIX9osUWvFaMSTRC0wvy5F6+hRex1hweH4ijzh6z6PGdVvyCcG
vLTb3RBHrXPMRV2KBm41/n6zOy3JbzIzXXPTKMZGTIuyOZMj1sVnY/lzwFStDWRr3+HGfWdynvGN
Te6twq5RoOGRvYi3+NupEW0McIYr6zU2GqMmZoAfqYaZ2BapxcTPoied3YSpTrcCEpVs6NTLTVYC
fRoO7jb/uzxugwNua2lIcxP5IBnXU8saUSHBs9hx729LjqmIOdJL7bqzttv8ua9zmWlLrRj4kDRO
Ro/sYtrsAlbGqZm7ugq1RTA2u8wKR4XRNKS3WSUUuNcVCILHgrGtezHGc2hEm0MNJ9Nkvg0oFynr
DUNjrv7S8vxmDKnzGy+9Gu7VZhpK5kpLHhRru0gYc+c64NzO7TFlJkKFh4oQsF7wWCV936VPGcTN
ntEjZH1xQ8Jg0FbAq1/flz8347OSZ+PVeHy4i+axzCBrH54K3lR/sMqfyh1z65DZ76dhzo3AC5a4
sR1QPmDs7Lp8Q+qNF72ZazGZt1C9JbVi+7pVEvf4cDu0tRu/soXB8UmI7cM8oFCaCGH1G7Wl6LKf
B7X2t8hho8gSgqCH6gKeRMyyc46xxV29G6TxA6nRhHkARTEVODGlWP0qcb5BQj2+XU5WseeL/Uq3
j0/SC/3EPVydfio9a8E5AX52yudzZe2QKQ6OvfPzkRiTpmNx/S0/+z5eEaKtpekQOioseK5mbPOy
ZXoK/TnPHkd9Kx4sLYSLRlATn/ccxOgDGr4C068cM8r0Xo6cQcVvYAWMWAskr6XLvSiMftzeiYmM
HCJ6zNrXyvJgRdc/DmIw8KVSD79JfnDjZZvIpBqzTD/n2WYgZrSnQcB/0y+tm6klw/6kUCOwMR4+
/TAj/Smkc2KMFuTZppLwoym7kyNw2cEWm6B5PU69G8UPtFQVEe8OSM/YDRoW7Vzz37nJm0Seioin
f5HgCn86w+N3ryU+br6Suk2cKGwXKtn07iE3KAU6YUSWjan97GRmmwJo2rVVK0/oKeT2z6xGPotc
OMnuUGJ2N6vOEgQLAhhUefv5XXw+yNHubTz5ytyBVdz9IOFh5NDEB/NBBt1pqjXqtotsJfcvrjs5
vSir+H9dB3MdGHSTQx8DoHDEZz6r9rXQUZoDq58qCuLQtun+cw1N5FjQVlxn3ucI/GuXRr8jPet7
PqUricGUpLHglpSwAkf4X9SGvGqYe7CzLGwk3NYnMCU9/oQ/LOavhz8u2fMN4qaR2OidDqK5Nb4J
0NtLLBpPSNlhxk41WcfO/Vxr9sh5DyVpNS7cbamS9Mwo57SKMUe0T5/hdujb96yp9q8S26jartn8
dshA1D6a7jW9gaNfXKYt9lmqVK9SCfm6CUt3rS9chVPuGMqQedAHN4rf1hhvhIdx1bggdgcytEAC
tnDhqfHHTsX4fOMc+35KFOK7NDCPq9EIOpWvVZMA2vH+1iLDh3DzBrXeCB6QAdJhvNbeUzWn1/Hb
4uVfjLaiwFmP/YBdSfMZjU47jhF0cnMGFcYW3R4GkFAnoWJaCUcFV2Wrn/pOIlJZ1Zo+9PuqcVY5
3+ge2SXK9aSx1K0MIMq4l381R/0ou+udLYgXCWz7DpVOuT5TXp66VJBxW0+w0aoSn1R9w+qX3GOv
utiFHmw0y6Ax7s+q2+STdM2aeJKEmk3bGSvQZF0nhTRzabOtvimWh8lbPPzzGWHV3UAno4ASbeVQ
N6w/U4x2VtrZ/w2nyB7LRcTO69I8GfZn4x8KzihStzBuuUcawB6nwgNWb7isNw2XmkrUFWZK14c4
r/R/QKVjGbHj1y69U0DkhKipKswR7Dk/iv9Rb4gMEIT5UkigrltiOnHfWo6KfjmA1PwjmZijSQum
n2oBdfFdHCIQMeBcuwg/SBQ5PaH2FQGRPZOr4VZsAm8Lee4k9zRzsaeh7izk5fkzDFiCVhpSkI/w
NGcI94PXrC1YvYrw9U6zKwb4jUWkyr5q8vmMPEs+OkH4YUCUDsNnQlpAiLIyF1hfQH6RwZRpZRW/
b7mrkGG2ouVv7WPhCouxNK2t3yBKbbp7rrGnJMR+NJ3VhHOw8JOUooWfFukefq5WqAZmOzWnS71c
ryxpIhxR+1S3IczJkCsAQXdM8i0xWM9E30X+tKYO0oBQ4/udv3dfaqftu+kbusadfam14jo5XWeV
au4v3QxSV4CaNbb/c4qgJI5nF+zzehGBoNEnF+lHKekP3iqRK3ER8G2TE2YvPiO8MFWOE6PT7SZA
q8c2b/emxBVhNpjBFC7nrA4/fSOUY8ZxvyWJvouvOr+wEdN3klEj13UvHmUaT8q/zLIjezJayN6D
hC/NDo+cdj+46xLaCviJ/ycoLObGBzvZ8RZGwWGg5SDv7KYXZPlYC7kF7K61Sn0PaG17n9C5LP/I
RByO85c4DJqqJbnRG6rVnZroSa9A0Dhionk12gvFrVvLDSS8YVd+Zf28uzoXTfPe7FLj1f2JxCI0
6eCUfnOEt2pitpU1aaKsarCbpKislohCLkJBF8/OYiqtntlkf3W4cJCEyU+DziDUob041FN8OGjl
hCIRiDeQMWLXVLzKxLAKUcwn8Bf4Ayi/kPttoa5wzlWfqXlH23smwHRZD3+m4GnYtW901uGSGTEf
G8vXZl+3AHGSPzNTc2THGWHgoX+ZIR5YHh+t5ha51zowSxrACqlv47N63H7d5qwYNt+s+m1QxlBl
q7aP2kWX7eHOzeDcJHbNzYLc+yusGqRU6SB8O4nnh0miBlqQQPv19YL5+6ySnWEUUQdiRFHJXfXi
8ak53MR4v0RdvQmn5JcpkzMWB8K+NkPaY7Ogi/emHneqrpHYCRMCOs1RUDNGO6Hm4A27dmt04sWz
z6bQYVUaOldr6qWQoJx2WPCqObUlSeqbEFvPTrbJcFeyn/LcQbPWxiqLrjRb2locFryWYSWQ+Z4F
5iG8m+WxFSoswql7zfPDSitRNsVHwJvtcNyQ8bzY2HvdSQqCdaOoT6+RQsmFpXHu6d1OF6An7Cen
OBOA3ISz+aHx3DFkavFC6T+ZQAVf1CyWqeMvxEm04PoH+GJzgDRntfRPZKvApG8+/9X3FeLGSijg
ojDWyxtLhYLp/BkuxF+2JtbMNTOfquvRSY+VyLlCkBbkNX4GXe1zNwwu4J24y5z2secUoYVzgwlm
te+xQ+0JF1imGU/GbZkfuSk4YxhIlLgiwmAmfcJTLASoHn/Qc0+mqAPa1KTpSUR5q0ZzWwL4LmIm
mBaZ1nUDUneChEquumPxJUIus8Vuh5uQHliWvH5BXOjixaV07AswDctgj0gf3l69du6pVNr/k/x8
N0XMRGCeCDZFBWZLRf1hUIwHgnBqkG/ciomkhYa4+/LweA+ZSVrJLFaJOVF4XLPmm8+YTD8+GCRW
3cbvCwoqSUW6uKBl+c5dBScA3BcJFLwO5gaycJg8WeTyGfMZiUcsYWzT5k6sWikjtbAb3gdauEDs
Jqukz3Ikaxbyco/SWESBNf3alWfbSP8Uvs6JXiLGMbJ2ajcyCn2k9EdjxHcV9M36da8MaXIM9dlY
8TqsoGu3NYPGdZ9g2AK69wSuiC/h8e/SpZem26NGhjO3UkDVbzsJNJj/dO1U8h0XyXG/KN+E/sW/
vbaxcbgQNi7tFWYYsqEvwOy7sOMH1tkOhrijxgwKG0yf2ElIAM04q33IYK/NDOF5uHN6FHRLNemt
b4NGIFwA11oBOWuuyzLeIah4lLDdXgEW40k/GowtiQFGrBY4FbYyQWF7qtNXWHdHK19aw448a58X
5O228mWFfn0xXPERaQvy9eUTIDDRxFPKr3JsV6aHWms60WH973bUJbv4oYRE3nT0JbbMmbyoqToi
cCqt5B6MMx+b0IrfpSNRGzQHKQfuXs6FWtSVbXr63hRiBVHabAYHEXiAlSgzYuVIlsRjfqwXhFxH
7OhiDRe52HK2XdtQAhwFMFWAgiIvuOl2iVmsvLKIRa5QNhNPazr5zHhqAai9tGkQuCxNHCZU/3pD
nqhsIiMxUlKB7MWnSSrtnMFAxB1V44IgP9a2YDATFqkngz8+DY+WSWsNI+TVg1VQEAqo7zEjpscU
mK4etUzsS69zM5ij/5YLuA0TCQRh4qUViBGYEUgA15i7BYtN2Q+3VBG5s9ozPDWfbr3CSUOUGH7C
59ihDX/U0TuP7aktcwvM5FGvbwxB9lxBX0hispE03F+Jl4Wkjluv3XBy0RrEIi+S9Onqb2wS7LTz
uy9yOJrqYZQVhA1m/zPacD66R/D+wea8ZKGJv5H0cbBd/ZbhfSNlbZdpQx24mm13YmJhvUbDFz2H
m3JL1pNS0N7+f7OHTFC6TJUn5Mi7aED/3Sp14Sglxg6QlGBex5v5Zj9pCJf180sCE9vGAhA0ZhFZ
q5R0T/N4O2e7XaFrXDv3RI2EgbEqfg+hgM+6RxOzy7FKkDj2chbld09otYfNdgsG/0d8M13foP4d
n9nij0+zW8LzSyVtE/fjN+hjFmbBaTbtE8YGR3H8TugBP1WIUweEnNBfXaDuSvVCEfhwFIhNnKuG
g4ETt7o1xqEAB1BX4dVLOizjtL3x6bdMBR0Ge/mgQ68jOqPYMR1jX+sqQ8+8ZKCIzys6dM0c0K47
x7vA3AVRdFyYiY2MBywUQ+883KRpjb1JpUUFzNcUs2KCohCynYF4GzOILlzDWpTttEDSdeCQ3Xmu
qtJCrDz9nZgQR5bnn1WDflbCiKEcvDPrD9+RJEmdverHQMzX5SLkXkFX/yMReGSs317+1iwWTZxG
ysCYgJQAGp1vHGQMvpt6q0p3PExToRE56UT9072TbRk9xxZninc26WZJDLEKCnDYkkraUeC63Cpf
jZOWcwTzzgdiAmhcsup4KTnYdDAte+mfQYEL/dwdKcQgmfop6btJ2JscXl4kmTYjAYBFzuVRxGTK
BmnWfrDVysoKuH7BE1U9+mIKPgR/O+uC40gvjKrYaLVPXqDOTS/Y1B7DTgxWATKN/hkn4FSHBHiU
voddO7VIa+jiCtMmT6bMvA5l/JyDE6MZ5odw6R+4ZTS7RWpvRyXch/4Pa8JHuW0ndTPSos7iSm3q
4L/l+t9q3RKm1JEmnPuGSfx/y+fH7QbjGvthI2obohHmRf0c4mcJPI4VKvP+skRLdj8PCBBiMQvp
X7jzrcp7nNb5thc8OHs/AG1V4oBClCWLORO8HL7mzV5+QLWZ7zoJNsJZ9LnneICPcfrXnmLMHuQQ
KcGpfJSZv69j2N6dM0pWlkK4JcnhIPnOmkvbE1hLig4PA0IlyF6SqXFRvaWFoofvbpdC/gPdn4iZ
OpOC6v7iabkuAVrxNvvQoodXpSieCkZcqoVF87GuRsy7I837yOlNFMyB/NbGzLpedRPr7aG7RFdw
TnuuFyEZ0nsXAlSFc/wFQnSNEtxOqjXYhTERV2aOmV0Q5SMWGiniXou3NMIcMLYjLFeeNQ8YHzYc
RO/LmtN06dCCVeTPAZqGwhFmQ6a6DvaAtc/4br/Ds0fH7Qw7nYHS30QYXxelc7U+Sm/wd7Q7WiKX
WZpsb88AwxLXVJ9uOeDD5x4tcFgLipwgMUxR+BR329tEjUZqjovuhyEK9ArNz334wS756idfahah
ypgEeLY4AmkVBiXzZHb/n4G5TghpVkqcO3A4jkQ03WJkw/CpJD68Pm6SoF/+QwnJW5r3tcEyC8Cx
APs7ZPpXFiQQYf89wb+sSoOTA6AV9ZZa7XHM9Y/Jt+4LlEH7XM61mI2+5HKQbAI422B91r8mvU4H
3YmNdNjBUr7lxmLTWFh/3+6SwV468GrcJO6r8AlE82jxvEqsB5GwRxJ07+GLNZZCr0NRdHrPjJ2V
D7UNuB9za2w2mL4pz3f10qkE3NDsSs6tafwICrnBsHPgNvX5HsvaDf7v1vGpP30qxuvDs7/Vi4YJ
DM7v59wkr16/fUSo1r0pCQ0Hlyz0M9Ew3ut9g62DWhUeVcdEuiHKhxK31bjQQ7ZdtpS3PTYGtsna
AcQo/+W5piX7WzBd1uDgN4TY13M713hJR9Z4IzfdNgMGQYBKbnzUh/DkcNYyJwMuQpLoIpbb2RzT
hQY6my378+pMXb2GhbF5uSDN+IpW008gEWdj5k4AfpJQgY7sC7Cg+m0sTKoajXBAOUW9jFyw5eAC
vgJEfTh+NTIC9Pc/aEVvEQx+0ZB3C0n+0AtqnVgzNu96bKcBGGGzy/+tgTGHKB8qMRgXfBOo42il
xdyWlSW/bx0NdeiRvaf8TY4fR1K6G2G0EDatY2DWVFaLUk15XLzpbrtNMORDrbmmRE+ZWxszW1D1
I7fg4dC1Ann/WNbZRFTz/oTD8qUOQDIS4/saJy3w2H8AW2FsRDzUpGf6rm3W7XbL22dva+QXo0iH
VYQtYOr2J0kKSgDkknU2yfmbgIc7DLhZExzZUVG7EkwpfFSJEaYrEyH6YJ8L017hi5gg6SDaYJb4
JrCoj0RULIcXSnmzC0FqXB7KuxfYcU0nhJgpYisb+9XIbo/M6vHuBGi2omd3/e75GhBnFBojYuzh
LPXvDllnZvo4ArdFfrgF0CS7tKvkWVHOVCjGyE1rgYxUKUinCk09mSQ9vf4SPIGoG5DXlhDG0RDd
U15B1wlHsCH/+MA4qIA0ONfrykREcLfvw0KKmHwf5ovCeOAshkBznJ3kQVzg6PQSE8M403A4UHsF
wOs7DbMUDXN5FixnSthAQn288aoa1LCy8yBcXANYxkC4Lf3e0sEQOWv3LvUx6bJMn4cSg04YRtvF
TFValDTzdtnbNJ4hg3A0KfdVfKYOTjIH8EDwfjNaJ8uXTzetzCf0EK0ScREf5M3q4cre2TpP75LX
QQn022DM+Ee9/oiAh9HupGQqkOrTR448j4VBc5ZfqzrTdaAeuSbfm/buFXcx0P+hX16j1TqB1eag
oDI0xb/Lmt8Z3ij9+dA/y4P56KOZKEi+3gJ0d1iJKvWRUPOzUVUUC8v0PRMru5VhpNB6qOrNcsUs
zNxFK3UfqbmMgaaZJpOBaF0P8WX5iDBp7C2L8u1NV9ks595WrQiJGYg01rJLEaQU81Elx6suAQOL
QZNbkqee/LFajtEqZUeKTQQJuEXaDgjR6sNHcStm8vUaFWywggkWtk9fwGRTCy0slOtjn25YOwY/
J/Nyvsm08/Rq99T9mMrMX+Ndywz4RHLUTkJm/+ooT2nCUJdY8pMF5rbfUbWvQnSwSZ4uQGm2MBDS
+0+ofP5XPfuyyXy+4f0t0/VOTEX4wOslHf50Smkq4GuZp6GXByxtxdAUfHQTWMQcK89rq6EX0IoL
truFcKCMiiIPv7Bz0YSbk2eUww2mxqUDYNHP5T1TufV6ECN2Y8hbk0cmr9bumHrJHuulUM8BxV9l
+pkcmx3eICBXjUNUthnofPQG87fRYHTS8HQFVoWE6gNZM4BGtBxszQ4mBRP0J05B6s5xxcXlROI7
990Kkz8vkwyJb9sRqLjhbIcOk7E3oW2O9qc/p7MuiTLTryLCkhdGLNThbsE5ThPuR7HYKI393Ub+
t5ielgUjVAO4tAZqONc5iA4X3FRJUgQXE30NSe1Lv+CLT6knkeQAxA46XHm4d8MSOkGtQWdOIXzM
OIZhOC0ygaOAdczyrtAKIaNTGeM14biMlDI3Mjmidvh+Xc8Dr6ak0TO3ciX1w02BeAqsGNn9L/zw
o3FvbPVPQST09+4C5J+yEWMd1Uqil/aib3gLru3WyE+hCXOqbuWRyFNsbjHZJJvGr7abOFigzO3k
8eJsRz/IyZvDzWIjoJON49ocatuCxk/v3kG/UiiWV7mJICCjQFX4Uid6LcgXELab2D3OPql81O7M
MLAsrgLLfCk1oXziBSl5xwXy2ik27jdED0MOpzP456yno6tWdTh/wG0eMD9VaqPvtZEIMGK3li2N
wdbowPVX5EmHCJN5YPxEfF87/bGsoVkmWeouYtErtV0WGeX71YsTEuWWFbSORbDuHyLdp5EJvl4E
mPVZjV7ARVCms3dGmZgwL+zahQsibR8xoM+kGQ5jmzWdcWaxXDfVLVw0yi2N5XR9SgU81OExfJ1h
2TMDXNVYnN5LE/cueW/6e5GW6v0XT6eLNJGkvUXZ/OZLcUlCHnzdM20zS7irTQlAHr/kdCNQDx2R
Rsx9X9Ii0mTc01af0tb2dgJ6cpWyyxPwrKvtWxN7hov8A30idyP6scfIGVPUy1UzYE2o4iIcleuP
BGdABUNHPRyDrARL5MdEj/LOxktf6WjnIcJ+0ZGuFzSTIKQALXHRbbki8Q6tWiH+CUQ5Ft3CfDJu
LIB7pjBaGwl4uQtAAdjCocjU4xfAS0KzQiMZW9g088H1cpnTP/mgzYWD2kQ2GXkSyWPvfgu2+i1n
DMYz3ro9XzlvDCYKi3mv/OaWmDmjMGBX2ajj3n5YYQPduWdwenkt3ua6UEL6yq4p3pmZTQuEiPVA
V2p5HYqJkaUOq737vYbi2Nfj+Nq1a88WfZnYGyOqq5N4HnNReZgFX4h5obobSiHfvemp4xD/OfuE
uGKqQeAJzIMS+R+CyQDJ3ctgEdxpLhPF7O0e6NZ2d9XLdvRQRy3he0K1twJxcLXJbnQuENFcdCZw
9NlVsH4kl474sp8i/6kDlj/FznjQ+c8WXP2832MCyfzHaa/zZx4tAOCrfWnkql6oMRpaAJlZ2m10
E6ttZYvS2qmlrFNPhe25cEb9bvW9/X28nl4h4PeM6EZR2EoXPbSQ5cUsN+hmyzau3eciUUTtUSH9
4nDU3lDLG/lPtO0ybxGDgOU6yKg4gVTS/P1V79YlDvjp3WgtHDjMo+I/HTS7U0FOwZoDLT+y1mjh
goyEyk7uINI59ehJyryooVZ9xZfNFWB0zoErhJdJtXIGjwdxvnuGK81fwBWGKPgdr6j39/CPZiOM
QqMdXF8sCWTeKGcrH00WwW8/0TroWw8WjKb6sbQEx/nPqxFpizOm6eRqBuEyLHyj93tjoo3c5rjU
Gc+QG8+n6S8E+qDFOmXTgwL1KgZldNonSnLp+LW+fisbFTPrAEnG1I3J6qRYxkykqn8nImU1jR5s
m8Ei/y2Qa7I6MDTnV1wiJkWW3trg8MIOLZVA7BV7X99Sba1S7rKZEDexiqQJn2mAMiy8p1bDul8p
KhvZXdLaPOPgrHQ/8Lnnx2xoeYaUAzu8uOwYGKaasgOpF2mVCOjYWnhHCy8xtc+9VVLtC31KqE0r
xhkzGRNfnh0Ik9Hz0QxCd38JuGtt0iVqIgb3HE5Sf7dw1v+TMJfNEPHJaKSwo0Lo2DIOitWoIsnl
VGYfe6/KhZo9KnciqWgBoPKiBixu3WP8931bDGiNAz23g67Qjcvn5llrxqbY6ojvrAhSUue/eY3F
q2fk93e1i0AYQalX4ZAuyWb5yFYEBgR/7hDukIycr5qCH6mBdcZT+oRtY9uSG454vuCzaywkAUPl
AflEgZj3TAnBoW9MbXrsB/OkJ9s3sJ8wGtDI1zJNNlpbKjeswkJPMx2RQbXGu2Z/MmbChXZtTjKo
FuNffBR+BUwDvXbG1fRQS1KzEBfl3Q+5dQRXQQtov9x/t/WoEStlm2JXoJyjTPPhQYswFiuMsD4S
Yqnpvj5l6vh0GSVMQ8C6bo1jEKSHDVJewLclvYdbtwqhL/MzF8UTxZOWR04puhkDcRhzQIBGhlIh
1ScbW8Z86bvidXp7OjjoU8Dgl3ZwCU/ElmDbcUa23Zj44NDZ8K6r+HuHakWzg77PiYYzooSznCsp
YrG12QqeCKeQWTBeuk1iuJDNJzeehv+Zrxtro7IrrFJ2qbsNFje5fol6sK7hTc2Fj04sexCN8TG2
f4UUDT6Sh1dmxyvmUfEa6DAwjWdzgTbK3uRXpCvunjtW6yzNUmgVXpHJior0ZBEhlP+T2F/I5mLx
ONlDKu63MaxsO7dPDD5PXvcnFyIcmiDN1QdY6M7C4ApAGJYNdH5jBlhnBiBXQja5XnAZn5l5YBeM
ITksldIsI2lSbtP/lqjAUtRExyMY2j3HvZaolRepfU1+mEP90IY3qNhVG8KnUVHNPpqQBkbQ2tnW
FoAVPw2/QBRNMfvEOZr9rd5sh6AaaFWnAnLkrNqRRAzIrv78cOz5o+SUETN6rkhP6Uhpc/GvXmvR
sV4W4lq95X4DjuQ8guDWOVphXQt52lFi+vjrEg1M4OPB17nYWjwVdAhzk+ucF22RWO0+Awr8gcUv
Z80V22T1BEVxJuXyBU3/gCfO9ce4QYea0/fCPEeLR/fhkiW20Lq7UokdeIHk2ksIVNBOk9sdrBv+
Uvvq8sDNXmt1uGauEq1drQkvWdjn7yGcQJYIjX7I0W58UDCd9yQEYZqs8z3RzafIfcEq6lP2e/mf
dd8djFp20aFnAAg+W2nCJoKhFnchuKT8mnWt36Pn6IeYs+fPFKp3cnNcaH6I1+bRkrrvZC0VyOv8
kfsw9o1XdBzHHk6daXRB0gNp1lOU5J0rHWNO74QGMIIwevKUq3kuRYxpwaw1LNRmMcjPzZZDQnbp
ria2Ol6cPP/xCfx+pgB40AaEbOKuASjrgbtoubY5YbsjHs9DKc/ZIpEsCFrx0ZATz/cse1an3826
hqfGtLvzcYdnqO3p/3F8rFitdzk0xhydGms9HaOz4jIiwQOvmfM+0N/Vy/c0bT/hFl8BiGdu1RNl
1OmYcp+1un3eD45Tqtl00qdGhs+k4ungMy9vXHTGgqOYZiKGfL4OKWPQJ5hceVh6LNQPgkKGXgtp
TmyN7nL4FacZXzphhYmrlsre5hkZ0p4gJVQ9n82eLm5Md5ku781F5VIARTRGH5qknrNYFP4bfxfr
+93XE3SMHK6+9JP5Rc5m7+l10PmDwNEBLf2nftl7H4tcjElZn6J0MAYYvMC7g9oGRgH6fY6aqn06
ZNz2IA4/ZxWwNw5CtW6N071bVfKB4PgrZ8Grn7McaUnK5XLqlX5ejmcgULnw3jWRWg1V1lo4VVZQ
c3j8qNnb/KVoW2UyXMDSibptfSdywo/8vFmXJfK63XiF2398l9Pd2ZGHMs328g4msmWbKf47j401
qjdjHzq/d8MmwvQ38Ml1hkzaqNUMMSTv3MYsS8cKQ/BT/iQC8ttCuWxJumkw5KltpAALnaKkLn+2
u9x70+H7iq8NInvyZiWFy2/UWNGpI6c5iOnCq5vkLCA+skiCQzoMIwmcGvjFwvbJFoVW/V8bzt6B
Y0jWO4QCk+bQj7rT8s3mXCttoPjSi7a86vaWQPlH4ylPSMyCoYk8PYHrCQdOzjGQDKjPaAfgoddV
XP3oHIphDKei/1ugYabOfiyYZANAuNNNYMwNFvAuJw9Z51tXPCvQKTaUBtjOJx+qUpWDUb3QlHqE
7UrdAMGzdzqu34RW+bnl/BAc/NAKJcI1gYe823P0225pme+9gBfTF3iGbkQiOYyeObMg/QAqpFnJ
t9z0qpZJ5sp9hDKtq0BUHPjYV3/efs9JglhAcw5rGYeLerYW42VDgM1THxIu9++6mR1f89hbfH9U
XCFbm9qsMSIv0p6Zu019DkSRGzy9heQP2iOWDIc2GclvQzly9B5M2kqVpvUAIw4Q1h9JkpZnM8YS
5/jOeS1VAFTsUEgnrIhn/jIwa4dsUQrtxuCwq2PQEHIa3KYSWo5ragdGdQP2iOks5P6wlwRsN4ou
4x6RJ6bQbj4wuUBqNwO7Jpm0N9t5S/th1kMMLuiTwTfljXCt4q1U+T6332XenzszQr0Ru5jUUGsV
d5CdCu4y6kgM5mNuxOJMlKa3YrhbIuR9bl3R9bKEWt++fhhNAd+empnDseDTaHM+Ip/u8iMmMlGA
KLDdBomy+4ZZwfypjrt0uH6D9MEByMv7PZTUeKUy+6LtsJHkPxlbUDBd0HkoTyLhHSptxphhJt0z
TJ1jI+VzeIqqSB9/dBQi7iJrpGsA1e0LgxMpx+L1zMdrBqndtU9i7GUfOT6fZmL8QzvgtDm5Sdjj
3vdKO9JyvQEQZrCpEeooFuJ+zyhuZLm3Oocc/xAN4YKQKkSzHDdWtoDPfJdXB/wYKl5ReyBs3AyU
p3t1YlrhSvkvYAQPr1c0ZUmHk3EmlQFPAqL6N5qYCPDlOO698NKEc99qw35fvEdIiVJJBBW/RNmd
M99nQQE6tpVZs+gTdodl32X7FSEvnWxVfUnRFnknTz0HZjaXohz+Gm7bFt76VlbP8WDd6i3LXajF
CxMT4kFecy9fKW6EmGao/LK97aYIlHzu/DMx2A7PkrWJWHLNBd486sBvZlXL+NdPiimUZidSOYod
oF/iSjofjV/bxZ0Rosd4Y1oBg5AD4RzifWkNjOXasQvfDQV5e1T7mlCXOxffb9tfhitFqjR5RJtC
7ENydM2MVTFZ/ogbLdvI2Slm6xXW2En+U2VsA3oDJOsSMRxBpE1iIEGkBIwbsPSjVUm1mNknkg86
ggBp3pP1f63IjWYIYFVb+CY/M0TABOdjGbSyx0uqJkqpTtXCCzytMWu//0RIn2+af61yCRkHxCmA
fetuu2+t4v5WWemJ4vJAZ7dEPEDsis+u6uSDMF9T4z6/YB1WCMCp6s1Mo/KpbB9lPSpHvxaDxL5d
QE/A5aABzkfkprvhdDDv6tGM+E4RkS9kZrYB+sAswu3KmoX8Og3EP950LkFVRchBFdBJ2ENe3nml
X9LxE2H3nCNfuT+aEDW44jvswQb4AyG5Z7xg5TNwbTi7lfEZmQpKq/JehdoCbuulpqHRcTnrs2p5
RgU8J5WFZJw1eYSOYvBs+USsmxdfHQMoPE8OY5E942/gkQY20xAKQc9PmydnU88iRx+Z27INtKy9
50YFjjdWyYzDJGJ4AIIfFo0uKAdf/B5CzVETHSSDnBN5zbW57rtiGC9YW9IgB4aF2pxuJIPgMX05
h4o86+1dp7gKXfSYqyjVLkyi6dyZJZcYtXWokhL9RfxWp32BDiwVcnUgsQAoxDmegUI9FebA/m5V
HePd0KaA3nQ12SYnVFMdglfQdCaFBHqvAGfCisiJWd/j+S/1gYrE5p3j82rD3TTzcverrTkCZXa7
X2TWso17ElUQWf1Ai3yKzcHQorAiKaUh1RstGHz1R2io6BJ2PETr0/x/wmSKq0tykvTJ8DPt2JxW
F9pQOEXg5WEQAr+pOecrXnE+nMnbJpdyfQ83EiGPSsncMInB6u6cOv6nXJM5ytLGaoZElwSVYuVy
TW1Srq7DLlx9uI1es6Kf2iTS+0KtSufvTxJ8xiquILmMFw0EcuIYiAYEO6n11DD0uKkhDC/C1DQs
aZoLMJmlsbvzrt5EdlCY9nHDblpy1hiymXoYxwSf42piJazTXJlIY6Vsj7xUQ/PHuRggBb2G8eDe
PcrlKLL7JlbP2hSf+TMpOR1appI6U4Ve8NQTHkfaS2AkuTA5NrGnYgjZiTCrgOV/QY+Xz0kPL50N
blJDJQeM/CXFOa2HIO7PMZmzcH3X14kVtINcnlI3bANOu9bJsLMGsNa/4dwK70VLKOCh4ajtig+z
onuko8brICjzMoUuP796eVE9j4e1+gJjRoEx9coIl5a44T+uK1FV4GiFyIhp1Wcimv8zLmBcA5lR
+bi5mIbmua1q9WuMeSoiLQ2+ur56rk9xO3+3ft5HiALs9k7tRIPhaoetsqSdh5hk7/5JPNh8OHrM
EDqMjanyJ6KJExTBl0JVuqXXIL17gYJk3brEfC4sPJks4Mir4ThqfDav7LDUc5W9bskKxd9i2Ng8
dk/KKlvxb9i3fFmcBwN3WJZUF/0CU71gCbzAaLCt+etCVWhVVCXacPzEB1GJcTX9Fkh3TNnBJVvM
/VkBTzx4aX07eDRD8NsMa7TkjUlzF82nTZX5D2QWMgUlRUd7yr8kfJyKgPQizlK67E3I4umcXpyQ
ZQs194duMerFQciz5p9Gr0U8dHjCOPwi1QelQHZKqtrhDd4trXYB798LKBTPx37K9VZdzJjzB2DM
deLPzveo91RWpCDcGGtkBbT6Ugh7J4JQI40dnkUXvA/BuebU4M+LYs87tneE5axvf2bP7EowXS/e
yxYy8x+ugW2eV19rZ667M1cCx34BQD2ofdXC+7OYGMGfs5P6lFpdq3IQM6PgOcTKGsLriKYnPhlx
RtlYxwIIMtbrlUH4ifYI4WCkyS7UIAi5AIF8qLwzy8pmJ9lc+o53q9uVZNCGKIHF4o2VAGDp/N+p
p1Ej8TOmCwSPHqi6Uir6Pc1MDSER/ONvFUBu/SaKe7VQkkonjqQ1Ng8ebNkcRjsk3WOvXrMluzuy
2CBxfzjJZG/6AMjJf/F+jxXWrSTBBm7F+YQGoqRH3LaQe2c3U/rVxOF4R7EYJyiXSTrJGHKXvl9Q
3RhqSTsOfDXZNUsg/zSYodJdqym2yLZO8mRUy4I3cmcYI15Ju6vL1Frc0qjO1bu0VcBQpQe7d8zw
GC1lpxRFNDJ83TAi2uB+B/viiA1xJaK/2eE9IymimYRrioDE71uE9nuoRvdW6Je5qtoJ2N6GASZd
xuT3c4jMcd/6sDCb9BJHqt+32tnUVa7t9p1w40+VI0bs9gTEsossuH2iaYL942H6U9zOjunEjNIP
wkGq7d8rqNfRn0SKZ249nYjfHVblGwcglTEr4rYCz3rAyawVRT+Bh3cOKZu8o98Fe61nrQMN6BRG
2UFknYDuKxlXmxqd/kh+6nQuEctFRwUBQo8MUfHARODUrueITgmC7rZJ0gFNEbct+9vd+rzegH9J
beo0+9Vjbiv4z/hflYMiKNhGZ1DpJAaE0Z3QBmpcaqgZYimb9BLkPBCL9q3QRSi/96Y8nEcHxTFZ
VE0TLjsuyUGXpErknmX+GGaz4JXfmaGY2CtilINrc1xv7AnpSRHQuM2wN3qlIHHIJvzc3ewwJ3EM
f832ZCXtAFMkc6aTORxQtKpo/8hccYZ+wZhoMGMTAq366VLbxoKhNqeE8VWIhMi3H8o+Ar7CWP+6
wg8swbaZIM2PtmYLLLSe+m+uoUDOSdeC0js/ps1XYZDhGPKrN14c6IjBYU+ZSMuii8RZCsT9GXEl
qHAalfZPiz4ijdUy0e+On49D/0O72QnN0q3b7N71Gr828ieMU65hrt5daCU0mzXOAZDvN4TH2YjT
bz0yGYQHT4SLqA4B2lj536pXJY7iqerMEDkHGdcEHBV2L09MWooe70FLviGdNXzc30NfuZDFxdxK
ni6jr1whfYA+ensN3UkGynItYiIN71+NGuPcGQd3bWwqbdEwZsyjhdHtpqyeCR8Hv5Jai0+bFZMW
mbPF+5A0dDB7Bla0jMcf/TX9CwtJepE9oC1Gdwmx6x5aUBj7+bqkcXWEpPUszYom22wBRez/KId5
q7Zxr8cF0sfUSgW+OkmhIUhUI/kNFhY9nvulMfcmyjPUBK7CpoDrIaxM1sEyHxhuE4PuOBRk92FH
6ensi3SaAgtyO3EmnX1M5xk1DPj0IoK/lAO866GvOXYfCa1lu3eNRb7GjubPVa8Yapf6luwdAkXh
uzyFVU+UFV5fVEzOiB25K/VBoicYqrSGIZfNGlMnvZJBGctnLsEApONiOwMIvKdVVPL6kif/Dkt8
EHMj/wDpB4KPK0WeEodmymzErQTW+nMRwtJCZh3a4SKUFCGYEXDczDT4QLS8cLu/KEgu/U5G3Abq
MHA7VXaGcgce1u2YRm/MES1pib0pACDkl44+AgCUlL3MEnFpg5wzdAI33tJR8XZ8cgWeL1vyPJjy
T1liohqhmL1StZ/eFXJvYq+vH8gxRBPQsDKEpYZyUruYTmXhGSDdsI48wai8lPVqEFFSP2RJgwFu
8lHKibiRI5JucmSSzP4AP6BJhjP+Dg8wHkpgWwM0qcm9IRtnzTk+M9Gv/GTJd1Y7PJxs4tbIUBvt
AsJcCRKH8wAp+sKJS5xTy5+ADRgYMQk+K/T6qHaYqIvOd50tVp2UXi9haANeywCRBNahm60JbfKr
uGW0Rfm3QZjhCvQu1XARhzJGtWYhsihEG1iJ2/ZxeE4G/Qoa96SoNvw6MK1K9RC2mkmIbS87ZI/Z
ZNnykclxbFST+xvrlSwL1t8pDCiFpnwyBdaeqFjAQJXAIdff3KE9dDG8UnID5Hrt4w2V8sWe1PkL
jJTFpkIO8gXcps4fbbtiJZxHwcERtFdbhmkFZAsPi4XUQoA2FfnUH/YXA51m2Utwlncp0EyHx8QW
r/36yTOkKmrTMjL8YzL5D9Ig3YT7roB2BtZU8LIOS0LE1/VqG23JneEywxXXhs82dKCHemq3+u08
sHUVDAmBq6cdDj6yhE5T/36IqaYxXmsmqIhdmDQougQSF8I+CsEWqh///JCswfKu0GdjKE3+wanB
psb6ARWz04FwscrqFrBfVcszqb55GBIoI4MmHs5S8Ma2L2Ky8u2VJkaqxCCV2lnVEhL6beQoMAd4
D2dysEJf8Fe12YsOpDoN26lTG7PxfRWsndmHfJ5lwLjIVLT3G3w+G3F1ZG+DftIvJuPfqYI6tpLA
oQEagyAoZR/ARMssX3AI93Tw9P6JySJpC0hRgkx4JtWNX0biJocxMHCm7lyZnIUqzxLGxhwdJ7Kj
Dv3TiEPFNZlFcdC6TWxL4DSth49kH7tEnwMsjPtkNcTvyg1ZhEGt5bdHN3LCB/vdpg68PRKfzKud
rjreuwSarvTyXsGCpVGSWfGC9sx/TF6+7mOtox1hteTjBe0KZeNZtNAEFqaUPn4eIJHaPIlLTvel
Nc3f4yGQTRiUUPYMEtHqAYakCClDaLjgqXV1E3fNTnC39AxZyN2OdQsFJmODWnpfYCCTptCdJi5h
XaULX1XAvmDl2oqYR+mDcDtB9UUGz/tBTlwPX9uD7MdbV7q/22K/j/0P+dJPONq0qpNUvJoUN7rX
aNPE1EaPINULYLzi/JYK5YZrOlyE9NfDWn78TxytfLoVd1LUZ+myNCKuvHURDBVbGRbylSqOygQU
m4Z6ls02xYp+YwyGx3C13thh+gGSIuaw7SCLxy0BE0PCAfWon6hBOUr4Ub+mM6UGMmxlQSX6bYDf
s7wabe8pV9wCDZkMrs1ePc+4hH5G2xKZJh8Vxjq3syFZcbHwQUN2UuWN33S7Io/YXeRyhr18ZhS6
qvi2obSZqCftikWqLGQLxgZ1YWO67d29pnE7fzgnkrgQPYBpPVFXMzEQeGTDo29TyzpjwN+1UBbP
d6YLGn4Z55VZfwzvylkL5KbG9v/MqzuyEjxzuDkTtgCWrvcOS8/CdCxZj1Bix/eUyEDNZgrgbsIt
7fOiLJBt+6O7t011+kuWG5KDWF8DCYKsVAqcVYGXWGpOZII2SnPJxw+sm+gxFUMXwRY7hWlypBq/
NlhbrohYZWCOrovrR2y1S2CWILnvcsMYRnFIAk/AqnxBDDmTx7p+p2t+Dq+CGjddcMK9obrs522o
TbkCuOhKvz/8+Z1udOl3ScWCvMWV/aEJ/Jz46vDS1f5+WIeHJXAzOmabI2B2v5c0Zh2sni5wjNFE
02DFJcCHQTNZOYWb9jiwT3KFBsX3jUEs5jSrjkZ9imWa/ZR4CynqkomIZaZmUIh5ffYvZcZnJzcs
2RbfcCSZrsdrSTKfzCGo8/NTxCzc+BDKfntll6jrUlK1EA9BfGvgoAwzyQ4vlpKEqObSZdmqNQ31
OwPqZzqxT3vfRKM3kufdONswClrKLTbZYR1HPbfROKZzoNk+bQgeSwHPv0p4gWTYY135G1xOmnF9
nUbP5X2dHhyhaWw1W01xxrwBNauKp3nsWLASiJJpw41U/5PKgf77z094cnzDYO0Hstp3DP0b0TDl
1TzOAQv3J2guOwbuj2Vfomr5RvZFUh+DaFKUEnZ6CmV6jQ2D47tUpr13ssK/EeR1hsj37r+NJ5Ye
aBVUqovFNYQIPuVWXiVyjs6Wlh/npPa/uwVhqvU+DBGOmgC969uyqqFJ/inXZgWYBlnHfKycj5ax
n3YMtq+rd0UNl7ccM9eYA2XQpIdNoZVdMiUpGl135TBCwWOz07RLcZz6BEMfnAkLUwlCrzAB1eQK
Ix/q344eC7pbGtChWuJmKQuYf9uwj0+BZ0uvOUWhDl4Wtucc7/FHrRrpDuUJ8jfhHfA2dO65bFS+
KdGA+Jmqvgk3ArxAi/Pm0tMlcx39L2xGr6+xeTRZUOBqjWs/T8ngfTp3Z8FyOM8vWiArDiRyw1fK
nL3O2VIzBpvlir8jHQmszd/HTDQovlV4vM45zheYZxHa8MenzCJewfllfMxlcpEz8AbPH66cv84Z
hPrTbcgu3QEhorYig1ReREljf1pEpPBXMa1tEJvwu66HdznTbc42dgXxw261s2RtHknN2uQ6/Sb5
NMoRG4Zyh+7+Mbpp2uuuY6rWrDar3cuK4bM3/YeTwDAubvYgm7xrlqbSTtivk8fiTV+WAeiUfP0O
EmAahdXpJQ88S3U2UMsfHqeovBPAV805P/sLcalqUwiP5aZvXUeuzMOqt5kb/0Y3OP4U5tzOrtlv
nMl0oQ9EoGfnOTECAKjvdkhsMe1E+dL8ceRNrv7wyXcZHOSyHNFx6Dy3a5tAzApBSlukBPMx11wx
2uBdoIDyPrbtpp3+wSRGq//ENOSnRWhfJBQDHm/7ou86xU38U/BQ6j31Cx0+gx7UaqSJXGIvGsCu
ZA9pKtlLGTTfKXbfPRqmxezMzkLwNqiN/oxXuSGQ41UbdZmZu7XVGtqvglUFCFPEWHmtH1eaBkJC
SellCP5ueC6PTM4GdBgN9wquhjkQUiG3b6D7jF2Yd2Q4LPT1DG8aYzdb9RPqlZUFmNu6nFpsLgwI
cbbZmFz3zsgCFirAlDwb5v67y3gUetqV2i1nhDkdXVrigAFM82Zg4SpKOd6TlfMwbpDx1JQjaap9
NonnkSgs8/zPLeDX+X0nJez3mltk2DCQ1QRZ578avqXMDQpky4TitDrEhjZLO1eZN0ceqH995M4O
5jokV26Wfa+vzHqQoJ74+ZmC+OdXjYA0NnMMYcShR93xnlbPal0RX5MX8/e064ViI2NY3dQokRFV
7aC3PsSjqbxAvVH8NbcWBm2dhQwBxfnceK/7/XXbePr9h0eSMo1iHcAvHWnYc00iJgkS4203TCTN
9vLsrAZalwCT+XECeLDqjduPDvuLfCXhVjGd9s0RuhZCq33mA9FQpVe++2UVdZEIqXOfyLshQWYp
eYcjXobl4ZjbqiT4QLYdKQqIG/bRTw4mIf+od2FzBYnqQgbvQh9x0ujWYqqq2bctFwRjFvfpgzkp
5kcqC2nCHjWBfOvfcpNjkXDpi0V/gM+gZJNf0LQ+BpIOJLjax1r6KLFZNWUy4W/ZcfT7+C7ppJtL
wm0LtXys/WDQAZrCsDXKdsah3C/nsQy/DuuklfM3hg4VK43BqZQ/bqsHNOIBpODMReLOoJ5gfbof
7beurPfrY2omgiSTV09C6FExHpGfwVYhpSCZ188OLbNtyHaR2EJwkpJL96HVvoomTiCBQDga1gZz
7mcy97AXBQDwgvvo2SElhpsgsRxxqefEg9qSYc9z6Ih6HZjN3uOV7OcrU/QTH5fum5Wr8EU+yJQR
XE3WKjvD17q/brcT0tl+UBRuXg5s/MPAJDLWX6IGXChQoN3vEXo6emPv2MWYM/V4UwJ53LP1TMIu
JXVF+5uq3zs9Mfi18ybGee9HzkzsZoLvihiknY1FWurwi8bHTIKTVWM2eBGODI2skTcVEM4ID4tb
xjB8PWbKJCtvQKR7/yUwHoOZDLsubxjj6pSGDamLOrv3EfFZg4p5COzLRBa8CZxs09UhDCdcWj71
7zIxnH03qgiQoPONyy5SU34+NhS1XWFA0y8jM7xeMCc+PnCE1caYy2NS9ai/ER028GdvRX56Ir0M
9/WQgGMeEdtRGCfg0VLYsPY2kN45mW/dg2ocPksQwsuGGuiQIaMDWRf+FASrTjEOPqlvbLRJKkiV
k0dj/i6bQ9srWJvn/cMnVgZmFEHIMek7quxxaa0oa4CkoY16ZYwtDMtQgHZ6PXlSqr1CcRHawbAk
x93LrZpFygbAg3KvGVK/yLU72VSw1/EKYVVwcJt3oOCmh1ew8f9N7Dwx3UlyO0dgsVNHWZ9ZPr5M
XHSfvX6dDauNRcdHcCJbaEettzAwVxWqp2Jx2UrNi23r1UJnMZnUU7LZeYEwKpBqhox7FVHldCG/
pAqIxNfjjL5MTFu+a+kpHqcAYHyaSdOGUYFcKcAa4RexiTUbnDcy5lPNHtSGJHf9I1ihdwTWVzmf
vomo4JSsHI+gRlqfOBO0YL89IfIHntPyy3eIRoFCBolEa7N7vPTdYA5RucUX3Ysep5bupqo11gC/
HwlTz7ulLEb5HH14LcBsjmjk8Oj5KSpYF7RBrAPeN7iTJ5hn1Pc7wJMRLN42ySD+JYP/8J5IjRQz
nlrjKKbNkZJVNGbuqZiAtIbfKpLbiGAAC2urinQ9d8czJVZM0uAeruMao0xp3K6rW6jWGuPLw1Ny
HHI7TQTSd9Pu7VV58TY30AJqOY2I13XyWw/lyeAJQbJ+S7Xsw/cub/0KqOxfjhunrgikBNpph/6e
iuH2TCRAYfJIP5CwY0mlzn46/EzczR0v7HC8oha+hUh0hUJ1SKOzr+jMxiL2bFWmzgxkgMhgjBfU
7uhnbKvxI5ZguQ01eR2nTEJv3phCjdkptHlbnpbQ9dDxho3jlqnWI8+/mAgOvxyE0KA58HBOB6tI
IW0sxCnxZWO89KpBUp204Fyv74wIygKRPtjix9g/DX0Ho+Nrkh60Zfej6vM/0r2rBFraZEXaZGvF
8n3x9jHYz58QYbZVOkXePrY3lT1g/eliIDWHxfTLcLGE5x0//6gj5Y0aemHacfSnX1dMeF/vF0+7
mBaxjhZw91E2OMPddF3n22f0WvDQm3TkqZ6I7fvu/eaJsSJFQYFrVVxW6y774H9g2OsSjefPQZri
LAqUnNaKhcwNj8cFnDumsYu45FUsDVnP0KzmkPJnE/GIhkZeVi6ixRMGlzmatnea40FANnGh+VoU
4flcKKuA0QADD64gDD8E6hKm2lCQNRb/v24hLKFxBjqAmmkf5nrRcpZcluxEY+b4MdNKIZZgYHyK
sAcsCXwJAqdXmdjM38F+UVgHosSYP8RSYAf+gTxa6RXEuE7ZMz+sM8LfroAjhs0e9aOhHAWT7k/F
4ud/ojxkv8gaFSIO+gcin15GPCBFitLgbGmGPAWTrYZW/QPD+r559hTjqMIDgckB8/JiPbwH3vnk
LwO1cDI7edrzk8Bvzlk2ivH5CHsTtXKAL9kriWadMCoIZoE2ndU0V8jyNekltOW4qICOBdrOfVF1
pEzoo1Fv2VBMK/M9yAEnnZI3wqPKWl8rSxsSqsQ98+VK4RVRmGdWhwBT8XrZppRbEdywzmqKPxTE
/F3S3x0qsKYQ75EYTl2TrErpiknTS4LtCMZv1vhqGBxSrt1r7sriiexjfU7Bo3FxH58wV+pwcqI+
Ks9+LYe2Ngb1fvQDtWpH10QMCbnZPKxVhU4fBqW8nP83tVy4rRDpPaLTBBDIQNwgFiU+YMpDGL0R
8ataBfTrdJjN/mNIls2yKS23dFl+b81W68Z84TqIbI7qSnyay6waQ4c8TYnmnKSO2X7aIZ3arN0b
3vpsl0dXbh4FyozIgKASFAzgyGHve4GIUr1LmUhPWzjPu/NcEZc/YQtOAgwmLMMNy0m+s6jXVm72
wmhosK1MeTuQfIlT5XGIpAi6tpDr5jfE+Uz+OGjvV2vdVeO2qQzmqQ1nHbpTcqEgSHF6ibcmwVZn
sSD5CTBCy/sjYGE8RAZxFq2DlmEWNDrgPJ1fGaNk0N8eTHxCmPGylOtU+4xjmoyGvV0J6jEUmK2t
wdFuH1lGGkWiN9gmv+WNAAcYzpwFDHsm5UpNDThb7wj/5s9MwL0pTyNmCIurxmIyI6PI9ozipXcz
4ZoFvh2qmVogEeicZhARaSCFtA3FkUXDEpjBXS0JuNqTz7r57aDARTfhEqD1+APiI5uxdaByzK59
GQpw7XjY+7GSrliqlFkcZgZ2Z1xF3EkPjO0R5t+VTKHs8/h6MgMQqQAWxIQfE0XYTrvVf/hMSKjN
fVKR8YQ6HUU14hICYqruwUTP+4DlC+F1FQex9sSWOJf08xTIxtzt/1UEtrBOpzB1bb6ynQF71nhE
wl/Bxsx5Rh+F5wGu0RNyNtr0dffnre4/EGag5y8mNNZJya6CNrxl1XdSRjJsqLGwGaZm4MofZ0s9
r3lS4qsktitqKcoqIugGRkd1dIJj6kYRUEHB1QXKltfVwfIXlI0HTnbMwUiO4L5cihQzWRLA0IFJ
VQKZLyy5BgyC46+8aSQifaaNlm0pWiG/t9nfDSAZ8/Pe04wRUcNSSvsArqnC4E6uXYBKHWtFgoRH
zfWazOI00rVTo3+RHKL+aT21OC9xXYVMTqrqKaCDruK3Gf13XVMwv626jbKO3W7ZfopPA79GjVBc
mobYt1OCFJMJ7AktgrBszsihLe63Gg/CA12gUGgxBvUS3uAIOIwFcZcfetSv6DWiw88xhqsXFyBo
K+ADw8Q4/ME+5BSOp6A6j8ztU/cFb4NnwWTsxNl3RrKei4BvRI6pt4zO1F++6Wrg1zKPGqC1910X
LoUUhwBHH/ZsJRiOtSJP1OXZSyxRan4PsTLRNWEztM4BCbQFECWeLNlpOYXaU/6di3yIQRkaDWyp
FvJmSPjSZ57Ef+wWGYrJpnRKFIyoyumvKmj6Ft6oantSE0z5BQVrLt9Mk8teYgNd+Gqw0Z2JxsbQ
nq4wcHtf+DjlZD+UhyKMVDkHMckO0peQEnurf4urPtnYJZag1MX92+XLtd/hHwuql2g8weHeUfcg
xcEV51efQds9Nr6tCw0ot/lN89R0cdT6AeM/uzuHVROPzCdl/fQS0xAkwifPM8TGk2HSrWSAZH/e
EI5WanEEGAQtMC7PL3eem5zAYbCJCfmdxSUGv4oBpceZP0E2wd6fTOhmGJ083DcCC9N/EjlTj39o
HVmBvEAO3xfHbnPQC/Beigsc2fWhdC13PLCOgbxJF+1RHL9qSNqbrtSwqPGJTHZmTl+ySgz+QhAr
ETHyfDQU2e0cOhazunqfO2Tz3QiXX8EfxZ3KtpySzfGahihU2AxTPy9Z2G6a70sFryXnfh5nrhDh
bNXQ+G/JqF6c/7vlQVS8l1sdSZSyLtOcRxJnE9x9Ctvc67DH9l8TMDECSq2Ozli4OQnTZTsl1oSg
Y8SIMpwmq0f44PjrnsaXz4o7asjpO728kGEIvXFxCNtFs96Nyb4NIlN+xH4dibA5g1XVysa6fZhW
fcTvROVbSIAlR6YYc1q0pSTiSGuj8WXBIVLmKoNv4LtPb5t6tonBMLaT6WjPD8jREByLZgStHU3f
e+gGoghsZ6oytiSLWgg67GBo3VBL/nvI8MYyBuQGNzGbdTHKiNnIvN+O9N5DIy7TaaEf9v1oQtkS
354zK5rYtDxdSySBC8AoQRDoHMKq5R2lGAgUuSxuG/rEdFpYXyA+56u9+vXi1xt3Ra6FJVI6yB/+
kXIo7ale0Twl4vCgWdbwedPgCRY309cML3WaSHPgPk8m3C0Lc6qTOIWfKQLzG4gWcqN9eLZYYhWn
2nNxasKHDce/StFeGlfe+RznKaMabWo6h0bUMYJkM0ogi8kVYtkHmPLSyj23YvvA/1kgKqmG/M4A
YcxixRbWSCfkR6+h+ni2QKPTQF+4lHjijwUxsf4gHvYfGtIsuMN+xu/yhi+nLXxJu+aZs5+s5+VD
SMLw9EiOhWAtHU7p5e0cn/IHBdyYz7CIJR+CftzXtjAEEy9KEv5JZKbBf1OGsS/xlOnURwCyd2Qq
fOheV9qWhBNQ+S/4UyAc/z1qDy3lS3KBkPJrE0amO8sLRcYqCcV/+JHexTS982LKn3ghyYHroWzX
XmIg1NZyLpiaD+18vHY+mPyZCe1yFm7EdhERb2tlSHMrBY96UU4RXZpD1K4FboGgsXjfYs5KkiHD
eTZ54xUOJspcI5ZGUYPnsgJf6SdUFIR/xEvAfpwtx5XCHeBnq7dKVuFuMM3yuheFrmsMrKvmI34Q
gc9LWAAqk05/Apdm46jo3Xy4PLd92MevdUrPmfFNPdrO+RhrpD20jW3fjvUMt4KLvBqGJIMZ6nBW
g/ci2a404yb9wNu7aYTKap4AqO4puVu7mOtQCkD7u7rTgwYktRCtA0lI4XiZzS/3LZAQkEIvU8GD
ymdnozr+oABx80jvEfWd0/awa8BclRRCTAwgqqnb6xyKD0z44HOZCfhTw07XuCmaIAyy+zxZTyqS
BiSWukL9ihUgHLvbzY98E3F2Q0TWQrwDhoJK2MeRHzabX7tItiZd9sXzNvCgyIB/aenKhhSVuvpW
btYyT07naUVxwzg6IBDkrUkbL/MM8kR1x1iS8f70kr9rMxhHbNc9NaD2RNOu4lEx6nALGRXEd7at
dOPCQF833o5LtWvnYb+kaapZwrnih3/Ods3YROMZqHmw47FwCOzclc+RpcDIFpTXXnAOakcKUCbM
CsGodPdqvo2y3WllmOjKT1d2rTklKjJ+Eaub/MwivbaXl3iwb/WL6+wWFwLxFLviozKRzBnyrooq
ow1U7oUUM8OKzRldUBXVUfK6GeMulU6wwA2U2UMU6875X4ezISjX+Up8GI+U2Y92xHZni0cl+++3
D7t6QzwAXyPi67cTFQO9WdExmr8AKggnJhjzOer7EdMC6lMDYFgQvkHAppqpH12QIUeSvKY2LDy6
RvumnaucjnmyKDhcSuZ8jpXEeU6bv8s1qdVs68q4PU8/RDRg6CmqmEY8V+LIWmbgbZ10ch5J/Sk+
b92oZi9wfCBw1z1Oh0nwvCGBUFQFXrHdy5AUn4yk3acWzguirJ5Lfb62OGza+i8nR0giXA0q9PPs
vr8smW/cJAk+mry3hpWtoSkAgWgrPSKy1CDavzJRA0b9F4KxyRAA8kTlZmCpag7Odlf+LbwtCCo/
8XGpXSuuo/vyTWv8BK6EjcgkK1FRZDBU6KaMgqOC2nioTuoANg0B5IvU6kFszdoxx9ML46FapEX3
fob3MuHo7RSAlE/bXRUP5ietVjRCayUUjHQLTrzZ29CWUhA3VADdm969lC3b1cQvNl35COV2yceZ
I7vLDB4fWrpYl0icli2yz3UmhgF4Z/sxPRhxwpNUWSCGqlyB1HTO1xpoobOVOjPTviYqRHaTfMiy
m9jbvfkdDUDZEbHdnhx6C2TOOWwE8BNacIvyS3OtuikMYqsAqOxRru7aYPsR5MwHlLK0Yts5xrVI
7N78rh0KWbsmfG6iFv2jDL6k14bhSIa1lh9Ozi6Lhhcf2kE2RLrjhFV3Kp8ZcpeKV5OgUUlmYEoo
QiRfOLxEqgS1IYOqQ353bonrzrLkJPSNPLKs4QFeynVm/hsnUOvw+KTcSjxC21mb+8GEF8XGlYvd
X7BZDVMR4oTAkt50kvKXgmnZexk/UjTfjFgn4cmNUKZb8rrmdFtRGcG+psVGPEAxfR94TO6OBBKa
PzTfIJeqAvrXEormO/yQxe/DQx/qMdj+c0tbIHa2/00ZTaRimNcfHHSvVe9G0BfQo6m94UNG+RV0
aLzqSqjNQ0q7v/j3tew5XF+ZJ77pnqkZ3fAHq1/KXBX+QuC+zRt4K0XbVLL2FmRuwEGtG4YU3OfQ
8MqXtjGT40lJ5HMm7L+GAK/Chc/HcDzGjKsADfdzbjE3nn/F9AV3L1vIO+Yadr3cmnESXrPbuK2c
iAfLFlMlciEvUzcfhBdJKQ10fXfDC/TCLaR23qF/YtGreSkfuw0ym9POG8VFuyuNB4HJIdAC950J
9VlypRgu/4f3JvE59RcDLXU6jFWRB7sFf993ahgXZP+SuhdSrka6lMGm/e3+A4sF824kCPi5l/os
m5sefpIOHqOy5m8ToaORJM1vYJrYw+RU5D4GgguoYlULRaPM0i6uMLN1oDrVAKxbsxleZbaD8dp0
aBn9hKvTi9pY1drOQRAMc7BkEzTO/fY3hB6PAqwCTMEKyQ+PecyweDG9jI78ueSiffXIYvNVlDL1
sOWxNTzF60hX6Dc4Omj5mXR5TIBm+8SJXmxaDiG6q8/2LFZwjmIGMBxviWaoi/Fc7xpP0YHKRu3R
ukd0oiC002eP+vrgz1sbh7HLqYH/SWvEbYlfdhXxJnpTPPTPSNJEviaZoBImFUsnSmQ7SGbr48Dk
VZDIrrRVBYQpGb0dgVE74VXiJ5j3hex/PFYciJ09TdK3wuJ9QWprgloO5HJiU+sN4hF4TN+QzgQG
3AWr/ShjoVBpj0OZzVqUy3FH1ia1KlmWPMoK9a8Nt+L2obcVPN7I7xS5JH2dTYeABn4f+zAKhzsz
KUstrv2L74Wdk8yxfhS9HyLb3Ybvs0+bUFf5mDt2/UuMhReMR4QQfr0utuigsKnSK50YQpUQM5E4
5LgqobeDzH3CMxJaqLlM7LXXuPqMZBYDSR5EoB5pFUkvM6KBBV1QtAQauZrYQbjI3r6xTH0QE21Q
DhylvOfecxWTC0bz3E7is7/KdVVFDfYGapZwl9eqH0lgMFvnDN/Ove/65Z1qKQ9VbvtCC4LBTVPa
7f+VNakqVxDH9g8fTNXdbebUnp9GtegDV3QDe+JPLvq/rl/uaAdqmt0JLS2UVjtXRjuCGqCEhFX4
WH94/eAFlp9xIeCFkyHiHKtMeRRqHu/472157qKM/RqFLHsdpCnmIOLmQj0yMGqXXratTku+XzIP
mc/XXgSH+iLFmr21oEoE039wXLKqt1DXCLreoEHyJEejtkyvn+iojRSLad4qvNA3rPl7BPJzyJG/
XuwSOAzTymcToBHVDaRGN/94NrNUAGfv1GO6rJX1+PwB7U/gSdNp1rWYLOt85+vHNmoZGyWUQc5k
axDz2GURYj5RHFDyklPqk9kHR9OhNktTea13sIProzWb0RiOrFEACttBANE7g0Anh9Q+izRecMK8
oCz4gTVzumwpYgqNDFl8zRdfwm5k29fLoKp2d8RlweuLzWSQjBKLxWS5CJGOU8HPGTi7FoXgWR8x
HRgG5i+gtCMHvF6xQ/PyC1Ux1wBwMeZVaxzuvOnXQ0MIAIeE0+SBuBKQ0s6g9aWqmDp+houp65O0
A+K1wSobDZiveOITdvFewNBkr4/QqS0x4WkxJ+UZiSx0vasmI78tClsZhZeNmwTgML/RLZbOoMYr
lg1roAn3y5k8mL6dhzjA15LrAgHNG3UwUAo+Ih0tw0RBBfne5giwiRE59xZ5xXhHxF0yXU84DrcI
SAlK5+TTaZ7JDUP2wnkTUqwmuxkyB1ejHERlCyoXPBxb1BHVOTdJ9eD6u7Z8Ef9LJSKT/RuPReJj
x0NWrVLRrw+wesKVLODf6a/+Wo58AtGmSe08By6kYHmX5XdPZqkkVeWBDs/ziOMjCkp5HMYZ1Ls/
iBbVAk+Qhn4lfsqw2w90ex32sKZNO6oMjY4y/Rktiv8NRz68TZL8tI5XHYdM+54B9SXe9lpvzYyB
FBNsyxJ+ZVMAIO+hrApbpmK6BXwXMbf0NEc+9dM2FG6sBbqQS0C7kDBzfD0P667PNQKl/5GLbNIV
nN9gxDdYmzGKWR6u9Md2Lc3WrEQMWCTfiKljqQCwWmvE5xATRO/XBZjWGjNSnrEufcpsD/Pk+TCO
/veOifkrIt/5bS7VtmW4FHG5uxIi0g0QpYm7qevWKMTB/zxL4eCPFLe0ju+iNhTYaIR1XR/ww6mu
tj+ogdCskmcpiWUbYBpfG1aIgsIPqGhhJQ4SxfoNKRuKejyAzMKrGvvzOKUMbUjbBsW0pDjEebLJ
qwAjsOWBGzWuxVzOhDmDsSxA/rO/RU9vK5G+Sej3DZ08ebchioTE2wzJD3GsmPvGfm8CK1ouczHH
QEMSd0r7TB4caE0lPsOaUW3mi1y3yI3CPLZIiFVCoUI9qMoHRbQMrgyIK88/u1AkBWqpT6rKQ0km
XZqraK+wnGUv38ox/COLJ+ZPcedEGhxXcxt8e3aoT1UAFNYLdXzoYbBszAX3qUuZf5TGl+uvinPR
Ar0p8/uZDEr2sKo6Rkg9pg18L+8DAD3dLqpThUJihwxtmgsA3gKSMtVDlG8OiesB3v5C2Lr0Xmkn
LofPyuSR0kuQq5RjsfAqAUAvwMz8BIkHvKlWpZxEV7HlTA+IUG9bwEZXT1xYJSNcIhu5kX7Ic92I
0DE/BgB6cv3g3TulsjCT2Qz7ov526NUGrCyWtdJvVqc4FmmmfnCbjs9vQilFki5lrGh8T1C2ulJn
RC+1GqreJdAEhjw/JmE9EY62Fcg7MAW1q1OPqcvlomAvIZh2+g1Uz5rbwmmz9QfXthB0AAQNihdW
nEgrb45o5pAswORDufeBYf6PlHpuZDkjfrYSm83zSQQNwq1oCzcKc6hVUjaenu6XpWdyU0XZjTaq
WICIgjM7W/msNA7Qz/9weauMy23W+SFNER059dbrLWYBz6YnVKLnqcx8Flsnkdu4zU2cp47p+dfK
7ZQWyVPrKnmr6M3zrRH5vjoru+Ldb/CGH+YO0C9vbqTy0ZmvVqnS6X0uN/b4dXZgJGk9c6zpOyrg
bCNjTX7kSzf9T3kvZeGyEO/GkI9cOStktmsKCOx3eH93759knmYiMsIvygYIt+b6H59iKTYKBiQI
4Qh6nZsohCt90onbvp/2se0TfVp3m9RBmIY2lizj9lndQpzHc8UTbpgrm1cGp0LYGPiKunWhzuwK
KpKDPyE3PuD4OCSuIrkyJgHcioleNO8u3E2ih+36gjIAXKoSZA8EPkq74Hkzw5JickkkhqsBYPtm
b5UVSSgKsjhHvVQvDS9suSRBR3g6rUhMcdG0LY1FzgSi3Arbcs7uU1P0ro1/3i+PLJe4yZef7q8b
s51xNmynnTd71Bd0X3M+QlkqyBbGrV2Soy1Nn4dBmZgBwoAjFf3SfZva885keaZaRGXEgTmmyqaq
/iJkCwA1eYxcA36GFRBWa3PbQnAnSsVavImHtWgGm4hVLYY3TjE+9pbfLpY0lP+jMfzFtkli7A2a
amXwdjJpsAW6wN9dmQTJP+i/RPfF1Iu7ObVGpYL75B4N4cf2i+/9uBJT3ZqYyboFDBVEt/zElehY
j37ITph/bBL6AV8NRxMvCse6vOm8+kXH9zmploX5xteez9DD66m+O8RYz9tVfrlk2MgW2TeVLJwE
5VDIsxOd/h8tBU/JyLty/0C+rDRDtoCrBAeVS4Otp9LjgwLZeedYWDEDljQd9sD6Cj5aRIg6NxFN
gVDAW9SvAIhBrdsG6rM4Qf+3GUhrukZdpGpt8fXfrYijHitun4PA+6sVEOM6J10dui/CoPpF6JAm
Hgc9ScXA1nH0EQdCnro7Ja1NL+gpO6nxqptNLKZnTKd14QQ3EbJO7wTBB2Rz8ZWh+tSMBdaxB408
TE+WMZt8fGrSxsGzTfPKlRkHWgLO0nTy51rTB5+giJiWi59EIgcopX2vYC/KilIMcnYOwcawzKon
gk2sJ+dvAVQZxXbGJZ9V3fcerqW4pX76ABXE/2J9DNKiGXXH32nB+jk6HiFjwJG3dzD3usOcig41
Madhsl2aCUXhRSH5H24RcpWg4ATc5ATv89csZ3HxVDWJM4fHre22WDG3pet62xBqEy0a/J9bIrUY
cOiBoGsNgvpLlXXpA5KvLBTvcS/esF07rIWlsTwoG5ED4ql9muw+0g2JHbIKW2PLSDb2Z/xSf1Oz
/08uU1ThdA8MIQWF9ua+6mbrlhsKJUAf+j7KC8cW2rZ5ixGKBCFvNuknjO8YTr8ZZfkR9++tgrHF
Xnn9XygD3ALiDOCHou7g0dTtLd5s7NC5i1K1xZ3B6xUvsdT0R8al0EIWHmk6qnLt7mtp26L6ruNV
2ey3L+/MB7P0oP2x5ZH7QXkjLNuJ3HsKCaFHl5/OEIULfmY4nV2qqph1KJOv1LHXTc5w3AdReKtS
8rv/nV321cUgMm0KLBlT1YTPYvgPFBRBuxVEBQPP45WM5/Jjvota4l0Y4rFbrViRH0mRDMOrg2QQ
dpAEB945MDgzNfflVYQuLuMmM8qlSdxHJJgzBAcrMIxR0i4lL5uDV4TfGBaCOXe+yDdKoU1QuXlr
zwWNOwmjd5ANMHA/o1eMMYP6xurpU6jDdL/rO/+CvvuikLMJAQILSxt0pp6I2E3SdhU9oNggsQT2
Q3btpmxHCk/IBzaAwfwv9RHHLT9w02BE6ouUOM4NDWxc9F3t/tsQoRMhTgcNNjn6QOU9Ck6fMTzb
fFY5j3JXqfdBGvjNKhq6GxRyiApF4fB6tqt99ER0kVaVScGJPkbgV9/Gzm2IDnlwkWnx55DwIXFS
urtBNPHIB1w0Nn/bWA5cCNLpN0L/lw1u22lDRkuzobsEGjepkG8w2yj2n2XemTRmgQIMULTPOjZc
k4f6BWe2EViTBZBSpoEw+81zrU2H2eevhieMTodcMWjNnNvXsZRciSSwKFXiz9qu7IixNVAjO2mp
zLeKuNgojv/ikt9nmnJnabUsM2HOOn+Q4jw4AIfCngF6OsnbYkpCEt+6x2eOYubRpD9dd13BiWA3
HKlXSGC0uTSQGpO+CJ24e3G1W+jdwp0SDP0xLmU45JDRJVryH4NKyLITHMeSG5nrZnn1dV5+P/hw
Y1BpZAG2GA6vTUJHCR7FYXnRmBhDJTOHWrlBqOXLoH44nMqfMbaaTGYhBALV+u90xwEyzn8M+4Gw
8sMTqn7GjI2fj8BN6eXPZ8XmwEbup6o//9rSMPlJgVLBHYFWRPNmCWYeV4b8ptWVMbYoOsJ7dCqE
5kqgYoa9Jm5/oEeNKSqskD4TIZZs05rseiKhjzKgOs/mqVr2Q6K+/kU/+M+ZfwL8T5QQKAMMJozq
wAzqP/0ftPXUnQwGzy7y4yD0Jca8Q0NVKJnQudHIaTojCwyFJoviIO2LlUnYHm56unHot6hT/Piy
n1rsWN/DkDLKwWYdrxthd4ajhIQp7khgosBSXWHK3myQogLNOxzagitRhruK9M3wzxZNjrhqTHQy
Bf/kXXZLNYOWAwHUn4IDmqSCPewn0NQGjryNBIsChWBdOlDRMnSO9KcAAkSTvJoI5FSUbuiUiJ2W
V7p77Lw0vBN3GAJThtCFKTWQNVdx+xCFsOhkEjKaB2hfxeXPV50Hb8GysQiS1D2Aw8NP5Wf6PVeg
IE955mQLXtbc3S89z4Kly0U/VBUyjVHvSIEH7zagmlma/zL4kmOcMdkeS62HXdrYE0zPLd43WeLy
xRbUZliPcwYkJQS8rFwD5nYRbtCJI4myXJd+opw/AN5EE9BeF5YgETKF+7lSVfHUh0IBULs2kvtQ
z4bctEX8K+yH4toTjFqElZPvXX/2n5vMGUukTKhhT46FI7aa8DnrTame364zGuIEZFWfHsWObqgJ
jWyJxq9B44E5OVp+3LU+jHBrEJ13LVYnFpQpIBCrVKO9MO3klYTQ2sm2BLcMmzczD/5V3cdxzZ41
+cnaI2X41rm7YZvaDHLRGxiFHPjfDZTlLN+Ob6AQO5hQ6BVycOhF4fzfrdP3b41LBoh6KAFxg6ky
wRr9l2utI39t5t1Z8ktciohCokwwvUmCRpUK3QP4aJ/FPOIQKux6DIrId0da/4IiPKPqbxG0aFy4
RFMrfDjDmfWSyL45g0JK1hZe6HvD09b8GC0DJbBS4T4bNmNrib63wv4h0mgpGm82c+pDKSdXGEo3
l56WOmDHInh9To43pTuqwPAIFxtdHCrqKRk3+rSrVNyjWQIwn4Ju7mSCV/Y6zlbR9yMohVmx4xhb
GZE6LmKesIOS+sWwoXwJWf0KKgDrBBq/6gV1nRHD5PX9p9nIQ6ANJq24cvORGOdS2V3Zsg7nLT+P
p74gGBic8fP9074Rd0PEi3m2VC9TCgNcuCxrBHe4HcY8Txza3wp7TYtWEUHSLiSA85o/4UBv+mId
/TvTVZtBpgf/JmjXyr6yW/PjEe2ZI9UjlJYL1E4lonb4BZKluOtht1jRLdZrd20k3MXY3ukiL6/U
Vqn9ONfMZN0ATAGyMmZQ2JC9dl8XSxW0R9Zi3P4eZRORKHPLR8iDLvAMvmly6prUKH8zC+jW8DpA
l8bfZqQ6HlXtJTK5fP0KEAt4Cp8qws0AGpdJ9Vbc0/aB1NH1g13VqFxC5LezDiJ1lZWmlECazLn3
s+eObyHfSfQqG8MvlPEeRQgHym5+teYJ1YvyG6+dr48K8ysFxL+us6M+fudpBCjH61y2PtRDQnid
73PXK37ZIrw5URhrnwq0Nzkq+mWkG6gmkQ7nVMkgD2bwJ5Ra5ZTUgixlWQts8yR1WYHeup7Clz33
jkk1SRislhzK9sZtLFmaint8+qhLh9Vc+jxj138H8IK74iG0UzcNE8UzgsGoktrfoZVidsfF2IYu
c5E4Oy71rkLr2qK4hOujIUwVS2bVNISbdpdvlFz6ehyDdWj+OPLZmtQ27VteS2r639oogddcSiAz
wGTJqxrQDp+N9Spq4s15Mwax/t5SzSrPofeOgWA/eykVjZRfq+fjdOb+fT8OWcRJXkHh/e8DWtXt
NzqxOOAHpSmrhhCZWmnI/I49chCL0NOG7n8WOaxNWWZlkF33L8uQlrfCISEAZv7p/x4MLQ1L6Vf0
WPyNJQOtCzRF0D+P7ASi7RoiM8KgKAihbAviRMPTE2Yo0RSQ8zRCya6bd7Gszn3rzF5MkdxfnMkA
MdY4ooqjbmAD5ad9c8utJOS8UWu+pMNpl9DcG6F8BfFvvlb8drOT0mHYDWwYBEjWQEgqGVfLdPMB
llLylDtpQ4hWVTqmql1k2+IgwVUbe0Ga++20U5uTJqLs0L6I5tDiqlShurfRXhrXoyjxQtRsLTlA
XzCGjZgD/uRZcRUI/HK4fNhy9HRhcO+HukE95o/bz2OAfIfuHISCF//wE8PpuV9QN1KEPB4J4Lij
V8JWvYvCN2lWoTwPSzXUO0p4i4qWpqVJYuSzXe+dzSNFyk3no9ffVCnrg2UCtXWJTXy815ptfrY8
DxpcUtky7b6678PN0OVmV3np/7Xgu0fgu7zz0R7bj1wHp7lv2Mw/WwmQpI4ejtrGpUNIZDDE+esV
ZHhsLI9u2ypcCl4JbuvMtmgTHgg2IzNsCczWEGzIYXwO09NLeuwJEYrSoYIgELey28rUajt1MAfZ
p1vKBgU8Jxn8nhH3L3zyTXw1NDBVgW96CzrYG9SsaqLtoWchcgK+iN0FdMMLcwBPQ3Dwy7G8WUb/
6+EDpKJI8q8xLRDzlnKfrf1ciIciS7FDvAMOvwAfbsrC7WlC+wM3rG0KcasvMPMYUrmkpuCFKe1o
TDvXhVu+JR1JAQiwCJ4CoaeVvDOQNFCEPutyiENpTiswNktUhN59oNjMKJAQ4b6rx5n50zXpO5Sr
dmmOTbODDosWkHhyJ8nVbIL7DM4YrVeyQruc7RRLqrKGVvK9isUC3sMICdV/UVo8gYepFA1B1OuW
S5sT5h1umqLsqm0D2s9Nh1qBafslt9RebkHc7suIxnbvAKigfSD2KAyt9vZlKYPZ2pTUypXcPKP4
Ygqg4RjqLZgeFXgtAEYQMsReVOdfq033vw1lJwu/nC5jz9aVwQJmiQhipZeLZFxMdDgKmSyypgB0
+u32jyJJ9kbFDO3VM5rYaBW5e5OP56e/WFSekOYK/u6EGHvFhvGWhZ2kKtUM3qiuUWMi/koVKWal
TM8sw4c2L4u/DuyH2uKcqiqvD/U91WvXl4xims225kGHoxxlhnE180c9+1OWO5M1947sEUWKaDoQ
UsGVpo4pp6+1HtCWcxiTZNZASWoiKMoVdHreUijBs8HzfUgVWsmtiDMCwojQBye5TI9pyr5pbUPX
KU3OvKb38We/xWq9/om7VEkgynjNPhLOnaGjoJrAh7Irvt/5RXwDfcAWFM2mr+JS/eQ7nMPgUlUT
m11t3J8NJ9M/bWBFfiejoDFqAfx+5DPdka+b6te4oe3qzBDiWVODmHEXwLNVYm3p4yLQOBdtIA2y
uIIaeID2elhqhgwQO1mVyDUxqYkPpk76nCo7lAWEEeXTSjm0hOAOtRhCMA/tUYEfqRdgI+eUYKZD
9zkG+F7K88SbjNTakoj6zsgvJNQqMYmJ9VDkgL6dTA2sdtFsA+WWee1S2sphWfOFq+/Tns6SoFoU
suq+w22ywaYsTvGBYiHocT6P3ro4KSUO/+sueHt19xAiXYA2yE/O1f/NFALtRPX7ILfKRwfw9VOh
JS2FUwI+eMCFmDdEw5zgriXBdB1lN4Jk9laAT8IeQVhtNxRoCROy91S2gYiLq4IWPbPpf4Fui5KR
MTpJVZmT24YaaOEjSN9eJ/TwTPxOq9+JiKohx82EZuOH3ZiTm8J6A9eOGuJs4lhBwiRhTVcy7+AT
zOc8msu+N4f6m0nQ+tXqK1hyqSgRIWco6Zobz5BOvGjM0R9nz7VAJBDCWuebS62DaI6DyKe2e8v5
cSzRYyGYjlXwWpJiayHoSPhIQsuKtzQsUPBw0yZz+Q3PF/tzF/jDE/nWS8VlfdjTp6BTKQqWMVx3
914EKdY6LvQhWrZ0ft/MJfJOeiNau5b6xkD07ZQOTNaQEHzD7WXkU/MeJ14novmI++dEIHsAMxMW
T8AoQF5DmNOHUnTs1S4mOuW7u8FeWcM+85im5bbPoEqz0hPUB/pJh9t1C4nRSRj/iMtTWwb0FLfE
mvz8Np0een1ecAQiuAmebFlR7QOwHBp+JqGH0lylJBGLjFVfwBsmPxu07x6S/83At2i6J6i/sZ/b
pCtwf4gkTKmubPJjZqQnhqYhSqqpR/0TD/rW5Gnwv+ZXyfrlG1tsUpsHaFPmv0k1BUpF6siIBpsM
YnJseXQu8uH1IQrMh/KRiADNHEAi7j39+iCRUB3UKN3x3jr5X5tUxJXe7P62zpVBU6i0657zwYZP
5BiULG1ehuh8rSE++XQvPmLe9mZUyGA/GuTrEFPbGFWlLqE4Buf6c9PuusjZpj7/zHLmJFHP/FOH
UvZ8YN9cG0sG/wTNHGlc8JWCBUNdw8T1mNZor0hnYlJnzkYvpuEf+Z0ieaKzF+JQNPPsquMKKXce
VIIhGqC5h3wMOIA93H6wUP5q5iX64B0uQrrbFCWx4T4AtVsjl1lUU4OK49lFRxwEH3SeZfuKoevt
lnxRTE4xiTKEYTJKEUU0Syu63x5oT/iQp3GHDfzyQDp09Eu/q/vRfQVU3ThVQZPvLO0zMm5K6ebb
9JP+NYcMRZuMndisOoNQEIDLmMCPu8lSevl37fiuu3jD/q8xCDwGpdnQGUZU8hq1QSFt+H9jKubD
e9mggxUcj7x1ua43ZRLb0jlbdUJnax8nqbqq0Tj1vcgNRG/stWcvlRWbIJSrrnKHiIWk2qpmzX8t
Rl/5kok5C5zQmTeQHK06WqQ0A1gs7CDkAYkcWBXIBJbs7rY/I5hWIZ2Djiwt1bo2MxefipvIhDmz
G5iLwcCpw+HjDDlEi6v9qBGXABdb+SJ1npJTh1hjg9FqQdMw184zDvN6T986iJXeZvHmCl46X2XP
R5PrjgT/8AcrWtl+Exk1p0b0XfwrhhJjU44ujHpXr3KHNeB1bzJioVdhks6bnhDwp+IqTaKYAHlF
7aE89kvim9MPbfqA8yiNoYnqCV0xGvQsvZ/Kt7MdI6oHD4Ke913QbGINAUjND6rgRU1weH1ADCKj
0mlnV7A6j7zrQ2QFniX8pTChZrZf7kj1dnMEUw7TpavaHJtp8ofaEOGUSMc3OQP2ipSsQOoG8Wd7
RX8cNdyDn2XsPxAaf2hEpTa32b/A5UV5kjhPaKcDkwDbuBfqpPs4HJ57oCpiFdWvyU22c6Zxm+t9
Quj+3eENsUSiJd8bIJlPk0RZpSMIQxnf8VjgTDF7vaROwgDQxLvFTEpSOB5VUU0hiEM8FM9eyfw1
xuZgJblLthBdtEya+5HNMorfuxjmI5vdZstCgPmS9Y7cwFhAOjploCUuU/Tinsj1TsYnTdjLHuqp
Rc2YRiKZPtmxjpQGuraW6CL6qWB/HtceIB5Lt60KRD7gpTafwvavCGLNt7vXDFaqB2R4cQOHArue
hWHssTWVz5TttlALuDDsQKD5ImSgWzrtLA9eXCyN0DwFs5ghW5ycocz/IHLFu6kE6566xVgJeoEO
PraAyf6/1hd5XJxfTA+0LvGaGCQHoI32siZxvYS0dXx6UBjcU9mDWBd9sgBygU5E4p8myobDEBPh
Q2ZqmqKyn9KdAmNb7mC26z3M9tqFoKihMOQpOonTTwtgC2efwtl8uBlEAFgxrIeHMQk7Il9pluC3
n7pGCkzAfh4+NHBw3qg4cs+FrT3osRksX/27yeNI64g6YzsharwOw09gl6eXkB55FoMtD9ZoUhaI
UGBG3nzkh4eEshRPjmF1OxykU0Zrt3XU7bFODHkTuvTiMDbREPmyScA/3MWWsqhSTFkCejpnCG0P
CYk9UWe+jCVSeq/M5izHdkRRlfN71Q8AGddqA9GcE/0zfBNFaCzCOWkaudNfGiqzt0v5G4uuyB2a
PKYqzKYKic3b1pRZrjDYw+X8CcWCE5OPWleDa2fxmU1tqcdSdHLXp9aMyEC95jRJw9RXgXMSWiYK
DOJjOSgiqg/w4jqDN+rTRX2NYsNw8the2qlefjSQjToStao7EROMF0WVMQvsNZpDqQ7NaeJbEh98
EaCIBZtyk/Raka1N689XxW8DT+Nayyr/gioFuz5Y+f1niFmTHN/cnIrlNGMvlnotpcpWzWa5gay5
gKDc5bOa/0Cke9FwB6NhveMlqQ/u5Pgc3U6REfX+Bv5zZH6aZPz3+NdtnpJDgroe1hILsLbJ5CiB
toEKDUXdQ8jbiYcOESK/VJGpB2yxO+XDl4x7lMycT6YSMZOacklaxBwKPTelMAxHnzcxKD7/OPAa
RRIkRoAGciCiK2mRaDIHErsugt1vUIx3Yo+qDHzHDgQfoeEqbgCFvdj43KjzMH2qX+7TkpmO5Yt/
g3GD+d40MERYJqx6/Z9flMs7/TyeYezSt/BqgIpc5DoEhATvydm6ltnZStklDytWVZPKA6VaKGYF
ZgJMEASn8b5JyJfZ1JWos7Yzq5hpJiPx/4Ex1dBpDdd/xGlyJEYjFib3H2gw5QooKmC2vPMnKv0w
v+l6yygUUKcotdfYI1uBK7sf/pOkjUeSCNDUYFp2ykN3nG/j2vc00W0pRkbrACzBotjbzB3KbAuO
sGV6KWJmp6JshTriXose2gkGXnkAJJt4QXV8xnhMOx05gI9FPVaRauQU+fkYiBqP72/LfN6UDCqg
zcCfYuU+/YIDPXk/7nqzMrZDVVLU4DUmsB1F1u6SEiaF99PwNOvwYRyl0sV7k+mJSD8NPy0MPhXX
pow1N3yp60Y0qWqEjgBiBtUb272J2dcGSiKdBSrwlcISLiOc/jy8akcU/63YN6b18n29poqcpf+i
+n+5cZjS9tEyU0PzYByrrPtftcLNAbAriOiq4xmpgNE94kuF0eJNyh4w1u3YmhDT0fg1RP5xMHa/
c9lqcH4X+CEl3Q5kdR3iLl1VfA87JsObuh6L3IMurS2WuD5R4jW8uaJRL/bM3VSHOMri+/GPeS37
l1byhFrq+MC9giMUN9ayobW2lpbRGD9Lxs1adizLWYqMoP7npEMTREJy0OeGOG7AvXFsNKd0zZRx
meDG0DXJsXPURcbzqN/epPBr1HbSIQrgVzvcv9u7i5f2SpFP7Uwxz8PuTU8rC8YGoROgMJcljDgs
8imYZY+eLETqNXeWc3qP3jqzKslJlmSu1/j6GSkk3Lt7T+wVaz7tWEPSA92iyl3co6J3Mc1LAFGS
OlUa4M5+d91mLnK013B+2Lz6UPOC3cJo2QQQ4cdURHbGGA5+QxAvfdcRKLKOWwzxcx1TpxUwVyO3
3WNhCtFz7D20Sg8tjJwoDxgarXgl8qkK4i3YQkiAIl+p0raGJhZpfT6fScYsHe9ObeaQI8xI2m/E
C98QZGt5JoqcihwSwvbN7XApHzEzmOnl7N3wx6+w1xDjPPSW10ehjHxZwiblTLAenuKkx+SC8coW
XuXxwKVhGBQWmxqEkgcJno1riiI2GpG3CWVy5H2svxOvKFrcpTUU9xOKxzlj3ucjr82kdcHK5A7g
1XHNIfWpBkRd8cnsH6SlDJ3fI//9llCHBFhY1kOVeqFNV3D64yfAGaypq6WFprDgBxfQJZyXbinm
xpI+OVJ1dafe0O4+WvHbPFcBpaW3dDttJMQ6uIV2ZX4JCBMWmDndbfAfu7QL0joJG0Ps4PqLxWEf
yZ+waigNtyooTQQifU2WQc+SGKiEqe9wf/qSQehdFs59lb+JZmW3sSQ3YsCMgt/cQD2hxNa0ydBi
5aUa9SRfunoy6FMxXJHXGduY03qvTSjdHjljS/SjLnyfjYaSiHVgGtJLgqVuXzH1jtx/LvsMvr+w
6foDYzOBBSjQ2mcWJAk9HIi21dQ//mJw65A5NqvuNBE0XEdJ4lZGVdtGHLLXewQ3Rs8LjED7I8n8
gqhlcvXUD7S8EHXJmxqE8abeAehHd50JCMaGYe3De7znlcKmYZFcUOc27AA4FCzkHfnSQuzDX2MW
SdE031irZtbhoFbowCsokUh0i0shpn64a1H4IfgZo8UPFNy6y4TG6OqgXu+udBcD3N975pk92mT7
ne4pxs8O5Z7K+N83ril1+L7re/3xFXDCEBjCdqI/r7Rc0u3HPGa3a9LPcRAZ2fRZUTmjOi6WUr73
YlrPPHS7mrM/C0HzH+/MPi4326rX8+VkggYUtIdfYmvsOfzh3YHK2t8NFHM9LiII7yWGKQcD8QFr
TIlKK/Gjb5r83S0HXAfFIUAV01J2Wc9SjqHviHR5DXdUSQoX81M0W9MD2wgpiPovng+680fVgAof
v+mKUF5y+l/r9o8R/4FjUwCNjDTxct48rQBS8zEKf0Vkt+wtJNFGb//x7p7D5SlGzHJx5sCZUrd6
9qiYEvJe6nVi3WcIZ0nPSYYU47dOGSLdTTTdSYwoj9VGbWHSofiCpG6H8uGK0uitZG5qt7Tt1CS1
k8t3eAKZP6tmtnJNKqZ/Gkru0CLpFo/ftVzJq5CvVuLHThs2JBM3UVS4CsKrzQuki1r9CfJXfZSx
FeBya3GJqdgfLFbawoR/q3y5ehnnFRnu62QzoQwc++PkK5Bgc0T/4sIwXdCCSWUdbJuLNmVFW/5e
XCyYdVgR2fPrNSmaIleMLdcPrVAqEbAumBkw6FgbZgrbzO8i1+aEA6qBsVBP7/KkOQbvdWf3X2c5
zGkt3SUXx8y3GZ2FBL7wlKaiZFrBUY8fFcizr0kc0sIJKmGJKh3/EpEwSdl4hpg/wHJtSsCoShNv
pG5B1YQkqwyVS5eJ3mujBGdKXKUV901mUEIJc96MaM7DPc+SJcqSvF8rvFoEsWA5oRUzHsUG1RSg
w9zmSk0tJ8zFyI+Wb5D8rol4RCm7eAleYYtMo5bEoHeQ7Jx1HBbG4bUYi8/XDjpZKUpD55moBr5d
931HU3mYrr6X9hqu4gdqjrzZ3GnPe8wCgK8Sr4yWm9tGNCNIJykfRuYsj0EegD4xoh6UdWUuwN0e
ujOEpnQAqoSokI09UkAoO9I200X2SnE2CJkilVQ+AE+c/HcSiiSIBJN4OQnL/4biC57H6mjyjyGM
ZLaFVUeGr4ymTcUDuAPyHa7kE9TMtxrixwyi4FxuBp8tndR/P2WfL5HvmXRI9wcqN1WTVZeUNcJQ
dG0pYedHufPuSvV/7RiBIuB6sBp1e2yW/t9CK+i3Cq3Re2WhzTwoXycG5BQ2e+ybMi8Bv7gNQ+IY
VDlbI9+DMU9ThyiyaOo+PQER1JACEHM5Ww1BtXRMknPMPzluiMMIU/e8YrUgyNXzMmlKvtEG3A/b
t98cnzFT/SObu6myy3Afq86R3aqDRykKYfip3iBDYWuXnEu1Rc+RcUxAtMuysYO0LYILvyBmaPcE
+9D8GdKIRuLf/uplXyDR3HbdwYoOpAkbTRkJ2wi5qy0qSUmoiGAi6Befp5ucV9mXLqNQIRsYo9ve
rU3xt32UBU8QYtkjerNlmxntSwEgDS4eyUqSBoM7aPAFar3fEzvZHj+bX8Z+oQY/3eZEjDe3t5fp
EbkaP/fGiz9+cSrXU7fq5XisqpTCgVeT/JMzH5XgGjPnj1rt4LtMt8D2munF3fLNkDm5c4qOTuw2
VMaHe/61ReajhEZI6k35LQ4HPbdYmeKueCzVjBoz+I2TlBBF48+1E0Foa88PN14/TOkoz57/FTVc
cmlbeQ/VSCJuMQPZMFaUM6w7sMIhCsf+7SsDuABi6BexVInn3qUV1Mk0m/eyVvDX8QeO8jXz1N6B
W8APmvVWAmwBp2LPvovk76ODguuqb/alEmtU/3OuTsRbzpYyInK6giIgrL24rwoCcUACt4ttH30a
fbSAAKuRRwEnKeHRbjz+EWyLk8hdhE4qTUmFezb1MsmyX1uNyuHGJ6uWTQ8clecwCWHMtZYCY1sO
FPaVLP8K7zrWq/iOkDMH4uiOWipKvxpaJJ3aaJckrVXr46NhUXvcioSbI2GaoKvdCr5hTrWdIDc3
BS8fuzqSevy6P+rMAYxKnD/1/JRaQYoSGAtxGSVPpH68QqKVYboTe236YimJA9XiHDDS2jQRq3zc
u/yE3zHtIs5cF5+uXjxQg5y8Vj4UnIq8YZcnCQ6ncUbM/BD5mLhVDDogCcOBO4XRblGbwH+P1EkX
sVRubhTEZmhYgzX9/6+GHBwIhknrKyqHrgByUDFe/XaasoYoPN6eIRj6mDzuo9uLvx+unBXnBrrc
1BbELTJfMMI9NZpoO5Lrg36yvSwbPfDknbLaY5PBED4JobniQhGnYPMVCGBYHP0UTFezEI8IhDcD
hkoEWY6UnhoU59mtVSvA2YCwK1EpwgBSEvMyv8p/PmCajeM5mpfb+DuzkDZNphVfNoSCh94Qvh2v
EomjRh95CXvYi/rhg46eMNBoscWlH3EEDsuB9daC7egdaVB9CxMq9B95/Y1ixjal+rESStzrhPTw
6sh9o6w7pTBqbNr4YwMVHaP/jbCWXGh5q3NxxctW3YX0wCEb8uGyHsOfD4DI7jgE8yeIPgVXZddm
OlTkcuU05WkOl1zaDSMGC+VyT2Qgbkwe2jBjyeB5CHtZyM1MFR3QgQ9Th3XVE+m+plHRjWQZD621
bY0gxpTuhvuthspbs79CSbaTeQMYsPtbAPdhRaGbEjYeteoFXdnG5lQBU6DrpL3R/PPAXNdyfnO4
L6Jmv5BgQyZpTIqnu5wKbj42jRn6Yxeh4WgtaflsjeFNq0FkVn2LgfW3dHnHF/ajI08IhnHWa42Z
/svp1eXNszO22ZOdWxBQfw5r0PqbY5OQcIWgSzkfwQJhQZhN4uqJ/tGSpFHHX4FEOmrYMZU3ZQiN
5cjc0gIThwaPCoUvPRFjEBhrdROKCFwKYMheH60yGiO8bX2afjKZw8Q3uxQOeZtSBCgzINJWFTW7
/B8jHerWxzLPUn/ByycNT6ZNIsUl2tJNducgFhnO7VAO7nqueZworIAUBtfVhPbj4qEibuPN4Lau
VxB0GyK6fXuOsorF5wGOWtE1imiWYlBL7ObURu/6XVZvUf1TMJJTYLoW51c/FVBpcdYLhfHNCrzN
wP6986WrnSF1tntCe20WWlgA8ASKSNQtmCGf3uowF8CTZIXxYwxH4TYHv8o9X1VtwpO3wIAA6i95
EKC/dVUMxzuOx2tb+4yd+NsDJcBVrsqstcMl8kjoee0j/OCXHdxGQeuNeKdGpxyNwwoly7tFfQ+x
n/iW9M9M96Dw1n+WderKFdVXD1KVVmMGIMm3dOtZhEV2iSqESMtGkRpGoE2WuIuQwJ1cfMtyxfCn
zGmoB/RqBS2ySTNM7zoRmqgqWn/uDXckk5T37vr1WAPsWzcUKZ21hvyT8TKabDgmL1Vi5Tq6MYM1
y6BC+ieDWnfuxMXryqAwi6FgqaJCtkjZBVYvCIn04ULyRUHUD60Z0pBG23Qr+W4hhntpZyhSdsrT
RYsPU3TkYzr8bOQvdgY/OTgI9LaWVLpRmHyZs5r7jUPY6IRUEbP8BA5Q6/IWH5KDcSeWEt2X9Bpx
+URCeRruW3ostIlElgtirSsL31ua/l3ETEjuq1GKwRY8+fc0D9XmOtYKNC/GotpW30jjMRDgTF9h
5dYkHRgsbmBtIjR67BryPZFSeVT5b2V9il2m8yMHBf2H92LtAAu/5+/Vv0Xtfi5bV7353XJCijWW
pP2cqLDqbUZz1goXLZAvvZTmmhFN804GTsKnHV6shyphXKMha5kp9MLFrju6P4K7fYqMCssKUNQT
zo6A/SCrgkJ3JCDHSkEpw6U9wVTjaiefnmdX64PEJOoOzhOs2y9D4i21pH1js/TVbhqZOgufMvW1
65hNc3SUfieR3CfNuPY7Z2e9Y1oLxMeJhYQlSPLiIZeO2wtnmS05643rV049bPm1SFchzTt6dLx7
nHZzEUs28c/rQ2/LIrBVqSymfegAa4Hq2ANGRhpQPasUw2NsBc3VjYEkGX7/sBTYz2EVR+oUf66V
/3LVwKeU5TmXxJrgb1EDvFyI4Bb3mcfGhrE7MOA5x6JVJisGzhdK0cgzU5ubgApzEJbXczCxfiD7
MwsAV/lOE9yogE1i0YFxcYs/C3RmhSBzcSY2qGzpc8I1Yua1ZvajEf6LuAE7iKvD+EYoGoq6HgvI
rqwvwXwtVQ+O4jKXtXD7BNeqsZguAyOMHozmZ2b3KSNgVPl0kF+V2U7duV54jmSY0fuf3AGZBgEp
5kLVtGhIOyW+OAJPLyZt3nnhmkOmR40VOsU9eRoyprP8ZRDNHSNn4yV/uQkxi2a8KHteShbbAYwT
t4AK8qagzrnDnMJHHC3E+jT8RSiJmDIE38D3SnLLQAZ3gUsyUqMUlLqOvrBtbVuDLBCORcGohTxM
YWch8ONXOHkO8jrDp9fOUEGMHmzQOS5g6ZZWLKoXvXxz1Z/hAGe1VV88+IPdEZhTeGXPehblEaxf
V5vhm9H9BiigcLtfTn69OelIz8ooLuSU5kWALhcMMBBjpxfgES5TEvI5+1lkOVVeJ7eVZRe6jvcY
n/+7mI8E6eZhqjNRJqJsrY5a9UM8XhXBUObt71JrXqmTy8bHznL5oV6+0BMxQfMsvkbAgxzsAGCO
nHb+wptMW5n1u4H7GBX7qca2+YqaJ1CFaw7jaul+6WvrAu97womcQwMgqsNat+qCIuXD/+wSHWwH
zS7zl93XraJyUPEPgrlwLfjkRubbfh6JBYZnhkcb5ZmfKcE735KVKa5jGjhXZRgzjh+P7eJfF5p6
qLpOAyJHQK3RO+iKaWyq2gtHKUGFhMUY9yL35F4vWv+iZqCHt5rhhMStKWBF1FB5iVm8FffFeebx
EUWoIPb6TvERV+Iwd7vGl5bCAJ7k3HQa9DED1+/AOHw87A/IWmUyVxDu3LQdxr1xKM4wsjRC6QED
nW+CqbjfB06UbPLeWCg1+l5/smNe4gUymlAWORk5Ymhl8MK344DSBl0bEh4h6+QVgJT7rzEbGKjT
37I0qMAZR0qamqRu3WnmNaxBvWyCzS2/lW41/lGwqbbjLlvLX8VfaLqht1mrAojdnYRFCW9GJrqG
ayUTgqDH1JKMte1o697ZiClksbgGA8kMstNQSnZwJL/0Jur9Ooy7MihhNduTpq+EccXSutIqJBNF
Md9ddQKprGvuVUqLy0VKkqeMQg4e+3XqBMWIvWm3Ygl7S73muf7rUN4Nk91bH7KcgyigOyGsvxYy
XJQpIXAyDBZjD1yTJ6GOt/7NSONV0z3b9DAPHi6JPz1qwl4XBzpqjkzjtuzoz+8eW6CPFnTv9Xsr
pFYhgpQxwOsAafj1PH+OugTQbAQuIsuBUTIuuYtq7M5Yx93OtE1dn8+Yn4+/l8xV7Cmr/u5PTJZN
fVKuyxvF6/fajvxiqgOI7g6gSBrGbITe9iS4aHkw7jLI6S4EB8+tclfXBxRdkbbcDkXBcOGu6+xr
jJuUkJPDsahQwBemdVMopY1DNMRiXG4lXCd8ZKyjjt47Mbs0S9+l4nXgYUb6LkSwpy68gU0JdkD0
Zny7CzTKr5NqvU1H/rb/vkybFtXhu4Uh8QBdo1UXdhOeQDx1EGkUBHmIl95OVk47k/16vrZxX/or
YOaxasTcPiAcFZgkrvGMI0/785/NrONA6UkIgwbc/ZdWAyJGjRwAFc6nLOo6Zqh5Bo0OQE6cO+PV
nm0VdzrWPTwlmMCWI+LMgCEv+gIDz4O6H8cXtWptclruyihwANI8c0HnRDh4A7GOGwxGgkJKNZaj
39gwd9Dd0uEnDUfcNoNOtzt6v2vQ2zbCyh+sD1npyYhP2v2nD5QVwU1zjRYxJk9TBQi3h+m1huB6
I3CCe1f/LjGJOZAXKUcY/xe/WDzvM/AIqsi9fdDRqaJromo9lvX6iXU84lvexS8Sg2aWryWHjLtI
xVLDaQdXal6jD5Fu6qHP3rXZTFrCLaRuN6ezx7Sj7natp91/98+N+2D130RJjiPVyKyaf9TqnrNl
yxMGpvz5o6SbSy//GRflX4RLZtfp5uv4dEjQjimhdP4b5iOb0EeyuNnHxMuUYYfj5GGMB0OqKnnT
TMOxWvhzVCR18Ld0QhQvcPiL2u6vcl4ne4L13pjtSu22vQ44LTnGGndxDgZ0/EDf1z9BzD31mdTG
yCmyH05wS7H71fHudAl0P9DY0kg90SaM7p0PuFhgGy86aA9W1+NhbqFBnDPriQK5n2XRyRWaSd2M
eftzwhlVWgPCbMWeIhjXo7JsUnaAXrKpbmd3fGR7n34W51nYwfd49pJ9qeXBA2dI5c5sr4Av57yo
jfEy/ocARMMuOCkPdQqEKY4Kt6AjfrQ80JcuBxk3GbstkSC4kX7yoZ337r2ao6CncujYOfy7gNFK
i2kyUQMgeO6TcduOr7rcrUGFDbXuYafva5Th5UrcXQbjf/l9XbYSePONFkoXhRyxX0uMENFsdzYp
L2tl55AWzExPI0J4oYBHjKdSUHr7Fw5q9a8G75Ucbh3twU1YAzm6JxIu3T3jDAQmFo39Yg6raxW0
ZiP0c1nIdUrzWWIPN5VS4ejj1gzz+qpSX0fC837IDioa4l581+19p+bpZHbVmipG35IFI90oKLsS
68uB92aPnQXb0WKH0PsypAGqyS1tcbq24rbGMRVutmuGMvCAsw73GP1iv9lNLR7ABm4JaKybEsqL
ZNQC6s4Y714ABYOBSp63NyhCRepxIWlC+/iJq2fRlHg8a8mSJYtIhJ2ztg22+yD/QrRq/MKy0N/s
x8DbRuPqbEuvkPAKjNBfZU3zDAZo+UPXXEmDrDreqpSk+CzCEn7V20llVkPKl5xrJIHGUzJOprR0
rSjWxZ4m62v2vGYo6Z08U+Y3K6SKZbTJAUBFagPlq5M6ALmLSr61y77eWl94aJr7bPlvKzhdRvZ1
3z/8S4yWgtVk99R7NimIsWFah92FVfAkhBZsGC6NlmlsaXG6RMBuxdClz2KWjpmmuFpriVbacmbS
u+wm4nWqGl21T5dW8YKQfDdxCqpF9NWj4tWROw0t+354x1AGVh/xkFomRivNvzc6sxk5kwCnah5N
nmXdc/W2OxsJ3wBOh4kH42WK90cl0/g7YQRws7K50MwQqCULH21j6GpBwBaq9uYWLrN+hblUI2QX
GpbUmrurEEXsuFJbrvf7X4KsEhaE0qBgn+xbswTMonaWCdzhiDXMtg+ndHk+7QzqUEVMoO++8XMC
+wrrS2IL6GEJUMciUp6D8mTqjVJd8ftsnsP1PpoDjffa8n0e7VqBzivKFe8V/+P33BeuTLVnAl9L
PYxfuHFmAkZTyxM8tR7NJI29wzAzh8Cmd0flurMl+Qvaog5YnmUSEwOge3jlU/1C6M8+4GK9EHgN
mY2sosSc+VxUXyR5YZkF7hAsI9GCvQiAgKOJRUjdbD6+EIcbxe819SWpquPesM56qkyt2z4Iu4ve
iIEsnMoWhFbK2/5d+LF2oCuBC2LfyaRGkwU4bpoeUtBmPXimpKXa3d+PzIKaxKXP1rd9FFFpXje1
9q1fFq428r4hYT/3LsTxvwTRM01hUwCG+atoilVnRnFCUSgzrd9wBxEs1zuABZloJlp8QYXc+E9I
V1evtxW/HxaUsmMRoQGsj9M5RyOE34v9R24/2XLVrJml67CZqJW0EMIoWmV0ey9yQT46L2Qi8oPl
Rx85oSHzYzThFMXhGouNpcpa69CH760EJ0gr/vKnYZEYSaLoKeEj/7A78BV+qcsGiGwKyiaM8FAx
xpYHGBAt0Qp0F83tnQ1FycUobxReOp+jD2seMAWs5BPqcICGbkjBMUu7ExtKhuXJH0GoEFYtG2KK
1bU7Oo7pauJVdp3Eli3wNwbEXiYnzkyHn+zkhJwespb7En7HEYd1t/CF/6eHG5jc31Q5iXxyPd3n
wZMYfvTJMriXHpixtedZLjXXi+e1T41Sw0M54H/ocLzTrjkrzG6EFOdCTfDNBeh+fpEly/Xdue1y
gPdH3V2CMXJQRjouZ6lcFm80YCeIrr78PXjN9L6ZUJHbVGI00qMH9uxTeC9xzdq5irqpPGdGzRHb
xEfqCbNbpP/wjndb1skpLul8bRsn9eAkN4VBXr48oWaaQaDdWOFtz8OouT5BP3IMr1/T2vISOUES
p+y5uR4dsm0zyB8lZpc9/VdL+W9azVuD2Vc+TJekWvJw2fhBnca2VA3GL4rV+pmPUb7sespW9lag
nMLrJV9Oh/ljBptJ3gj0rcB7cJ4mu9NW1z7qQvSYxWl4/+QKLOEFElZnC1qkt5x0gm1G5HrxIvoR
KsaioV8++1yK6qHwZr/ZGA6qn9KOUj8IW8nwSZrnOD0wmkII2n6a+jWdhLMMwUlJ0lKpD/JPCUGU
ePTBhUyWYNrYdbqDCbcOB/sykDUhMrhJZxBT/wssYG0DQeL+dGM9HfWOfcAWe6h1dHjVNu3yoULt
Hw7KpGwAhKMyQIpxlEipMkRySd/27IIBXTQLTAzoLI3jUoK/iAmBpuyqmzpH5VOp9eiCvg50KpfU
LFQlNG2zeqE0Dh3F2euDyhFuZmiXITZNGghJakAfjjmdnwSyNIcNFYyz7kNGN6rP979LN/75Q8jy
2KWNkELtJA2ggctWLCThLvMAqyEiiSiom2FPU4y/eAwPXxqaMLvbbi0kltmMRWCQWNtSiXmDSWK4
3s2pQ4PP+jyGv2N1/CkrCCK9CcQu2QwGdG8ZuhDwfPuN7jI5pD3hObIF6MzlLaOWv7Ex1ScxbCj9
REYQfe8a6w3z+NW0I55hXMA9mOlwvxkSxmPB3S5aGj5eE4O5sK7LwuD3n5+BQYTUAUX1PJraozKT
lmSuBIa/SO8y5oLe9Pt348de5yPv9Vpfv2mJPEz/m2k9azzBIaYQopZlRfV33z/29azFX86doygx
xSJEq0U/PS+zNOlCds/fw2A+ANh2KWMHzt10ilI0sq05O38hx274Gc0SZyoT1EnKkEdqGAFq/IX1
yruFi8GU+y17w905JQXpBtY3OXzghTYe9N6B+aihmsPDLgOJOweEuepuZpDqm9kYe43LkhhyuyO1
hGnTJkb7wnWjTLE+PSkmR0xs/L71nK7uHRNwFm5S4DfFD6rLeZ6bCYorNcVn2HBKUyuk7119vMw+
AG92ns3M2peuQp4oKWL22oPwmEPZOVFFPMpfFM+lt6emA5loUkyQ00FoYcGuSnGSKHdQgSzs+QqZ
QeIjATb/7RMIRqjH+qk3nr+sEVlr7zBvtBYfrx/MkfttvfDt72hOu8UH5LQa724tlVADulcWcnTh
mfkQwOmSOhSUM9ois+9dCgyTIb+8KYxoc40VqjcEzMc7Zf0E4JjjV9npo5P5IhL+7CVCGnewUtYr
bp5oxzR1Fq1FlWiC/uI38ykh5HVlt+7GQjx4kxac3TmAOLzXPYUyeSv6XI0Mg/GRKWIcI6CTGSEJ
mtYa7rYBv2+9RYZcT9UmQPC0Ied06DbuGhCyTzNAtmO5B5QDhAhuw/3HyB7NFCY33FSNdo6Xdz/k
qeOLmIcDv75KVYJDpC239blSzyvRKAVPf6mkH9wqewrkAfl/py+MGGBPrH01Yxi2h9FPrXZujFu7
tKFj1LNfqUqQ6FDmfnwR86hLhltXNks35IlooBTiB/04SNfWtNFEl9dxukIkWSWb7RCZ2DUJ+odH
eDBRM9mpt3/w8D4s1qjUrIJSG4xiu1mkHYVxfozmks26uRMZiEx7ExipqCLwqZ/wRD0B4mrufCt6
SmmGlhUWPGeapHh8iBKEvnM9oJJCJTyJodHgrfyT4FdBO0dJ11hbWZXwB4hYiPXPe9EGPY0ziFC8
+0goP+UiZRsf0exr/kTIygyk/9GrBtBWS7UJ9H+NOr7MO3cSl2w1sqm9VNy7KcpUY01LebaK+VgF
9Z7qCNqqXD1Wy0XANUjepPzkoW7OkhLuGsIwqvo24yq5vF26gD+RaJl/OC3ltCu1Tn+LLhxZFwPW
0Kt3ZxzaBYxYzPIhtK+I4CuVJCSWfpp7yMD3mQ9h0vDnywuHJBoDWHby1T/K9wmCb2h4MsgxaWWa
H2ropuYb2tcXgwBoT4uW8VFox+a17ivKwTIrEztKZ7/5HuSzJxKYwD7y6z7/LhBxq1HIvGLw53vY
cpJ33JEqFEgVoSRnH/eKLN3/yIqfeJgWSolMy1Vr5WNq/TXeS7GPOtYuaJ+0ba5r3BtUecqNtnko
Wo2mzbv3pjYxJVbyTDsMEMKXQq3CJ6GKUnBSxGOtLAHw5MnT+K5bNRIqg4+eOxE3rirzM+nhGtwo
LezQR3lxe7jVwToPwb6HDqgEwdnbzWW/ae601Gr9WNTxkXge6Vk3f99+9/5lWLzSxeRZ+LF7asLA
MtS1E7UoiIbrkqyHtlDv/PQR9WdiP9pk/pzCN6xNJG/ggAI2dBOcixbvYgW+2fxkTZsl3QRs+C/5
qlfdKhZoGL4HDCXVtQa8QGaXh79gQucOaGWpvhBx8Vvha9vOBk5GAKknmDBdCNwmDyAXSujGvFqV
iMAXxYOOTs9dCAH8eF8C3f1aySIye4uqBhFvfOOJbA0aQvgUw6ENYkoBQKUtN1RUPEKMEBYVWJhe
efRDJF9bGPPc0p+lzXq43lr+Pw84nZe9rx5v4SMRU6llYGD0u1PycSScP0cmII7/9hP7lCDPg56C
x70YoyZ5445tX9H2uuU0kEVbFCcoh3iTTo94+c+YJP2Dx45yXq8FdpE0iPXZBoHInJhCFDsWvVHs
cnEb/VrJfxruus8M94lUk/6Ij8Zpc/jU2xamarqKaMjfFRZ1aYMMA6/eovqKxNtTYrkyHRUa8Riy
XtwSXLuv95M5kHv1D5XIG5hodQr4V+KNL+fokQ5nGCNg0RH7FQuBQKj9YbmmRu7rYI4JX1OsRA7T
OixeTIAYRieNr5115rJB/cdQc0BcH/LcUek7oXlZcFWkTFsSq7Ypk+2j2rg+AYu8DpqLXCa0d1As
EZCYSHYd2RXFCmG76uIrjD65Ypnbp4qkzdHj+Te2VmGA7OPL2FHFljtqP61H4TDuehd3O6qKmYAR
hjJSXali/OOhQlYx678AeN5mjGMWCGk4QqgdVtBNaUiLEnKqVRHlXQrztxUdER9OFdaSG/VT2p57
yowvYX486pIC5uWaDLVsDKbyNbSlbvVXhJ/gdB5BQwlOZelurYpRc8gu5AHWQlto1Uu9ef03MWIo
yJskR6LAGK2sPWsQfZXyYZFaObqQPoav7tJtGsvL6YG7prcIomTXXMqxRNGBzjqfwFNVVH5/c4kP
PpYnNrqtPg94KHctNMTFT7xFK9XWviZ/WF6Fdqmg5B8P214ksuwt/2fwPHF/5BR6Rme809gCbXmY
/RdmSi3xprxA7pmZIjDv+lrdPlBM3ZjnbLJSaKPI/9OpyDWPxDoxiZs84OVUOzHvZMTR9q33xaEI
GPYKrsg9Eoe7/IlUgNJbmjITLHjXUWUE6foDNPp1Xd0QbQCvIi7QauP/dhi98tJXFnlx1h+xd+oI
sTUw/bvNpRS6gTrKsQzA9kOcIc9cvFbI+NdZg0Ue80tfOWEhb8b8GeGZZ/BqMcHtoHUAFYDoDEs0
sueZxzHfi6ek4/Cs9FadOl2ZwDOk4FWKawHdDnIZ530Bkp11yyFUi9YSLEl/BegnVsOAAwRa9meJ
urNvuoMkQXdH9ojUkeHgJrXHgNCEQOvY4Q10XCRGyus2H4+KLyH/L17GPp54j/UU+cLaRDHcWMLH
2mS0+LszegwHvBEGzSs/aItw1MOUJPEb7SZGYfSvBV3Ae7k9ftwW3jbOJexyllcIM2Tp86TnaixR
IAxVSuKycrwddHK6trNTI0MNBG4JnflPpr9qFjtQ2FEHMOC7PSJAu2Omfa9ZA51Vj9FCRPX6gA5o
IpGOwCODyxCCkfBZ+F2jbINPdUIQRWFTUzDnBD71HaA00r8rfbQQON8AWPIc7bAgP5yjZvChz9eF
QLZwpRvnHRwiYcIPwlFhsoHHYM/ND8lrXX+xdlgNCN1RUYJJrNWeg6rxZ0JOUxKYyedsVpLRMf9a
CIhQBngS6vAUFByhm6818EU0wtL2DJ1h/lSVi4+hSk7sZ0C5m+0arQvDqRyHqMBzoleYRgpQIr1G
iEUm+azcWAjA6bN8yAb+pYC97WIIfLtztD9WA/LJxRo9pNUbILnQzlguDzuxNdOLMvHlFnV80HHE
bksV6Hu3rDfmQQTkKel4fROj/13tHvBRl49CfeNOCHYhJn5jjSkuVyYWZL6lLhRkC4oVQ8Znk6Ux
0IlkoDoHFZsBbo5ggQYQegn2ZzcIwNtCyrSi/A2QPSB8QLbdwIDvWkciITUV4SZoW5fa2glT1NPO
7gZeHPlU+Wf5bCN6y6Ho2EvNRsgSuu4jfdM7mQlQwrJuvl/OhvHforeHKS1OyQtQ8Jq3wXFIUDMy
abfgp+HEao8b9sylqnygl9sv049a2e1lqTRiVqzr6y3Ix+j8naI54wuSra3ipy3qTwL8omrLHSfd
MoK4IyqNMRWILMxIRMK5ruQLJHAGdSiwWZ0uJVGqE22fxbM1BCbm0cuNcqyHMkLug5Rf0ueUOPsB
uzLi9MYuhMU8YS2w8kr7mTQuR7p1U0YXRgaolDLxIIQ6h/smNiPvDmMG736OT9GMQ+9QpDD3OmWG
QZ/7kt7hBDW63DYtWt/yrROrkRSy/VRpsRTtdBvhWN19FSPcNcLbdLSbRizS+jtMxBBuEq/dfe6U
ekZGz1r1HkeMOhJB5TKU7pHUC5C3zoIcalGfXGhOH5XcscNhxPe00ZYRlgsQIFqkps/fcTUU2/XM
PnGbybegrg+gyG4WzMYKPl6oooX1n++WwznLicgvHQYB4DI4GX/8amKzsc2qN/0q4csfFHGzwFiX
/ILZCad058sX7RveaAlBSDAO248F3gxNN+jOhE07bvhXBeAAaKeunLzFwEKnCblnePE5H/X7qJPt
Dpe9G66Rg8xgYZUlxezABIA8nNegizBv4LHjCVF09Lr4cMP1SsMNk04ZL/65Z8Qllp4zftcXVJAE
51Z+whk1lAAIY0PX7trQlftpT8KWhLpXPcbgLvNAsDQFmHYbKcP9My13KkH48+8SpKJSrX7jAWwD
CRilP62iC4v0NkSyu2HChD35I+1O6LwGmSFuCL7Adqa2pB2boWDedKZ2dTohxCr4Afk+CnW+g0jH
Y4I0vQvKgQQM2Ez1atMwpJPEYpjwB1rE3K8fNQtk3H2aU/OypPdNRuom6++Um5uDb9mmwKwtayyj
T9Mb7kyZ0In6AOhBSqbQfxD+WBgMM8Vtr6XERpeV1KdnNprF6H0k+u1YpIgUXI0ypE0Sm2uA6/b+
hgHgEH24mx9AL654sygTlB9RJI/HiczhJkOZ0AoZp6Q78CGCaGVVWVFrQ6H74ESLPThCzS+SyNqD
IsmJev9YHAxopF2PUJshwBbnaGEA11HSZ+KhJQGT0CxTRji0yScwi5LzNkrIMK1jfaYcoln8lJ58
1xVoZG6EZsinnqaQpO21aKPrvcir0X4sgFl1GUGI1EoJlY7Cxj5fUT+iHPBgQxgdbdoomNRcNIHt
jYhxxtQDZpmQNC+2d2yLSQVV1VP6QxxD3/9p35id8IuIHk0TyW+8iSD5+SOj2KhvnJtrcX3ZIN3I
Mc33naPgl4fzAJhnJ9LJDXgf2M6n0E7PXrjvIUNYDpNQ5E7LbkfiPaZlGLV5JF2z0S2Z5MFyOfrC
ZDegqQ/IVLWglhTCp2q+V84ua/QYnOP7QkTVSRdYxNUqFJAV5/FSyrdLwXkbN8IULgqYXWTZu4aQ
3u0dp0oRN//y6vZKTchTr77r0k9pa7yUulbGcsUAfk0mZRjB77r/nnVeNBG+zvC4JZblLg8MWeRw
i5gsS0mLac/CN/qKxJ2nCHHFxn8K3YHAOsorm2dNrPrlZBwfVyKteCkEs4eh8D8w6FI1x4H8X/Ja
z3jc/TgZy8wV93pCgZuZtpkWBuouaCLf5GmFAoyZtIkPCH3XjOCa6jTZEcWv1thdVkVZwKnWwgCk
03VD249UJb/mMwKFtnyg2dVB27KLPv7kgfXlWUte7oL0fw6Hc26+GjC/VUDHOMef70W3UNVVY6uN
DJY794c6HPUSaLa5KEYFAVJC7mXaWJS3uEAldR3nUbjKI0NRyuSo3d5utGl6wvll72xuok0Skj0J
LK8YfDCqCQo7C4dCaz3BkyC/5I6ICqeobMF2B95QnFzwQ4imZz/IJXADY6n9AAMjjRbAfgHCqEDK
kDg+Nr/a7/gf7sKfXMoONl/aVrpNJ1qL8l+qTx+JZttkHllFCunp2t7bzN0kXTP1dP3s/iBIHxar
9sljyxiT5XUDYePBfQpfgbN3vpa7kXNtiYOiDVcZWP08MSp1NucomlWvCxJOT2t/yP/j/5tnzpua
UIcYgDu/u9g5uMRXdMmHAqBkIRL1jpMjZHazB6qIEyiQCvugVaQAwB29nBmhd/jzpoTdN4XGgtbl
UofgQpyoUpBf7AO+oJU5zqHffFS8XbLjG5gFYUvsl/mQuKw3vo4OSXi90Wn245jUllAK8IMcbvLV
TLr0dyMD8+Fva1GE3nImxuVKFJMsqt88bm9HXYCBElpJmCt+3Ut+9Uz0P4Noo/2fwXfcynX4Pi7O
08Pp6LFDDcHME2BLFDtCXmDA+LlpcQvv8RgS0WexVntbzUzRIlYy/zXIorBQQ06K1jU8flEpHGHl
hbHvakgRDONzwwZZl+5q5zkZWkRsoTKfBPSLJlAJM1PsWZF8qT371si9QBzl1+QShseErVrzFLSL
Bb+RcfPCPUdfl9SPX8SutCafQw59f8zJQNrvhkhuj0QXClJNcuUEuMwiUVeTRZL1/pY0uV0VTJ9Z
H3yCbkKX/0y4ZYSRNCURgJUt/1gm63YOvXlmGCduyLS80JLCEBPrRcS1bURqqVqdGFn2NaTZe58n
r56TbEhutzLR8rbsjZ/V6GlnSMprrfwQJxGxUVPnNs+IEe4ivtS5qpMHZtq9FsWwsJMh8mIsvtiN
ppFPMu/Xvr/27mlnusqgPSmoAu3UBpPG9KLn0MpFXReRp+9iq2txiIHxQJqsBL81o2mV0/etA509
orPccvXxc1pGGR4xDEBR/wrMKndsWB9PAxMLWIdFA//u0lXljSV4w5BgritOqqkiixlIjVC2KTxH
qSPD7U7NG8vH5kmH0pOydX1y/gTBRuVh1tuv2p2QWboYSwGYYXvf/Dh+RdvCSCJRw63IG9KYLXtW
gv0SxQnGRtcedzzI5VnRPoAj8XXVYotdJeeO08wkW3i8bwKHGPaRC3iFhhXE12hZmg5ITQDahw6X
cupmh/xZ8zounXuZRk7HhJ5VCGbRybZZBK1y0h14A/YtLRYpXG6zBhdnbqbtRqXk7usrNJeo+eEQ
mOW5JQKox0UsHqEnx/+WHfj3eXzKpTyhLYXUeiNKCF395uU00IiafSznUYxFDtXo3HcaKlGfqJio
JANi6kWE2VEcbyPn1d03isoOMT3i25N/QK+jM0etemTFPufQ6kQw5UVqkQtFlQGOcPzziIYbF++v
oRuAIHwp4uMRKnsdYcCFW+bb67vnzvNFBhIVQ/Itodcz5gOYPkH049TIK5DVm1+HtESruGqETuS1
66GtyMMd2wkNh5mxltbXE+DX2oq0lbx+hm9l2dR53QpH4jfD831P5yDTQvvnI5o2Og6QuRe+/uxD
meqN+MG0mCXr8hEoy+gNDhtwRUvX4sPlXF1TQLdpvuPflnWMb/G8QK+8/babJOez5i3lnX6nXmHM
KpQIJOF7lNodF2e0dHGj6llpMqzUGE1zFHZf8Jo3ujHnF4DoQ6nZV9rxyeoUaxfQGC5k+1/2VKpB
2IoPO/wyLFbHehTmdSRXOAQvygGg00iimdl16R4AyoK5uwbnsoissGrPyUKK38p11L69gTj7cNyR
synqvsjt1WCBXJ33vJI+pPTUdauhfj2rFTdBn6fM2JcGL38Oc26Cc43nLRs8togU8Y1ZmoJGkf3l
xrdOrRmpHiU0EVGlfnEfC/f2CBGOXBLnCv+Puv6ZDn8ZA4XlIBnvFU/5BOZvB/goZkfcS5hYVqvJ
WUP70kRuG9c/O8iXocWA4nOe6LaOntAIQZ9nGhgcq1ocSH2RwW4jMVqL9QDA29gq1hB96Ambb+oM
+BilOJpKvM+ihylh/g1WZJv8ciLXbXtDypQKX2qTz2akh8hVZJFwE7Y4TElTHt6vZfET+JjxcvDI
G8Dt6lRV9PyryQYzBIXNSW91THW2Zsi3nlZtaW8yj8MPGEXNrcDZj+SM6iFkYdOTJOarOFnH6eCP
+6WyUJfxixn9AM6iqIPyQufwtV1Uo433QGbI5k+H6G0qL3u0A3o2yu2F2Rf+tCmdc5AvIgZYu30X
RY6GHJfND8O1n2goTc7CL8QOf+x8SEWgEr1khITjE7/CzQzYuDGMRcyFCE9uxDgbotg8T3/pYtji
l+bhcMnFYsbKnGLmcu4d5UEUuv0hqhttSoc7jNYd/xz7GHJcklVBpvp6CgS1t56CpT0wQWr6MZgl
jdEAgka2a/OkcnWSHcc6mxOMXveoFt8G33UFkABEntdJ2gwOQTRbkzHfRXe37hKXVPoRhHUROpeT
6Bl3vWeMNQbP0zLsy4aubxqQ6sEPzoQ6PSeZTR9PDeLgoxZ8VOhbychd1/jBCwyXhtrFBO0xcBox
3PY8ymHoDNL/fgy8xORBCkKL2qXGQB9fWnO9sygRwFh1W/bNlZJtMA79nuHgsGUt4FNCkzfsz/58
uEFQLrNaACsUegtAbJksD6zoZE3Mp67a7nc8m7O5v4ANZD4/vsR+8YyZh/B71D4jSD3V0Nv7MY6b
ofPGLAhXhN7PjIXf+r75XyYsytDuBCxDr88eqZlWgCTHgPlV0J1r8TI/lrMkCOlvsmf2ozT4/UMc
MluTnajGRzVRB+ctzleIOfC/aSnqOFjwrrfraXFkpZEARset3J06hLwK4t2yzEilNB69L/XGMzOd
iynvKFpMyQC2ucJrknmVyPRoZixWU57xgJKHJ6GvmIBAb5PCyGTviWAq3thV8kAISU+xJhNJJj8i
IPy6WZ2PdDeUYcRzUCrukiro2aok/C8XpxiEx1J6D2iI96d6wa6dyc2DCKJRXze/q4OmEB0Yy8uv
G4o1kRonKreSOBjeTHCTVoPBLtAp6EwzP6tJ89kTpScZRWnZaamVFZp8q4rWtJdbSWK3spmiV7Oz
m77LDZ1exeWcwTt8Uyfn0wfsr8NxNATCIonMpgdTXq8UpyAyVTtMJqTnpqR5anNQhyHzvqiq/ac8
Q8hUSUALj5ZbzR5wt7aw2+Ct8ll8vRp4/3kQFmPo/QWpYwktVwwZmGgQXpUiGKii1me6H0zvyZVR
mrO8So2Vp1kWvvTssni6b4tIbtk5hvEMsdObI+/gH7K6g4omWPPGwmRvUgNsm9rIL600k4KviSci
R74xO6gnMbpxW4PrLcBKdbbZux8f2ryMCXoYzjXJYnUNbozhNuCMk2zndpCYjOKBCzNThhFEO7i9
s5PYevt4SZ034fLsTeRKA6vBKBlamDdqicYvLy3sNwqarv8veh556XV1M1N6jy2xFmBEHA5iNsq0
KneA0AZJ0VBV2RQnynrfEi2QPZ9NSA09S/lQNlBZbbe5uyCMskxK7FFieJ8lCgpRHoZTJCKpcUoP
kul0tFdk4aNBiB954dsZGqv433ru/49c3+PnCrf+4u4600bcLHkMw3RZuB6UD+IdPknMOSxnkal/
msK5PEJJ/vnqHMd2bL4mlOnkZP71wbiyVOs+ODYGY/6sYBOnvSHGEXXBU8NxAh4Wg6/QPlrOEUwD
8wrai6GmOLKhhRLfbAnqEI9DnclHCxYlBZVOD7xSAQnAxKDlURAHoJW9KDqrs6OsKh4xCO81U4w/
5HbNgeeRfwNs1pVU7YOn+hbqbBZY78+Skc2st6H561gTYxJ6rMfknPTUT/4QUsrKsCazrL8UKYBy
RGuBrPDnV6zUJJ2dGEE/tvQB7rM0cT8XCWE3c7HLeGBssMcXxX2awwR2onW9tRiVeDts5CvFrqLj
zgP8ucNCghsEwWaK4UrgjPB/ciwGYrFuV4WW4N1W1jVe6j6iHzTUavhDcOE9vEwScEmMUmTmuJuG
ZwohHI/mpcsfbHBrGVb/4ZoftCc+GF3PGVN5yHfehQjJ0SEyK4YHHKueeQB6vuWFq+jcJtQlZPbn
NpJZmFWmNsWqMGI1IeWX8ynUXOor2KJYU4OyJBa8BbtLMUD1VqqvZaOjMsm778wmkVJMu5fQ1y+a
2KJx3TVzy2s1LtnE9eP9j72XHiLEGSVZKu5P4uAc4HkcXh273tTojCILWH9fMDVOwh1qxk2ga2/Q
rmg73EyLL2nsmRAlcbM2i4EhXf2hSRnxZcsw28+uYgmTJ+OmmPtSSZzY+tNlbB+yC3+n2VZNUuH4
5B53A9p7AGO4Oqp9KhwRexHesg4BMKAqF3C5uv+sZY2iIGnjQNGM/+MrAumVUHz89rYaUFJvFKsn
6J/TfNRTtctE+bESUhoWO/0c8Hq4pSFWEuzCGdZZ1Bm4PP3DJb/j5Wfti2jdmIDMF60hGyIqHq4m
9Zylsys8WRx7dJnsvR4wxhWgRC0vPAShRsl48qauSyHAoEuStHfLXQx8MQhXWhZB8VZw3SFZcwP1
uXjUMUQJUw12WGBRlN4dlK+TiTKG2DX+nlwiAlXY46fGrkSOfuXxBj72tIBNXOWn1Qs08QBfDt3P
HkfIAaAenxx62HwLLckqwq01K69wlXV03wXgNt9S0LxOf6utuFXmTMgJrjS9ho56L6LVnQDMV7/6
6AO9KJBo8BG8CWYLOtcxMloDVt/1TUfUDhunSl029dThVlwp2s35Q4IWlk5lFN+sjAy7bSdOsFpP
OS32bfYEdJYUu3GAAZXycFMYFqN+F0y9IzfI6zDWimULZ9sJiLag17JPTPyEs6jKlKIIeFamQV8G
d1cKUvNeNzs0WQUWP8QrrlCQVztJVpDoZDclGP5SRZfCC8dAU8uqAJfC4xw2Of/7RRaUjbjQQT/K
1I9OC3NDHHvyd9tqzRArNrXslMkfuugxo8L/B+pzdnDgS3ekwRjaNvT/AqCmvGCMHR811IkKA1ic
4Dhf+jLnMHlN3uhFQnH/WziOWkb9lRfnTlS/uwtsrHOZ0XBCQ/jx0uz2ZcQl03+ZwULdPE6FhC3b
E4+1ePGdQYmZKnsaIVN2a3RGY1WyjxQYwolSbgHhDwLbJfhjG+HFSEy9Z1Zc6LsQtS8Y8F/nUm8/
y+bQRfhkEIlE3UY9BWkHvJGZbLQNOtOcxc3j74M2pcrVQZnedBaAddkOmeI00i31o0FouNLJRWSW
jfw8/FzDtwSI/MMpNoDFlJPnUxFQ8Ey+WZebMj7mCuWNbk7XQHNBVtQlGPSGTd4r+bNv+v+sX749
jr/dWh2pKTM6zWuEVt2gZa1z9BpcpQsliEJsFpGE7QbyuLMoyRPr1di510GL8ze+yNm/YbEUIvGX
RtJa6EkfKg4NTiwSyN7U/sBRhEPbjQZ3CJ6YKMMtvBnrtvm1YEJM/hCceVr5uOJ4Df4AKnrwtyxx
/89lIr7SdNsvems2IlU0hwbNOv83Mmvyxu/NcIuj9Nlc1FBZi/qQRiRrvnzkl3Mbjzt5c2ez1ufB
QSXV2ZDL3tB6VAp9/NHlQ3bKmC/T37RuI3ihLC80CP9FUeYyLqCkULArcCkywY3pfSeSxmBQ738K
D/SPDNo/7+dhaoRhYTXrpF8yjqoX/Gd9WyaKmVp4hW14alEfo7eQXLVvrEikht7mYLfvo4f0j3hy
CwtpUqMKmPCvw2+OrXFjOoW0dcXJb/eNk7e3LK5lgkFVOf6VdZh8pMSGkijGtpCzaJLAIQbSS+Qh
rNpuUMYd2hlRP1Gnef6/XXcpzixOYeRiXvXV2kBtR58ZwGzsNmHlCwRLJDqgh8Okghp88+HFyjbh
s03WkxqKexQ+t0+Sc1TyVZibuVe7+noYf+fIHb7OyjecpZTllupyAxlVpARskzHHEhAcTohQBl9S
n1YhnKklfVMHyOguOG0bai8LmpJe43GgwTEPBRdQzMY/xmCLc9YfhGf1Kf0ZlE8pLPCjX2gVrKa0
VPCoDeOaLUTRui87RXPMDvVv9f4lOVMyeGbJ6FsU4tPJtWeNLFvoa1VbuUAzWCSmBNXEY/p1Xhg9
n69LIAsTd8k2Z6OiZDBh2ElrsP/0rhTSb4Uhr6x6bfTihFiOylSHdfGO/Jo8KrZc8oVotk67NiNP
UupBL0UBGejO8mPbcXCYgzQWHMPLA6dHhm71C1Q5SOVrK50trNPWqz0+efSVt52BNLNqP970jBSp
HupnrLB502/PO/NOBWs3VwlqsifKQso62l2vT5AO2FYJXhdsk3HuggdQDNzfWoVWUTO2aHQHVztD
4RqfQoZMwSq1fpsu+H64JMdVIe/QKYONwkmNHegnKXRDB5vPZkCF4mC+nKeB2scOv4sWoRJzzbbX
zYlzhstE/Mjg3DtL4bZZ3EBgMpvVMeIwHM1GTYWmm4yondyvE4aE8DxWV3Q3HLICxYV/5D/XBu3C
7bb3yx707nPSX6L2nlLTLnqMg/35SovfVjjZ+6z5rrIzFf/GFrUyz45tVpXGN2WaW0czY6SJ7JnF
NVLIEilpjEFOX2DLPHzCYVtdxHm2+dVXuaOQU0m7GUij/tYkOgjZEN1aRZLn+WBG2IbbqhpCtK1c
w9P+JQiJw5fVvjTV3q4EyLn8kw8F6I23Od5Msp8nXVn/LfdSlcTDucmqO9WQhWWQVn2eN5Oizgpe
sII+3GxNQ4N8nMg0qcLVFFso9RegxYBr4r6qYyYdHD3z+sJIKBRfekh6k29LYJkr42xiSbZxD07o
BUFY+PL1Obdv+RXhXNXkOj317xEWg8BRoWIbuspZRa0zlw5+kVRxtxpRYhUIDjOISrprLFt0uyVw
93Y4mdMn/e8Jg818FeeyPLIb9bjbObRGcMQAytjh20v8Nc9Iz/qtgl1UkmdLWCHS21ur134ln+nh
YEjYMsRTB4P5A0BMPsPMkjvtwCGc5J5sVFdvoAWWSyM08F5akKNPW+0uOEOtyzgOgHJ0k2NY/Yl5
2l3ko2KemfnPTKXnd+WHxDkKgNIpHIDbP7n/W7Ezz0d9ddVeCKckt242y/I6va8YZ1+tPeVpCiT7
uN0UHlJJxtXvhv0rIHuRfpYlkf54Ik3V49Tyc2160fP18ZXsKN1NCxO/5HOV6xd9Tii6JJ2wox3t
yuW1iICWnqYYWW1qfNFTXXpjaI7IqJ2RS+tBYkXdyJVUAqrh5SCHOhnlRw7KBCWp2XQQBAy+vV0X
fADEJzSp5dabWYahkpc7e+fQSKsayv9MQijNv83JX7Epr5mzmSBrBLjzE9W97BGH8cMd1LfvEokd
hyFkjQfCo9R7tdVFUOYRxn1N5HzjD74bKSe+O/1FA0arWwKJHWKstItuFLbMtGMjh8RkA663qS7k
aFpvbtyzW7KG/bf5d/hknRqD2QN3bx3nAhAhT/IIS4o0kVebvebjDGNBUnCYCk2Sb3Jd0XhprQv/
1bwGGsyPsvSb6UeF7LoPIAym1zO0zcaGzH8qd/7EhOaLEW66nAEHSL40pFpSKaAIeY9xkrOzOBS2
npL0na27z4YGXzmVetFA+AKtuK/DC7ev8BD8sna4yNsWyJ8MwIRIi2JnKTUXwOJicDVUXv+xYWuZ
mjvxj45qh3a9rQ9vOaWqbK6duiDPXtOV7ybEApEXBBVV7O/TNdblHm7vVTVKxTgTwShuc6CiUhfc
dr7R9IGpz4uw3OBxst1fsz1aP8+lhEZsMpE4tw23aAd5U7i14ipwDDYwN371XSWEi0W231wYvaN1
4IJFpFAKcvAHbsNTBnkbYrxTBvAh7R6DrwZYynLUg4MySyFDqqlBcQtc6o9xVyxX3bLQnXECnWkZ
Q2pvLJTO9DHQfnF6Ju0+edGrHmqrMgjqny0XXFlhEyR7DLSnWsBwiW44MPilI0KxJ4jeglFgu2I2
LbPiVJJWwCWWUy0yxgkZ296Sa8jNYex0BqIdzRr5UlsI2gPxSQcEmQWpmGxMZ8fgijxYxFPDBUCo
sxIbEiV08h4kRkBvua8vcPa05N20Ri7jz3m6k8eSYHlh4FcrXiLyFcI9Vl7WJzNY1p6j6vC87ojC
ZfRSOXmXUUu2GwFV9fFbo2pxNG6KtOoykygLS/lCvo5RLideemU52TCEA+AtWbRk2meOlI1ybrQn
QRgsNj/oWneOESQON7CRZpigr4zUQ79mBM4KMZdyRM5FNtml7upjTH7GBLIt9svmgQLEQFq9pF1Z
2ihz1ut8fe7rhUoWHY8TLRiUiHG62i6nrut8fDVzerJjAAwFZMZ3Snm7KIvQwtQwTdaVMSwacU2Z
Xef90hmlP6BjksqpA+VGcTwx9kwmNr13pSNilSyXcsEm7RDSrwbJD7uHJqZ5xLWYHGiOGQuHkBZa
KVi6gKykGasRAu9W58GnHP42UmL/lMzjHd76SiAIGID2c7R0aHR6lXtLqMYjGvURo39pql/JvP+r
UQzSYTOegpc9dBMFMZOXRx/mpsUC6UMt4Hh+1y/FmviX2O+8c5FTxj2Vg48KwvGL2bSE4E/szgBd
xuogInAPbxMcdqCMn1ZQUYL8tEmGeBWbSsglkpruZkvMUNMxlRAN08Stxnf+BdnxFEQSrd2abiQC
iAD+brgWD3VhAsAQ67DQE+P9d2yYpoC0xs25N8GY0p8x8M2UsczfCiLT5osX1YBDSdyar1zEdHz1
ahGyYG9/Pq0BVvyhVW8OtZ8SRXT4HQghjH189DKBaku89Sb0LyD4gRqv7Z0tQ/mQVksPu+x0TYPr
sbWXnPNZGY0C5TenDYuWbaGOnhdwPKbqOOLnPXRLx5B5WPPKf+ZfwiES9J4WmBGLjBVk5KkhJv8N
nkotHjZo1/tQvtjs64/F5FsaI9dWGlD3ZA0Q/NTUAm7iKZsmMujvsVoWsBD1GPSGd4WtDtZtweL1
blPZtVoGcrc0IOg42bXRNyBURs4HfzH99AIy07gOhzsWve20YuqZQsrTCTC8PXdVZLhIWAp5pP35
yyur9VkWWiFr9iVX3WiwKhLkPU2W0cj/W7rf9QrvWaJ9qBk1xZW7CA8/25m6iBkT1l7to/H58Msh
iJfZM9S7k1TYFaqofOcqyScaS+gaMCpZNUY3Ygs8NUtqwNl84x6Cd/mg4CfmTA8MaDhpO4g8MjH8
TfwEWgb8OCbn4zLCRajKlxSgPwG19nDVwWqY2vsfpd37BqvZ7EXpYd1vycrXr9nHUZ2ORCkMTHZR
FO/veidYEGwGUbspd7TY2ErDiaDVi/2nrMpYTDiAMu69vzgr8PvW64cFQ7ZUM7b5VCE9EeAST51Y
BLttFWZSMY/lWMxocnxRAV+A0ObTMjPdy0k8mnraK0lcQoSFkiCNOF6rtlWKORAo/pkYj0hy/aWz
aAU/SJ+L+CJW4Diix/zEC7tCYryIIfAPivhbBmfxklgSaQ3BhTVtZgS7EBwhOue0nG9kLtfZY8GN
CFv3syEdoRROnfeVhossyKnoIjqmc3H8dLHXr3k3zwBklNLQzNGvXpnA9r3+gUcnfi0TSj+WfUOq
agliSiLyul1L/rfc8Snr6XUYh5J4XncsSvvDtX8OnzztjOZyoBEYLwjFvcx2wPq2II76w1fiHJRy
7TQyD2J11ov/fJp6F33MXDz0u9SLCw7pi1qCKTO1DBApnTHaulKkc6diN06ITKGNFr73eKiB4QLc
7BD44Ae/1/zub78ZoekUE+Lzl2xqGBMkMVs6sl/xuQVPTcXOpHWadjQ0P5o3t8eJAAAlyDGBWOyl
63Ett0+bHFpKNWoTXVt/734ThIXYXbJ3QeiFl7G7oFRCnGpi2kpbi99DxdCHrr7uuhOrsYJa7Uyl
KTDj3hT90vW80JIoK1PsuaaHb+B95pXqFwwWEMpFB+0SklmVcGpAu6Xtb1p+YOmIcZ1Pp4nEyjlz
plxD0VtiYismw+BNDcs+OEIB9mL86DRW70RM7iXhiIJtwtjFE8IV4BHO9HEL/OveuEVe8Hal3WMn
qVyXBwCt+CrXT9R9ciQ7zNOooIh6YSY/tjYhj6LFuIEKrVGNP1rDWtnlWaNJ/8BVlS3BUVkdR9BG
sU9epCXYh2XmdlvtpEvrOiqjgxTXT67tlqURhUUqj8qgx+k+4AqXoYvMaex8hoQnUYi6JheOxGh3
X8nIpHZE/7eO0+oa7Z7P+XtmH9VVLf8+RcMZqHDhgxoEz8CqwNrD95SSN/x0GSy5A2GPFVWwjvgQ
d3OxShOcNKYvJWHbu99MHt3sJ+SycJh1YQeztjf7ykyUcQ7hblK5Z5oDu7QUHpblV3AxMt24+Q0G
1EE/Os7P7SknNw2TuMf59f2y3nLCPdSqdWezD5NMETaG1SylwWc3C99R3IFbTaiutTJF3YACx6yG
e2oTIEPwQ/YNL0cDsRIEwMC/h7qp6LQUQTN7d6ZJulH+6pHMbd/G9y4dNLnlZAcn+A+EFdb+aGo0
4QUR6TACb9Aka23a3G099AZRYFNxsejGZcuTCtJXCtcmTAt06mxYGvC8HIywxXKwDtg/0tODoQcm
wlghd/6XTZFIUDqsAsj2ETbF/vFSr4/RSPX6ioTse7lRUScz/rjBL/7xbbPialIv2Tb0x5cN4jsN
dPuJQ+0XhJtHsfnoUxIkck79A4RQLy9zpI6YIGmmltVW5V2sv9GWO/mslgWlB/i7xFxL00bIDLQq
h1x/PXka2cC+6n7Q905R18IUWjc+xKXoPj5tESpShP6ET3JVo9aIEjgDw8u/YZp5JiUxWKR3z/tq
2SkkCo5HVWHDWoQYDsBqNrvie8fdK4dCMiBkg8/IHSQHUQdiINbDd17oT3jWOy3HN+gseHCoH90R
NoHepctyisO2ETWH9BfIQyCQV2+b8ira5XDur++Rkt2i42U2lyfI7kEetvjqpgfkCq2CsArJRH39
M1Ns8jLY6MxJypofkLbn5U4SpK/Jx0KVUfdxOv+TJvHAJWeHsOCSbjx7FjsAtPJ0PwAwC++D5r3c
Ja3wgWd3JaxOAqDCSgC4jVJmD08Hxinpnq0/4e+7/wQnlUnpBAws/xLUBvAPbEXzGNaB/VpLmQIC
huahuOZ0mjS3qC3RfFVxmIURVPyw/w+OCM4n+/K07PUAJxhxJfpOC2uQoqogjUM8casesoGhlumP
gWXVpNt6oxtHeZNpFpC8TnYOe+Jt76pKNlNKKMSx8Fuuz9n0RS4P3EiY0NWllzHPFEZcRxiRkyBI
jaSb7vrTD+FsVWfpUN3IbbavlAq5oXmVPZxHtHyqkAEmiCIJYrciUP/g9Z0HPSQhThvervyX4i1Q
Om6Qog0aNkDb0DoR56QjMnf3QXTMiPI8uwtlt+NanNCxUDYn7RMjEEVxoPr2fRrSRF6sYpc59F0z
7dU7ROd3nSU3nMahxL3cOVkLTJbEi+jC1jmiyCHcQkOQwEoS2WZt3rpu+7molD4ZfLu8yxJDdnCq
fUaEQpMKFvmSAZH3F+yoy1JjdVmklcrd7k7QagoKKiiWG7D96MTbDl/jvCx4W9ADkVNcPZDAxsKc
rlz+pVxLT/yPdslipMM8+0X/+TDTMjVA5wb4fJAOuk6FLS9VS1OcHTFl6OfG7zOuJW1QK5BQ5SAx
fcJXsUtakhfUrOmsPBdPirpgUByzJo3wxaYJiaDoGgFcLwOCeolTiT1TV5ZI+5d8026/CXXEv+Ds
IIYhWKr8uFGYMWKXBXKToaS8+hQgDrqs8247YVB6wQ85KLKel3KmucDpjgzDs8hJNboOliQEagtV
e1CyyanAYCcNN/kfCcIhxY4cp6euFGcfp+I385Q0hsT4+h/nht5wlBXl7+HTpaG2L2l+JTZ6ms4n
S1nvcXcjqrOTs/QS6boXtcQMdjpw5iBBxZP5+ZiMY3OTpMEJ6zDw0fIUh54LFguNuh2vwtCm8ILh
bFI7kFZzryUYDGVoUg3HY0ArRqtwuZAmJILOQT2h5skaZGn9BZbX8iaCf0XDQ2NnF4hvYBX00GMW
0WRKUbAHEjoZSpaYLCWyaRzUbxd9HRIsRp2rPoa/q2p6SIBeu4e0bDYEegCjQsUVDBOgkjc7CrX8
zHCNDTzQbCJfBtWlBYaLX+DhP3X1cLJcvel9jY1vXHzkUplQbIUKpkaxiOAEZEiR6bQQPAUHHlWx
m9D0piZOOxnR/r9MV2ukryyeWiLCefVYCovmBfhsZ5wUWUWpkVplsrvNC1+W2REejdsN4UiS5PP5
kH+yPivaoZb6KBKLlX15zhgilYPNZY/Dje6IcvTAcsv9bV9SwsPSvhWavWCP71Q69eq2WRH/I15T
CXQkSJvthOmu/GjkuYougz2+F653+vhGjSC7qAyn6572oFzraY4x/VHYWiykc3F1y3KoVEp6ZUw3
kbmj9zyTxoryVKd8wpcdifeHZZ8hF6DSMjRYA2DlBcPE8msuXY19BZAoZG+lZH+TzbhY8M3zAkAa
DbT3hH6cCVZLGKC1jdhVfmjYHc1sjjZxcbSnJRvSPSDefLfGZjjXsSCXRjYaOmcvAPLZQkty20QP
J9FhUXd8Yhmdt8Okza/jlRfT3aHRuTMh+bFvO5iA4MIc95XdqoVOgm36StYhqA0PlU0WP6utxIxT
6eJQpG97BThVlAUT19iZEmPov85pNBG7tBTbvv/i1nKlEgFUznj4ORHGUKAFNGB0NVCkT+ApyPNH
Wkk/vB2gzyoH/ZNHFqMXpC+VsbApAOAtWZGyPZeFxXbVL8H5DOY9txxwS2NcJS/2Fa/CBQQYguVR
QrWNMkTFbN9BbeSARfrV6QlBdu5k+gFrW/X9fuCllsBwCDREdes4BDDtukmSykIpNpbXd9kLi/wP
wb1gAEpuxz5WJniW2sEN32uTya9BF22HhoNVgnHpBbZe5B76gUS+cbv4tbF5gLf9kZSLzQSzhim0
A16oMzDvUL5Dd2KONGSEkumZ+j33EnnSBZ8XQ2SCXic6b/rHSB7A1RvUdwciq8AOFLSeCQZBdJ2i
MXb5NgZSdv6q287S4/bIESCahdDv9YUk8v5O3rFBiMLCRbeaFNvaDVQl542Nj4mDkw7vkGq73ogc
0O91SQO8asgIq3F5NDXqq4W8no5LUR66GIrBM2ZlBGL+nHzP8Y//3mRCyiMGekJFZ6G0PiWVEzIz
9SIfrss+fndVBmC8CpxnVEXAPMedIyMgyl6d67yqL4DQ22F0FdOjwodPyWqQ6ZKy5YhveSsFDYld
t9t9cOLJpwAa1VTTYZJk+SiBqUIodPWuhfGiJVgx8IBqzxWWtEypEW6b3lm8bmzNeFdoBGG2bilM
aN/Yx4zc9gytmeKHY3vby6E/dUpY2O30r6lVyO70hGcPcNfVtKUaMZ6Tdjxu1r0X1xKq3l1mBqA9
qDZ/PATDvzFTLpNTOPtQyNG2osSMY1jkrMY8xSZ2g1k3GZcLa3eZ3ymZ6o82C6R0FOXILYBO13zS
vYEcdzvOTsjkrcI2KM6SND40vMrqsocdpiPLghRpuRKc3muEWuzovlPtlL7VuQ9Q7FBXCxICj3MN
kFAqHSXa8ah/spEB9QNmaQy0JHjPPL/4nM/f7yW1hN1ZUvh6Q7riPlgdKkYeeGb2Wg+16LZbQtFU
2C0JK/180MA3AoLQUXtGRRYq6+0sZbTO/9HijEhGfLCzvj469WrJIPmUTSK70nPRoDN6zk4rw9MS
Qb3vFy854YVfj7ZmhEToLkKKVtlpUBHEUbeQ+y4GR5JLnGJFcSr3dYW1qyTBbtY66JsXvkwQ5NI9
nJ4tUygQmIcrZxWYvcU+Rs4omQok8qsqFOHut1hKmTR05BHeHQY1jYZTe0QlQ/au65h1r6Q46qLA
sDz+0MzXHKtDDs0mKqrGTmsKD21lg+Kb25691JVK5/y2z1+vSgibN9KPLwoV4i/WtH3AGLeWlwKV
ZCcjhwmHGpNWREfTjTAjf68m8lKb9TCK1wtUV7q+V9mv+3mA5LZcV0h3RG+n/CD9djf5DhqZ4i23
ky5lPhyoVejQzK1xG8eCyIuhJsPV0AXO6BCGndRdS9YCuZh0PANzgTe7impYXyu+Yuw+c/Q4coVh
Ju4jM1kWvfxMOZbPMxTsBpsc2oQafOyBXAwm6UDUXml4YOO3Y3eTCivEHKddTYrGgrYacDZqqhll
8P+hmBuXMhviAF0+sBjgIR/7CAxCcrCLXV3is5wOFgtYPuwZ8FBI0mlXPmy8TwCY3nkghPYij84w
+HIFP+utTuQfpeZgl6TuOfclZAEGYZYBJMsLc90ijs6d7Eq0jtkAHEE5/0JJBmGZV//xFmuCam5p
I1LnI7tyqSeKFsQ8y5A0WD2F6kXifxjTRHQi+ALATLxIzFeS4OMa3e+sS8TNN73/FpcOdgnrJPbr
EMprROzdBWHISKPfGW90AzcrLJzYvONaZSdzGk8PWHoZepKRW3/bv8QXE7bEAkwN3Wptl4nMIwdB
99AKFc8/Y5voQUURvkQy9wgaQn7qko1dXHG+IVNnhhdIpPvHWWHTUP4KLr4lpQLRvlQqN7RbYXIP
qG4gel7hkWD0WvKR2fELGMWZiJ0YwvGPGBMEVFKmVBVpLopR20IsPolhuPmVMXZCCfmf2XJZiYVm
VEm0eEbQJWKhG/cxHGqbkvAdiSjE80N44FW/T0LxvuLj+jxMzPTk9DKfu4DWwF20CPS1XQNbfvUN
fYvx4rdO3r0rO+BuR0z/vHZ94B1THpGmJu0CPzIWdGPdAAdU0T7BR7b0kAbiATnQ9Fp+lBX/GQGN
IRHer4R/htBEOg/vIPWyfKUvy6iieF4wzYUYZWjKZxZrlXQ7PBAGUHbCegu2qubI9BQQdDE966J/
0KceNFnKxsl0Lc9wyliIVIslSBs/iyRLlNSoS7jdCD68p1IoqkKbm50O2WKtzzAxEd1v0s63lild
QpxZNfYNKDQT2ZdO5ab8U408wl4PS8zpIaWRAsI1/UyY7wrlCq2ThCAqSFTUj582FjmuwZHCeqUB
s7/25d0vT1VJIAXNfUFhXnWMV68bqvWT8w2HwPqes7csakQfcd23OF3yC3yfA7PjOOjc4SLRs0ly
/X/OkUYgqxs8RsRM8XiOqjjwmsvHQyzjAVDKhxns5Doz3phhBGGb6+Giw2OgXJXSEVYQ8yxBEThX
FMP+Q1hjW0UA/nejPUgnOY1C6wG7wRgNBbKRhnw0LkQ3Admpr88AbWbx/Q/mn4Sm6EM4RMlANaHn
Ya0GcL0RuRW95H7GcQ==
`protect end_protected
