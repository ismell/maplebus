`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9qS3t+34Adw3J7tzEF6mdxJrAFan02fIUr/4xjQbFxJztYO8Ss8efJfcKuFdSM+KgMwDxzut0r7
7wUKes/G3A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D0xSMGVp1kA364gfEeBgZ2Tu6iS7kfQ4zOA/16+EvBEEf9d4urc39zBLLeFYyI+kO+GefLswguDl
LrFagcSf5vM8HJcQXy6nYClvbBVol6lGSl6JttTC7gD4/KAPOJ9yJjmDse6Pp0VQLeNYVJxO2de1
Qg6YvPIP0TmB27TZpAk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pa3K+4uLLYd/JDdKM4dKTIzHVhp55BgjObW0d2aXf8oi+A6zi0d9p/h9InG96DGGV6OGmaF63M5r
D/ZvbKf4SK4g2ygA+6wzuS6HnosV8Mhi9DEghG41GRMMmBiZ50GzzC8q6+Zqvd36tXHRGp/XJ5OG
9UuHwOAfHyJYfZW+670RVCanD8JOUK3zfJGORgc738FPH2ObEHJqWarl+/7UazVnUXaAqPgtVZKX
AUGFmiTmYaBHnHOBTywp1a2T3SOGrs0lMoktS5ia63W+4QHt5bQNGaWhQyyYf2qW3xwAe3RcZYhz
iarzMT5YkN3/AiuDsWYW1nyJQFQ8RsGMhksSMA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSCz+VtGXT44NsvPvXV/l048m+nIHbFkEqlytyRY56VQ5UwFwh0Hq7ptMEPECN4YBKpjlQaTv9fX
VPkJAqzm6fQ35ymXEJsK91Rt7JTjNeSC54vRUR3yaSVnwF5gCDaisyPpXt2LhaTTxLVX3QW7Tq5X
ATruKUzAJXwuE8GFWg0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zg+/is1koS4fIUk7L++MHC6v5WLMmMP8ErlAst+jLhMPnoUEx9yPd8id58awwI/b626nA22mGWMY
Kl+7LuXpSSz33I6sf6J668LCCwgloJXoM4d88YCwfHS3jBFOxAnx0N3jjSieb2lxDgO//zri8e0G
RJTduyYmXbdelOjUXLV13VxxOTYMxwoHAYlRD0p3dozFYgddWp2OHVngKhVWR/jpijxUT+A/buTi
lmKCpTNllXIQAjIBAPMlQYJfCDaSSPZyvRWbfgPgNqAzGuNReZ3Bjjpk2Zx5yZV+xTXQJlwo1q/L
JL/5jIhwY21gO5b/QHaYV4ciSjKfcSuU2KDxBA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
0/4fBZsdE2xh9wJ13KHLYL1nla34IpfgL55KmCEOb9cRaM8gVmfCmm8qKh9im4zapCjdIoJBUeA9
DwAid7OwQCw+x6NopLmry2GP2Wf82NgpOIFSHF0Qo8mrm/q0ZXr6H/gDHn78Ix755tuLis8xbM5R
9IjVtYqSkk8Bg7/k4lN3h7AUca05+D1VgUQH9mQUt4HttTLkJUAnZ82nmhfkWKqPSbMI0GxWopoO
3h5Yfem/9zWYtMcWAv/SpoAjtFOJKeLvvVMR8KBpHdxr+fGgoQV5c+RxxUaaggS6BhnAL4/b+yRD
ELClaYyFMVj1YKAYs2WGi4WjVnGue/XiHhkr+njtzb8nCPOrC1m3n8WTNTld3xpJ95CD7ywTtBzs
neLoBBQ3Fh3xxuQ2IOQNPPEmOR3bhkApOYmlxL/TD9VuB6zdbo8CreHf7tOg7YdN0DfemrMEbZ/j
PMVMA1RmA+jRnvXOeRhAV4pCg2QoQoElKTBOP4sfN6v4aQMjvEm0wCr267mAl2xCR4+ghpblsXIU
WKEERhY9k/UQExwSmoDXUj1ACD5EyhAto3tTG1OUplpgqS0t08Zoq8ypxhuzk+l6tc7+KRxDU464
pNBxcASlDHXYpNX/qzZMb96i05kbnSyaeRljOtUaY+7uAmjC362VRrlIbQahVTAVyLKpxbZ38pHd
LMZAu2pBnGAmuXxEzHMfY76uBChwab4S4pQPzgjhw412OYZfl8xJTieYa38xZV43R2Lr3A+ZKvbK
KV+San71V3TnREFagiWONdmB4LEjAR+3ql6Bcv3h2YpHfgc3i3hs/D2LnlJdM4EhZVIOi6RVdRvo
A1gFSMmjOIQ/4GOzJtOEd4unQvTD42IyydLylohgADyKNFzUP51hHsWKec0BtsAW52LBd3z58Wel
WpI8ExcSryyqPQ3GObRuxSa46sYLI6tZrMul1Gjig1JEzpUY/L1vnVGFqulbBRaxLMgR/AL6382r
UgC4t+1Tdmfjv3DMoPWQUQl1ebVAGcAZotSi2W9Bn7W2hhz/bNCIKlLlKfh03cl5Gkn19D2ogHgM
FZe/Cr5p7DDlsl9RlvoAkXalQKDSRCNNUkGltiPI/4dFHuEqGRM6qs20cRtq+CW8fFGT5C9wKtwL
rRFD9TSVBD3JrfRQv3KUBPDbuZr+rCwH/yZQOhGiyrN1DbyOiltxvtfMoRtMeas7UxcPV2eD/jl2
o4QngUu3M/+0yppDeFg4YKd2kcmwCCVa3Y2AoBdifqF0E1C3Dj7OyRb/EwRO8gEcrVDU4dBYc4AL
ns8TG5uFg18uxQHuITF72pkJZFApZDfrCV1FSPxn/b/eAf8lbR0yzYWJoMgBMuOd7nRxqHI5Qln7
u+ancQRDvFeVOvOZzYJuZ8qwtCMnfEsOM+6UBVDduOG5gKcLLTb/nPP06+kja01gBZZ/vhY3xFNH
FubvmWA3xfzUmD/ppM8M+GcAfiWjvC2XK21fKxqps2gHZCeKTheATKC2afbIB3RbAWtzaH95cEae
QR/Neq8uf4OYBmzh7MXSrBWxlsxw4llA3YT/OnbKVoyVkXzM7YaMQ+ZBtiP4sBMby4vJ4S2FTa8g
D1Ms8PXZn9+3nIlJQX51WeU68ciV2O+3y4p9u0D6E0da8o1bvfGt0mHkEPVNhaKMDFm67K5uQKBL
6dlgkOmqeI5bzkoHUeHt2wTwWx0EPFtvPM4TWAX3buTRLkmXyACU/zZGwx9RToKQnkHTi8Z03nWb
Tdfp3VgmZ7Jj+gpnOiBnqVTkdOoqmGWDICS9+mme+AZgpeh0XV7hy9Vjzr6Cw9tM9lST/JV941Yh
CixtC6gbXqfq6KfA0q7tpfogQb5Zeu9PKUFh//odw1jOFS2VspMwHSUbrFn8wsXdlnNUwYvvjU2W
LyyUhsc+IFeZnn49Fs8wgtHa5Zo6ZUjbMqg05tl4qaSeTYTeXOeq0IE+22DI+YbK6XFF2UUt+34M
rNVSJ8svykfjMBXloUwNWDB8VI5JCaujpYcSzNy4vPYPDOBRiV3EXhnX7sN0vRAK7NwNF3of32zU
7Sgf2GJ/DMvzbZ2TZqMET/2E2+3p3R/HpRbpjR/6HIvt+fnmAVUf9KKSIazFCFTOXKhyLy7E+7zl
gcLss3iNx/VeoeySUNVQNpi6rKTQpLAEXNm/r9ZWj1YTXPscX/WY1xsTdlOXpa5Wk6pVSZhrGjt+
MP3zfm983DAC6kMmZExI5nak5ax6UZDrxfM2pU7ncwnzFlVFvPJYZ/0WFQ4G6rjZy6o7D66/SVei
B2Jdx/xOaHqcLBYfkipDB5j9IX7V8qbxRx/RJjunIdbduTzejOalqbT9hJUgk+ebvTos6gK6rLhY
Hg/e4Dn/gYzWiXbwtpsXlXTsz6dS8qFmGfOnBff8CYlkTG4lyfpguWn0W2+qDf/I38QlDw/OLlRa
m1flLIztcuOQfWLuL2dllpqqB0OURG5BgmEXOk3prELxrhAjPsqbQefV+eXhXLyn3m1GB9V8lhqd
RBaFbv/DFNDAM7WR2uoCSzJfE5962EFilbeet+JTbz4W/WtcjDTt0d/g124lRtYj9IXhR/fgk0sp
7Z3PNKE4lIi8tnzY6tbzTzWkwVDhaZITSz7I0nyt9elBM6FE7nLRVwFmGPur/xu4XRZnOErkaztk
3EH+p/Jg1A9iHQLz66yjuYISw9aXLM4d8MnvIr9rjfwcIyEukWmIWDlhLFZ7/aGYY4EuK0A6WmxX
y2CGboa2V2UeCgYjoNnosAp33Xu2W/y6YWUR71RgNuhtPTofRrhCTVazp9tx55YgmOM0OQ1Z/dJQ
8DgSZLqhArXmItX2gnJqT7EteSPeYxzOUReLg3Gvvwr3c2hsOSaaXbiDPeuXpGCJVgepwm9s6QIQ
ZXly9IprSgAP+27IzFR/CMN672Tsy1MlWnoS068Ur3kmvYMQgCfjKN+/8Z15uAaFly72+iJUaub+
2+b2ntm+oxem4W0wuciEPHIKWNX1iFVHcTv08Sdn6K2mAV8P3/uVSLesiK898UbV2EIY9z6I86xG
VqwWJmqE4NCzRO1/NFxDYgWcc38W94PDVg6AgYCrIdAeCPt79UsLv68jZrJTfZ569n12l2gDefTJ
QO8/u7lCt8Jj4Ia8QciIC8eyNgljEUmgsGk4GaJVJ8sUkKZbfeshm6/m+e87zQqbWjecTl94rI43
Uil1rSHdJUFOCVGXN6Ip0rdMB4sAiSHf7WxaUFESLN8ftklVsCWXdRolXZ/LTiCvQwjjzcZ3jdHd
LcGssCvCIySyTntgkaw+DMlZfafoHWgaDDQwG3+Z7109G4/JoTI3Gv424xKJ6IO0GnL7568il26g
OVfsfBMQnPKySJfDO9U72qzHxaFZveg3a0qJZQjpYGCMrhENl9ogGOuFZEGUwMQk9hz5O9Z60GKi
WOskm995mnbPubKlv8BrN6xiRg6rTs+eljhCcolpyqTeqLxQ8mP1SsjFU7e+EOcQdgbf4ZPTOxgA
g/QWT/EPF9Af0yLnLXiwsnKYq6du+2B0AooyoPFj3l+enDcBAVr4WCOJTTqTu+yhKxv9QqsF2ENn
9GfJ1du9MC0qQeHvD2rfKEQ4rqRYmVCtgxnHxdg2QxrqUPTCSFwpWJNq4h411gnMK6VBNYOUcdFt
Pyegg9xzaF+1K0coXtDObOh01I/Jg1DgeZ780u2BwQacQQ/xEUj5zcQsgwxIrUb9fx5XGxzmaj9s
N6T/Q2YA1v25A5N4jbR3LkLuTgR5P7cU4cB9s4YwPLyuSQ3CJaaAXaqesZo10u3MWbl7RTCCO2/s
F0/xSwL9cUxPWxkp9VTXdfrrV9WaVHX9SBrXjICHzhgRCCxeAeYAJki7fsa+9TBDN12beaKUI+XX
GttForFuhecDJwahltq8d057sCS5QVtFIMgdk1qLycgoRW2IbTDlNaSmySYvlCmFr//mifvessZs
uI/POjXCI8fW4nc4SfuUeoIhe6zL3+DLFp7CfQC8zV63X2kt6agORy1jz0HH5lInEXJgqtuLnTlk
W/5+zDla63ZRhFziAoWFZrVfPi6vsmwmJOXyhCFRJnyEka4YzGc7Y8CjmBJP2Xibm+NQ5IOLyvMe
JVn43X+DwCE1NfWNpfLcmO7/ocG4x3CWOAUyb7xs4LWhiXnwWmooxGhrWeya449x82ihXlPDLmKG
rm+Hz8M7Jyk9kSzpAoyvFNvhsh0JBVDi2wAalkHwe7bNyYe20CbO8gynr82DxsDbXuOsXIOrwKb7
0OC2kIN75LlHnkwp4keQy1teduP//JCjXXVzDcUvPHVec6Ar3iNPqCcxKxVMqh67gtIqYI4WyURh
quUxVOF4J2xcJ70ker78ual2EUTqDsCBM3E3sgYNiFe6YePg33zkqThnweYd60ddyWU6fZxRmwZZ
BBk/vDQQTMiJazOhbFjeh4sIEvfuDfwJIGaa//0NYbwnd6DhurlSF/JRv2Vvp8qG8g1hi+1BwDVE
zJtt621NoNR5ZWMQq+x3cS6euZl193Uizo1veAoYg3AhY+MJfVirneis2l0XPEqFRKXL2j/My9aC
UTvrZVykl+PGrEi8/t7c1831+kv1L9dNUtCR85migT9/hT/y+f+2TMW2RFf2ZTSHnM7t0DzL3vg5
71K8QjIEp2jCgTV4TiEsOeXTX0x9hqvkM0n7Tefg/mI2/ikqrELZSlsCkVVtRu4PERg3GCgsuv26
CjI0kBXg7/IN9JatsTiybRWknpx0dGZIs3eiyDmDp5Mev1NVlqLN8JxcPsSagA4N+GD5TGe29bX9
1dDvsghZIID1n3GKDI7B+aRMvlSei1xiqfPejpKq40r5R+Xj1bdhUcZXGRU6pLl3ZkRtH6yjSQah
+o3MM65kcHynYs010/rW0U5pxRoqcFAOBj0xrLQj4RmxbXOAoMyn9kl6dIYTU3pW3t3Amm6PKdtz
z4BT17ckoVDuW8RArUn7Gd//dxMVbNFUVrWZ0jSL7+3GhNayPb1dvZD1eHvtdkrsi9k1G2Y7yp89
y1iPYy/BkTotxx3p3aEgLmYtVcuFdN7ZuYNqyhbdYeGJk5qyB4AAdC7pTDl26hgrbRSzQfaruznr
fcfOSOFkSIjm3UqCCcrzFwFtaYnpgqPMvVOyME0Kmxczf0V6yXW10SDN2z69PE2lvpAlAJV11oMd
MNNTb4bqUH7b6DNv/K2rfy6TtTVahFINhFRG/BwoIoJk1Kxn1ovqCKNyfTPpzgn+dtnbbCwp+U/U
13WOvIjJdnz9qXtYrOlBhzG2TLpSW8Q03iTvvqfQ84oRg3ZS6i38zD0sUXbgrM4gnkKYwz5TyIf0
OfwJgR9vqi92BV92YVGs6w/7RCeHzXNFpVsc/cHVlkTufV+RxpuOgiZvwOV5mlrzQ2UpBn7owsSg
w6jNg2CB8pAInwvPaBRc07jZrYEu68ZS4INFSEcZUTBAxNlitJQ/kvpBJPMHjVASbCjhCMnZqa9s
nfQ3JDdY5KZtltqDuROmzRgcDMIbTVGJvp5YW+VTaxHSQVjzqaoY/JKNEG+SLvp9WGIKsLaJ6brb
7nDKsm/b3wDE423jEgev2RwZcOi/3+9BO4P8GllUmnAcpi/f2grKKbZQnzfhglbvUzBVsFvDNyoH
Jj55Ce1EVpqiv2U/da/D0qeAnU+/8pq3TGzhL2uw1Q6GadsIifMo1h0j+UVJuX/Zhy2NUAcCzq9D
ttjM+3LDGnY8C/ieYZc32QBA/cwvlsXcH3Lk5eirYD2y0q7LxcRJePTNTPA+LPTdgGDtWTOL+0Qc
pnzMZ31a5K5DQbOhkx+uSxCdiamH5/6HYn14zuaYQPnsNvxEJLFvA0l9eJ3Y5nkIKdTnUx+wlEJo
AocnodJiPYxFU2To086NvVi/vN39JtPf6QoGaL/ekQDEQwXawkUzAvxtzKKFV9zFVjl4IOEBtTqv
MU2J+gZlw9zJ/Ciw4DYMkoPxcjYAVPO1o6qGi+NAidlse8HJ7k4LGXDb80xIulWA7UQDsj4Uo9WP
Byh1OVTBIoBIcVNOLqh4ic3swAQ+LJXNHsMuJMkx44SYpYejYkxW0q8D2/DFobsBYiqgfxNDJLdJ
ygadg4urUF7sdEdwPpmTjfBRkkO0jZBt3xB8NaAanfbBuEzE9Av5oAQumt0E2CZJw8QVM79kXAsU
QfruUp+41SzymaiBCoq4W//zTImn6ZpRv2a67S9CC2TV2Th8Rtgw3MeN8xsEP0glZaJpy3bN1WbW
kpitPqdYwtbetBk/GwkocQCs3K1V+PwGXPNco+PXSRSXByixFVQDUI7asBfQcTBd7rO4ZqMXuN39
BOgUZtMEEu0bkxaSJTd4xfYdauZpn2SZ1PSFV0ighih5xbov6ExbHeOqvz5mVDkTd0eOzAWUfTTg
UMeHDtDzmYkUqJIKuw5Pke7OQ0xG6LTcrUYG8FR9ctjKmqUrrjOZK8p/sNtCqjQg3IAjHWtqOxLv
FDafuu4g4fwgGeHp6YsMxuANnlx3dRgNaCMzmpzDNaLhKBaEym8FIHi1MSHaRTQEYZq47dmUvz9s
po6ySRfBREcdh0PC4t+5Pw3CBSgpvMepZivY3XCye+tURCkxCDazUG8cJm/5GSwF53cgs5ecjeR1
tGGgLWNkAWJvem4Yu5mgsqgXOsSzK/3hPnvVgW5KM+de0k0jvfiwLeMB4/FiZFg1g18FwLXtK1Jy
GNiX/sSS1/KZSo3jwnTwU4tkHd8WXZdLx2JBe0eHupOB8T9fiTJGUhxFRAjKgKW/ol7RGS8Cvjc7
plpAncerS234vrEe8FoIKFefTp8AycTKkyfL1QJq2gHR1V5vEFCb5c28Tdwk8kGKBHX6C5DRSzNF
bS7283gAchNGFlKRaA0SU0yoDfB+l3Uo3oECoCEIhCnY1g8NM1h5iuYW/G/O7Cbkizr8XHX6NA2W
uPZjliHj5ud/DgR+6Ul4LSDiy2kfeUsfhpKxms4+d8T8v2lXgkhZxlVvp2SBXh+NiePAt54MiwB8
fkNnQthsYbnpJo/Nu/81Hz97bD3GDkoyUoEz9Q7Sm2o84cSJA3YG/oSvnb3uJD+8uznTJxcr5pta
RMqGsdt4QU6gzewf4Amwhjwuxt37vLy7/sZRkLqLKAhhk5T/uM+Aa9CU1vKwY9ZLH8M2iJAm/oev
nNlTHEi1diT2Yfmr3hjmDjQ66+HzXxZEsU56AW18R+xv2a4yun0QWZ3xW0rIM1SVGrQWwpuuGTSx
EWgkTrP2Ma7KTStmRfoh8nawLBOv28gCCK6PHXw07OwVHWtpsG59CXbCSTFpF/eiru6i4IWKH1Mj
FjIu36xXnD1ixm7wvm1m1l/8i2AIoh0GjcvovTLSjVEEVLvYHfRl8xVHegTbtjOMeIX2QSO+1fRH
JbVBpv1JjgLvIDWsE0JhGJBK+aCV/2ZoHB0gmSCDxVo5jrM6pimpJo2h6RcfBfs01769eJeT9+US
X1wXdJuo4IT6mw7Ii2oCf8YFRwVzx3UVZdUMP16m+OWe7m07x63z4nA+0xCeHTEddRm1DkBO8tuR
7D2haQva49eZpWayEAZIBzJLQHzZIeKM7G+sbslsiTZihDQdVQ2TQEIqkgqTWrR5BguW/ANmNmlp
eBeoIzsXERru3Gq282aheOPXmaKOmxQvPzWYFL7dPUetOf3tUQ8OAQ3U+j7Eg0ZkDOI9bRywY6gw
zEbr0grM2xcFVgfjX+vo0pqbjbcKSJltg4NM36Lf/WLosuzqlUmuOgfYkP3RabYXJ4fPxAHLYOiI
Ts/GjGbiSWuQs279M844yTMohOzrvzyVbLeyiVMCL5kRFrzILzEyRBL+cpBOBP1FxFCU1f7rRraq
NqmKB0hxPuEn8ecN54BoU4Z50EWg32dbHUZEZB0qUJGyfjIqv/+6cwepBT1xg1lrmijD4FffhcPa
uD4EZJA2pE1dZ5ENdXp4H6IdwRhLUWRzb0DE7XXjh+yykLeyYFrTfOSpR+upSnQKfvBtWc8eZTaC
rOhQCgdqPOn3hXQHVx20zeypJ6b14bRcAt4pT54shQibcAIK9z74CprmkYTzMUfQRNDFaMsegQFD
EvfvGOdQE40PFbGM4JL/ZvY9vgHvSPiSUDTHb2XQ9Xb3srEFu+O3I5PHUZxtYSJT+ebd95InQqbd
BYrfdwnTWXdD418LFYAw4P8r9Umy0MMZNse7g9lhPy8gRPDJcYCz737rA+xB9N3kfGY4YRcnzzwn
Se4cSGGprVMBPZuycvUBawEdsRZO9Ceqh8aellAAHE8DvSClqnPD4Rim+wwDq7J0yu9lklJMNuNO
poheM678wvAW0FBemZiapBk8rzGDT5TseMgbb0VIaIwvbQLIYNlDs9lyx3YxIzfopd6FBJ3SaK/P
xHTSNqQJA+pcIi9Z6GBVKAEm0svdsU74B6+QnzjtyQNpMCB3yGzDLu6j0Zj8TcH+SkI4hCVCKcV8
MG9D0dIKHpdgbwwcpEMVMJxAyNaz26ltUf9jmQ/ORDSFz4M4itsAy0Lhsue34vG6ITPIzmUen7UB
aKVdSVz2MjQ6G4gytOr3vvhcAQNj1IMroPvT0I7APfhqWcRJeNwkzLRX+UWKWXWO1O47ZUbPktIc
1eS8KUMEv1OCsssAeG2et60qSb4GnPMGmgIU55x+DRPMkVCd9sK5+zy77PyQAb9NcQjp96WOolo4
9IHcS6ix/9Acx5cYG9YwVje/Ovc6KxsJGUlbOODg2VIFE45BcjOVDIgQL/BBQbXzrN+AYu4YFrZt
gYkwRo8EYIGoZG8bDCPrJmIs4RUAvbtAJmLFNbq+/XajW8lC3sMUSEQ/PhKvoOPt5KhS7b/f4euQ
Pj1Rp2JlSzLxw4zFA3JjeNarb+RBKfpFCSLcvwnOr/wrlDjG/pV3lwHWMWB23ETVYDqOsvnwtsMI
/eniKO8s0/VYlcrwsYw0gS2xRI4KzyFs/J9ss4scMR17OtQgGwIYR+w3wGCg5vN4Vc8euUTiVl2Q
Fmp6BwvSDiF7mgxY7EuplpApMLXr7k9ilTYejm6MMNlI8rQsZ3Rzt+w6pAEDrdlP9C8J+xij2hbL
TutPg/DyjVJQbh6OseEMynbIzoMX0PNbfn2G+zzjqFKGk+2rpf1nKTJPfOqXFlERDDK8l/poi1JP
HraRciYnlFzMdDkHYah7YW704VUtK5L3A6+liTszgEPElKePGSKhavGY1CP9NUTLkt1/I0TIUEKl
Frh36JsjPZZCRpTZUswxc2QgmR1VuoK8V/vdRid6kY1M+40WXWKKZK/QyQXjgqCM34X1kZgQwrEF
bb9feQTN0E+ycSuixVDhoNdfNVXoNtabyLoEkPC+JxpE+QiJxDcDxQSLeTRItpoq7c49XxGb+y3D
04r87zBdacfWKemxqL2mctftFU0aJDFOU76t2FjvlfI+NoQ1rHpGUU8MwaEM9qEOb8c/DLe2lHXh
XEnjSMEIcCPoCgzBc/l26VzGS71xJHrGyCYn2cJ5vtGpnypBoCUHZADZTHaqE/d9FUMBSz3e6jOl
f7wx0qlme2kY3gr9gR1m+Ad7iJMFj0KqyAq9v29KJj2Mm5Bqe4iN+k61gnjvHt9cX4IaS7SJzfJC
JCQJbHkuJYvcruJ5mJSJA04yw7ex2NKL4FtQ/yacK2fAjc8saMV+3Fmb+Xl7iJ0IozLf/fdQOqeh
JmsKZdtjuyz6RioTkXlqtPtPzxlQC1ykdmI3BdhTmawjgDwuDDPU1dFaC9kVvxyrz81qhgeR2ah5
LpAIps3FllYgvPrc/Mpy6MXAj1KKTaueCylOOGcVYdrsaMcjvVXVogWeG/TeuLLAvtW5Uotq8pP4
6YE44gLISwjzVma3rxWh7riMgnBXGGn256DYjr/ZYtKRn0nSl82onXh33VotmpZfisRwwekiqtuc
bWrWOy+olboD3F6J9sWUIJhAzy/85xcS0IxmKyX9xPwcjWmuY/QuckofLEfp7B+WcNIlj8LX7lI7
rAiPVZZUlv0B5AkNOeWf4WgCnibLOqpqQgdwZqHplFx9VK0iHWLtQovB7XqlVR/5tYLesNcBWdNz
EzZfWSWm9jxVqhF1Q4bP3eu7WR6dexHptydqPIf0sF2XJEMezWZ8Vpsk2IKYjsBQvMEVa12zLC2N
q1T3C0dNBWqz3rzrn1LyJ8CuypW8mEEe12VRWxzizfr3I6XmSB7a1LdloFFen7o3pMne
`protect end_protected
