`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SYrTT8vRVlz4UcbcwKgJ/U2zcY0Gw+2M2xSPd1pCai5wVCAHUg1U7EY/KACUq4fVXVxbAR+6kD91
+7bt9SIT/w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SrkE43E0DHSeNJItWd7ftK0x9usmjrS5g/8t5TOe5u9NX+OZBrNZKow6mNsFzQJyBhPtb5HpJwCJ
gdALQI4luG7aLmleMTOilyx6bkrkmMvLcQB1pvf/hf/Pb8VJRBoc2sO2Y77lbCDxRHIAci+oou6q
qPNzbkg0P9G4nlYiDV0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hVbmY8XUxCZkcX+QFvZWdwniOnOI887VPdjJOihjNGombqL4NOu2IQDAFjsRZRVsJ7GJAwUYdtIl
vHuSnCeSwExj+7HFTf5qUMR924i+ZamuuTEu0/7bt01+Fale4VAEvHFh2dE/ZCb5jiS+FSIeI0AZ
NW+0U/NA63QMYepLe1j+TpK/hDn1IHfFsvTP/KUq23ntTs/2Bw/CECwhlnmnL8VS5RmPx1YTT7sz
PiNT36ft+DgOmrLp7LoXDRDWt4sKbbQTO3vWxGVMDxvz9+jea6S4w+g1o+zthF37N+X93TVe+JRH
HVyN856chxJZxOFJbmsuW05ivQxfoPS8lvl4Kg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fZ6/SYhW8TG8yxkmGHpw9sbSg7zzri3DOGB9q0SdOXhya3Mioz6gmHnbrV2ebXufk63R39HqzCBf
wKTDvfKqegBEdFT4ZJ1+bgC1VYJDxHjyNeTx7rQYko2recj18a6bZaVbH7lL5ua1Yd+2Is+zHcTK
ZiCtnFlDaWZRrKmfjlo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F0obLtODuPglv4OWUeueqwSWpOtsiwy5TNdPfzLpejVjWZjuW3LuakjFNh0Rff3e3Ve23Qea2tJ4
BitB9zJkp75pwzMxjG3OgSPouZbZ2Hft4GW2OlsldBUfOBdSfFaS3OUi8SRAkaCUttngZMD7Za3v
7cWS5g3qnIMfMu/RfSKF7IQLhO5IadoRInOhBxEOgT6UlQOILJvHj0X9p05gWcIzZkXhc71N2/qZ
TENjfk7pS3FlvlxspcNx7+iqPHEgvTaSTORvjbvp/ARyHr9cUDR1X+TZHnADA6b6QarADp1yeEsw
2S/qjtcGcabE6Z5Jrv/Bapia/oKVPbETNu1Uxw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16944)
`protect data_block
pcN12pC4aGPN73n+MnBWYO6P+NEHtuBzDkl8If00SYsVP9RMvFu4sUVmMmoXlVbtPHH+p5mDLmEz
HZt6CkcpYxazPJO5aCtXJUXAA/nl3RcfJwwgGkl+JVChzKWjOEOW83EWSJs29rp5wjZHpSrb8SAs
hjfWUWvnIBybSY7SpLeQlQKPugwrky9EZw034lAZEXkwEtOqQ1IcrqcFr0hH8pv7hHcC7c2wWQjr
2ocNrIaj8QkotxfMhE46umweN/MipYB5paFKwHlxJk20VBImpG+IYaYY+eCwv5BJxjaLZfYWTK9w
84rZ4l7qiw4kliewyIC9ZmtQ7p80yHkXLoPFB8xipY37G9c13FUMqwGB92uTHYNphz/3thkVoyYn
CUdukqBWF+ZNjHxIhUn3/0gmVw3OvqORmgYGXx1uuS29WGEsK+pR/UUwHDIEZJmx0d+xFph9fVmF
rK/QC60Y0JTW4Oo3WGVJN/2cEkJl3LNPZyG0FPbQs/JqzOPU9ipGXSCxyArC6owvWjB8LOSHVUQ1
tXdk6ilfH4tU47XMTJ3wnScs1wRamrcBmqytjiiSEnXG9Exke3fTihhBW2FfKmupoiO7gw7Ip3VK
mn1F+8Z+sljxoYGX4Jw3X3DdPclry6gkWxX8ICT0x/Fpzgep4Eipnwr37KsrLn7xLk+WfVlg1u7N
MznOy3mKts3crdIw+SfKFbJ+6nclV2GfN5z2oBxUrcmAt4mtkINXUyOPtkGEd/ex0Xr6oAEk1k+r
wzeoxi9v36exla9q8eIbI4TrO90Iwqp/mSYWM9aNIgGxSvJNbyqpxu2eb2tDm6OGHhmJ8JODsVdc
DRxadOpoRELwmhjWl/2BkBbtdClgZK+ybPpQFBmTLPjYZPTe3EAzBPU4bNakaqM58cKNkQcqjCEc
SGn1yGOQa0AMHpv94cKyTuPs0mHBBVhzfkIlrEJXgA2yDQqG1oTD/gVyHzr1lTY3iWNykE6IDAsQ
fsXQXs5cKTqf6HHfZ/s5gfbGLpNOVmCOkSwPm9KzCVxQp7zl7p31sWWB960QM2o8tRondbr4XRBp
q6l2d3pfv3UmJ7Ck8yBLa959gsoB8kGjwSdz8jwQr+vIzek8T9HHgU56CT8PXvmzff++fBVlgopE
GRIFk27WU15LQHy9bUlWGH/PNqiQgFsMUGKOCPTI4bUk0v5ApjVr/G+02zuJLbdJ3ogi/rtmoTBz
IbfKz/3q9/qalvBS2GOqyK1zErUP+WldugOhPM/VhZK1XAKwftJg4HA/n8fG4w7QkuUqC2PUeQeI
AfrOSRL6h98yU4wQXyGQMN/j2ITKkn4HQLh33JS/hTp44C1alq5SGl8OgD4VdJA3YmKQBuzc/Pim
AA2SM6ejIfvT8e0TcZA8cobMb7ChKWcpbeZCdyVkE377KLdWa76EQ9vpHBEvwEaivPYWi4BsMTsF
UkWqXLPlRs39QQTQWGP7QJ7dNyjfcPgxaUSW5bj6GI2vYDNwM34dDcmfX76c/OgMn5l7shaIVrk7
w3d9jezTy5uQgoTgUSTw7Vpkn8YYrP41FEyZdlRsisA3dmcL5vbZaWEjjIFflk7QD+7NrwgRqZJZ
GCfio6IVUwyaGV5UG4YnhLeBKr/0Xf/KeVZeajQJAlvKqdVMWe/ce1EyrWti+aCXcmQgF3ZIXHcS
C9NbjTXvdUtNrv5k2dDaEdlx1Myz/CTmi+a9cp5eeI2Z31a/ukRKjDkvcbcclSBnPOc9/xMYq3H8
zUeJ0xJ+MqOIZdlipEyCiqc9mMEM/aYZR7XO5xxRWguTnCvGTkGVziIFmIcVZbWJHQaRTTuPletH
D4dqatUvO3G/xZBuHHHznxb5i+meEd/8SGLoEt00xM9VuddELfPiGR9vB2+kyor3syIwvlkNxv9z
9r0ks2bwTG09eVBZGYvKnqEbz29x6XUHh2RRGdk3DpU6DI9ihjnPvq9zsujYbMS7j7aqoKW9GUy+
ui0yKJx5rdBjjcJ1uUF4Q9hI9s0Z4Yx23WfWkw3t/Y6HGQUtvbNj2y3Xw9V6kvi/nVhHMNTBeSF1
igKWMeTj5wykWhy/z8zgCOqCOgs16Bti11TjuznJD7rm1O9ho+uc5AYmlFaXyTYhjLigieIaOTQC
jQbd4DDzRuH4WghZFIQR6Cw2xDAoyBGqSzjkkWS6OTc9CHeoNSG+weFcR1VDULGDpGDvY3lR791/
DwMdoa1XET7zdscoI33w+7KgJ5cTY/fQvJmeHIvHlWiVPnQjKTS0+I9j9ctSROKNPm7mSBQpkuHw
3j5aQAYiYhn3YY5w938gwvkNq04jjMgguSEBfTj/AEpMVrj9+892MdGZ8dOMnBIHxOBsiivQnRva
0OMzn9HPqHZbff/nC3C5yRW5zzUz9Ac8CYeD2nQdXGLMV+mfa+K+ZbRhjM58lchMIrdjsyfhv9UD
aji3LImuV+0S9x0j+ZL7ubVvT/LfLVYkc//X3oLnNiooxwDvWNREYEy7NAVceNqbQp1iWSiazWcT
iMIckKxWxvO1Kv4XQLTHH2bf0cSHEz1oWSF27d+P36NfE4bBJiqghsQtYXxoNBEdhP2Xo7kIJKml
8JwAuj3lfX/pt+B0Dv0QLAM1FgKh9ycWvIJiGBQRRtlDA1XbiN4gDFdIwONGyZgvOxIjDsdNy5nB
6ptfBcAcCmQ0XPfQlggz45euZ75mP8v4xYtVz18e1M/FK2jkfaXCseXojN9VuYxm6TDaacEsY2Nf
3EdQTEvm20gB7Bp7ZIepRsbUVju1IUXScgrYarG2AdeGgap+jqvc8mUpwWjgklIkDKbxi1BLZsCH
EPrSznxsWVLbVP7YC+OIM6bTll6TIjhXGUd7O/NfhFRxq3i16OyPTAktRa5Y02V7n5FY8ZHzQZYR
ELFityriaLOzF5tVMK9Q9bHwGMnmLf7TRvDNnko/zyah/ZqiLB1Oq+m7mP7mJA5R2nNL88RPyE1t
E2AUfO0nrJAL8EAFWEy1X/rgvKnbk0IPxe6V42tBFjbPxQ7srRjMgX6C92keCjCgnQuh2rPFpGbj
kCUrkOxdouIpdWfP6JZdWloRf3e8nPHC7XDefFOBqW4EeaC4yj7zGkEgoea6xUbx44ofTZKZor80
cSFn7vbe3elGiEk5JfakbD/xKU7/0Sl+J0hgYgL8S2TLxrXgq8vn89fB936fXTaNUuBMe6BhTRH2
j6Es2kPCXqKsgTU3pKyxWm06jkk4RgENyE4M9Px9j7t+A4EYOGm1NOysgLFAWX1IlWRbtjUd8BZO
BjL33c3uSp4mIWAq5tFZcmm59c2s2kn8RWXeJysX8e3S6vycSzG5DS31+VqfLDM3qOEaDkOqfh7g
x55KDYgGNMgY/9coRTm+IIUxQ9bYCsv5f6oSkQMDX48XBrSR68gYbMN+7Fk1cwr/2IDQrnDD9Keb
r7SiU6P3wdG0qjHrmmLRDLaTB/SLMDv6GXV+rJASltK8BpJpQdSM05mdXmy9DGpWxSWryhCkTL9q
zNj4g1xRAiVEH0B4Rf4R6zA4eLcXZXrHDpKB9OhzlFZUCbbnklQVl/8FEttizueW36nUA1d9bZJq
krhpT8boBEnTIreyvqbl8Mfpb/ZH9KA+sNXwOn/fN/pNsdcWepUrvu2ParAjuHY/TWCGvzM3ypOg
/Yt+hXXTbi2zz2BwfsywdA5vXesvKilFQSxRQbIo8C4FxGTAO7YKMTCHiyqIYMnhSWrYW4ZRZkSi
aL05fvJcfLg8kptUDm3dNP7dgr7yxeNhap0Q1Zf0doUu9CGIvUhzUP2qfLPzOsxwh5NDTg7FDL40
FstJPpUhehLBuWlg67F2WMdPmqe+g78eAzyvS6gRJNRl1LEA6tO7IMKc/D4R9/R/CmjGCNlsUVlC
oCSny5w659TBiadEf3e9Kplu4ALbT4QCePmSKMF/saxGXDr+D/8HaF8vohir33O+f1as8Z7v+mTt
EXg79e9XsppLkGE5cWoL6uwxXbAbjjkh5pNUp2tWWI7lJGr8zI7CTfK5OVxlIaBrWuEWEvo1Mlib
TSIVZkLHm66VCNdAwAwb7xLhBNY1Yac0f/L1yyDBCOjCl696ISoUFGqKdR4JiI9bLgLG6X6zDJyH
8qxsfNGUtXstplM1thQqZVoJ8SKDgoYIrjsrHy1TMpTd9RDCBgFRZJqEEgt8tlWPZVcebHEZ6kpC
nLWUHyAHA+ppZsB3R/KZxSxSRQADOodtXjnJ5KXQhOvzGqYvh12j1GAaudHA2uTq0plOUheETjlq
oQh9iebVguxxlDAQJpOuDh0SJwbnZEh/LAgZZvj8MqL4lz/4ZExV+1NN74wl0Faw7MELZ3//mXBZ
4j42YAh2UOMUAVz/8BKnitbAxCiC24uLSVaj4MX8nZlpVvyausF5VZENND4zbBRjakw9fc96SSg8
572FFbjwRDIE56rVZfZWaRLxh3UfhpZxf4h30zrH8zolLQpJyxxoj16ig+u3nmnGZ4R3oPvEH34+
LOjfHvWuahK/lPp96Irz49lDpUoxqophIU8EL/gsRwD12DiKgSHyvKopkmp2LHKLVqpHiGkqq/dv
NssJhxp5NCODRNHNO2yzHXn1rjUhbc4Dlwj9g9uSAIEoMNJFZsc1KgEqB0s4oOS/ZHbNysOi1eOk
kUeAFFclBpACWIfHX6k33+63eIMFLyt8eWZpwL3t5/VDJB/Wc+/DEsJN/Lz1PfMbcoLOQc6PumQ2
6m/gQ7uYvh7/7GHqOIazQvrW/4mgN1nykSfu2TaTCJwNknN5F6MV7i/BjkMSGX6S+MXUv/xp4Avr
ToT5IcRWX9kRU+fJzEMXzOs/jofFpzNKn5O5p94xIZppTEt1e+uRN8v6BS1r1tKEfZbKrD+xyejB
jKG4VXX1lTZo27ezaDbOJDDbLj6wVs/85u45IvF3Cg35qHSEmg5EwZUSRezPEYr2sOpF0jVmBZC2
B8Ft5C0kN2LOEYyrjB2LS4xBFSSSqdApWrQd2Ic/agonqf6uYvFm1VkHtV4LvlGNuiFZW3yx8hyz
dj6NE4bG++ni6FAP8iBwJ/xL1GrEpq9Pz3aS7LM/D2HlolTTPpwb1AkwZSTB7rANruKRPfw1UREk
2lCY4Fb+RVBe+XCHJATQPJ2tW2d64xKqlqTkWjCDxoNFJEBRIK93cFbDJd+HauALYzDdAbO1KKD+
bMmtUljOUwnYWgRBhgU4ESfZsfyKTJTYHiQB51rcqqnNww8oK7ejMz+SrX44bA+L/GzXNQndoAq4
dJ3Jwfvbrl80JZFN33osnQ0wmyjrGRFco8TfEGtKPoaoA9mXbDk5sgao5F8n0lIZk8qWmla29f9n
hABk57apcnpvHElVCVmrAAMsjTxneJFRFSmCwY4615P0bbu26sQ5NWNHELuf9vq2mj6FjnLNeWwI
bbZtw/3uPURfZttAVL/ZVgHF6yP9Wb4jaGauRVRU7bIk26lrRDQX2pqGvuBbq5rC09NvV86pI9cc
AjjO32ZYYlSJ4KyWXIhhGMLg6vRUFP9Cld+lv8R9/+UsT5U6ElITRVKMVwjsOBD5o7Qz0imgNKyO
Fcq7fBugKInWuvH6aGYx5DyqEaiJ5SPu52vyRmePwtRghgN99mih6RkXJmDM75jG3egbkYSKi39L
Jmd4Wt1EzPGN+1JIg5H0s6ewzq/PsMRLFhcFiWVBKupoe9pD6CenIQ95ZpMCOfVaDUCsegGFuC94
3iiQ8hpnaoB6U08LTiYH+RYhCrUHlhVRKcxW5gWuJRg90XA6p01l2lvmVmFqmgyWo402yoocEnck
mX/kKpOdXKxj/Wd9NysMMTTTIVvEHuQUZAAnSuF2Lv0hoKICorYWPYgo4BEYqVCnP9gWyrPKHtqI
EVpTe0ARobVWjwRAfNL1v2c+ta/3zfFkE0mgGLfMQeG+S1HB+7f5MbH5mGwyPN2y8j+btlo9skXA
9E/96Qmoqdv3HqGCTzXqjd1A3pHg9osvAKTNEtmblx8tudBxNH9tqBb3yak1szU6uvEXofy/4Vm3
Esb9seDBm/u9prscg1hEONwmfP4lOJOjkd9B82P9OtRAgVSlxu+0aZ7nuk/6FCUMTeRAHxnyt+Fh
xrKulS82qq4MbPdAEdpjUyFEhJ2djPqvaZRFo/PnrmQM32l/A21HyeYWJM0op9vKoYB5LOu7zgVx
ULpkbH6Ff83/KSqw8DWYAtLjhFOq01mNVvZ1rzHa1/Ql3DcwfceWWhr31cXwBZli6eHJBQgbyffV
zO8MXRN7KGg6kKYtpWTnAJeoT4SgHgYSXzJmI1b1WiUoWeArQB+70coW1vaUvAhWATyoZnwIjyG3
OaVUrt2UcPk5eP5AMVEUqkqLpfxBV74F3kpAZAOFXawEqwZ/cqk3yIdK69rM4472IUxVgxVU0eVy
6Mw/bToNnqytfbCDF0ZlMIsi+CBjLLB09K/KJq38/s+Rc/Wyz8OGMCD9+03fwi+4Z47hA2SCxOIa
/HrntLyKpwYCXQ5tAZiGn5KqpJIe97LwlgFlk3Z5hF+BqKq5vCjUN7mU6b1I/+iMhLtDL4mvn07i
FZsPKGKIvhUdQER/kRyCGP1KmvzRM0XeLaFpL+kPdS2UdSCaVJOuwMh+FOh0niJkbJgiyKtDSIH7
hwDefALfIQgHzErKAiH9ahK2jh3GWLOR/PZrI+VofEi2XieVGsNzYnQmSfDBRfXPhWQR4dMy3Gf6
0daa0NVazwsElj1Ljf7vwchY3ha/6d5jLEIvx/yKfMlW6+Qlapjko4pW6PU69kwsLM1umv9TC+py
Am1FSbH1hetZ6mVlT7PG2s3Uyc8fh7ak5QtTdbwFM7nCdthvyfKl+/clbtdVOD6ekKKW6iS2MC+8
+YvB/WjfSJQozGoJ3B6nTHpS9HyKbZqGwxUdr4HMye3eeyx2PrVkWWFT/BiKExJhB6Skx7arjMuX
lsNEiumv5iq9wqp7Im6HGfpc+9U6kWe5cyf8gA4blWsX6quZ2TpQ1WqNjpe3623KgvOJgz0Kjvr5
RUyeGgNxphs5gTgASn2E4qcWrTnjjDt70ssoWsuS+q5Vm/9LaAsT1qLWZ1Fe9p6xre2sbj+oHLzs
/X4BXkXqjhi4ANrIrd7ZWR3EO4MR8im83y3F5oYZUUqH83AoptLykWppSZ5StruMyWUHukwt1RHd
rdlzr3spGe6ebVRW6iJfCK7/05wDLRJeP0q0NQ7hr5inu9fxTWgsWIucMXpW6Bki9npQ5qXFJZWU
Lo1uUqSJB37gxurlPQPQgwibkbuzP+WR5V2lXZ3bm7V9tSnAtCZrFaqkq+CLixb9Kjfhy7K6/j6k
MmJK0BGuKY05ruHXsqdAXCX5pqwl27GS4RT21FGQAl8kpyoXaDZbaxbvS36JdpH4vJ4WSDXVlesA
3255La5ndZI4LCH63SGxjs5j+UIN45bK4iE19ifKjjXxC18bA902CPfJAYkFGjt/txGCgSJq61vw
DsSGDBIxLdDqcX1Pa8Ia2XaVB+C3KFoqsf8l8Q3kjMOCXpHVUg649l4i0Kn8jV14gawzeFmxKPgL
hsu5vn9cO2tP3kUDCHmhEcypCxymmYC9oaI9LZ7Y/i2NjophXgi4FzPWjaL0mq/CWuwQtdKpRlwF
exMRIrKgdvClrLGA0i6MmCyIb4SkOdCG/nZxPSwBiGhD66zy+9TobNeTZW1cWQhLyWXFE6nnGwSV
Wj4xLAehUvlH+AzqhHyzEiVTS5mPq/m5DkMCPqHoEYsCpbc+ksY5dfFCgxtKKFyg8X2eLGR04Z8v
REHn6pq2CJ7Z7iD6cFih7ranE0p9KqDo4U2zXYbMoLw4036/qtApTDzQmBJ73WnvQvRNGVHOgF3Q
cQ/OxCorK/AjvB4VW2F5Qr5PFh2luAaP5/qfJFsZBSh1lrmswHZRNEqFU8b14YDsQe49ny7ql3dk
Ho5+OzXT6Dpo4SLrctNLvdu7ICALQjNRu5tiJ+4BX7pcdfIXI8l0ADp/Kr6HQFIWV7kU7nEL/hiM
RjUzyz9zcw2MCZZ2KM7Hg/YC+e8vzz3tEmmfDm1QQsGkuaT1Oxd00shVAvdj8o+DUO7N5rr2986q
K3V5RA1nmxXn/jg6m1EAqSDqWQm4DtkRfeIb9pp4CsJpPXAA+tmtIe8sQNy/p8vRP5NpFlxVU/eY
zLqB2aVp1sE0pk0KbAvcd/2PLDOFBeThi2b642uxD47gd/JnJg9r4RXPAkviiPbQrpuTMa2n3IdR
uNJAQ0tpEetz3hSicRWpTtBY6v7HYYTss88jmtUmPq0NZoBasG9QOmcb7mcYFJp9lW9lrM4dlCSt
2ULt6aZqluYegwruxqJ7sy9crnlF7HvD9iTdJzRki6ADoL/27vssG5nwKOCUcekoFv+K9+mMYyVv
9wk2q3Nj3D3CJhMzQfaGXAg05EGvLGby/nz8AYfgQWObKC7o9lkJ5ksamlmAiJZHMBbLi6y+7FW8
Z89msrAZTvwBe+F7GUTZajl3vSvme95YomVtBVNDWLqo3gnOcuPxnKo95exNmI3g7ZaVbKtFVQXC
9wNWq2fwW3QPD/usEI5udB6L3fw+KVOutpxQiulKxIS1T5CJAAzKKLZNa6jBxBHdJMQNwUVkfBMl
a4nL46BHNjYLl+j84Gga3jTukBr2zOKedY0SVmdr8dyiwy950EmkBTBQks4tlaqFAnjuWQXqSyRX
dVs7tIpOA+cTgYbFjSNEWD+LMlL+jV6cllS7hrioxCPN6OeO9afHuJwFH5ROlENY2zdE18HpQqSY
kdCBjlN5ex+IkXbZZ0KRWIJsNIcTnmMwmQh6CzNKki4BkZHRj5i4O3qWgM4vp/1bsm0qAQanjjqX
i8YNIA1eAbxJ6bsy65w1UtG1l+islgGK2sogQ+EOizZHJsrVs0BLsxYdTNU/xW370WT+k5Blhnmd
orkkCZiA1RZ4q830fqRxOSP5uT+xVY55DU65i75hE/6S8LihMjkEEla5azFbwQelVq+qDx8NESt5
ShkfKG8khNMEU/9beMp/rOBeZnFDr4i5nM/ntiFyEhdiebnFNuolzghnsImOJntlNAuZF9jeCfXZ
4lRQAmSW7tZp8NdHpEqZWjTTgXil2Jk+VDaJ3i9Z61Klsxh2FReu+31tavojTEhvQXktpHEEt91Z
29W2o0XsSSkGh3W+LN9hIoQAtP375A6EsgFIC0OEP1fLYVuyZRwtg8cE4D+F/xwM+5bz8FDDzbVu
3pf5asOzo2KvOBxhKXzq9Tb7S4MWUlU0VvbBzpmy8g+22p4Bu/MMHwza4rCkiTh6a0ipF8ir0xkr
v+VJVY8DSbHoLKtLdG5wcSKDjTZ++CT6ZcNhkHmKIFxFu9QoqbyKVaCqh/UpuZeoL1xXs7D0fXNc
afonh5smCaXuRbohgQo3dxn25AvGkCVyay0+reqFXXKuQQuUtRYoty+o6i+q29w83pH5dL7To8ij
K4tgB0PFS72e4RubuN3VPvQKPyxM5o7I23SRdr5wG6H4L4iqXAJtjUJQvXEiN8/vukS4wCL/+32q
HuAYJfuUcus2Pag6nt290ubYoLqpe9o1JVnG4dnzn7loaw7gjB7qPi0yxKEDk8kkiRJWTSR6nWPB
gfW5xpJQdsjRURkNn5qZ/2WsdvWconP9lgpCmkktMExeTe1xNosSYBgJL+hpiovDcPk7g0VImm6d
si2npoMpeyPmya3ElTXa3zrT+2vTmacGYm51aJ4usha9wUeVsGLR4HLWxEoHcK/z1+qhjcaD0L6R
OCbWMaF9KyE95ygXiZQg2siM+ohLMTkEpOUPLMlmJdAxe2abhUybYO/VdVXMGGyzh6bmPyz6Km/3
3ev7W62ii1br7lHdhYaovSSVJTT9FJpP0+GJt97QwHnX/SFk8xQcuX/ehIypAxe604qx3cFeawVr
WHMZ3rj5dKCTeuZE303Va6TmCH17V16La22xRR+Q5DsfdspJld7ltDn3IH8LF24rscXLKyfRUtNm
Ne7lynwtQ8/GkYMJSzx6FrjNgdxafxx9xDEL4KXslp/a12N9i1UdCO9k6RdZR/gL8dSabTX9jSoX
+DWreGV2uOoqv0+U4V3s7van3Sk2qzSDiIZcdhkEzuXwcELTiILkd8IbEbfqPecast3Cav6VcXfy
j/I4SofqeMsgj3OhdwT3a3dvlX3TkJGOWothod7Fkx12ZLqCn35QK8R0GtGVqf4skolpapiSsxjO
Mo0R62/O7oT5dShZ2/vEbShiLI06iI196m/7lgqZnTM2nZ7wYkVhGrOClUcUIj3DUPFBYJ3Bn1Jx
qDmSUAZcNZdKOzPuK12YVI7/JE01201B0jANFFN/NqT+H6hkqw8pWWz1zObIuL76i/41bb6Fk27s
iUjfJ/9gvWT4QnUKmb5VJIwu2NtY209jaU3Z+WtE7y4C8kS71NGV6C+GhSuq6YYvz5HycK6RiyPt
emMPmFc+iXhsTTMogotsVCwJEtiLbc7SFpc5LlBiRdnh6fp5i11IlWwS+cOwAlrwu+iicPZR3Og/
HTdAdYEPaKk36X7tZVSbUj13M7GMcF1IdTVe3RjmrAukXNj1K8ZeyKW283vQ1kd/3zXWhZu7vLli
itr59wxOqdiesgxB7M6QeVDJJWowCloD4Yj4CxANaC85fkK8ETg4KDWl+zfxMisTw5RkQdLji44D
7iab6O7NrkgCuZ8XFf9mOlBgn1TZT0KLyVqqItKiFkfz9ORvvSk1P+kNc6YeYgSf3TPEHZ6vCbdR
G3Ita4REedzJukeol5ub932gU63PdxA318R1TwZ+jMYCAfrP4kaqJE+sTkSGH3dRYXJorqpDPpVH
L2jSEQiAmigNp2S8qc0NEvJWWxKmn+UYYsmZV8D5REi6LZJgCZPFPTZr7i/p0/ordqHp0nI5ar0h
fezGkusIC3YNWdMS72w7ngLHMQUjfNO6kBbcbYUcp+Oora/xEJ+hmt9VBlaoOkJQfjj33ggHPqxh
+hwsUVbS6PKVmMe9im9ZKAdIdhldQknmZ0uZtM91NyTqsqZ6QPpgACeViu0UFIqBfthTOSMIJEp0
T1KCyKw1rDNaiy5/nnN1bvGXJaOdcGAdDewVEih+ovw59Nk17I5r9z8PBo8yKdepRKdPxsHIkrWy
H54Aq0EXfXDEf+8I5JmO7HtpDaLqgkvT3+uTLznas4jyo92ukukIb0IX4X+SyBo/aHctC1BOM+N6
YAkjTFhHvbwFZNpRtyv5OptJvHFIIjhnsVE6BuvmPnP4ET2EQPfO1GGqbsXPiGHRu34EqZhaxmwz
HR6DMBDdng7otEi3/vUct745mP04xCcnxRy4c1/ws/pHh6ll93btEnV7fA8lGrMiLpvC04WQP+FF
URKlP9mgbqS/Vh4moSYW9Nism5EYcrbEij+8+dVeo3Xni5VJArnkJ+MzSLRkrMgz66AxiEje2jVU
B+Ny2ivP7gXWvknaH/PZVf+02/i6SSJCEZssKQoJ5Uupfv3gNKLouZcKNpa2C2U4XDH5kmigA/lK
C5x7DFHNizNAk0oFCAkcJB70szxPRivsO/itPeOybkqIjHKLe7LnNz9i9rFoyQkUvqw/9GzLDG9t
h7aYClFTVVSIhwNpCVtnAwEaP3HldiMg8h0GgDycOA6Kh3WdvFkXABEMK2F5lRLP3TzXtytnjS4b
+2s2dtJ0rGI3Sqh8+sFZo/P3GKCpCFhWkAKZC/iEWTrl2O7hqmLtcI3+5Sgvng+9X4M7rP6ndoCv
TgarkWoZen/v6r3/5RnXTaNr2GNIQr+zCKqqSyXrPWE0mAabjkZqgFiih1qC6CNVugLRiFILPaNh
TJhZSu9GZhVFVnLT9F3oxL7okJ8P0/KMKjrS+Zcd2OKE014c87TNHZhnPDLIpa+8lPLGZhhZXmLF
svu7h3zWk16frhbqfuApV1YFIca9axhhQfxKv+yRin7V15laCMUrdleuOKa8wFDcWVUBmxC34eVt
S2w1uJwyedDXHxBfv+sVoFzCa6z8AJ5u2iasWI4a7jXd6C35OdHMMYnhSHzJxIDuezVMk9P8fz7O
mwTxKzVEfK/Q6EauLNTIxnpdtqj3fhBshhoA1TnEDdx5JrB/DsmWjCbEfEMndMjGyE/2omNmSifX
ZfHu3sGOf5kuSfi2HmEOmaHBLlhaJuucl6U+To9fFtSfG7i1dngHC7nTMCx4wGylWyZ3WElF2Aa3
TSpcM5mRKCk4JzHxARNuTAv/YfuzRlqbJ/jmu0bC4Pp9A0IOsoTI2ITBjsoDTwQU17B7U4MzTBg1
ndL98XyQth97C6nPEduITPCBMNJlc6kCEYKo8PBJFYutI6vq3RgqQeZ1KMvEJENCohTCWg+e+ZTz
CrpWtN8AY+YvrW1Tsk3dSare5LiuZ/L8cYsmlBzQbis9NGIO9LQ++ZdGJqOiJHjwIjPLNlGT6KLE
XFmHzO4tDBFv6/nA5oiRZ2b40KM2S4iZ+yrsMeUovGnP2SIRINs65ox5uddP0l4yIWf/cu3EbyAB
19LxDByPa3btIc5nfSsfFXzX6BzLjpklNjAHSEoDah75ori9+BC9IWRjioI2emBDarAr84IiuzYw
dhVH62EHmO2n/W7zIi8IIF/4/pJd7iASF97FkeRwSqcMx6IxVxm7uLEUGASfnRyxpATwA57RCPlC
ywdhEPJT7ptaLcaqT08dBOo61llPVboIQTd3N5ztYUw/xDyim+MFQ1FSG+Pq8gNWNvdOG5ompiLN
K06VbLtzb+jAVLcPVRI/bk8JHh0CI0Eg4w8KZ9d8x+LygdSR+xvSovPhd8iGXWC2nnwtGl5lz6d/
I4tgMzVetDi5YlquHSoxv1yoZqEl3AFrWft/NV057kgIT63GLASSe+Go8R8W4vxB3dPpBkB20oS4
jqr4SNroADqu1Us8ITpw0j2TCtIVyFbcm51Rudc5Kdcpm3bclGrKlt/muWYJB6/87j/amx0t9pBj
D1xjX8PZZWA7qacy/Nru6Y/OCKwdNTSrNbODDVmJsWONK1UPpK3Wk+s8T5KNNk/NHiFKp7UipT/r
2ihtdGTSvdsf/VBqVJ8ZFNQq2uzl+Ksz5ij7FOSnpf1sks3HBfdY8kfVUvWlQg87erCBIHX6AtkJ
Y6p49DTQGIRvSNfiw06fgg0zJwv2Zzx0uXMK1V1LWo6l//B7S5n7JxheH5JO49CcOLZQmypCacUg
iE4FKMSZQiuSUz2jBjl7mT6cObZojRieGB9p5P3Yh4AusPr4+c1SSYaIdC/7M+DBW4zBN12CsupF
Z137USvcGnj5T3XMchUd5sLh+OWkJDA4Yo+a/WLl7iR9Pb57iXK0zaMES/0zQaheGNs9tAOyxX6R
WpdqT99k0hv6DvZiuBaeZHFvlZD/MK3ujNcCPqx3n0qBMgjXy1gDwZI27CE3fpEF0NaKiT6n/Ps+
wzVVCrSSS7CCt8ufwXfeLJ0FbkOiGPcC4Vl9DQPcIVQm49qL2asptNskFr9hIy3EjJp+LBGiytA9
oT/pVq9WZ4EV2B1kjTVCk22Ix+lFPrGoZUL9/H9BTpBP0KETdEZLhgBqe55q+6NuH6SITI1k45RR
lakwPUniJLZqinx6yNaJZ4g5xC2blm0kjKPj+Xv8/oJOPcYmGt61R0/qFm3Q2HY4VNTSQNjvD8gp
MZHw9xYYu1ELPD/Ogh2cv0ir1TQ6L/8ZgsqhWPm00t0z8HtWOpaL+h+ra8/Z/HGun9yRDd2RxD6/
KvHmcvslil1AcfCH+UGPegFnYXQ7fuA9jkkOnKbbc4bLeSQaPDkGXvyC5sZDfGkBLmumDOJofQDX
Sl6YsXp8oaA+YYTchPgqbVdGlJk4kOSKQ/d96UkVWAn63E7lOxJzxiVGo2SFA0E8cuQIQdZBogCK
klq3qeVSsCrhL8O2tMkHXlknnTG1tqam/+6amI2wr1pVRXvZkY12BU3OgxgFCqjyrL52zHnz70kO
/u05IMNZaKj/vz7VvwXFJJVvZda8P8BOShhORPR9VrRNSf/ZylNsFqIK5r6Xt0QbtEznUgWK+4SA
HlUsIq6HuN3PdFEgVGLT3sqT/W7/qOm9rLnqCSBS3cqG3J9wiGfb9bRwJ1ilxCpF7X5Z7MJnS96E
cwUE4r2uhX4xOmJAETWn+mMJreyVLb5Qpl78rAHHQua36WCC6UAfyTh8OALR1JROtrFxqzsSwGSy
npci2NIjt+Ov3dVRLboVOtnTzadFAlyjttf6bBj/Cy2aQFdMQtafBEDLRg86iXnOLzZbhE5Tg4IP
f2C3FIAK/1XFg2k7ZKKGy9FvYYdVmNnrgdRb+ZiyZpAy2MOJgrmWCjzGyTjEXTpNDVxyrUfNPYtT
azhDnsHWWGIIaJhcWJNN0u7VVWECwlqakdIV59GK+RTvuzn98t/16EBFSfLshRtYgFMq7TilDid3
zThp6qGLVx3tAPdOe2N08v7iRHJoUlhrPUyRzeHpKyVSYSTgCvZzAjzb6Kg4VaR77wbZ7q7QQUHJ
cljtgupVHAvRT197XKoQwT0gKCHTVOfod7913sWtvDNRA49ucv4fL2gn2285cN4FWuj2//T+AurY
DevNbxJzd3wztT+7/0/b8tGbvbRsTpKz/Bwn5BCqJhDDLOO0lT2aMXF93Y9ExJ1UQBZcZ0WpxArQ
JiMs6Y65Nmf8n6QeZxpWgLJNLjZpS7+O19QqLQbR6w3fhceCEYePmWOq2GVmfO8zIBGoXaWSOjbS
NTjS/0Wua0WC8Zt/wN1tRBXHc+hlKX8D4sWBIWKo4f6kRGUhigOZkw3saHRYctfaAgIjBra531Z6
ER8irYnm1znMG4oSo5Xc1xPNwTGUko2mfUf1H9A32oSRtOuQpYWSsg/AGgSk56inK76OUSejRhEZ
QUUFvd2bv0nKuMStsNsqsFrtAFgotzVnl4jDCWokxvvPabru0bsPobBYKUSYu8cU0ibE1tsv22yt
bQbWXZDhKA2CXUyY/HXfDbmazEhVA7FafoP1kBwlMl2N2xwUf7l8tMiehEwfqbHv4IQoTNv+VBBW
tUMBDdIhCW1vAA4WYuKL733pPrwuo2Oxa+7MM76bJrrqVAmWbTL5Udr9tNBHhC82n/B487nx3PUV
+C3ciTKtT+K4mwgS2FERvHkmdKiDU0+msE6ngnnfO0nAEK1IBPOh377gn8m2l35IF3uahi/e1ygx
EYkGyOJzm9N8nXERNFLXN+gW3z2D82a9gJZifqrcXnz/cEaneuOxDoPRF5EmtlluAIHRN6AqLEGd
wYhQRLoir2h37fuXlV60cHtbQZ/6RD+1RvAs+6Z79axsZiOgfhUx8n6cXnFLfU27qEG2ZHv1aqOO
DeDgTNmCHaQIar3fRhBkXUA3WWhGYM4l9Yy5yFQAwo5g547D5uBJwZGeF9P6n2etI3Lpy5efCZaI
lun9CmMgIqpV/OW8iAhAkJVNEdTZtJNDO8pW5Q8PwApytZpbc0gkh1lxFZNhyuEGCTUjidGI9TRP
8pAzSBYBrYHcapyIphdyZQv568HinSXYvEvYSVp1FNTpDs48XBxcFqQhqmH4qzw6Cdro+UWZncqa
QPI0wAPWdfElllyQcqyIkQK22CJziHyfoNz+fBsdEmjOytRPVONh4NiV/HGLSoH6LpyeZRplKcJ0
hdEdQAwdiH/TseA0Lmn/d6ZXo70KZlSjROnvojVt3AkZa0twC1qGVvbC+e1VkTfdKtxsQ0SiaysK
wYw1bKjbIlZTufMPdgx0PXIZi0i0J8lPduI2ofjBQsSHWCpq5zYed75AEBmmTMVGV5o/HqC4y2cu
+znjXZE7HA6xhItiF/ofmH58fgYB3VcerIghz3mFa5JwR+jurgdYTOJLUjhlFVQirToQp3B5FcTI
xvIvUVfKV6qKFgoIojfB1H4k2JGDnRDX2xMhbdybVhzW7B9LjKLFBAAdtewsuytrT4yCN3FWfiNM
f2/qdXjMYjAvkrzUZ0HcqMwmGMLJqSvnoWuy2xgxHDfLf2YGcP7bescIoQuBKRpv/2eEsDWxrl8K
ztfy0RZHKan+4TKzQaYVVX5y1rfp8fhJsScqAPp4sEEjzyY+/KuEqP4ntlSXEaR/T25hIMvrFtYe
cNe8kF0/1iVv96aCw/R3ff7OA0AJIU/Nb1Tyov7etMSQxMMzBV0vlbj4vuZPPHE/6PNFps42M1IL
qMzv7kNVrui8Z+JDqK9mpjvRPsmq1EB1juo6lJTc73BAxp/aqiQiuDPRBiICwo74XRPZR4KC4G6S
AJEDsK5jNVEUgKlber/st1FTMb4F02iuekIyl3QUFZe4Xij31bojHm4FZRtXZftEqXzLUvhZTQjH
4vNth46bvYsFDZNXhOpE6QZ3SuH+lX+8oW3f0lVeeT1lJ683osIimbBVyJeTGo9KcZfVjYNkYrCT
vGrW/KxkcMkKyIVXbv2/pEQOXhQ6wgYfiIoG5I/Gn1VF9QoHco7qoIsE5iSs8eu/j+Nb+Hg0Uwmk
Tc008Ji4M6r02qcMTBS/6Epo6+q7FyOAPTSRzKlJiALmso3ZoeJfHmXSbQHHsolhAPV2iukZKuIU
z4Q1alLTeFZMkLYzkM+y6J7OOC8K21gGjCbSLkAVpki2nG85R/++Agv8j2No1xc9PDIHZf0xsPWu
h6YqEcnZdPNJNI9gb4baKCld4E0Pwo6lQvm77lp4MuQ8mwmFMpA/d1ZCArb3tRUcvGGAz38R2Ejt
swgaJ8zDPTxknAnShdz7kX2AI1y/wqD/3sf6VD9sAViXKg117lLu7tZ9ygAcdb91H6QcHXt7BUa2
+vjl8Xs+bfB7CjaLOtWM3+pibsEuerbMieHS3KkUMVzNbamojTo8wSjZMnYHdjqbAraF7IBDZxgn
zsi3tiFiHuD5RzNIfHbtcPC2bnyDRZHHKlGPho5rs/PywBXX0ULrlPKgHSnBbTX21huBqArbZJDD
tbOLYDFIwH2H2t/rSurrgjKsYLUlGvvQTFMKbRui84FNASCvDCSVFIcb+V0J0lztkjWlQyrheQAT
4uoXQd7+N6/p1hTPgVH46BAgOhJwdyyw5Yz4eQ1tznC7LxX0unQ0cVjiduCcsfnpKzLpeV/o/Vjt
wMC33cetIeC4iftjCtFh8icJcfJGvPrivuncAlMeMQ1xF846OJz/xCMqtLUesvZY4Qv0qRef4A2o
bRRuYCbGChG24dHTYRyeENfKbvHUEYxtzfoD3g+yNRfcq5EgLrN6YZJGjhT3EcTwBvOoPicQHjxZ
k2QbfRmLs9ZObu4QJ9evkxNDhwnhL7nn399AwKp0ybr86+w5Lqk94eV/zYYV2bRtTqaAbnEBwGzx
H0E8ioErmWCrhiLtkRxvW0hu7PSdd8j/EtbmERcXMRp7nF7sRVWnhmncd8wJV9N/TvMVFhg6pCp7
H1o3Yrj/vMNtGI8pbhUYaNLO/BUOIc4Tvkn3bgVMMIhB6VwSVvZfLZHIySmPQ0z16E0bCM8QIaoH
imX3ztp8CVqnGJqpkNVdoSXkxQ/x7sMr8cubveNb+3keBzPBRY2X8UK2qlEmpXv9ew8Vad+7qpgO
MksBI45MOEJLATyjZIoAd0HdrCgSDRybViSKeUUg5waWsrMOcYtX60u8rgIr/LHJaPNf5ACxJr4C
BbQ2LH6+w+ZEDXWzbb7HBA5BIJk949iE92gs3MB8vJWCosb6k9MdPrHsimk66psjU1E16+Jf1ch6
dg+379MdJXZFWVvzmYFcsD3b9cXBnrwF/Si6GVFEdvRHO6MhlYdGoIE/ALo+396zUfPydu+raYWC
FGQyXL+ukRjyQjduhaGIcoCi40aX1Zv1/pNNsQf2lMDDADGlILBY+KUIJRFR3jlzR06U7B0S/7jt
VX9BJpQ0JgYyWvvcUm57pwnXvkfGFVCvuPqigTolw6cosr065SBuqi/ohE8pmNcZQPQiJClKdsOI
gWcIKyPjboCdlPo5H3G0oBRrBbi2d6xb4Gr5/vH1RzP/+iq/QORFZ44sfVQbsiWzrdeDLG4qjSzV
10tDJ7b1QJ6gJhYTa0GquvPJH/ceSeSHTGN5f54e9N7mdplj3IXSFwF7+T5yJKiRbK7Al+7MFDdL
Kx4ps+kUl/CgK/CQPU5sAMwIR/yE++baYVekMDHWXu8rtSoydurAJKfbBXVJmqiG/bF03mgJDaDE
WyiBSVKB1CDlpmS64q3OEJF7Q3wTmxjqTDmQQIOOJ2Aa6zeO3cRQqExAp3sIRdjRd0C6xAutGlKR
hhl5yjbai4GViAe2te698GFzlcLoIJfQrMZcCWExocVm8rD9Oum5xUUxNzpGjro234Me5CNM/3EO
oCGOSEAVzviEDVXdm1ZqG7QxMeBdLcfDPtuIT04HvCm/bOaHOeSY08Y+4MxZ/nP+yJVRW9omrBIu
WUoNWt3ivjBoockcDNkiW/dLqRv4fpshHSZOp15MapSIJQbLqgle5droXw+5KRk0GFrzQTcnV+z2
Bygc6S50MGICW+c51n6kX5jFpdvxl/2kun/H6FpH5yQpYbqYh5P/DtMS7JteLOHG7sazWxxAY21z
B74E3gh2/sAbgqgaBZiNDrf8SyG3PkNDgXYLg86tZN+NMFCczhW+BVo/AX92WWXVvgTtiOPOb4K0
gZ9lY4wZm8e5uRtWFqy4YPuo0JLtcwEURVbf8sWQnhyx3WM2zhgy75kvZCdbeGyxnc3dYv827K4i
M3KizGsHqjKYpb7MZmF4ZOZvYu7VTepeN+QkUjbcE4gPcMQMAqOpisBf25uWqwNhJx8EsmaIxJLn
Dint9YURjvwyqzEwi/mwS11e6sso+LSsHsxm5ZzFA1msM+e4yOc3qGGje9Hjv8McPjCrtWRvM8pN
0qUxVVQYPV/jb92rItyrvleBOUgxbNwO4G6Fwu3nXSBErBwycYxYf32kxa/98gKiBY94yBte8QZm
LQxNjtLIgCVjqj1q+vGR4GyhrLLqcCx8deaUac0irq3ZMH6YU5pi88lcAcFoN3RHXgiuK2nIuQwY
QjChvglfoZ841FgX0GmG4wrOZJnO9WNjldPRsaWT5R6zkx+Qa8hivV78py3X7gth7ye6hWW74Sbp
rDW531ie6ugPmtAJiLTKUnE0mqaWrZPH7tgpK2O/2KGy7l8jSnQ4Kzf5jwCXroXD9nbfh57nbkmP
d6FsdWrUZUqhHuWCOMmPIRZ9v7MzWUWtFmdyWs2ngqdavjeJVgpre7SNuZMpS8dh5XihAZqtRUBI
3Gpm/VWSpGGzJnGj63Y19LeBIgsUJ7N965pTiFIJLk/jSJ5qaxRllne9VB2niy4x5zlU93EJsvBa
Rf6qSJcBCmyNSLpzwNEx5FD0Y0EKOLqktU6CFXJ3i82zb+47148YQUM31pj1kHJzBh/FpWDfKqXm
tuDg/9dCJOZx/E4oqT62cEEavO8h5lD3pORHQhyAJleZxv3JDay+NAW9uGUzKXgecgpo6wZS1iEc
P0NRmkNEp7cRYBqBOwhwTnbxbl2TQBe/egtRo4iDdFeM03qrPhA4T+CArFwbCCh4BmoR9YIneM3D
zTPJpll6u3rnH12UoSkQR4iKKYRYA5s2FuKXDkd6cPIOYnc3d37U+v8hJdCNGCMEkQ0EKNEoIoHz
5TF3HwtmKEE4IlYWmfvWDtG3wMjXZz56zOd5gHW5xzc0RyXvSKTMiNNShYpGcFTip94I/g1TGQ41
pIVIHgdtQBMGshYF7MejBKMyZwU0cB6YTnDbFNZmX3m4t/NHSzwPFPO3JdyVHTJ5O+pEz4fgoEnf
FU89+1S+2v42P8Wdu7LOGl23Vfdn7xFvOdZ4AHs2AzCk/xiQP0hp/tCPR4R+C8MVtaWUHYkrJDTD
WYx4D10nRKTVOR/g/hIhXbulCD6ZwVPKzt81WqmWmApQhYdXNrRJ1AdxcaCkKzOYKuyN1fCbYlxy
GUrofv7OPz3myRnmwWyzcl68INQAoPvOkYPJugB/98MkdcaG6dD1wuQwMfRZSWpKejqxVXrdM1WF
5mI/y9/+DuA/oqSntFd3Kha7wbpxBXQ15FRsHK407cdxzmwPlwZ2/eszgkKqArOqnRm9W6KujmDG
3mUTX7YjNWwQ0DbUN3YaWAHa51FWzJ93peQyswvci7k8Dyd9h0YwNza5yFO7WjTEGggMHHKhl2K9
snAa/MnQJ02Xj+Ljl2WWQieAfD8mk5IlaA6LjfzJAMqyCva81+d6+VluZyFtzSUgVURqW+CbK9Qd
AGCLnOCkWsTw2NawPUKT7pk7lX77Mnx/anod4gsvck7KzDhuFtwO/ox9nNnrbQ7d68f16rRPIgHE
4055ZZEO4Behqw7jRWgtwUMF1Vp+DUoSZfr5TDK6IkwJwuTAld/fPKDZBBnFGdOucC0hJ/gHGERX
4dYwSINdcQNumf+xGx5vnVlvZUrNTvROsvFt0pth//zAF5mEgAlo8LekDbzQeGnLk5Yyb0QvmWqT
ke++0mKCfE+Oogo6iaGL5ysiZJjAVCiBvc8bjFOoNcyq2KbbAHht/LkrchhGBaYVB/KqTOyuFoxg
20WAts7zOnxOeTWi2ImqVAl8PI6G7HIjpiEdNRh6zIPy3TohbrRpGMJgzg+wmoEQiV+laBCDY642
qER0UZZriiZBdP+pyb2UJ8ly2y5n+YLV1kBsXQAKeeAUCrpbfhxwbTE+ZHMH9PE0hvwnmFBQm3m8
1alrYven9KiaZriZke2YckaHeM6Pvpfs/JnvL8ApeGQwVTkPVYlkaL/2vJkFOXA/h6PdGxqSsjlN
cMrg09lDI5DYiNnmyv3DgqaJc94R2ATN2h9HcCfQhRSJftcvlRGDTEF+MnaQmMv0irAWQEYN0GXR
SXpq7S6KPn0Bg9vA14/R2ALzkEtbfy86S5oMxjP47Wv3E+aX7cOw5j/qh45OghY0XNQbFWz5zMsm
pkkohMCu5iu+bZrUBe5EONQZgI2+V6O6k60oIdYsqQ80otwN5YNTiCLJ+Qb67OrHD69onuXCofE5
v9ETlbjtCg8SsfnwbeuclGt0BLQMr3it1VxMgA9G7PjLkOapi/47H8fed/HCSgRI2aiNph1p+Uvt
v5H3CPIkY0usGHih0f27OzuQYkigi04iRQfRUCcjaGHbWEdLyUw08JxgQorr6WhVYDOLmBfPiiKC
hMTgcQTVdv1zgRIkNvdImBvomIaFiGWQuLY1Q0zmpWEk96HjgP8roinClN74iPue/izoHZ6AU8AE
FcHHgL7GNn/UHOh2ZAbAxB4WRfNrfEGkwPfUkcOHoAO5w9pbSd7pRaQ2b9qLMgk9D/has2FR0IsV
htH8EDc361UZ0q0bc7FR8Dkdt4DBVcDF9OWMxPGRjGJ6ufMPwUgCCtPKTyJi5UgRlvuPsSR4eDaC
kzZuMuZrNa/qn6p86y0mGv73CcuQVWCjGIfu/ba/pBkm+L98ob0mC9299eAPy0lEic//nddfs3Kn
3GMkHM2MWnkSuOcrufD0S2elHFFhH1f7jeueC1bZ3qafOlXEqfTYo1d7VFJsLKbiApNRyGYAzBMY
JycB/0uCHwKHSNFH+iclt25YYQ66bThTfBSu3L0aSp+SdzoX0rvQTsHN0siKNDc/aTBJEB9pJ3sz
FCeC9rBD04AZSd/2qXyohIE64FsCUSMSYTN1eFoBRqWEbtXVPS0Vf56cTnSfqSgfD4oRZ1Z1MlhQ
aoD3ryt1808PE5GA9KTgv0CfzHdELhvWMgacFwexEp9ssw9rYboTmhTzOy4oRTKidOK6l9vnTuBd
WtpJGjYYA3h1J4M0JXIEQbM5UOvFXL9cFVzVXk8iM8nbtXwaN4AN9hQIDDcsLg1QfNubcyMcRmXc
bw8JshnU7h/UwXHIFHI9HmonOZIx4H9kpgf+hrxignPYisER11AouSQNszrB1D/qAPDwjNBlBRsX
QYlbW3yfROSe5MCxwYG9GMv7eIvhJ5DnqzLIHCUspvTHWM6zSUbPjaiVjjX0KTJYWYfY2z3XHM2y
/U2Y/ruzAotAsXZ52gmvN+vhEaKC2NPy0Zs7uEIsc428BdcNTWOh1tsXjLIbS2SSwFDk98amM6Ob
HjBIL/UvxtEy0PfN0Nzd0uxKS1E8LUAQlIYHWfglr6agM94fZeVgZfNHpdXIha510hobTgRVppet
XWKGu8P8hyxjGnbKgdy3e4WB1rN+rS8T0NLsvCyhzH5cfj8JQ/bDt6/69GP2e00d2jT9o6s1etdE
gjaJsdxAZs8os00AbvMO+z7oCugSS68dGRME/a0lP5lIRh9+4FhRd9hWhIc5ZzdbHMDLFH/DnzwN
o5IwZzgwLx6txxVfJSZLrlu8iJdkthuHkSRB5EOh+cCjHNEtVcm+yFrr2EnyHe5Wxd0mIj9fpUjo
i9EeF9CrnfzTV2YRxG9sQeQVTv/OdRraxNfvc0t8YhQ0S0aypg+jFKsq1SB0iSVtYUWoGszYB6QG
BPlWRKA3rYjYvpM5WDIkBooMddLV/TCK40CHMMrMPggTpemSSbHfmvAMtql0SqQvNv6rSoumIw2S
6whlscv4zYW7HGo+fZ2M12YVblJkjUU9Y3CEx/l6xGpg3P/DgZm8urWWqHxjBeiBdxbNmGvWSEfI
e2hocvdXyyi9m++jhSpbygpzqyewRsjOV0T0MwQ7ZsQzauGlsfZ7m1SbHr8BM1Cjg0uFsnUsk0T2
GtSAyMriTKLzVABa2tni
`protect end_protected
