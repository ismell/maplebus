`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
maPvl9UcQIXB7Dt0/Du7rmaEhkJs8Kra0+gGs0DJ+Udci22VN0hKj2v1ClDXftYzfDw5OZNsMBzA
CdcWjA59MA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mj/yVYoKfTlS9Fs1l4FDAeHWtjrinclJCnOydiP6iGWrG8GH/4ni5qHXF7a1dwAgYBrPbhM4Z2tT
XyM9crnlGmV1p2DJKkdar91DlKXbVFEGKQLqxnvvCTnRkNaOMoG+rlULDhmaMDMvmRxh+8tw2M40
1za/g4BXzsDB5iF42Xw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UZB7T1GVHARV3upN0hardeFXwiATAM6i0qchKfIvGXgdcD28P+qkPUkEXS41c0titPluLdGSwZUe
y0AXOJTw/6vCUxrHvRMcErOveQLhLePIJhO2EkYGirpR2fgMV+SK5FHEAAfOTuYmw+oZc4giXEEY
VsrXDol4awmrD7A4GSce+K9yt2HRmKXH59u2inmVu7r6shfr1h3R+am0Epl7aIaqAbkY0Ng6avsn
wHGJ32G1Asao0eSnyxUXyUik3mOmuiCKTu7RghEphHuefoXwTt8Yt4SdT2mSZmYsjz1WpjoV4L5u
lfXFFP0vkCxPwc605xloTY0rKLRltpIPQWKq+A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n7D8zZePoA4bijdSCd3owbHZwgXC0fsqk7FzmqDgN3je7hGvKGAkDQlJv4gtO64L/rUE2qNTnLS1
WBMdtV5y956RrGxLKjDQbj34oHqYybdaCFs5S+qqTqZF2uSbESEb9CGOUv+jQxsqVZjP1K0BWaJB
GTcVIa7g4A7Uxruq4e0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CNGEITwolhW5MFruCbG5o3vaYmdFFXEZ3sAb3zOvh8tFpD8oB6IFnXva8qN/CGhY7Mzz+ukgWIAf
sWZk/J4zIHnipOqXgbPFoBvCvgauQvac2NvBvjb+dmsxzyTF0tZlr95JTI9Btt0bJMOH1nQCdFbu
tNdQFEmqIkKL1bPiNpbLSr3cLONBoiN9iFHWOWMIR8ygBt+8ssWjuUznXkVLial1HfZJ9yVJlC04
tv2aLCh91+OWMc+8hmxXOU+/dBHQKTjJiXpZ8vt9Sc5v2NyAfEJNUXG2TEL86WNQiUMbdK0OiQ6q
8in7tFDFlUTKsULz5YHgcDhQGflwA5WNE364+Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13008)
`protect data_block
XegsziPiQDmkXqECFdtfJp8UVUfNvzprvyv65SpQwkExqB5XuZWNP1hmAq2YymbMDgIZrG9h2uPR
FAtTwWAphpb9xKq+Fuu/QnazsYHTLyzVpGYlUFjqOAi1mBrJe3ECSsKFLIiVF3eDR15a1hc+qiEZ
xQ0tw5MQuKGnRrYWSIqjOxX5dqui/FvrYN7XNnwMUbPz1fLKzWTIWqrtBtPn/sq29q9SJt1aTmiZ
xF3ut/yY1/Zv+Ub0Yo9P0ybGIx9FhGhViQuYD96zKHtm8UTuS8oTz2W2ZRvEXiimNRMQm1ZQQ/1T
SQkdshb3aE9nzm+jkb8swm+KXdxIsF706tIa9+pmlh/R3dZrl8itZe8A2j6zmI2Rq66JjzV42ylN
ZuNkU7SycJPH9gknPOViRVs2gRN6PO2/eoLoWuvU+DoCd0mvd5BG2zITaIY4cKE7i7VDNJ2F+Dbz
C3fyPEX5flSkjxKKYSOzuMfS1X5repRanHQc1BCrC43ZWPGY/5OpAjLHsSyj6IEYyyMt6iqKP8Sh
5x+qM27tCYbCT6O64ZQ7OuxlU02QdAwLEOMkLioJ5CO6rV86wLfBuCPkM97cIDfi9pwGRuqxvCGy
T3DroPr9NemxwBC9F7JkzVquooAp5skd82JCSPlAWiSar1BMff65YBzhxNp+Jc3x1ZpRA2GlDSWH
jeN1TnXIkgxkk/h17rGQd3Ju36rGjWr0Iymn40olM1zUoB2oRjDc8zUEcXZUji8r8OHKzdi7aTOQ
QC1NPl1tyDKsNHt7kN00f8awhYtqMGenPEQgjhnr6x3nVG0ZZXlcZRbgNg2gSYFzn9V0iJFfgG9y
Sifs/Fo75RpSr64+hBvUX1f25geuBwSRD/lYN51OVWMA754s05o5+Osa11eGP4wLG/Pw3YXMkAjj
Y4arc4PbMqYb2W7f9En091qazW4SfY9zvXiwRq3TnWq+Vzn7eIfzX5zEQyb7QYgipfH7mZluNG40
XHxWLYZ6F2I5wWkbKveapUgodM7XqxCyorJgqjTFAUF2+3u01+jtMYezDk0XOsXvHArjuNn2UZj0
9KSuG+mQdLaJLm/N7ckHBmHG+lBRn4LcCWCIpB3geH3QmvnYcN90h9b7OHFTrlX2CgwVXgOqAA4c
U3SBqrIiZqHenHcrp0/Dseex63DStGvLMNvJ57n0lw50lJLfc8sQMoF4JZPxjWQoX//eaAJSziS2
tKK7Tq2g66cBNLblCoXnWL7Qcxp4kvfrfOCct5RFm12++pR7TIwor5q0E2zBksCrwybVwOzlnM4+
VJJBAGY0gXpK4KlQKYlEzlgjINfkM7w2M1fd21zA6ZgMDSrVWkEgCMfxoCRAfY18tdjyqt+sPABr
MnQp0sAaBTiqZ36lhGB321b4yoVDDyoI0HMEE0H3iIrfokZhfKV82uI1WRiSccAwU3h9yFyv9vQb
50r8uE+d8lj+5ynyvZK8c5rhgxmfDgIJ0SuLUDGkKEffJ+j4uZKjzB677Hf2WcKisv3wHpiiDX6D
soi9b8uFfnu4oRJy5GiWxtGwZn47rqNk8jd7W1CeDi+/qaWxDoQQDon170T9im2HObuOnCWzfTY0
iIZtSM2Wjd+q5PuQnmxnfF3lXgItiA9ByALsyJRinWtE5iTXhnN3utTvBMOJdrivMINcgn09o98u
nRxwVR3wmLr40rJfxPPWNizvkP/8hQihnGqkOsN8aHa1RxYwiu6Y7XbC52OTV8aZvAs8bKrLKaCn
EqvwaQ5McuYeztn9gpNAct89QZ0WR0DCxCdqow8ySdHekr+sSY5XVz+HjNPRdoa0T7uLxuCDibcm
A9zb7z+Y4H1+LbeA8kchQO8DIcMgk8Km4qO7+FTpuJGrfBm2GG6BfudB30OU8l9LUhlKfI+ogioa
QeQKR1GaqrCFtY8X7BRhoauGWkHexBdasUdR9OK4mjksAKhrm4yZg31BnxZFpB8hETTKU8HfdEAO
8DeN7Mc/CXLncebmCw3lWY+CTIsmMdTEvNnN36cogHbYJLfvn7K7j+gNU6btJkgk8zuecqr5DImv
Gg5gLL333pGl+Nu86MVcwRB+LLM1jwYbm3spwPvn8rCHtYlvpzwVmP3N3TdVakmBrOVqe64t5Y5e
aJ281WKK11i7mW0ajvmIv5r4ag4UnG5y0uCnZOFPl123otZxnXIsZw2zbnMjAvcZ6gF1BD7WTTME
jkkVcf8VegO/dxbul+h9I4Srj2ix9jF2XNSxXFzZWrrx51l9Whpn982PjoRfMBt/uhotz2ooLgqw
+IHZHWyyQMB5gGi2itngnbemY2ztJxaiQdH/mjwYCC+fhN16UmqfPA213+F+iELO0QmHz8uDZUU5
hqnC72tIjyFVvMQb93hT4LV2OPkmhG1PmDQOQSCWmz74/9S9wOAEAwyGFRxFENVAmiJOtR3G91vn
JkPY7kJch4di9pkNRweNIlL+svzZy04LT3HbCuQ1kC27hJI5lByk/jQosFBSXOu5qLBWokhah+yQ
coB9jZIgoONg5SADTT+vVtBxUIIjxQGsV3YexXIwpOJ0AHkZOXfpvpqRo9M4IRZC3vDueGUJGagx
8+sS2GVwMkuyeZJpNytMK7ZvtTowdc/FKCOkgvECs1ytmnoahXlT6pVHpJK5vHAKt4C3vBy1CrQ4
pAXLOnwjxtrmTnzBK4Q6eiUtOpyef4jHvCqScbrM/6Y1KCbP1TzG/TUbpm+4xcyEYeLHXRLTEVNp
FJoJflLBmR3WL7QVHiaUaz9n+XFvfZdTuiSv9nR3Ol+ZpdEC1ZUxZjYDq4HAWDhqzWpiwrNBVDPt
MORTwGG0PLa0IFLzCiR7pLJQcHZYkuAGQFzC+HJil88fQnTPG5XkVzLKYNBEOVzyi/qjZvkfHx5y
qkmcyzJI3SWO/dA+GuuV0N5sEdc0OHWqSRJyrza6TlCyBeP/toky1ThOzjhuUW3eeR1Zi+WBCCaa
/ik4j33oK3UP2EIuQWx/NlxaFTfH4STNNdQqRfIPLwNC8i3raEXhS7dJWviQGGtjUA7BnEo4cApJ
b1MA7YfqwjYmy3Rk8ANfWC4gqLwk8gyTE/NGueLOZOuYKYb3qGIPlGpGx5OjVIRhCc6kaO/yOyQD
krOM5OUkq6w50mE0ymaNAtDpT4sz6Pv5bdxxuF4WhQwx8/BVu5mwr2wXSLumQ+QZxF2ZHwbxjAeo
HrUuAf/lBLnqZo278fPAYlGNoV+kV8VD7YMyrvn4oAmop/5mo4PT0H1ghFTCw5ZRZZ7rpQyGgtme
YXA10k4htPNjdUW9MKUaxvcaw3rxiS+Fkkom2YzuoLL+KLQM7v5bDvfUu+XQo28ntEgwiw7WUfxV
+sTwc6cRJklXHT+XXRXuwk7DLqcKHu/2OebyFXaGTdjSHxzMJ8aS65/toV/ltctSsMDt0covxxKc
vU0xTfdBMd7/JoKkN6FdzUXgaQm5FkRSzAVQxfActorWYqmNChjN+bmVVjTGYqn23jv+r+KMbWFg
3tQ27+rFKQYoZHhrsGdJJSL6vc9ffKgJZDdrILS7HeR+IuyqR/+ypC+RNpa9IQJl/Rz5s5EPuMvz
2rpt8x/MmOFjR6FpZcAs+G2+CfhaiGOn6f2A5Ww1BhYBg8j2MbjDUoS1B7ZFlPH9twYwqt+24SnV
5WteygrXc0OCOXGfeXEOiKp+mSNgycLFST6/BrP10hgaTEINCsGjv3MnwvtGpvvOHAw5quS+F8tM
PXjGN/Auyf8C1DOG1maElz19HcmOY+jABXeYDAamzuvonP2bJ0IKBR/rKA7sIPRlEcArUGyKzQ0W
6aiJiR4NecMpmcB56qir04UdBi7Avdi2oOEoYKl4B0Cq5HVGLwdmi9iY9g+O6c0eps097TCD2bg1
LvtVGucM+QgGmKpjmiEROXq/8xW+GZZwuH3BOIuu54ocytI8a3wJ6dXuXD8S+DPVU2wnQlQ/iNQn
TXoTGNC5GSbAEzB+lXreXNz4EPz2ogrUec2YIai6Fm1MsNSVFZwlGTa7q2pSnQ4YcJMIqgtrcPEb
IFKecDGomn5wMnmEzuRVizqGQNAZ9mB+bywQv8atnFc1PqsgzzjF0+OPr3PALrYsZhLQ8RvsSL7H
psmyr1UoZg1HoLIMQgUFPy18uVVXnuAA3Iz99ssDM4FTkmRLnfY3gL/TX3D3lgjRg0JD8SeBbq2b
rwrqbgakumz7ZJ+5OcToD+CWSXe8UD1Yw4vhPjFppfNhDm0JNrRzFGHmPX/D/tZC8wAhDoZhlJyx
ptsX+BIBbV6zz2NFYYf/KP5fIgUHHYU07nDy+41/h3wmCOKU9z0N31d437N0iHaKKaCNJAiyU7mO
QcXUNT4UW4DDHJ1WT9py8qvmYAEhs4/u/McJd5I8mEaSzt7IX1L/qLERBWTRWys5mFhSDuepa2I6
TkkmGF6l/HXdU4nMpwOwWm3EQDyYmOs4kAgCIy2P/729R7cOeA+a82BATMZr1nBzhOB21Dx8J2PO
psSm9CcPIhUvaTLhl3Xg33Xkwk/LCNiK/G8iuTQ/bVjAhER8eGpj7yE8YDngzk56j71j7DWx1Lnf
8f+y9B60AfXH3ZG5jqRWg/GO4V2aauwnS5yBCEg/V9uWahVUTyAOtl2Sg6d656hJIEoAO/VTkHtS
Yuzr7DhnmUvvw1/1Rmh1mnxKTJRbhba1mOJQwbWOnFICVOaNrTWdBENDELzK+BuPGtT62dCPXHQO
I/cyyK5Ev0rRWLetojOKmTdBjsY5HGecjH3J4qUBFeWZ0QIHtSUvj3bIefDzz+aLPQVbTTXeSjwv
spCdZWB8hmQvi0/L4TGxPeuoeejr/d0hRDAa7JVTczoW338u+mjlaDEaV9xYwdtWQ8yh9+R7BwWf
NTTEwCDqGtrjjBwNWURvlrKGB2PFJTrNZ97HK3ZkTwYwmAwEbasdao1N0Glxk7eZ+sUqGIIIAm6q
iGaqhl/vHGRrqy2mnJaXkAHUixa14t7CTQwMereH5J1Sy9gkr68djfGeSfJTCM/BLNJe61ePrfqy
7eUT8CgoJCi/sX52bWahjZf45OPThh9uBmyrThjEGjtbM0jFURp7ODmPjQGpLLVXEO/Oq3vPEZxB
aChxbwYSrkVUpUxm2x9vGK655huIdAnJO8amhdeC41L5Q9TXx+7MT5h9RHjoZo44e26hZrOD5uO1
RIglI0oS23qX1P1g7mQCxY2a7hgUS4PoU/7EyGZ5K9ZOZbQ16cwFcfYMkVB6ruPccY8WuzPp8Jgl
qCd0jG8PCGbLuOQybnQiEG+CQZoj1Op12ZzlnL6RHy7gy3ZU6o5Z52jjEgc4mkNcDJKT73EScbl5
bvuvLADm4iJEVtos+ybsvPTdmTCVBDe2qZSbzCx4AWX4iJqIuotiMyRZKeohO3NuZJXN2EyQn5UC
rWUJDUAYFU3JWACn0SIMfISinZxwe+fWTxhuFkc6ubzXAWeTmin72jY9tBUMP3wnrrfB247NkWJ4
UexYp/7UbloOZaxsFL2yxdPLT4U7FksAmEQfsE14oJ0xSPvUmEr7aSBGUS03RkwoLdo5t05u9iUq
HGG6Yn1F9kJRuz5CXOWSNa8WHv5x60YbI3Bqj2Vy0Wr4FXHLhmElJ6Oxx142lmGQKaTxZr+z4hL3
h1aVKrdzxhHgR18HrBP6GSNhZs002iEn3q83RAPKCfG3x5sKQGcZIv5GX0rXHwpn6h7BDV3Iqifi
mgWZK1RpF7PFlOofg6ThP7DHc/OVZHKphtsNWtWNuvunvkXpRAfHrZ9QoCtfhqE6hbYxD7wJrCa3
3n5QzECeUUpJ4zJI9D9RqYrHdeIL81hoOV20hvVyZb26HOIsovSw+yaAm7J4z8gngm9PJZCXgmL0
AfMTBsQV+oOyWFf54u78LG9L2AA66qYorXl6TA3+BpnRnNMxigDYzP+aAu5DboVV2W1h/23IHF/n
G5/0r9mx2dJOg+JHd5ldoy0uO093GZQzxuKjfy97ADdeT7LBAqUhU/qXqwAJGYjoCKMf4eX7SRp2
tSud6CG0npocVBiAcpFbvNUwY7n5bzInZI/1swfj7Ae4w9YyIhKWwWwWV/Ysu3rWsiEDEW0a+g1j
vICFtkJcvrD+D5IeckMu0tiOQAruSioJLYqgbiaAHZTgiwVSqfc05htEwtSL6h7dNm8BxDRwgXyg
jpOCq/jtHe0Y02LNlhzt4cKCS4qRU3R3V3zEHV/7+iuon7mz7pbL8SKSutKWIAdBHS1vRLhs+65W
pO41C8AdchtuVVF4QPxb8hvcdT9ZqSVVANH0WiCAFiNrdxSawddEw6nsWEmXhlhbxJiyu45Jbhup
ah9OHFIugTX91zv66VRqvLFH3Jf/271oEaWOBiY1wB57GbVMIV6wbwaj+WQDZYFyW/SSL4Hj929C
XPUQrNAUKiHSx/BY95fhQz000z1q9a+4FLRcv0F+inVar8JefLYFoMMgoACWQccUqNt6VGwJbU5D
DjMiRi2cowD8jfh8GIbQbMI4vqvrtT0UPx84kMymXfD1oEsqLt3Ruk1n1R9q89MlFTfnlT76TITr
a2rQwvYDurDSyCRTca8URBWgXDtFBQ74ROauOEyHSKpIaNlodFCWNOif86sdQYTyp5Uyvxw3QO/S
Cm3rKkTxbZwMwqPUcxxcSXLRtZLbGc2EGbEKAUVmhnThWCfQk/hyqKg8MwCwWuOVt4X7jgxN86MO
SZBq9TL3Nw35oDkVxrtS5wmg432bL3aMmgxlVG6NBvnYCw0ILaMjCOXcDTjgPzrjcTzad2QFGs66
+NAa7UuHbX2MaHBMAJHCoMLo/7K9KmjjFI4mcMQS85dDkH78gGL2w9OhAe0fEYOEQhHpwcwlwDaN
9/8b3p8yd0kGd3NNxgBIOrzlzIU/9OqcCGNCDTXBOOFkPP2wvhgMybXLVSj4IilzrDUIqWpaozfq
RJuPD5PwO3WlwGgPFFOOPakK9liWAyMjFepHj8exn5UkTLyUQOmjFsKP85kMAtc4nxDGUT8GiyL7
wFLCVnh/V2kJJICjLhEZL1LTEqen5j5v5cPMBJ+N1r76NeqGSocKEgpULzzYYaLMg6J08I2+jGI0
kLGPZvyVB2ty/qe4w6uXCKatOKdTafgjNSq8K+3Ts9c51FcckKy6QrnRoKYn38h7oFvm8RC05/vA
P6L1EECv3UPSEa3g+h4gjaVMwArQ+NHcTRE2xXC+HJTwoXLjrNg33XlifsVKDuHODoMmC4KGZvRE
3erlRfzPMQ+1ub3tBNrD622KbmhcWZswuvo8meMXjMHD302Nopcn61jObPaZtCcgvuSEGTQUN2PI
gVVdVRZKJHS9L6gcmp0wz61C7lc6zIFhLHxvQ9TxIdRNQoaqYvj7kLOZrDhjCdAjSgT9sPjb2iy1
3YVZNmg58M99zsOa1OKnafS1NvJrNW/IOgg4a2Xm0CmtxYM2KSy2cS3F4cf+Fa8Oh8SiRUf4weT3
NQkGKEQVOq2Q2qBxzCyiBy13xXpGg6ZDelEeicKTNJT9+n8Qpg41da+YTOYK6UCM+2NANnRFIyRP
TSB8fKQTGz/YYjEtC1/2l2Q0mz7NS5KfS5LjpaF+rYOsfZaB1TlfPweJpkO2XHTz0oUqbXQNnFrT
PRR/9U7n1CGVU5PWRl1Gq/iIe1AhEBsVHgj1fRIqnF7cY0o2+VwtmfxhHbZLJeZMqIye+Lj+jvB1
o3rlsTsFrQOs+N/Gkygs8KF35kN7j9/q7vjQlogrc89GRvgxBit2Bg3i2kLY7g//hTkMjBwrFnAs
0Pp4Dq6LuLTqB7kEo4pX02esfFR8/Q4IO8X1sWxU+kbP8tYOCwe4rtwjJZpHtWPhTL9UuwwaGcZg
pf5fxphs0eN8GQyhW0/B2hstILkjQ6FeRMchdtipOm2fD5PjZ2zvoRQ13elt9yEYFQ3igbjtFZPh
1b/bjioLCfjKfsBKsI1Yk64i+iYFXz6MHbqGfuQSfE1QEFoU3j+hpqridqIo2uD9ropE7LKnxHHd
oFwqf630yNeuIE0J25WJKaT/LuiJv+wi8b144Lod499oZD32+XBxsmZnMMZ+14+ZqorAG9MjEW//
UCDEVVKhs7WEyl6BgZugkMcoLdypafH3G7S8LBs6upOPgcEXoz4YVmjF7YaXs4t+BkCoEpcQi+Zu
3MgZoxgEf5tO4MIo+6CVaTQk3N2HoqZC7/VFfC3cCYjXFpP+Wqd5Sqah+Fix86TFeJ+SFwrkFKex
9Vuu0ohfn3mJYUWLlQ1pJDJJ1sFcfb15dRx2XhxyBqrTSLQPKK8+rHRr8QS1z8EsjHztKTYV5YRB
Ye4mHcsY8UUXL8M9YBFb21xqcAdtLoMfk7JBmoICiaEzKIIc7A0h3fq7EJoSLEAyidRmQzzxgG77
K8AJriLRlvTuLO+P0/naBj5f9GAQ78UYW0/MJgz74HwAf8g0gz8n0DQQAkKd2D0THxVeNGHh/pO8
OmQD+2nnUwPQa4HGL/H7Or2zy1MCKNm4wDn+GlCmWtgs78VIsd+lsBXQw4O5MlhGgbOXQsTAkz+U
PK0Uo6hnxpVqPNwLRc4hzyAwKmFq52Ei+LT2Rew/m+iqgU9GB1uzQaQH6461hPwF5h3aNo6qHuZ7
GVAz9O0xuqbujGQyxo3+lSGg3FVNPCj9knQPKyNjRYctiI58ReT/kbTBKwIUsvMfd/tYtQCSMa9A
rIOtxL+KKa9XiKJ45T35nhdXTPsFiw5iWwCdMcLTwcNB5ds4RZeT287LrzKGBMrZ+iJsyUF8L1iM
ThbyIFE/WIMQKbH9YSVpiRdAm7QUw+wLTR4Gug1a+IJW3rAfxngP8AiHhiLweuX45p0dHEdkgP0x
ikq3ApCYQu7ZoNH7KctUs73wD2RONitlL+RMpgufXxQbapBGetW01Qh00Zc6pI45iMHOKoGLjXgx
fvokafZh6iZzXYld3yCSb6CqXpMGYhtMKqZQ8mO6tLu4e9r63GXl6qAt5HERc6WcS6ECIZxy9rex
Zujv0M7qiU2NmYDWsgU1Mnq+zM/Yt2wcoHxK8mdbQJTcsKaSs8mUaQRxk+G0gFC3WH4GoysZNZJR
UKTJhuMDJE/84MbIh9gWvSchM+VN8Sj84kOVmNOhBj3bWI6afhiM9LBsofPhHyiyhoteejBu3RnC
gUvx/qG/XiP5TKP0XHNGvOlaLq7oArsFSx19H7c0tG7rbd3y01pQTZkMHglUkVwUykpq0AFlREJ+
j9MQSwe240Sk7Es+UufcnGrRb0dbaNlMa2RHgInr40f0hDcni8kVrqDdGNXpIoH3XqowV9WnZDcb
lm/uMiBD4FB3T/SKIZBjwpJ4FgofzoAzH7nT8Zc5TFyjN9NnrdG7S+/l0I7YGyF/tyZcxts7ziQn
Z5BhND15Rg121rvh6la67FYba3/HzKaTolgesSA9/B6SOGFBndAuv7QUc8Rtd7YByA195ydYYrND
2S5ulfdd03RMNCgbZFtVQmrRqKmSMOrhBK84YAS0/fRLJmh3F3yvpRMlyvdT94WFTuoqn7TgUYmq
kpznc3W2tHmcqrJWVZvFCEI0nsxIAMZLAUKCydrzSQNCLC9gb45hzaS5g2EFBovKfsgmIgfbl9WG
H0qWy2DMo8Uopjq2053mLJIn/eKk9fKwUaao6q5914pELhH22G+wTXwoyVczSkmSEzxQL14kn9Zs
ke1GjifNP3uLQPN/odUT5VjMceK+V6gmaw6P0dx8V2WdG4TJrtwVbQKjZ2FzFh73aIky6VqE/8qd
gZjLbhHNyMOITYQwDxAIUgPkFJAI5ES6rTKgr/tHgfFEKT3sCsepV+MYmOJacIfQlQ7fqhSHWxyA
quC4mr5z56dlyePTB8y3X62Aatn6zAMiyF+n4yGg8PE0JEpkwSw/2rUPTPhxByf3HAWApiruMC4Y
ctHPfaSD4yX2Y6tCnK7dWKdD7loMaR5sylLzoNDNpzvFtBQl+sjK00ObRtTZfaXAjkQSY0ln+uW6
B1h7WhNMbqFoF7HamrRA7Cfn4k7FMsLfQf+XoQ3ZSIvQVDxrFbLhbyz6G6V2eHMGD9lxU7zsx7DY
9gmT9jLJV45yF97IJDaXDq3yvdSfxfo1A0S50PrwakPc1sh369gFU9i1xNSl/8XCrrTR1830vCQn
1M6hgvOJQ2D4saEcQOaNJzuBtNRObt1xbfyMJkzLf6Rtb5/Y5xSwY+bKWy7sHncPjdqX9RMU9itY
nFYlPMiub0jDdKbvNfHf5cwjwq69poeAUeXAMd1t/fkhAUxZQu4o9PbfiRd2ip+w+wO3slz634/u
RpVF6gtZxa+iqTBB8DKb4OnjmempqNR5mOYmU8fuHL+NqYOsvPrecOcnbXrAOU1DBUrj8aNF2q5z
xvJ/cxJ0Lzsq6aBfgxQdkUoEgApa7qwx//oOvV+fZrxvU4soPV91Dh62yxTqlo9gfpqYNYlb17qs
rZfYRXu295mkC/el51uZu8tir3jFTjEgbIgeqVD7E9mK3FLNjKU47ySd83R+I3b0ddGskMnrNG83
uYtJe6rCfvnTBbpE8AAeiB0vA/JA94IR1/eOhcE7KftsoAxoTShPl0WKkQVOBPmN5A+w5QSzrD/L
s0NvSuzR9abJ+prLDaUjH60yug6kj+W9q2orVLR2in2DFWMswcEzD12hwu5CsbQtRbX/rY9r4oiy
4q40j8dq/dhzJ+9yrIU8E3iWZbgyr1p0MJ+pt9RjF19aWdxo/Vc1gAwL518g69LT1FjOG9VnlpUl
4qWmSQXIEKvJOgAM4nzv9x/fpxNWalwKASgt2qbzmD7aw8TWXLErdLdbQ30tpHOxmkAxRvteuU3Q
LeYNWQxkShPTFCDLLwu2T+MMbNBa3QrjTT2sJaLr5js+7ncLPBETb5zWHAWCk1Igy7FMAagHU+AL
A08/wArwzRm5O2QBDdgP0e/dtDbUHvPHvhyO4nwdf8TGwDJc5wb3cq6/O+UXLfLmyeR4S4Fipbuu
3ARTSjugkzarJ+rpKNDN8cyG4OFc0FhtrHTbhzZgca3V7G16WwNxhfM/TkBzMwpsn5hObIq7OsSN
ndN4I7R564z/CIaEO1lS6VdUoNKsQOyEE3Pa8TcFQVTHmNxwegRHrqbFMSNqh6JZiL/g9k3xzmNR
6rjCaIXr+Hy8gvSWD9oeeD/48p7xYbf+PlTegRZfH2m080OsP9hLc9mRSDlauKPdOk6+fu5AuNEh
xdepopbRLKi2zo5PL/06vLvlcas2OYkeMB5rEpcPWA1NbQxe9Mb/wTfpGEM+5eswM47QNTL5PmMw
1f3IdvsKA4x2Q/GcEPfYhvX27nRr06ovurqIm/pb8GLn8X1rnJXbEREvW8KxQFe+umkmeemYU5/u
7w5+Wawm5Ny3dF33uIhKR+ebpMGkLcdPqohjPCBJsKn4peImEpmSJ7E5FTbtx24ubeoLt1SjcnzY
UKax69D64WyseSzBCI2eAzQTZ0OVRESwgZTeWcHQ6C/fSBZM1JbVEq3CXXkpFMmy6zNIzTe1BBh1
0+LY6BakqWrHWqLdbZFkXFu+01XofvlfxvuAC4PKPKXGAEb/ajo9ZgwJniB4bRgUfzC0803TjVsL
qseMMNLrzEX91NrMeiu+fFWiPd+BvLqMa+SVEeDH0e6CzR/h+VgCRQqZltMXBPIvMgOKZv8UuKhZ
7xg0pHc6LgzqzSCGRK2qFIu19mcPGGHa7x4VHWagMTFFXcQwhPx9GNiQMBgRhhESDFKnQ9hu9lGZ
4/TfcCPKGceLY4mP9rQqmu5dULDiP8MHSDnnyNsdbudm39YW7KtxAlPGgsOdda/VNqBZow14Sxhk
/MiSpUynWEVMoRGlux6Bj3gqAppn3yPbHoW3EIXizGXQiOakbfu+TY7Jh1pjZKCLvieP/Vl1X0mf
pL2o8gtgvqJlvSyw5AwXyf4qYgT8I9YvTFdo90bxzdGonp8EtQDs36dvWAFmkdGWOriHUBMDMY3a
o56vwY8cV5MuZ5+Bi/UTqhscefTaylxmtXPKKHhkclSo7uGmu/I9SIzt2dCyWSkdkgnep0Ndhi0o
6xDYJwb/9wLSeYS3ZpuKq+1QVUZDBj9kt9gSPov3nS9TmN7afyQcemoZZQ9c/1KuZTViBjMAriLr
AjGHyH8MUM3jn94q3Bd8f8oOm2MoW3h/2Kndubn1OuCEWoFJwJQiAbUJgLgHclS3w9h+vvA11ZdM
4noymx7opHolXzwveog3cPORalQHL8P+OP2xyRAIxTE/PHSr8L89qUrqptANO3MheYbkJg0hvnP6
sFST3Aon/EhrY9QnimY7FkZzTYY8CT8b6XPP772m5DCNMXFSLsfT9wu8lehhJfSwSdv1/QzRnY0W
DEBVuTr9+IqjVqvcrAAxN9f4kazohRcDXkHwur4bpjGjRUlDWkNRmhBhKOJPSEu89XW/PUwW4ZNE
nUNJD+sW5n8yKBlbpyx/o9hoiJSZQitPbxuUd/MhT/BBy50Unfk4HpNepjj5P/DVve3jk1tFa+Rz
xSDvIaAtdS216McDitNNI/kM23aBkZia/3vb/ARSwx7m0V6DJ4oPz/g4//EhZL1n+B9LDEYAWuth
Id+r027GT3tR7EwvpGsgMiqK/NlVGQxKM0wOUx2Adp15Db1F0bs/L2YlqL9lTCKX8sEIJJYEM5E+
RzvqXxuA6+W3jRdfSk2vdHb5l18iejKEZwpIqz41u97iBW7duV0dnT3zZPzJZZI5rFAk9YLBA+6Z
0NP2pZc953glQjGLdq52SrWKIIfxWuNHbUH7F/i+LyyifTt4I+pVMJFTzLB+mKO/yOGQVYVNx0eZ
MfOdErB/aak8mBRYvE/DeC8MWO2+0RUPRuNxeq+zQ1hGfYXSh+y9JHI340/ZykkuY4Pkz9rdSEKH
iCID13hl57ryKLzOtZn0WgX7tSV+qOqtiI+08VqebgJarZdBFIunr0dI7SmA6V50WuEpfWOgrSio
YgDvR7JlXxgRppxkCT6d+rT0c7EUWsyoWxPTWfEk6e4cz2kCYPAAlV1HVIAXYdnqbxPhlRkyTvbD
exBuHYo0vT+avURjyFUBTxylVwc3D5IrVa7A9gDN9BKT8usCNe+c9VlFaLZ2cJJ0Dcytt75VhZBB
5NQclqlsxKbU7tF2QfEB/1P0tUMuYQEhPFdYlNszycw2fqwONAt9ifwax2vhjusgjZqTGUP+3NBk
t0CLbaDj296+DL1rvbUrJZqj+tdFS+mIBeyuQMmceWZ6a95BV8nJUulXs0cowAKgVltT/HivLvU4
iLuXxzOnN/KcERm9SBoyZMh6eWPE8irmfOt/4g/E3RC+BBpxpOe2q9M/nShbms8Ys9FP9CJoB4tz
FophNeHMFV76808crm6UVY8kZw5UmcTV/AYWo1pLDbS2PqHVUM/biF9Q3y3nTsHqaTpb4PPudzaj
QnA+7eNaPpMXssREgTQw4Vw0aPd9xeOAVlJpgmGiZpHCJ/Ekw96Qnn1eaHNNhva9IC9ndtLtJXso
cPsFLnE3lY2hihwL0ZHfOOIaXoQGCsydUT4jNR9BysSM1O/VeNdnVWxDbUXDhYwaxrTUucfvSZJ7
JX7Yu8RRwwl2vTnK/myUOV2Bh0if17kHcL1TLARAJCcZEWbQgbkL9Mr07VCnW/jhsvOTZcKdy1Tw
E+6rSYAowshCNHXFH7DYbL8AoAsF3oj/OtjqpywXVQhAzFHESMa6+mXyxSQwZobY8cMoZiqgeuxz
FS+FDBZmDs8FvH1WYD3dgA8S+eC/CKDqAPpnRfWh8Pl0iglR6iRSZmmbJENSyFqnoSmr9hOC8XBB
YoXDuAT+/U+GMW44tg3zcMjMei1yrTIjYBF6yQcdR4rhtgoS+GWnfrp8YyP1jSy7ld4jmHvQSVRR
BAfCaoCtCuEvGkFrF7CZRU2Ha/FsAPpS/GCwFx9Bakohg0alpd3IGF/Q8zd1ZGG8oWJSJ6SSFDJC
r+VlorlZS8wNJlx/upCXgOQyLcyVTKl/eRYDUwCIT+pYF/+070zfD26taLUsp7Od6qIyFKzb+Ry2
IUuevwPfa/g1LDk3Y1lyUV5vqzzHVn4SIOyN4g+Gp2se9kYAcQDNyYN56+L9Wyo8gyBY3Wx+jJep
T8mymM+GI2H2EYDYUJLtAA8AMbSO5fzYwZ1suYvfwNT9NOnmO28FhIn/BsalaaQznA1pdUFP89V5
vprCZsmMLukOoZ2XZ4di1lb0YdCAJKxhRYUXCR0GGN5tDs+cnH6DWstYN5FUzzAeOVURCdb7pGOV
N9MNNIxpVn8I35hEZIZerGEVwn2+JsRMTF0bzpdbVdwIhdwg/Uu2Zz5sJ7jDOQSf8EhMyDZZweDU
t0SJ1Si5GPOhQ1EiWbWhDheUxCxIwA+CaZgeUEizyK61TXpkJzYMQdpY/mIFjb7sdHDUPU27lqdO
ZWaqF33ZnV3bkITGsG50f+BRdz5ddCty7JLOKcczCtnAhj2Yw9eiseOHoR+MCFG02cDs02HDUoYW
aDPXOFXSLulYvJsS9iS9oINfC5k1g2488ACJdx3cBZ5QXkEDJM/r5mClRES/PHOy+4DcfjgD3c5B
JV17W2a8RTH4xExOESNENk2X1D9Z3Z7hfm/i7tuY03/FT/cLVMqC1nYtt9vgdUvBV7FL+8A603IF
Jp465pWDiSqSNygMOJw9JZ4TDcWwpNF6D6iC3fwH+b3zg7tv/6wimdVO35zgSzAQBNzYfu0MUw61
0eZsiSyqpplVuoaGp/dsNMqZ1wLzEUz0njlNxjtqJBJLRkqW1qX4gzTm4i0zgicKYQNjCpZBE0v5
jbHhG9TJ9uaLApasDphiRidBI9h0hbEHgUpgjN5NZd/7FTolKy0N+796QhOmD0wyh9pKBj0wjMxB
IRFJhie5aRzHoZ++plAAxZEa0gvo4JxlrqVpfBM+r51RpGXy0d3va7smJwjJXi9t5//zup71IfDw
NDgm9QjFnfQ59wt2D2tLoMtyj06LS4OMzEvA46hnzznU4MUoW9yhIS5nioK3u8Hob/nBCcWzT55g
TMborgmymurAZi++ObNz9ofE2p38zA7H9tU0U4h8Pia050eMK60FVBlnSLhES+RCrwysZ2u6v8mI
zt5KuOr8/8c+dHAFYedwOaZEH7+04Uzh5T4n7wk0qZFacY49x1LRFe3w9FM2sKzP5u9Txs1ZvHUF
GFI0yOgWUFkZyz7p0Dsf5h/30lKsqG7UFXHsR+/Cpwu5b6VMmoCk6EJgt+AtpvzogT5oho/B+W7R
1/+bY24NC4KKT5o7uFITijIAKzLak7Ev6uXILVetUtJotqxChQt0sul//IU5CRrRHOLys8cJCEDR
kyHlFCd21x02+tk9I0oVGV0HVqPtxxkDVHn9tB+Ns8BwDRwNoJakiCa+GJLzwGSYmrNCx4jdAoxe
4J7l4GsZXuxqjpRNIB4/HGSwuCuvlRamESSHzd1YD3p5jYuNczuvIfSiPKLd4APnsqSOudvBXx09
2JPqG+Hjnu5QzZHEvXCb3+udxeyMnIBLKtFsAOau3X7gad1hUSYh2JU1vvJ5zre8DbVJYtFhEh4H
RnQZwKSB5Hs34onSWbX9wARAMjmRAvjzY7jRXkZ9NVLUnHfofQNZLk6J36awXAI+OnFJNT6K5MjJ
ZLIVf7uCOKB/eltoup0mfSuXIMQplNG2CXBQHtr62AW5P+qi2ov96g7ZKXiM4aZvgRIvNjKXcJIp
I3iYZsmK1EWJWhzlqAVebQ5vsP1H+JFJyjrXCnkcT431XXF8KACdi4VglqFUstc9P/Mvb/1vh56D
ycgO60LexuVqaM+qhnkV9RDccS0S10LTO0UQ3IV7hYoWdOTJRwIKD+r0mDcqaGIZhTbWF+4wKRMf
7LP7VDlMdeqe7n2suEE7J+/ejHWdxFXcoJoKN8d6w+CZjWuw3RCesoYpE7YXcg+iil+Ppi/zzpc9
3OPyO36a4d/vtaakwVLDieV3o8ZFa0QBOzsmOL8wbU6ORM5N80KVnZDmbeZije7syMwTTjYgaS54
0Q98A9AAOMOJYCmRcLEcn09ZMWcX2Z6hPKelK13LHbkl3vhFhercX78cqf2W2UOPNHcEdg2i+E2+
MIewPR0x8jL009Xd8ud45YtEtybH/C5+zdi30LMGrVrYDqY29vyryA2W6nAyd4Mrr8ogfOVI/1hC
ZzIOtq77rZhyvFy9xS1iIy+8C7Rpi5Z8gZQgpi1tLb02VCeA5m5uT5O6Mt9iqbHge1fXcZtps8Rw
SVOCMcheIOPkAOotQ02JPMScXZ5saRbzZLpyp4DGWGAjOgAVn8p8xknnRw9EWHq9KjEwybM4SLmR
ZSAQR0jMlsqwTXTwL5PNJlmrPH+N0q3eXEqdhgjySO8BZYLZzCQ9EjxPTIlmJJGKnU/Y9SNze7eG
betHh4WW5QS5Ke+WpjGv6ednHaE3uqG3BaDstsXET+jUyYWEc1tK39KPV6KsqwpPwCWu4OEwQJoK
40DBU3ei9vVd+vdvOUNEC6fVMBGaIzGP01duVSep5IUb57RRT0yHhxdtGs75Cil0Y8ZvYdP8t9tx
nqiJuGyPwyMU47Clvw0tkbmE4Vge7WkhKc31/ynXKSyTKGYuVFEUaFczbR5wsm31BYqGfI8ika1R
moS4MXK8kKW5mO87oq3Zc65GWwmNWOUvUY2HvKBgSsF3B9TS+IV9YzL18NVcxsvn42uIXfJW4k6h
lauNaDvldpuuOhMy1LWZZULs3f3sIwGapV3GY0tUnQ1Lg68i9rl+S0Y/VdB3Z1GtdpqEItTQ+wNC
fJvtXbo1eq6KvwxMaYkHdfrvFOwb973rU3Eg1I9jY53adNqjXIUF2IeUnjiDIe2RsfgPzjyv2tBW
eiIzA3FB222TKxSm5myZzcblgxzukj5VeCff2Io96aQ7XhYECko0XtFGX1asv7q29eyecXVy+1GA
I9OjaVMQi516YDjxM7Z7ngvueVaibJb9uWWpCkk0q0qrcVVL5vZRdWaUEOWsLi+Le7/6/8Sclnrf
pPiGT6XVQpTW+iROSGN2oQ7I3edB5TQnyGIyl+Djf2v2FVo2w+66zMKmrKntuDe88MQlg7T6MWEq
/U5sWk1JnJj5lfEvL4gX37p+3zenCn1tg6pbyh0/oD7A8djR3izbjBR7U3xoQ7vwMk8mtZsoqfLC
eZdKPGa1s5+WUm95kp5n277/m9HXc4lsR+KN2gs34agrSECMIKPhM5yEwiItytJi/WznN2bEdzXF
umAxJLsoEEYDKx8WFw+D4OP7Va8C2gi96s/cKvGWaIdhOvBShaK7+HS/k0kkU6APdXVdU5FyDX+K
9GHGAmzJBCEhUihhbFFRGjuKPc+4IYpU+yYsAq2vKeBJfpPVteN5kxb1T8VD1yBUU1T1lLjc5Sf6
WpNuUSlF2UBDefC8
`protect end_protected
