`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UQrVVx0Ki+S9hN4EA0XVMDwAsr5N33/CSVu2kBhaJOhzSXT0t2B9E1Ngy23ilekqSUwemUvC3J/l
wqO5cWTVJg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gq3Svtc1Qc59vccEJ0VGC+Y56URSwJvkyotD4yYAy8fMPsPnXM1Gi/yAAk/a+ioarn1g4AVf9cSf
JBiWcZgk+/R9frQKH/bjFbrlhNeiXUtt851AiG2NHUZhTis7R27xCAYEcTQC/ughB7GqQ4/ZslcN
39hccKvcc3cXnmd6Gb0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YdWaco8NbCBv9Qh7Oqv/ziUUS1qViC8CM2agQKWL9a4Sbaesq9OXhuQYuzYuC+cW535ljhhsaEar
HPzVXFHeyXDZ3yCXzpAKAEKoILgm5Vv2UEorrMelt7kdRTsTg+LArFsX7rRuoQ7oZ0oSmruUl8UX
otFtXb4D5gaIem2Cq2v16fEfgvMajmuWkmnr1OMT59evXymKgPP81ricdC1uORESygSCiGCjKsPd
uzsavEzh+U0h1OPpDaqmYmD3ma7RKq32cNw3v7vbKiiCQoUSHdSaD+lo2pqnOuZqH8V8Zn5eVrk5
Fxjd2MVswJTYQnrRuNGGWfSqwo/gm+NV0U1/VA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYr4RXzxhcg4OpTxxqArhwoCZhbC3Lfl2TJJZpMZYRdWTBMHodFFiDntg3f/p+r0z4iGArJ7wL4P
tcA6C0BNTGqYMXmphSkLDdfoCgPxKJZ+K1JXO6wkEO15mF4C36Z17fW+pZjt/imMxvQQDqkYmboS
BygNczRG2swS89VUrns=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jIr+NNJ0cz+3MbFTjfgtXaGeWxsjFiGIMbU15l0Cd0jrd90lVxPylhSPGhfZae45PB0D1RVjG9+f
Lw8MkaSbePKxTRoetZ8sv0p5uM+ShaHWq9WqBjl7d8agXNuB0eA6JI/GzpFIKOBc7vkD3gctbtHw
Eja1O9iRmGww1ku5nKleGWcds+387T/vyyeTXThjNEf60J2H/gQy/4jKrIj7DB+qDRn9e56N7+iR
eibZo378M1mg80Q4/GoBfZSFi0Sf0QUHyQay4u0hbJapFMXRQ7b7OPYQhmGCfELzn5DNusM2LL6f
fduFcbzoCL3+14NM8Jk6/PEcKrzI4+GHLLDUXg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66960)
`protect data_block
2bxeJKhBYI34JW26YLLnikJ9st32jw8igEN6bTeZvyUUXZW/53c1unyRrKBtdjzuuYOas0+lc6Tk
rQo3o/yr35etQ8/gUPEWH/Yan4HaYwuGQJ/KGCLOjfApBDUz6J3Nnf1jC+pn773sP4suY4J1NZLw
UIN85zOFQovoEZB/6aYDjJQk9CzftdIY0pwp6lg98UfUEsrrGpTsMhqzkTOVyiSCc6q9hZzEgCBE
ishUh4OTWAH0bQzTReUgRv6OJDz5nNG3zudiErWTGDhAKbsNuTDJrcu9VRPRnDNjIhMIsc0U4vvI
itMbZP+bPRgU7p733M67KBngJDT4JspxVRvi47/hw2uo/Me0NhBCRok/AdpF/ELshfoRivI2kzlO
WyVhToT+G4S9jYHBcXINe1ZK8kaz1NDcQ8m8uYvuVVMTmpAKQHLwD0WJ3ldNXeOEBfYKY1suqbMp
0GtDdOWmJ0GKGXJvKvFzdshBdZUZXkVGJoLzbONiMX8b5r+NKxtr+vfza1h8Jy1PCEYZE/JCqqqd
8MzY5edCijK2yA2o1sUoBBHONkhlqPXzDuXqO9Tfnjo80I1ysujPSEVGNYtY9N1hu1UlPK+PjoOU
wjT8s02dao9A/qkBa6Y/EQOkv7tVTWu6RhTYdX/ayBaWJWYECmWfXhjFxY9YQExFizdx4nelBC7J
pk/m/Qjhic+8ZY+cDQ6OAMoDYi8R12qHLhWxXBr96GFjIVGYtyFSw6Jzt1kF4PhOR5Hu2ceIRuEP
zZpuXf1ivGtgidlAt3JY79nECss3W9wQOyBDlAYlwfo0Spnsh4FONxGyiY55duwiaKjogOIRPlE7
UEAXiBbwbgwymiWnbP4dz/rGsRUsBH37rP+X6kQ9gewOJ7CWGH3kPva+9Alo80Lbu0TI1Vez5S83
5fnb9dsKXdx6y0HYXw40VIvcYjYUnOG7VFutXis7Ux39fX4Y3tQueZsEr7bh5W2idsFHSCdkB05d
TGU+qRKj8GrJYbHWZ+ChyS0j025iwbjU6NrYvnArE0d5HHgVl3LKzbsy+jJln22yROPAcOEN9SAd
XTw7l3tgEu/oHvlpu/pej/c8gwjHFpF6rgekPO0srcGJkx8RHt/634RoEfOgWWX4F7xXFW5A6EuA
ozgdgYKIQFzl4zOad8RVl+FDuz+BP1Lp82Z3JdrekvWgAHVrT1khZPG6r+G4XLih3qNBqPGtvuC/
08uA6iAPxyH7HVwPihkaPO78Z1CqkP9VONrOXb7PE+EU5jIzS/E44cdcYqZc0c7O3lCLlOJYptzA
auAMfce1zKEpB+Txigj32+mewXuPBQfFqs2EfUOSlk2d//O8UhHW9h4OI3zKJ3UxVzs+nondOlst
DkLiEdh3OuGE8vJ8E8wks6NXauug7Z74NDI7RMCt9I2Ts8ylNxoiCx7wqvtXn6bZ8QhCnLY0Pi7f
mOKDfbEVI/5sjjiGDeD3/jT4uwgcaYMlulXuksp+u3lkrGP1UXT+HIWmbpqM/OLhZe3Idd4H8KyR
eBCzru0kAPB+nAeICLjh+0+6nBtiNwWu3rrMsJ8uRL0x9buwkoZoOKl61QbyEQLiYOmqEBiuGCKj
BoxShQR6wdbAor0hxM/qXX09PFcPfMe3tlz1llFwXlovtcI4u0dYvz45ChTLHAMMWCbu32C2RPq7
joBCWb93IIkePzIpPsA4L7k5S9UJoBZdqtEviiwB5yT84frKhpIEN4ZR9ABnPMBc3/IFEivtUaFx
B/D9vPQoU2IdMHbR0NvuX8qxXq4M8T2IMQd8+P3OThmxZFTC5qYXvTqrNM2bzIaTQvd+vjjRwt5V
JK2URAYblH0t/2Fena/Na0p3kySl37xf2v0PdKfhEo6kSzWjCst3zDKqsyN4gS3vROWEUjl2yE4e
gP6Ja4n22nDfhylMOcnfKPgZDyVt8emMtt3FcL48BZxTx5fThksQKY+yveNToAskb5nPhkoP8Q3z
XNMo6BHZi8spDpaYWVYIcV483w9vg8xzDxPD5/kkCMd6gkr+2c0q6Pmh/Mg6eggZYyM1oHJeadZh
tZFwy7nUXQhbM1IULiiD3PcCoo72xsRispqAwmmVGRaoUST7XePklOUnu2bPthS4MdygVzNiv5br
ht0EDcdmySw4b8dNfcPD0QG5H32dh5BI0+v8gKelV0I24ybDsvDhzv69/YMNDxYprDYLa7yd3WTG
gixXNTwnV3bzoSFCyDJm/Ywrj+V+19Mc1e11eziXZ9zTlnxpHc1LE5Zje6iCQzET1HFBLJG87Qx4
ZoH/QnaOc5ZUhb1AOeNi6z+IJKZ+33s/tfurZNd6jUl2TDJNaockM9vZT9w6uz6lr0EoE2x4gR3+
6BNN0uq+VHhg44XqccfdxAbSZpRk04hm5gxYKkeMOUwDAA6VifBHIm7XX4f0At3hP19wsA68WqQT
7OUNPhkXHlmB2g1sl3j5kXICk1jNKHSNinDhqBd+EpaAqbHT0qWkQRhxNL8MgZUkfndhR29JI7tb
aNhElt1+CRFAy8p91joKlvaPReXml2pWrqdwrm8EX6gbL5Zplq6egSQeybCD0EE5OMvnMLPuMUOq
V2ZxYcmwlgD5XJxl4UXpGDB+TREmtkf793ijtUF1z/b3vXD0jqrmaIY/1m5Qz0OGrD3t2TE6cKzH
k/1H1kRapzjQYW0dqJxK7Lvq6x/LtC7ku2Uep2eEYRM3cYGJg1RIN/QA76hIuglYZEkPsUkbLDfe
VT3RTl8n4UD33xbU7mob5/AwwI1Dr5IQ4G3vkZQKoy2JNMwNxLcBuSwgqLUmIoP7KxRC/HeLHGlA
9S2T15J8vP/RBWECq9ZqIG6xuO8/S8wsl4YgtLYJxZvaLDQZ+rtPE05XpkV0KYk7bXSbud+mMzur
B8ppK4CvKWYcUuKuHHQzAjn8TzFs/gy8s0kZ9BX/EMVbaOGTQDtXRJO+rGNLwkyz1UWhvj+v0Fjt
/maRjmv2rxcr8avTAwnCQkDE5Am5aGIwPy3a1HF+xayV4u+Cxd4MLGi/zR9r6kwgrYmG1xH29vF4
Cf1MjctdOWq501lBbbtw7o11UubGJQ12Vkzij7O5NN/mn3HE5J0nNgLn9zAb1mfks9PFz3fRm6TC
avlf95TGIuh9LDwMdTPPn8Y036ke8asdAo7mNdbknKK21Wv6V9p1l22dCfuX6grjbeQT7mTrVqty
Pb1IjoaYwKki4m8+sNeWWkaitBKCoJcCRqC/XXTTtmMJG6RTcXbbYNPPg71MK9Pyy5eGLcy8ICVM
mIPTlcg6V6kztAKrmG36ntRQfDrkiWzGu0WdxnTfAvdLuPOzKa3zcNKseKMQNK6wBNQ3kr9VOINv
22i8CnNepJuevSwgophVyN6UlU42pJOVpzkqhJ30MigntvIQKHq9g9Rek9xuLW8x2EOIb4EBv48a
JRTwVuNi/ecRA65BXsykymp5FdbiMsK31aJYojcadqwdpD9XvIsng4FkayLmTLntebsrEGrrscva
l94pOYVJSD+yI96HjYdn267EhSmaAS+VjeVu+06O33ITafeW2W3sHBw6rnjC7k2gHSrgBLvwqjfm
rU0HL/l21bXZs3gAy+ibwAii+DSoTsAtC9MmSefjW76+5ie0aQG6ocyIVdG6QU/pvwgB8nN0o7Qe
krFrGlu5Cm957OGxbksGK93iAM8Gss1qddhZMPleYmvCstQTaPSVmGlCKyAAeaXhP8QBiUNNNEps
C+BmtTpNNnsm57qtBTlr5VkXtLtqNGR1CncEqW/5Y7VGPXPetgr3TDkpxcc/FknlvqtNj7OOk1cD
CkKCMpYRkoa4yCD8P+5cZWMJzx/jHJUVUp2kJXpE+bR3F80i+wWBgUGUdZvHgY3Tx8rBgWRe2Pqd
PUSf8Xk395yuhticH3JJfEoiVUg8ENCHx5s8bAHFyRvG95v2Dvej+M3nOpUHamtnaVQgaIIFar91
y4LS8fe1saA8S7J66wWJdp9Y7zRuuvSfmGLIZrtmyYsSXK2PK4vJCh9BXce2QEHJ7TGmK+uyJ9JA
ENOXEPZopK5TNUZgyTzETkQSHMQvyX2r2sZxuK2MIoFMH9xz++TlArCG5SScnFbWxC6fBT/NGjqK
dFbQaRTPl593jCV+NN/WURfWPbe5V2PCV9Kj2aPramQChYWior6m47hPY4mDaZxdmtc5cIyoWrH2
zP3fDAKfIkrHgkIY2rqF//OyODn2WV0oHda4uiULzhykXHJNJu1G1yUNYyM5guZvb6USRaRrtVyQ
f6x2n6OnsOeNB3sWMiolFselgMLWoafwzY+KYlUyVzR9bbFmDlUvWQFrlI2WlDtWCiONCHUKBjmf
cQnIuPQzhkG37JVWpEY07sA2U+scDPyWRNWTgY/pmJNCbnnAO1c5Ksu0xfEWezq4oCFPaKZocv4R
Wg3/1vo92TA/GbGdw9p9gHUm4nIzMftnlw7OHs06MCOukHECPi9rzx/Qp704HmXc+dby3lc6YHDF
gsEUIE3Nx+Ue454GIgt2TSquUbc5XX0EbflJslrigP7erYtejA++uh3PXiPM21apNMkT8CxpNO6I
lBy5EmEGG6ic924TDunXJv0mFv1CfxzP/XbShBB28OmOOtFWfyeDoXoaRUsR2AhkU/C++2WMFsZG
5G22W34r+g8UKvWHsd/7Z/4iepQIEbu81NRYqhIQzgE///lz+Vau5ld/69mdPg6/E962lQ8Qoxtj
PXTl+JK8oneWStLzbkNdc3hL/r/qTexACuQU37snY5j9SxFWfqaX4TyfOEu/dLp+mMkES6qp8Xxw
nV7yd77vOG9zYVAUpIqX2P43duDsWLIbuDcIKirBoKybpyHEa91ogv8Y6zk7uzq2lIU4kPuarc4o
fEgLfRB0Z5JpziaXzzRtqaCZqASOtx4OAo8LXgM6Yf2J/6dpTCI+rRRY+qUFct+zyCXAaknVMJHR
fFVLXEYkB6jga7RaGaHxsufmr6RYSiDDGtf3Si/bfsr233EsC3p6qr8I2MGga8SowwyllvD/7BWU
nvyHKyD8HDtLVjzC9BwdHcb4Ri2D79Gh58Q+RgaWs99JX+1+pGL/O0Ir3jgE9y/k0uQz08A01COW
cop6dVI+Y2N2HOgkEnm6hHjLEP9sYe5AZyBiW/AB0i4/JOo7iRu5Myiasm3VuO3Ood0qSgURCFGJ
v9ZYXt36FLbwmXbIm7ovuBm7toeR1aqlWWGdhTjlxdIajKJp+p9rcIwwMZaOjB1e8a/RPj1snRyu
INxtVcnuAUS0Pxj5LaPsdK74bW50lc0wCOqY5mgIs/dRRRAZF79swoE1AnMtz3VnwyPJ2mEvfM0I
YPWHRMYsue2gctXE1kxHjV5cXt9zXV5XhjULMX0m0eoiqfo0LAVerOowXzyKXD0o+AFme0RVPRYY
9AMQFFG/lwMB6bP5jqtsoRcMiuMmtOH5X441y2lPT3NjkeSAa6N3ZakdHYtDtl2M5vEFgXKMqIjz
gHLFmukBHKIbFnh3JYQcaqpzQgd6uZEef5dcHura0OlnGP2aZaAYj8zHyaH17xLfsIw4ti/PMebr
a2r2F6X75Eh4yT/MCQMj66UP9ulp7CwTYCK2ue9I+tXElFKSanPc4nrvop/Q/SfbB5cqTtU967JU
TWVRVFoHgkLG/ZlGpys0cgIWbQHkpRYEqwz4B8wpZCkmzimBdy+p7+kIRJGIbAo4ffnXaln676Z8
TdfT6hQg0jFDJzjA68rHF1bFV5RX3LRsurZXnRCKAdn8nRsJ3ipPWPPQztVmkKKmBw/M8MvhDHSS
pze0GCbNmfVIqTm1CNDsPu1yFiJTVcHqMpcD/WHAeDh1m9lQvubU+WGB7Od3x392W6j4J1at7ytz
Du+HToeL/Fu0HnbaNHc1hfTDRlEv2kMPAvoqxIMN1Hh4UumaAjt3Q/O2Iwsuik4pQnZ5c+a9INed
VsyEW2EfR+T1ToNiAKa9anZ1HaSgs8mbPPqqx74Lke6aHd1NeUWMCIShPLMb/t3/HimNw9vuX68w
qfC/SBV0HJiXUSmiM97OlU/fryBrbkVaU6C8lH+uStrC7GqSjYHvzFObX52XAcr3y0D86mioVFbo
cAdX6kl6/++45UkmA8aQ12H4+BDcuf9ZhJ3QOzzZd/Mlb08ifktsaQNMJz77JcrYC53+b3g+75Mj
XKKH7f5bUCJP3Yhsm3baO2c06hdyCStR6Ftk/miMQHsLk7QTdE6hnCQSkP4tX/7ioNFVHIKlscsP
4qSmDFJ4FOCnGlVkBmklhU+TegxLA/T1ENdPUR5gLoF99Fl4cp2FJrq/ez3hwehbbdFcSncL441m
UePhxi9K5ECvOVMj/pG5xM3N+VONXY+U7PZz6N/5qxwZ8RYXBnr8sW9OmQ81X0uaUIIIRU2NjLVo
TneR8gnKaJxc3MCFmCxrT2HaTzL64sTYtcSMe/L6m9Pj7QPBGvbvkik9wtojqomDDDvNMwRe0tPY
CXLUDbUHcYJRWDkI3x2JYPuqDld8uDdwVmjcFzcpIWRNjCIrdIf3c4rOT4gKyqjoIZQ/J2BASpiB
NNGuxmT8WEt0n56tM7ldjpT/V9UPbuoofSkM4wugHpNBY7zsf1JsnYcWVTtLUP277H9Y2adjmiI/
NADkPsixcs0nkid5JWlbWnR70BuhJKYtBndV/CIEufy7JCDVUWUyUrW2WWdylAZ7plZNp5/OEeYQ
ADJU4EFmaK7EEMYY8paq09EQW+XX1NdZefPapT3VrXl0GJKyS51p/zN3JG7BMlPi/0jzT//LBS3w
fp9H7OvIvCWeVreGZ3/eQfCcV430L9m2vjvDuJWPRy1Zs+2ouZLpG75LpihwFLrlGmJjL+jSC+Bn
qcJen51m4yBiEuMSRCKBFyBf4oez7YOvmbfdFDILreFZowoPnX432RmoVIABaNJ6FfUBBntJjvcX
WqOiy7QOHeOfaPIOXHYdtAnn8LEvQPXgVpHcBMjIBOMM9qHHyURm/RLClAEsu9RgrpHahwXLuv7l
D6K2IErCCm4wFERkpSVTpT5ZXLahOLNf0NYg85Px+7co6khbt8NLaBBhsrom+e90LldXMp+pHuJ2
iQC4KMKRz1EbYIFd5GgiORRdVm7RpvLtGP/i2UbBbvwzGOZtoght4ei8IV2RI3R2BDe/CZC28NfE
GJTjWH3i/1PFZFDUwQ0vU97ePf5Qv7cbDQeX0+mY+EUIS5HJ3Zjt8h62g3tmUbEuM4xdx6snTPhA
pXLzgZ5Q8HVoDjkR1ezu6DAo9ne28tsiwd/1zL3Kwdc2Ar9iRmAnLQ85Fg76/xragYCqS/fOHhHS
x4+yZ+/R4XrRggsnbfI2Aywdp0s5iPLD6I+k1GBNnqbdhLXDO5L0CqDddswOp1RiOeDqTyMPMHcQ
Y/nyvxkLz34mRl/W+uqD8JJziKL9e2/3PaJRCEo5bN9l3MbBSE6lB+HBi+UPn2VO1vsDXfM7CH8e
+QYyEp4MRlGAGs5GChpP0gEnU7htipPaBHNXxOw1AzYefNHauatPeYooXnt9vfAS15YzhUkyYAnj
KJlpSYvHVDx9UaIqdVVnaY5mfdV8YCqALsSy2n3Q1RmkmIP3WRTWpgH4cVP+SUv0RPpkLTRSjqqU
Ib4SJiihctH7h7sZz6gI/7GHY4wy+dATtYQ636z7u6qJp/mUGpyEGJTYtWyDtPPtSWfuIVzvA8i9
GExJrKjbw9zLUelR54R6OXEyFs7Gm7qfjieXpHkFCaALbNxnpvfAThwSLyyh6up3w+oJ+VB1zvmm
XveMUiaY4ttTgCCwnxRFiaOz4PFkWwAcZjyx2+mPnNBkdnLQjbA5mbU6ITLn/mI+CFtZLHqYqx6n
rhajTmAuenj66RJh4wts5ISdaJ+ngWb8dKk5JcpUDWrNt7TH12wQKjsyE3VidlHbC3Jt0JN1C1GX
nozDdwb/7ZOUv/kV3Od6oyd9Um/FdGKcFBln8/UTj07vCbwxwxO+3GoNwXrNnFdrq/nxl/M0FNNv
c22f1cvaw+YCCm2/WtWBBZOXmWgMN3ytX5swjE4OwympbO6a6wPbJ7YqORiN5KAWgC30ZXhI1K4a
WYDeyKUJlRJxb9027EXrRk/b0qRaDS1A41FXWpCMAuHsnzTJpY3E46MishTZLI8e41yDdsYc3/9l
9ZyjXD6BfbfAV/nswAoY5o11xUEUicToXqB2Ofqu/u8Bfd8vrttZZL4sX0RJuMhX7dch3VMlvVPO
8o5EZgtfFv5HzJVJnln8xtyZ96fwTdBaAU0j97ymHe1HURjELgMYtsmWlVzlFs9eMdfiMl0EatGv
W4Dp/jttpO0JT8G7JMRGDyEtXVCFOP/YH9BYcDBrXN+eQl/aeINgXz/ebeD6QmUuKNypDmU6rrZ2
7vK2OL2r82ZmpsMEEMbz/YUxHFF7HIiaajDB1i1BM9CwbCarnzFUJHojSJeBBuq9vW6s8g1Yq6dO
hYtZ3HTnhVRnssFjoFWbCfXoROqbcM5XKUx/q3ZAAWic32mXHfJ490JbiggVcBSnGKCpVKSr1D7K
rNFcJyEe/GVW9VnpH+3kyk+SSWLF38fiVBpQnvugRfgDIVIj643WIFjK7rN76+WIwphhhYVyH/3z
S6GoawLwtVPWv8BgHff4KpXVOIo+m5G7g+TB01ZEdt+t0vmfDXsyodTOV7zHW6eaG1y6VHgQqQcS
FtT+NyheEfVkykJjbBXgvRwROlE52b4iFe44WZqOPJpbHbMqh7aY/cixydvUQgee3z5KrxuhzHrC
ZW5abqdwinP5E6UJHBXWQGFsTApYPr1tP/UV2ZWBVb2n0UpeOiv+sK7QgALWWdjfMnlStEmsaXau
AKRl50HIuikjqHy1dAy58mzC10+RoAnz6aZ8U2CQGEBIa4IvZPlofW2ZJ8NrAUxr3QgXAMXj9tHN
4Kyvhq1qRZc0ObvbDu8n5wd9CxaxNkuEnLpRHERmk/MJhmfuXpQqTpQ0eM7F1uLtl4KzlS0mZtlM
PlDvtRSkAFa/Y3ZdUZiWKzN70nM46FjKOakMTOTWgpiPyUdtnzHeJiFB8Gj+fj7SNLUTA4dZXdzF
QWaiETJ70amns+OLfe6I+1yzhKWvzW/vi0RaPqz783wUKCJSCpk817fh5YPoPO3RaGdYBZROyMpc
uJnBVOAVa2CtEw8nn6fx0G3waw24sl050TkQic5GyMhD9kMwY/xRkArusB9KQkT0hAnHeTI516Y4
nNCk/FdWPjaRh4f2o4MGXugiKfcDgl8nYpzIC5QfFuJa589TvzR1OyfmAsTODSIdijrA6JMI3VDo
91df3Ae7kq0f7QzBRKWblV23qdTEXwJkaW4lrsgFPrQY7s53gBi8KV1mpTZoJDFOUT4FMuJQyrrs
N+cOyvf2gEDx+lURqdpQSajfKAFm/dGTsJFEkAKhVW/Wk3DC7CrAH/3EyHZlh0+7VLoSipGw8AI+
XMEix8g7t2zk84RcxiJEFqvw6M071GW8FsjcDIFTyMJWsIiqGR+A8H7tLbMQ2UxfFFUkexvu5VEw
dUOxKFcslh77sS6Bw71j9pk5xFjZdfscfMR2I/alMGg24gEh66b39VjgymqLS6OUwVpH7t06fgsw
VJR2p3vcCfpW3Tp/u8L3OTy5OVMNOk7BQuFpxEjYEI5QdtZtTj62P/4EadmGa5JpyuCDgdIIrhrY
P6kwbKDKYbe99aG+tJodat0zsYl1ZUa5dwVhq1zBxGGHeW0U8aDVEVozRCjVB69iuO3DTSX7+BYd
u2zthQb9VtxKLzSQX99tq0D0vXJ1hEjvCJPX/HsQo/ve0aWVqVK23Nso5O+TKjGHBsV3jau0lZzQ
AIc+qCLBKPHn3zoMAGCMpsfzy7C+E+UhmRZq1muumAKR2aCgNCIMJKDSyImi1+8r/8sP8wXg2zRe
98ftVoS9d6Y33wqc+cvK5ZqC6DDLuo5frrf0O2AuoaZrbafAdaw6LmwW5mES0vGQouxra3mx1GRw
0hvC68Gx/UIiqxnCu3EVUPwVTJu31CxNlds68YoAGBRJupeKvS/rU7NrUY927YhCiR0fOzZ6XNNA
XJG6nexRCIIgadOMU46s/K5UGutMKSFHVnKzpALFSV47eLneNJKPi+KmAAeklq2wSzSHdgKmztuS
N6Cgf6PXu3fL+sNxEXpHMM2RQ3bIKsr9kflx9NnTFQ9Cb62XM4IR8L9KS/k1XVXhMYgoAHH4WJaZ
2MOAanNpshIHlfPEBDP50VA12m+23wNiY2jankNedDwQnx1XV4yvQTNFLcQUQlqtG7GntCu9WkLV
WDV3k2zD8JIAe8D8DZ4zxt3UdMHPJlz3BAiAKzA9cjAEkqSE2kvKaplOkeS99VeU/EQ0J+Sc26sS
9kYWRXhdweMvZKXDW6dNvc1Jl5Ora4i/IL/aL27xoEti5a/oEO7db1OADXNHLzmGWLwtCY/GXJv8
KOS5xHFLGx17R8COOGtnbhJSKo/FGENIglB/56N8xO+oEaQFUoirv0MqWIrjbx+vyZYSGNHjw4AK
CtR2qT0gzV94Uqf/W9rZUAROq+1CMQfC8+Xx3hGCsOtHPd2a5b+v4a3qKgvAXlJVtUapioFXkwPq
XyX+jzeqgMIXC9j9MCO+JyT0kBDUi7mliEnbH1gKnA//IVWz+CWRXD+36XYSSpeweVouiYyB3F7B
YqQJcnSDz5VjTqc/NtE7C5TGIDCfMDMkzmqaBXjGGSfuYsn0494Vf3jTlhRkTpRVzkvJIpQq02xi
qUR0MFLcsjPqqzBa1PLSdI3NDmYmsZvU/f8KTk7IHLDbCwxpSc1/PvNJ4yhDSvr5GbJZqm5TNBQq
yP3n9/R7QzUwRN/EeVHG/BTQ8vjS75RKzqrrhBxRJbsVOXtiXZL/XjG8HA0YBfoHzNJWXAJwV/P5
kZz/U7nWe5UkC7dsZGMrEfQqlL2N40q8omzy+f1xPxdehFHiy9VS74+tmpzyZbdQ2lZxRjfkS7BZ
uZUBgS2pNCRMVofSy2kzTmDh6EGhJov5sgwUeLYJ0C/EMn9MgnwK3JJXxYdvO/tZlTUhUOtShC49
LFpMxYzucI9QxLLHnaKg0vxs+C8sbwgWGL7cuEhHKfF57JSc5DE0CG+fGSE+M7IYCXqsQLYIqkkm
eH7EKQvT1qbxPg2XSf8Pqzq7qt50/Q4s/rish0PqCyUSGc0/u+IaRSWn8o6FX2+8MuJWVxFCdHS9
ofbaLMqWqf5ltHixYmNaBfsnwtO0L0inKeWIKmbKZrar25EnQ/nan1UdMpL8iHIrh5YbP0ddXtp4
jGEai1XUjk0FLinqiqG8QCCZZUTo0YDUEJ9BFg7HbnJH6jmQIS886qKogyFxJQ31i5fGWlzuaWQx
IB3cNwmjUIdAcnW07ckJA/m6UchNg1NYaGNSVmAw4pxwxz5s4WjHD2HM+wXZcYxcWBsVzsAfoBki
3peUkBnWRawMps/rMsgI9P1fvQCid4Fd/r8hlOy1pTIfeOlBbios6egGvHy/kuvkv86fyIRGmY5J
Chzc3rgsZD0w6ThnOLrEEyZ7X1Bh51i4LbJmONuGugmK+MvndKcy63ma7Bg0g/IaI07vr9k8+E+W
op/l0Zg/DE2vEdJX+vElrU36ZBThZtfEiFVAR50eLZLDFntLjzNp/8UJ2LaOVQB1mKxNZPJOdq+Y
ujacb4VSFpPGrUIohv/RwyY7iEqFh1qbREMeusDP9w09oOFsfxyv3KF77nglM/iqhK2n22zZcZH1
8itCEPUAJJO9LVUMgMBBw9zyuC3fnIolVR2WrTFdvLKy6crT0+RoRvCMeokl+KNscMwt9+Qihjr6
vjsXKpLDU6YGYgHhVqf7+luEOCrDlU21DWFpRTqG+54OvP1tN8T/jzZTTeVY9GOKB4Se7adjNkhm
6GyrQuLqMHRXtunsFhrdmL6ZCTs11MjKcYOQR01NEsK1VoiDLnc7wAPenvXHj5WtZ8ceQUjcbwu/
+m4kUuykXVbag982Czc/AOKp2hpkmTuMD6ds7tIelq8FQgpo63cAeuC7oiloVMYheU2fva0s9Nsn
9SNxv1E/laQboLsqjzDWh7t6jwi46ie0gcvHPZWpDjYbq3XS/BS0IJM25btZ8z45coPMtC3oiB6I
G6r6ufPNxavMx26cKj/2ISNBAMgZK7hz03aqi8WncJAmnoMQV/OCMEf3IgG4PY+kpJEiFqzecXyj
AJn4/Ni3JXSACsp38hyX/+Oio5Za2M6vg1McuCcT1+6WIqnnfAbEZHCk3gk9mDziWYxxPcnSi8SD
t4TU4X6ohrYEoobC6+xH6ZM+AneGnhsr+B90/ndUTGgddKeIYX6TSuDaOch8ycOKmTyoRrbyjuw5
8fhHdyd/eg2bNV2Nb+wesypZaPE0hOc9JMg9OjraH4jNyfkTfLF4R/RgFY/AQ/uyaOCPPtDoN+TF
mEbUNsTFU6oo7SfmoSQgMIY3OTrkFgvlXLq1UJD40u12U084FuXNoeqVonGtllvsbTIDzGMXPkOh
KzJgIpnbWc+GVZe/wI1ncEAWPShLxZ9JkF2J9JcSs0fyH4YwSXuzWmK7TXUASQkA7fL/CA8gTS7x
Cum18OObhIJo3sAQHVt8SBtmt0ixcdyICzL42MZG717RbJ6MQxecDqeDgvCZ/llGQ4A8LAKhUKq+
WGReZ6MisYzWyZAgxJBhm/fA4W+jChmGj4OjdkBhe8fi305+DzlQha+UCVr9Q2IVEWUurjQJHrkY
yzAUsoCdX73HOMYsF8yjKWeA9w0LfaWCr6ffTTL9pVxu9RhQYrshhpuvaQWX2KXR9GuUnHkUKk+v
X2362pA0tf4j2RFyp2XElFGyHmRuQvVNTnZfC0pqaRVGyXzeFU5KXGrpKcbuTp2kgORCiYyRIXHe
er1mwoY5cm6knLpApBTbhip2iifs8dKFt09p5RfxuH12N3KGyvNOPi250NJdN8nMRf83P+uvxgEz
bWW2K+fdAlNBtIJ7Mui17u8yqVNbguIziX/WKrNlgh1LZOW+vaSSi3ihC+okdxCUGp3OCt8brEkD
Tzoy6uSdDqmmuUJ7OJyRya7XrOEJ7fUrU63bXSeMmmxUkEnRcGUk0HbpTG6kLda8mloC0iG6K0VD
vKLQEejqfrzU6mR52Srh/7j2cem8kuFKhnuXo4exxCjoCC2JYnshEgOclNPPHB5dt0E4I3+basjK
J1ga/7/zcNavVpwB9MYA8S7QzhiBkMKd2+lebbug/++PYO4FXoIM/xeJd2MAlq9nN4tqXs3STwlz
469DCRN7PSddGbh9Puwv3eF+c0IpHKOOna0a5CdkYJ/5Pt6CpA3ROaHOtA0IEkF5wA5zqip+EPAn
jlPq9bBWYFimvcTrhLf5LE5D+i3ANvccK1kR4toNggqPeAgpeC9EByv5MfxfBSjwJBpWVfZ1gwDy
q2eqA1atTguoWaEl/O8L1/iVKHNSrL/NyFjfJZp6stdBtyB8HQy4KDna7uPFpt2pQbknuGvleW3D
9e9lAaPzLKhaQJlXSCc+LFz+NP+6LUhMkC9jgALsXXKjU2trtlru9C4COO7iSPbAb6EQKSC9+nDU
PX2JXz2a8aGc7lXfqV82gx0V7AIBYVb7WsLjJq2Nwot5UbwQPnAtF/7MmBoRULlSeIroXvTRIH/q
7lYtkZ7ldk3pgxbPRetaZivkl5oMS1azfOnwCtF4c7bFXR1mGJB4B49faFB1ioQ3X2U5P0sPoC0K
zYy1aAuFVb1YXXAcHxJ8rw6a3ep6NB0s/DodlcCihQn5Uh3tPS2sIYv+wwtImdyXx/lWRFfgqCY2
FejICtbARfBzojHDYzBrXVptU6E1SByDk1tUGoz+OTsZQWiLQZXbtByelq2VmZ6PtoEdVTD0CzvP
KBS3iqQeLJsUr/Rx2koS+7XnjdOUDPo3JCNM/JI8h1eDYaDHC00PiWHc39lA4XJMqNuOoKogZZqY
dvHxafw8c6DsHWYjl2AVEZAabPALe8mVadCsMtmhOCejjlZ+HuwYpRyczp9du1/zouwVqTBM1QrX
kKJgDnjVX4oY4aYi1iDld1pt4RGzOSnD5pbO/lBYA+/Bi0ZbEmv0PeNem1KL2AxxuO+Y35gHnuGC
kwq52TmQv/iAyQ8Ai9dvkUYrkqlEa5xqyqGc66U3U2xwhZLXfOwLE6XzKv2J5jsLTBvkwdPPfVMx
Nlx1PpSSf/rLMjoL5JnYUfsgBC9S9Nt13DPN32aX2M1RDJvCIlKT4aGSPdgsyV4U8Lmth+JWQLT4
lBcjE//nIDxJDFs8FKRriJnP4l+/kix2FQ9FVMoaF7CUmB+NFoZuTGZu19/s0U9jeAGtRnHlgFTi
WQ5BtTtlF2o3Fpd/db0D7LNwyUvmxSJPgl4bCC97ApJM6wjOBgoHNJXby4H327MvcRugS10JJqqx
u4j+ALICLB7avala0nPPPeGfvbgrHr3Dqm9XQjt45rfQ1cqQX7luV065OpEpbcO+5+iON0QIqEWi
DF9QvJ6epEek7nqu2aV1mRmiB6mpWNx/facUUIb9Iw2oeyIECiDHxeQ9w6I0/JCrdWXDOUTtuxEs
MMQ5zcWk46g7RVwkMvzvs3Cwjf5HdBhdtQN0+AT08cCAodPph4ZYgmuTNezm+jA0xSbUr3cIw/eH
te17tuzwodEXz880nhC7+R/nv2qss1vB9M8hqdWvQ7BpzijFT93IGOQcyIisxKXD+eYu9X3EkLbQ
bUFHGKPNIziXjl48cySGA8mhipVXs6T0RfDRp6mHZAeo/bWsIyILwx20kIhKFYjrd/89ktrIUimW
nmAt1Jh70nQ947uw1tRwAIIaN7oiZpcALwoVBFEL+agXDaKzHuly9WmZjMVSVaSoLU0qG6nAXG4R
Rd0oRhMJghpJpxrgQMOnwcTWaPCcpeaTpEQEdAB/PSTzWTYgldRydoQxlJCHL9EV4ngXSNkLr2N0
CbrSrFFRlcvqgNZxRjq2VR7FVur8F2ufUP/M8IstPOjweW1JMsUk0bdO/kdstFMBJsYUvTHo/kDi
gaePbN8fGoTnw7u/faIw2rQ3XTVsNdINO6OTfmjinir+OsfGcme8QANIcPndoXkWQ9tkbfrwYypw
z9wPN+sL1w/Ygg4129drMtW6n/fQGAEFQ+bmNQJlWmgzWhoZoXGneBUnPMwLCxu4g0FZt0YwYpsr
pa9NvmtqHC6qiZMqvJ0TZMqvP1YBogHE6iKno9bnLmL174M4pRM8TWzphtZzNpBk2GqOhjX9XROt
xFMVyUu7Cex9eAsp/JY6CPqIv4hRt2VdKpDl6OfY1tzamyBJiu4ewH53Nm4+I3TM9h3T87QGD1+h
1004NyF2UlHyZt70G7e7evwhh+vHeKOUfGhdj2ReEyPvstBNI87uedvsSCitMrL1vTwpg0dXIxaK
UnPPhTpEzQ6Xs99lxwlJouozVzYxDn5OetII/TZcFB/zhhELZ2Hf3KuO4QoW87I27+H00hb5z6cc
KUXgQ12GqP0LEcpCnvRvXmENhwre5jVLT1aX1jrrUaqoyUF487Z+puIjTKtqkTGTuxJNdJMVThik
88EM2r26Ng8fr+c4O076XayYmy4tdUF+2ArC+WB4Yw1NV9liTDHW+sAZWI3GgZC17qGnSahwf/A1
a97pgHfPFoJJCAY+hqfeyn5N/8992/+jlyyLwhe4KSm7dsO0l2O5OSKTuwmFeH+/4SxhneabDLwQ
dEMm8FybTnrJ3gpAyWPaZSe59FybtQbARJTY+z4gY+Gkl3bQssaBw+PtzHxd0tk2+ZlnggSkXdwv
gzsSKweeqep0dmN4r3ZNy5tzEsJowxw1CFdEfQkZZecx8bkvzoivvCD+Q7hh8zn+ABDsvyujveu8
wt1WROIIzl0P+dnDva9+WtEFLuJfaUdaeTTXB21p91F7yfjLPT/OSJ6Pnf9u5dOWScFSgUfcWUzz
HD1OTZCZZJevShyTMXTK8y4kj/dgIeaR8aDTWy6KThXhyC64f2c6DHaeZ8l+ZHK+I19+47Bnxrpf
ZVB703MTeK07lTRwmdEqNIny4E+D5XgUVL5HWJkwJf2/RmJX76asR2Lu/tokYBPDbcXZYypgGlNh
sx9O1IpbeC8dpG7q/ZTPwzda+EeQO4lD6iZBegElw0alZQ1zDejbffrth+hDh6+KgDqkRwN9Q7mR
yHh8C5GWCpbB56QXYhsZURQKcSuOWNviVu6nyBZ1KMm0oRhHRqDbkU2xA1OD0mrDTersIz6GCXlY
RmdIJvZZ4VMmuHHAAulCTfoxZQQOZWgqAiTnLCUWi2v4DHwtVOFbJiNFCP4BDzwjE61T1noZe36A
g7b45jJZEsHPmfBTSBAyyV/PfNuFdwhxOevtDOBKHBYl/3SbEqrkai/xAtjDFg4b99cEdmPDjt7T
MpnnBBl+gts89tZ2O2KTuRtGnfXtfZE3Q+H7Jl1uUfN8GaLmvX1vvB6fUMFCMkpOHIzRwqFCsHuK
23qncfVPPO2CdmYD0fieo+LO3FXEbiGpU3PNZW88bct/boWiywJ89Em1ocSlucyn5++s78Oq20h8
LitNAxpq2sLeiiXwAyzai9tKsoHi03nkMl2YEViTjLaNh8EBxCPkNYw8tBhOPHDIoUNpmiP964xh
MwZz3TMb/eifrwCh86GpmOYDaYjWWTGVsvT3YCBAiGPAw6CvrXmm05rewiKhWAMR8xrX62VxIF0a
/BHGXheULo4Yf+Xt3jVdVM06R7IpBNpJu4yOtGHC3JD6R/U/Ygr0Egapr2RDLY3IOCJATOLof9DW
QoEBvQoHpH4vdkbWeiV6bQ4RwRelp1Pe8F5kc5fUEEQOZdDaptpoCa5S8P2pUHPTGcjlK3AaZGT+
OjxZI8yLezq/VSBIUdOnCN71KOOLmMCaF4viRwMDroiFGEgDP8bfEv/tgd8obnYYzOYBBqm689lL
fQyF1N2lCTA7+L8q6c/iB3SbqNzqAmwdDwa1g8TQrbz8fGJ76N15ZmlYZmVACy2dd1h0+dijyMMA
m7Lvc8uuCcbzn52xZE9zTg49ugrB5UFMSOdyoU12bsTOj12B2yC9FFWADn2SPIgKix5US7enyI/9
TvsOMH7UahT5rT6aU0VrrTs9XxyrVN8TK1omHkw6lgPPRgpDn/epyY46Urpl3CXfENW4g29D+G0r
p7QWylp1jOF/jlLRb8mAYnaKpPG6cL06BVio3e2yz0WWcgb62iNdDwxos/EvkqwcbWBdeTh7Gz5H
ozIrOf2iG7va9J2FkOsVcdnYCKEL3gNW0yG/HvzBnvqJpjTHjIE4ejYX8M3UkX/5kPxm3ivvFO7N
WupuHX25CYeHsitGZLfgL9/9bYtlhXCRrbMDM9Jo0rP8MFfJNmsbhijJpZWNaMSs4wJRt6AuaNrR
bQFC4Ty+MTr/kp53/pfUv2BuLfb5sWA2Wr7Peo2/mn6bLYhIETFZx0mkwLSVdvn20bT9/PpuD3Rd
GSUPonMBxqbM6nWuSDnomBZC8c5iJkBjBa9xLKu0dZd9LlK+YSlXnx3/nxpOmuPrQgwxkBwIMywo
ym6lkal4FYVTTjM2TgF+8GrK8HFNe37m2AmxeFzrGfGxePEOLpA2Kqz/wuWOaFBnb6IBG6SICdX2
Dld2PfKKlD8hk8Bws0FmqE2Y8kdS+vTxereE+7q1pT2sNNx5tk1IN5ChK0LNjWZN/B0LdYwElWGF
dIX7MzRrKLKXCWRGC9AUdsucVYTmZiUG0/rt1EvLOXiO04gBnw/Cni09GK3lKsCPrDKaN9Jd5yt0
EDDzBw4Hwb+gCSd9uJDiTxtsPkjYaMR8+6DBnEs3VtXhGJ6w4yVcavPvaQthGiAXfaE5I+RwgrfZ
pxw6Rf07uS8xq1WRCGBhKxuZZRI7fBgn7lrIfy858tn9+6NNN6UE6MKu7KDhilqtkg2nzybJs5LS
B0sDVLtGfzNbbjovuT8tR6NLsap2pFmE6mXG3o10HGHm2HIjq687aG71rlkqqi0Gjq11s10CJVbr
8AGVxqTeELnPRI6/Q+U4z0ls4h1ZrGPjHjZ+vbWg67Fdh7A8E6JEMfhYAghgb6kz1izFyqc5W0GP
81ZWqY/J3PdT4f6Y5RrivPeXtet5y1ltvKf/BLoQF/c4B0Jeoc8cMckIgoZ6uCWNc26G4PxIbekU
bl+qwakZNCkdJs/OYYPOkxj43TezGyzQGLnmW+HTYMgjcnqs6ol3Dbd0pkHNFUboH7fUG0bE8/2P
b0rXeXiBpdDLmu2FwPe4nVg03/OOM7AzB/LKh7YAybMaxzLAc0Em2zG9+QFru5WMovMqAyOBU7ne
wm8iBtJnbIBtnCrNwMhGrjv6x2Xo4y7yyAHwaV+Pyitwf1T71+MfCE7QoaBOiIJtdrVrsLAzNTgC
9WFwydv5Y/j+NOYAn4NgwhmiewUQp8KuseJ1VQ6anfk+2UR46hJrtY3Vc5eGbhupo19kPCwUsKYa
SY8hGAKZkdKh994NcjsON1+hL+Ij6VsONvgGE2O4iJ7n/Z98xL21xZQG5OwipkDs/arEbwoj/kPw
Pywe9KO8GeseKC2/GVnbExy1yU0ZRxURqQOb3AG4B7sTx4MlVUKgA++MQhVSXXVIMSXis97VIA+p
MnHxGqSCkzqhiCAPy/e5Kf87c9ihqhNdcHEGW4zvgiWfEXuA8GQpGctyMbE4VlMU3vz63fMtb5oX
9nC8etrTtZOxzOXdG5gTl3XsWPx/ic/1Vx7SGJOdvUoG1UGb1Hh90dCEsi2DZEJw02CHHhrd+mTy
LlNv6M11TL2HQFTGQVcbtUQauEjVW5DwiGTOPBd3sB/fr2eB+ZXqKgkHrDFG+5fjMMkqx2RsIJKO
TrOPxg1f+SzoAiCXFQuoT3DB9FQ1omtIEDufAd6FSudGdrwP9pGp5o1HZApcwxmvgID9HmlHtokS
efVyy/doWHAR6RyIJvLuqgPgOpzu/7qHRxJ7f4N1XmPVyxxz2mxs2GaeL710kKZBTHKzh3JaUbSy
aRLsQ1eeOQ5PkB2D/VnDQueSKFkss/8AD7ol372tNCNrfDx4vg+eCVci//STvlXCwVNaWmUS/5dB
H3G4+olUcKIRoDsBnMUfgi9DENPVZkpX+jY7pdQT6LYHyevf+iwqhQGqzgPM4UdzF70nTRZxk5Jv
dU4/EBQPdH6+jiKqhmbm4/FnvY5vXuTN7P+mGQFgIkyyRS1bIlsBU4B4K+wG6zaow+y7T5PJFk/f
GdObylR1TtapMdTyHM+ADF4qmcds0Cl+avS0Dk+RDPkl1zulhtQhWWAVJBFHKCAaMMBe3Dr9gy0F
FZSTpWG4fTMWT8QDRN1eOosEeG9mQYjEW8FYPzAzTI+EeY6Iqaw17VaVfKoxGLz4h9qiSPsAdkVZ
mGSEX+Ow4UTT52lPwArPNbjSTsT4fUg3YWnTFvPTCjlk0wUGcmSFc3y2y14QVOwMLPBD1Sd9A4DP
aDCBzta7NU19hqR9XilLp/3fymbZ1DebYZ88e2ANcCowX/zK99KL7ESogtHC9naAufN9zfTmO650
VGoAs+Clfl4QP7+SncfN4XgRloKKRz8fvpamRrM5Je7gYccHIJPcQqP4etrwWO6RGkxtU57YPIBM
Tm88+H6glHdE/hzF3vbYQTA3kYWZ6ebt0bx6jEwowFK5oxLsdrpBxVYPnkOvVztYK3nHdKGbtz61
laqw9IvIYDxtuv/vDJ44gfF0Fyi2lfMfOT65RY5PZh5Ei3/a3BAyrdZJHgRBhIGkel9uIOm6duUy
+2Y5+n9XoLPdNzv805RFU3YRA22g7G5z16Cz1q4V5evDFjFUlEUOv/3VLXY6mvxVb6M3s2mNQyWM
ly4+tB2QbIF6pRpxgWzfsfFgkOVhUe7BYagqCwYs1KJnNMzU6r9Jz4TUuX0WG4/rJh8tF0G/jqXD
ufk79+RaMsH2musbZWBQ77dbIH/mzz/v3wty6QhWki2cFFXbCIyTT73RZ4Es8MBHik7dKhXRM7pF
QG1ZgPPWv4Ne4CskEg3l3PmMbmbDOW0yTj41TOtQcEuRG81+bl0zzVjr7HxXSV0IiRtqld96ucnn
G/FE98OVq9c8r/olArGK8+KsgrEm6InyN1A8eO7z+OF6M4xNSPCN4v9/EUkALQLGVJUo07UxULaR
nN5ncDNjPvBZNRS2KiJtQLJgz/CHZkIYj9cBrZqkw0EidzEtVXqZT0oJE8ZM6nYQYIdqJ4GPqU6U
qJb3M9FcXeRY37wh5fAx4Y+X8k/DZZFSZeN9f5ytqrLQqDwB5n3xmkvp+fu8AYsKlf9XnWHi3ABI
cU1Ru1gAd3vBsN3imE7LyQ0WS0PrHnkRg7DnPo6dvHY5chjroApxFCCELUjQsC0XhhDrTUvsClwU
N29APLqRZMpb14VN3fgrzHvHGOqy/UyEv7J1nr5RdwrPBARiAbc8aD7Ju3fSa4wEWUXZHUu88gRI
v95mwnH4cJmlDYidO847cf3ONUpR9ZYoRSMVXHcLOc7Cdg35xvcEi6tGipkh+1y6UZnHt9FOQc7W
ku+dzWZpJNWUQXGkNpiwhIMLgoDlNgOkzZDcokhyj5SZ3jv9a0aP5UjOQWJdJgpdJ+n72E29i9/W
pvhNNvvixQwadbgEXjRCQulH8wQXyTdSFugZaBfOBrOlb9/Y5ZtfYRYKnrGw2SNui3tQ8oAfq4C1
5wgNnrCVqZBjixDNGh20/Lz4Ls/+uTBLHHUqO+fMBI/N/RfLzyVgmslnDrOSf+Ur9K7CrYAWcL87
vq+Z9FVQLM7TDEq79QEwhvsuV/xu3yyq2k2eN++DhQ2/Wyy621B9M4vn8WC+OJWH7jkeqR3oQXD+
RJ3foBOuuIzOeg1MIF3Rhd409x/bEu8FHgGXLuP1tY8nYU1Fkc5hTarmqthq2O49RJvtGd2JsEDU
DTpzkScWo2lWJvXVfAYTGzIdsDcNg6J5eFLHhBrysMOIhwZbHknikXwyZOR7V1ne7eBjLvpmEja5
8sjnm9UXmJUrlDKpyThiE/7XmllViuL8f/E1zLETjTDsKqZIogAl1dmSkv8hJqZ9uxbs7zzgaYfI
xWD/wACUor3Fkb9Ct0Pa8KIuVdkdJDqDCcHY+wHJxe9gbZRdTRIxgA+9Kmc1JyoVoYTPG7xk2rdG
9MgKlhdRdQU6hBWiJjNO/hzqfy9xJ8xGsXuIRzB1Uf6BTMh/Ij/aIKf7nAe1e6g6xTzKEl3zW/YU
yVlOUbpr6+GeINdNnv5ioTKQPT39btkatgI4vK2+AvWFnuCMfOnCheO1uWb8fcHKoYeiKKzhxQ/t
jEbAmc/7k75iucx54wzBQzSau7XYBubBSpoQZM06p4AOtquks7I5U8aAkCkvoUuS79cLxRFlItgJ
KxlzT2TtKqMwMYxeIGPo4Hv51JpyXvDmWCnem3FBtvNRxLx1KlFcBkpw4CEOR15lNg9ONZLsh9bF
jaqx7vFUL3lYVOobyMEo7KcpRqwa5JWSKR9bVeeCrvA0/oq88WXGLvpXJWIzgVdOqN/O0cgHp4eA
dbTgIWL5P4Co7qFf+DCkXo1hv059ffqnFHGlYgH6Uw/xRZL3J6GDN3pRblhUb/r3tDxiu2bzw6B3
KYJJwhZ/xvd2T3RZTo3LAOxomdNpbEkIJzki8/8DgBNbuMq1qwWPZcaB+NLQKdQaedMMXRKfvtmj
VcuXrY7fTkK9eqpU7bXGyD/loscg+tAlHObzAQO0jz4fYl1EOjZaUXQLvoPMXF8AoVwoo0LU1qbg
idg3JN5Aqd1VV/i7R93WnTIJlda+lmDOC8j+vxCDwO87ij7nZnFCHSVJbK+Qx+/8ddahu3iLXwVA
2DfurzSBHBGFHYbwjzAwXxhAEnFqaH4E4tnOVttcqTjxLhA6Iwcaas2fTIoZAtvZtNPgZ4XK4nnk
i8JbadJnc26gVKbHBZZnIZxaFtFXPLjeUP0ZOGFVyFIhofmET6ifuwD7dBqeoPO3mM2QpWX1lXnk
B8Xwb35kfwPS+DiTJ5siW1nb2WP/dtEQuRXQ2B4MVvPSp9PWhr8vMr7b9YxwHTRyIhgjnZ54Secz
HHbSUpsf+GIbcRY/iMsSjcRa4CLgmMNBTVpyyFAdi4cuwemN08nxxxB4E+xEB1Ye9/463P/m0G9c
oJTXgKcgcBc1F51sJHk0SJmHey5f/8TIUb8FewYsRYYxelMMMrh0BDWl5FHB4ICNpXAomvKGoZ+5
4XfcDWAwpMynFiqszcMHh0MRi3kKtxLvq9Ctr9b+I+KQBeIFuicc5FLeIMCMLwl7wcIQ3Cbnlk+7
xRjwRKmyCl1bLwITRgPmQEh83CPepnlZ1eGNJDNPFWZuui1wR2YOR0cCIvKs0mXiy6wQ8ptOBMoq
8gW6vlHjqHsvmMODYy5PyqDRDUo7aY8vvXLYOp56Av+yV/+o3YsAK7lH4QUFhwCLhQBcP81zZ+Rn
+loOIUYWsiyPdWpNi2kqG1UdYVk0vslX/cXOUOv8Y8dznyHeABCrbJhvlOcqB8eKTWHmMl8LeU8C
JWy9Zuj7rRXXbuFs+uHAiRyX1OGQE7qZzHY3YT0w6P2yZ26MFoUP34nKJ3o+cwTEX7gNNzzQvrNp
t+6iLFJUvoMzW35mnd5swndHp51tNqcWl4r7ZqYiHrL9x7kNxgtk5RvEhti8YF5QQ30oG3om5+Dk
J+eEulO6ZaM9mV8YCE1qzJN0DsbMnzfixdbvDeiGOy56Se5b3JbG1lWtfxg0Uf0HzRWQUG+HURfh
t9B5P29AMWmzTD+CoCXc5KT1umP53OqvWpQzeRHnkc3Af8kDxBCejFCjzlNTo24lZ9bRcXbgLxvU
OcKSLacIoDPnyISLRdZd9mb/YS3aRuABbXtQMCl9RgL3NUeKQdYQ01SZ+u40KeR8Jw21qzq1ABjN
Idj1jbvuvWzmHY0InM4clCBakmaAIRd1L+c4hgxyV8QQeB3Awh2/zto2Er1OapOZP6gMaJQwT/7+
iYf3bbzSyC4a2PnUzTC37oPoOe3bsxn+QJtXCGh6DqX/uz+2q9GYyuxw+vfXbgxrOv4TTwyuGuj6
7wN/A+63XipZX/lgnd3gqa1jYhAST7xQ0UWyAXQb3Y6k9xoQzZsMWvLZc3AUqcAyZEBlEsb00WWP
6vP9f+TGtBwB7LNEorkaVXgejpzTW2fGU06QguyEqJuEwMZ7A8vHZpQPrjAd72FkuJZTu5TWUb6y
7WgseMARdcIhVRaoK6voY0SNoRRFqAqHXbwoDQcR6/toWr5MK9uTyNhcpXi3wrFDcqT5r0ALanC+
556wfz0SWxvctygnzaZVGR4JojINUCCgpPkz/SUoz3u3mOKVQDtG8E31aA46VvSR16gh9tJkauYv
eUDlbZ6TStTiYvLMFULIEBSlZKN786s6sS/GiJo4BM2FHh9hzhMhRP9+i0NqdNEvs7JWfB6tKZFq
4uLKTXPyOZ7L+9X75IefrsNLXDmXwEXdOfTPrjVxlyvfIU/rH1pJzlSxCUtN88/w5/GLlFSS0rcO
GAM7FJbFRIeFKaVOWX72jlPfepHy8YzAuOk+G6T3kfGH49byiphnd+ZMnGRiS6cdkFyY5Pfin7YB
dFwmC839AmOr0TXR5y7fCm5hx0qUZwDA9NOxxgjUkn1/DY472yt6al463BWWcxKbXKjM8jOa0GAX
zr1MGaUGeq8wl5OuiZyCFyy8o/iPowt7y5jMrVihl2Bn/vnIs+N76NrMZ/e/Lmuso4Tf1kDMN99/
0G+qQd0A+K21o9fyJQrsNODZe7bNsFkwuVE1Ie02gqvmj2upVT4kMML/FgL2N1AxxOQ6/jgdi198
A6tpFZLpWqaijsRHisuWI6k+CLM8cM4/T+juh1n0EEEvcrvKhBTospTMnqF/WlB5uAJK3EdglB7q
6nZeZI2YU9mFf0x3q5e7nPIrmg3T9wKvG4A7aqrdOypt9Eni+AjclHTOcu6dd6TwuiZ76roSh3fQ
Rivdb8XocFLwoKWXM/dafhMP1ImahNeXk8m8vHA41f2WV95lEPP6PPfehwE4O66lVtbtWKQ679it
brIsmJehagylWfEz8uW/58gfxIvZJCrqaqCVONL2bMyJaU3/EnRe2kUjJrDlWRrcfKh8UFPm34sM
uqyCmlZcKccEoWOqsIPIv1KF+PqU+CS7uwJOJpuqAk1QjRk8ZT8PKW2FXJl5m1ERmiCEOADTJwlC
yd0ap0AXxfzN+EgiEkuXdaeCZTRkuFEyYN+geZ3Hb/lzPDw1OZGyJNNgQEZsblAiEJDJAk5pvnMP
fTzQXsBOTpqI5eZNuGhJCcSyAPMsmZByU2RyYXkOTqSx4fFMGbqISxjyXMlj5M/Zpfm2gUgwnLO4
WpC3Xf26k/7yd9RMM6fP7iPPO3LvmrWwWPS61Ts1vkHSvwk4eORLByUF2J1XVjP8qHcEAfPGo+AV
tOnYsmMoWT5+ZhmqP02qtUIspYGXhgSXTr3hDlU008+rqmyVilUig/Cx/fEqrDLb+eFkZeTnOzgu
vflmDUcDxu9IWRinXKVfkLKBYerdCCPusUv6XueyqQxYZkN410IOU6oaVOkLyIKK/ylfx2e+ErBD
ETfo6rtyhgRbUI2s7aHDjdz1XjK4/UG78xXOetfYzcPzI08AWjCzZw1ZZG7jyYq2LpWUVCQmXs6L
wlWgr3Ef+ldfNC5TnSqoyZHtgNgV9rF9+HTYT45RGJk5kHgYZgox/0luqCvXJg8AgNwJWqQVFlMu
CfbTiuvgNVePhtOkVmk4HRt1W0KY/SD3XW+61XcXW4TA64rtjGQMhRL2v9yZHQsOQ7PW2LzLKXXF
Y9f26MGGmz8rDHj1SEJSXHGhHiJWg9O7tTuYmnejMcD42+RRLv4d6KaH+WEM08PwCN7fcOaY2uLd
1PaRPI+WgTRY/NOK0gIrJKehET9aJJt/gF3ARHpM9vw0z+CMtx+CFOGu1a9p7Zi7h9dTaqj3oo2V
LZ5a44uy3YxXtf22SsMktglkkSDsSTHGIto/XWSg/fttxBw361ojQ2cBaTzsLRqoiXP/MHbh8Ovq
L6bFQgjjFxKxdQISL7texa7hHjdArv4+StT8Y6fyl46IUMv7rQcK+HrsbjPENcl8Th47f2E1KdOe
3I+S90IK/n+4AQ+5T8I5Nvz4y2NDvP7I9YxQuTAJwhyhfSHEb7nQDqqjH5Jp5JfrACPfpfANT7/f
LqQJbC/rsI5TjnCsOk4Vy67Nytfqb7uaTICF/tywYHfE6E0vDA6aTaTvWd1GtZ5/zLQTUq4gu4tW
h7DLC/ojcIJFScX8A9xKYOJjaDTR3J+GY+YCtnlRFuWT/pkemjRl6sV7qxI069k/mwOFy2IAvauE
v5Sv/dn4gTljba3sJ53rMJS7Xjy2jVfeUQu9OQ3qitPftu4Pz4CmNuDyv4GU/a/nV1909c6CGraK
Ogy+L/NxUMfUZqDtyz84iqyJewARWmsGT8taGJ7ZPl+OuL/NibQKLTDUE/0iv5UKFgb1BDuZDhDV
ksextoleOQDcNKYr5Xb1Sx7Uxe+4ZyrB4utq/whWdDNrGv/AlUNyaAQ2lQEstJB4UcxBN/yZAO45
+wL5cILvR3ddo/zcCZhFfBzRZ50jkCO30LLI8upvuxYv81qAl5Z5eFX+mgS309igQ5hD2nQ3rQvR
i0c3KjYiEZ9XfdFPqEA4O2xsNr4Gdb5biQFRCj6UP/dt7eW6ZsO47OnoKooCWiM/z0UxVijk3YkN
Nw1KHvCQwpW7Cxd3+POwKpnd2/wDTx5OL8RDQY/i959ev3edLLf+S0KzrhFu9SGmbdOOqfFF0Wy4
SPU/cOFVpfPKU2NeZlaxPFioLA8ezyVxbJox2e9OL79sVdmMZvFauGOdD5uHTfh/dfzBhw7m/vCV
WWBzbqI944Gj0fnZEZhQ3cNzzExRCfb6fITnaI+6IdFQG5EiWSLEqkEB2b5tbrmcbsKF9WLIPQEo
vtxwJCKuL/58wE4P0v9W2SUjbBWDTHoMD8dOrW9P9j678C2AnVn+4Fv4573EXPV3+G5z3MwxKc0k
fTY6zZv43Oh8c+EBD/vnQR2MYqdP5aoxQJYmtUJdKMNCqor7x2e02mo7vcet7F8v5hEDHWGWqVAP
bBMKqw1Im3jjURDVZ+ArO6mNcrokdb5Q3SgSXcpLxmNkVqYaztWgM7YwdF093c74uQ3/IXLsK4KK
Cj2itcERmvNBUXuukn318L9qBes8PrO230+F/EOmH4iDQ2kR/5Tb35ZJNUw0M8UUFydlRvs+XThA
3apeTsoVb4JfE4IFF6uXwsx5j9TNMcmZ0Eg7eH3TsMwwxVuyXKcPsJgmHZ930WpO9tQ4UcJSncDS
jiq7H4UoanlMzTqbFBHdRUURFI15fye6lbgNcekuewhYa1uutOwYA7sbZmYfagYtycfeR8zeCVBW
tTEfM2lkUY7bgkulVTKLCXPti+3bgp379YegOB+q2XZIdvUc7ZWN0kDuykn7qKJ6J4Ie4t5ViOKF
mFe4trnqZmIHL/o1vEANMFhqWdZJLb/cW8Q7R2RpCiWN8MpJFgXT2qyfhRUpCt1DtiBeO2DU8ZLi
Bt9uKlK87XlSMcEYVwfwMnwHRew9qyumQp8hzsoryZU34fjj4jjGvIiexNMxhxk7CuuSpB8hCW2O
OUDFOtgnD38f0inbDDWsRdvRwusTFn2kVbG3WXwEJzWTywJN89LvXoaSUgIQU+0HchoNv4We+zKK
m7PoSgUDUg4YvajJd8YPjb7C4oobjP2Uoa45HMQlHn3cAYjICwnF+CXRtIfcyAEzIU7GcuftxOMw
K8mPsrNvDaBJ7gVMib69A8TOn5PiFJipDqkNE+QvF0Bz55ma1P6tat8WnZAMr/cyeG3AE79qBXx1
Uwr0se7IVOcN0A2M/6DcKxqXyBtoEvaf32Gc+asTr3MmFc0bOLnuPnKZUxrrymwpNhxg+WmqGqTP
pT1r9QPUprf7sPetmBOkp8I+6H2d31ExXqJYNyA7eXm+skjmv+2d70AHFI+5FcQ84lXaPW2OG+uv
6PYecCnyCjaZHwGh282uSLuR4dKGNE/b8R95yivQJG4P1OM3/OiDShTy13sfswh4gp8CKHA6xq+p
C39npffRGjjaEF0FH0oQdmlWUd4+S2svNWym5KTXpJTajXoSD+SXx63R54KG8ybknoqh7/aamrWC
wupNOpWu5EXnFFGwwybf2m/b0B57JERcq9DUkkSQT87+lWitAZmv6zWbS58lxxRZDmMbVLiwNuPS
DhwFfYRuvmWinR8BgovS5WltiZWn/vuLe1pwBSjz8bzdBeA5WUcg/H+3B7nmwzX/g5QFi6W6tZHu
IghtgqcKwf8axvVYxXKOrmVjF79DBQUDTwfjdgv48pSOXxRrmf6YZmaUFpJRsaXipm0Ey8yzZSiu
kMd88gP/GOA7B79AlBhzJgHzXsRepaPWqigM9hOSM+aG3FXjtqE8SQc/ITDd7lr6DAQp78AsNNnk
7LMcXOZb026fEeGUwuFL6YpqLFSshC8z069qzspJGcOq+H8QbvQaozBY0Z8cbcNjyMMcHr1RcDRa
MMd55dOu9YFfqYPJlsnJR0fp02Y7qlBawi0L5u8tYAtv6w3NOept/YoQsmWdYZu+1HAxyyhjit5z
ZRhT8NGtuXaUVpTr1V6E+17QubOoPaLQfHB3jv2xTSQ0DRTdlDRtD7CiXtbGvCoABmQCKIPNaNbf
Vj7eVoE45Ugl4+fLD5FF+mklGFGqB5+2xJa956bhcC/euPKL+QOj0Jz7MX0cZNmeBOeJj4Xsvcf6
aJZjfnM6XjBiIbBiCHsmLoUHnvzkb3T/aoWG2lENnZCBAoA0FtNS31miygz/pgaYgkWX0xPvsltN
ADW+UDOC0Nv/W1TyUuMdWGIBYOLj86J3cznzDxBvxmzAQET+dae1J0GHPRvTtMnCqOb1rfL6nji8
bCsbNGNFMsMkyAKTuVN+Zv+3MGlJNB1dcdlCfRGyv3DFG+iBfi3Ifo/oJ8YwGqOjf7bAaqv8R4Ij
JeleghDc9+clEItxcsGfYrYDIgTYvU+BLv6ZtLmIP2f/H2eHRZvP0+yCnZ1N7ONTJaBGgg3EyibB
/TYQ9uokMudgVXv1OAoCEu16mQgvRfNvNd54nZo6fNFebkxSOfwkHcnuHtCFlcUqgeMFKisV6reU
UaMYfk6T0N36tl3GgKtEkF/iW48rPXG+ptbfL0Aq1p5ieUkEeLT3omUJCVyjYXbmudk7rhm9xsim
fPgbZQ9hoZ/clpJzGsah6s7w/QYHaqmiqqbQ4FE3DoDSxURriTnF/9dYEJwfsT+UcDUNTVZH+3/b
M0EvDdS8PHvcaxqMkefyKo+/0MOD1iNnBQWE9hsGuVxgzZuXwANtf0WUjpjL/TF1alunYog/PSJX
v6LdQLGet2Rk6y/TutF4oVrJ8w+bldW3ASmUubzSVSRlyvDXKspIiKLB1UC/aemb5tetBof0Oa0C
rNLW87WuAE8Gg9Q6qlOpU8yCs+2y4G+uQv+/wG+BgcYRVHlDMaAzsd6lhxd3c5o7d2yMGUbGRCFU
gDKm7iYt/UtL/v21oMkGkiuiATs1DuFwn2sFuL3vTZ76JSSiCMM4SA/ZZHA1rpCMLuoJzmgWRQtS
zfgajjnyL14P5UvU7bwhNRar7hhN+ZLR91pOk06mzvv7G4c4D17y6OHGVWrPbxXfgV4uy/Evd5C/
vnUevRtaMMLvrQNEXgVJGu9ixAI3p/FcwYnKnAoSFgMWPlu/aEQOqNiZel52qhVWTPo64WhBk9wN
Gun5ETvHoCta/+tHWpzN7c0Anu/I51hmMKfdXh6oF0zq3F1rdrkhI1T8IGDgC8vlO5qHjcmxotQK
wBI/K9wZrEnfBVSLGWCa9CEb4FaaD1Q2g6Nj4aeM27M3q74NTRJQLhBu6mwhEL2LnjgqrcCp6mfk
SQYVMi4ZydcOudvGVDSzO3N6Kph1525JWPyF1npC2UwnHYq8gMc083E3tZCoIHWSMxbcL9NTUgl5
N6s0fBuGM9y11m2JVrfE+NV8JoDPJd/sFcDSYeHjOFpmdem0s1fvlAQjBD9q+2RVI1ppMmMUFjB0
x/z9SpgvBFbRFqTmZCv7qw9Tn0kR04CiY7B/dAgieUCoJFgpTKl+G8LRfSyduV/3DPDvQRN6eLAv
4yN0valf34e5x72cUZnpm4s39CrKX7v3N3L8VfOdZYwDCaugAsJM50v60klemf/fMbnFKFLQU178
9y9oXDA8E772mb84eqjPmAf6DCWfd5/zStLMIDcaUTuALz0UcAuncRyGxFnFjFWgsqecjvII4xeG
bRySwiI+12jA572OmtdfcZ6jXRlLiSgzryVn6UNVytUswkT51Po3r4Gug9dN/t/4HlPoq2xxzmJ7
PyNYyA8mfJb1OCU+5UqbC+fGxFU5XVUJoTkTYPs3uJ3/yx7WvKekknztgUgIO4uoIV+CNitA0m/t
ue2AuEfkW8ZNv/WX+3KU1N05ASIoDFw6OWhj5O44rvh1XV8K2B/srbi8s3O+F1cU7mt/3JvKKZd4
Gde/WkHDQj+FaQ4H6eaAQqVR54bI4XwXxf+5rF/niyj3WVBgjJIFcsGO+Ro6c4dmNoIjbuRqWpYx
N38DNaxz+TUgRhItp0cLDqYs9ND5JsToQw8WnH3C5J74gtVu7XtHj9fpumq78HS9PgvkR2suaGiM
Lo8CNxr7aKx/ZucASSSn1ahSaFaBxgFsXMNokhk7jSsAqqcoPmymHGBKoGYJF3sgUF7PnClTsk/i
yOaMxiyBWDyEpX6ywc2y6tNIr1s1/llo2C7n/qGWumpDe6Gk8pI4mA73DQGZU7iwjH7pNKlg0HJf
CWjAfTuCeUpChEmCs5antEmA0j4B17JVyTAPU9hsbX7hwi6T3amjhY3hLs6P9ls6K5btCxnbJPFx
G7ZceYXje5OXav+Om+6dLv6rp+Vr1Iq88v20FH+rx2JcAqQw9fOESu4kYOsrKInzfR5AVaHc6S8S
3BZcjTX+U5reaM5GfqmVm3R6zbMIG0V1EFqNvFUuBXbFCA1R19P4HGa3n0X7O3toOoXgSVI8IniU
9pCEwP9iN01iZLE3/XBhnLrDm4oTfSHF6+loh0YUw+Omu/c5RL8d5OAXcMJLJ0OYDoStxBvzqmxe
QV0V4iVTrEluRszea/2KN4URFaCgGTMZ3br0CPR7bZ/NZ6+hRIRTfn/s+Y/6VkgOh4lAakXNyK+o
pg4B5VwdmrH2+W0jO71Uz8T2F1LuxdtRsgLSgPlc271Nl7qTwaM5l9aKd7Sz/KBXCcKHTH2JLKVe
Sn544FI3OfejU8uU6AYHdMtNII1dFeAGYyZyt2oEipg9/HnoibZ07ikIJScV5zurVH6aXx7OHiAy
wB92Vd/SwtSWKvZqT64KBvNuKlP7NTlf9FH+vqEUmzZjVSWEe4ZqFKpGqqwZThSntMpxR+ItPFsl
a7hoD1Kpfwfe65Wva0ukTu6Kp4nHfGmrkpog5HA/1taN1fVGPwSr5siiaKM2U0F9c3QLgAPH7TAU
Araq/7jzSm9BdHGcxpREEVTJ9aYeERBMfx8rMzUtIjhBdWnU20nTpNzPKhCg65T+ocWCnjEN2+UE
T5tUVoiuVDN1eT4yqbrtJXMOBtBd19KZDh6AtIAYyFT6lFuvuBiQemVKI1DjKido+tq5R76V8w7T
Fx4OmA4lU5t16XEdhYH0pCcTSvW525QApx3Yi0Sxb/cuyJoQLFEiYtnoQaQf9ZVyDBEKFCtHFoZj
yvuf6H3ZiWGdvSG8G3YczdflErStj3osmsDD96xjozQVxogxu5SgdRDdeIla2ym8E9xvYWrZ5LL9
YaB25kOjk44RSibxNDpUXV5l4tcQn4WSdaLBz9+cQfXKmH6z2eMF5LE3KpuKUWUVa3+s0zGywIqr
QVG31t+YdY3knj0qPmPggB77nbaz53fIQJG5gAKMBxGG2uBV8UnQeo7bbROJ4nmW2WL7xeC6S2h0
1aJw+FPE+UJxECOGm7LqcL9d48cn79aDmSWgEI3FXEhdRUq75qrITKxIsfYTrAGjLRAfYHqSX4bo
IoBbRPXKgLRH8bcujJPw9+Ns6FIG448Xjtakz3AhW/KB04j8RZwRwatTjHlqu4dSw59OwhruzAlT
J3O6vwVhyM1sYUSj7L1HuMSJJJQzpGdqnezPFhENN/RzD6id2YHRbYeB+YPlf3htdw1lRPvDXtLd
Gg2uE4tgeVrg9rOwmmMkE73CTnhgMxUmUYccVXuxelRY9fCorrEHKCnXZAxk2AWmjYyyUIvaOLFz
BU/ZiVLyaimlC5c/pcR1yFBtfIefr46jSGNhEqVnTivWQeb+jaU7DWSLJbF0kr0hDJo84Y9ruWGy
hCDMZscdvcWy3AAQUzV58RFC0MUCE+VHuamrSDav24PbkQOvXmHIw8hCSK/Jcii2ZfqWGbGoobhF
7Kel4g8UGQFvbt8+sHCnaA7nWoxnTZq7FPx3ahHTobY8YjMcqlqlUa0kl/+wFYGLAX+M9hPx4D+y
m0JMm0lHEUB/1sI+9x1vUNfA79H6Q9W6+mtrA9fkHsRz/NbjVjoqJr70ZUK6013xeCWQDnYx8YrT
QpZa5sYxjaiPkMaAChXjJ7PXZ9Vm8HJtddPo4ITiy0rxFk12Mbghm0F0y4U58JXnuMWwknF+5RVI
dKX88S18tKBjGIE3gixnDwpw0pRdeRSedIsXTkA3dKKFn6HSOeiiHZlNZc7CB0E+j2s2Khr5ugsV
oRRGxv7pmj7SinLOd/J/XRxQDRrZPceFAbKaarJFS4Ke8AGyeHcGVDe3FjHIECyVBC3HpxoIOUN8
IQA0oLf9SXRGIKC2ZSASeXtC/kV7+HCQ+BNlPS0OYkzpB7N1q0Vq3yCLETWFbYaxncaaiZ/C7uhu
oCrHf26MhCaQzc8heisP35EdET8UnTCwneBVge21Rq86o9Lv2FDVJnIco3D/qSBlQ+iTGFyM39eX
O+0Yug7uRpOA4CQRXOchtIKK2Hv5sIJ3kFigx1zE9hbcbNdQFjvqxx/FG9VivGzY5yTttsgqKUiP
Hqtt2X2Bfw6ws/f6sSLG6RA6mhVtu80b9RwHjXNcMtufs5nL7B+xivHOmzWs4OQODYEC7Qh+zHdr
ixYyQ2YevNkR+nQkShpQYj9UVqm71lWqlgth9zFrdkovOHigHMfCT3Ye8BBBUpJwhR4qYCBlPyil
z2UaMQugr5bS3bI9KgWocXiYvIIQJlC4t2gQ6mRJfm28zMyiw36c+np2SLx48rBQMoTjacxK4TGz
bYZE9wYg2WQ0BxE6CIByBruWx/DR+N6a28WHBDbmwIOIOdhAKLV0e2jDHnZ+8srXKuNJtDl4J4eD
1aQyCZOrsaEhgG6DrAinKebdMb95tfpYmI0i+HVblD5ODilllvWd01YNr0TpU5l+pHVm+SeKwZZE
wuqY1zoCVAJlDPyC6H3Px2HKkzyl26R4Bt01ol7M9aW9G69fCe8wf9f1uQ4ASR5OsI2ZEWD159SY
1YsGQPEPy4cwhcQXQf3VnnGVOAIXQaUqFoD9heGXKVy6Ot6bNWF+Atl2413pSnPIRku4TDao52LZ
SLLdhp5biWIKV5dGNY9dB/pT9edEvY2lg3SbY3S71WxxMtDO+KxlTjyJ0PrQ/N3U5l5rCCA4+z96
BDNOHKTZxSfgX3fGZ0YJFtOL7PP8IGJAzpGOpIYUHi7Io6ZANl7c2bnYM+XY7sf3hkdroxOfYYLj
GgDpxpi+oH6aRnOeQ2mLD7jN/wRKvXWARP//AHW5orYhFWZTiEPAKqIjWA6kBHMfPCec8ExT272h
vpsbzZ1yN9HtYHDoWLoNb5ZbCd1R97+UtKTR5Nmmpp2DJ4Buv50lWjJ1zRYQTejB6OuBrAcq4ziy
PXYB4v8lN1S4MBFSH/8oLtN6VDQhgNMQ88fDd/q99IjbzDKoo4PWeSGsHX/Zf+nmPs7TmerqneN0
hxca1UEfeDVUyn9JDPMoUHUezp+qopl5/TRZjjsUW3xDRYm1UUfLKwq2578+1Qu01jEVehgPcsC4
wSitprSS1nakWpJegc507mAJPSaihata373yEpxzGPy3ANXQHD88otOSQYEBM0tSUU0KNsi7lREJ
A9QDTPZV0M+ZhM2AXbdGADcwS7WfcfTbcw7wcRX26G0nBfrPrhvlagCQOnPyFTbVPvPbFX6y9a6G
ta8OWD9E75jy8aQ2amZzUN6FZg+ObPr55twxiIVcn5vX8THq1zH31i9PuE1hX0c2Sdu4pPFYOKP9
M4yezxlTJyAUVc8L0vqJxF4+1JWo6eG9xZknzO6Y5zCecGXgXW3uOy5qVnlddtqYXOM5SfVelaed
exCNrcOnt9lJQ8Tqf8ZRBvEdPQ+LQeaNVui7h639/RIUyL6k0QQqm3ndTAb0R9IeOkxAymxSFlRG
Tff6LIXTNfl07fcDV89iBgcdQpi/32ol70bUJrehgmUUsWt1ypgihl2fHWtvpjH/otIYIR7UkPgG
nBK4EzvD0MXN1fNSAfjbw/d0MQQrbpwpOTpgO+QXv9ThsdwMbGsO4QlqjFbcmoSKHJhmPLPGE6mC
jpTLXgemDepqU5Xt4hkZnLIEAbvSXRJAx/qyhbMZjUG9zmkMbSc33NPEC5wt8u4/yCgguasFam5S
1kJhh6rXbs7jV2XFrrml+l9noBYG3oDHLx2kGoD+ahLWY6Cq/PgEmtzuGEZx7r3LIz6tr8CTgeUX
ECZejfJuKEPpoQYvw7/BgTQ99Kr9Wvx+nYla6whLhlCzoQchPaqB76MS4QvtwHvzHWzzLT4jjDIP
S6s0su4I51Yx1MgYdaKZCvwlGfESlRoJVdVtucQSyvRJnu2fmo3GROX3csMMMrPSlpyJkDSY0RUN
tuh+yX3VTPbec6TRVcu54sfYl5yG3R9iAV5v+8bv1IVLLfZUO0C+svBHwDFSSQZznuGgo0fG00eo
1a/zGRDURkBaDBr9doURUPxeY7N5HTur7FIbRnSyNmusBbfX9uToNI9r9POY7G54exqAiY8xTzyW
oC7XqOUBXFFWyJas9niV7pgDbnGIrAk+/ciP0exJvABDht1JDuS3fZQqMdTagYnWUusBoWlnngfM
WUwTQ/se0ZqHWuxQi9xScr0N36N2F5/idXZrDoi6X9JsffGgvfTUfyuFTCx0wigUuXrSd6DvT6QQ
D9GLQH4EpBIYL7YhYQQdWzvLNgncS0lhe8pVU9Hh6BCHq/WLLo+Ad8UOcbo6B8GMTzJpD1BR0HIY
h3sEuP8X5if+FW0yVliR+QGk2ykn88FC3uAvnAkE5JPxwE5WXukaqdGNFIdkSYXTGE0P6oW0liN+
MXqcainlzwmfij6NzGN79Ubk0/AljqNJ2Rz4JRZsNpnaFqdmvyKNUHule8o/z+yVxdj/kZEh/+Sh
fPle414iRU/Nw1TUGZv9V3ytB3sGAlXeXSz1BoLIYRyNp+NEjlxEWCSVVkvBcvWGxCv7aInDoM65
lQtunyRoW9FOFg+wMiYpS5kcevcGvDE57BPlYQZxyoi+crGRSX7HYwzCwv4xwAYFWPSXyAR80/S3
jZXrhwjqGYDRjjZust1tr/UBA+2DzPUHrgV6nTbgAiURF2X06COcR1wD95rhobGC8c7maPbkKHey
BqCjG+ICmbKFFu6Lqfpg09pCLYALZPdkBoBXK/MW8vWaZ7WZlKh01tL+lbpP6WdI+PHyEK8vYwPi
SR/K5rl1WK9xdBqnaEe+tv0MQrU2KGTCRwFKNDvInqDsPcA4yiFkgjyAvr5LJv1j+JtirMnvSimK
Z5dh1JerVmXyEmhacMkgNjFigVnQahi0UnG0/jHU+HCc+uyeSpwcO57J07+nrbVogB5p5Q/XsxSd
r9B2hIEqr78WY2bZuLtCY62GERUGC9llg/09YlBUY65K4LC1racA9UTJjSBa4Ig+CxBGFlqfop2B
q8P9DmIA7qBH4z6h90N/okGqOdfi9ctVW3oAWYqsYsz3SBFVAualqJIRCjUZYO+rXeSctvDJl0rn
lE0Bfqoq76GfkMyEtLKZp32XrTkOLswEDvJTi4oKUHqlQ+U/f8+Gm6SkZXMth8vqPEvE91s7EA8V
Dg6gktu7nreJrKOj3k28TQKBPmWn3AzXQMiW7jIZSjY9u0DZzRlQYl/k5UwNA3DAUwkl8z1XZCh8
pKEpOAiTewxeog+eKOHkWEpgFuuwY8O+7/iOlgANAg9XhMtejVMwYemygcoW72yOt0vtbT8hKDn1
bhdXkumIdT2vRZqY3kJboSfPi8jdGQuERHKF1aAOq6yo8jUtK7muTH1kNQkXn36sqJLygoYEnxO8
AnGcVbeWZfbG2z+7MK2pSr5JC0f3eB6GA6be0kIrzi0dd5cQ12km7lvnn0Mzyq84/54Swqa0pmD8
Mhr1cL40SBORAEYEc6xryJ7WkttcWXUKA2rKZuUISgzAwcDfTkMShm+JgxcV2c8Qt434V+nCGbXf
LrwO+UClqd2xXmRNMGj3ryblFvvCRGQ7eCuc5DfW9Sn8a9qQ4+9NVk0c8fvxGUW9phmg/Zv5jTXS
IYeyBaKZTJDwaO1oRENJMPn6QeO5pMExM8UhOCRVsZJZx1cmh5gulHjWztY+tlXhpOc8vhictgX+
o2/YpLKTTnk8sRMsZbP04DKF17H16euRhb47HFGl4pLjWdKR9o/Qn1Oa65JIB+YRuOufa9QQBUjX
S6A0e2cCB+qIgOrDcxFmyU/64c8qVumMjbTxDj7QKKUMmPWD6rhR+gaOl3mcXcHOeDeX7Lu9BKu/
7LkeIVtARycwsV4gPGO6osqZJa6IjvUn2eSWbK3ZDjy20eppM9cxsqszijwX+/cG8ZHJQyyy8ksA
rTa91VmSY2fkKq/3kIbW5fdSu/rQuc0ZHA5H3fFwWcmnl34bxYS3he6+2h9MCJbMTsIYP3+1reGX
MEslMvmM2z4OZvvgK5kH3JQrO2ICKMGG6+CEEWaPf1EIvRxiUvBXd9gK2UOK7LHRWBltICo12YbN
z2+8NLQnsC+hL/W/17WXS1oG5PXMaHNGaYR8kS7EKU6NYCXR3YNNsyUgnx7SELIc/o18yL5lwewl
JgboEjbSdB7JgFxfqL+dBsEWT3A5VsgDO+us6YU06macclosh2iCJjXFiBAmDnZDLCc0l/t6RIXz
QCDtf53eeEHyGa2Qy7RUAJcv5ItQrd59ZR2QVNx37P8OItUakbAdj0qXg5Hf3WzGzGGypyli7mG4
H5xpGbIraat6xgWaEEJ7BaxfwR3rWfOy23nA75oA3+1BpfaqnzB41KMGu5tCL5YNNuILqtNiFy1Y
55f6sRuLNDBDR6n0+swQWX8+jplECQ6nvBcXlu2tgvf9VVjzZecULM6PjoqK2oc+YNPQnKj/MZ9Q
r4wSLZjGP6NAtXv286FLs9Qz074Aj3AEXEfBqQ5B2yIytphz5Dw4My8sBTKKZlc+RS752zb0dZ8c
95vHKDP4jydc3K1EFYe3EaXR5EjrKt2XT823Bw6DJfcUSrq39I6fo9Z8SOMPHdP3aWRboNC42AHl
AoSmN5ezffGHxnxEgW6IxwPkcCdC/bc0r+LlvwATUYNAICpcd9dsAUyG625+dyeF1RvIsBu/k3xp
oQxUHIcRL1DxQkaD7wpcADLiS+/7/8kKmuy4CXw2DbAQNCjBuZnsC4+8n+7lIucE0VE8vZlStK/d
m6ve3mMRH3OQHIcx3qGzwbZ9hsl+CON/Jfu6I6ujwOe53jqDuFP54TjXKm2IsfrVtIaIh/BjreAg
DXqO6yGQNP8ja9XgJUd/1MfBPUauKchoc3BvUKSNfvKJH4079MXGXk9d1pzlAwXVQhaKx9AmmGIo
jhiRBuHVNv9cs4NQoiPF8JTv1nFEl/sjIHNeGQNCBjRFcy94AQymgv6Q2c1Es8q0rJuWberk6H1S
sFRmy/usJ57CUBIH4GnbuNMOLBe9rbiFMkWotztwPI/0LM6kpBwOEa6XBnvbdIlbfV8MumyvpzHk
7mZHsfVHU7Zv8ISXXMgL+tw28xBHn/2gxwFCJ1jqV0Cijghd75CnNMy4PoyXn0HivY72xPag2oDv
M1XJteF8qbp+TdPw7LnEjv6JFCldk2ujS33FkEz2MCSz7bQnTtF0DUVi14MYOWnyH6i1g2AfqEwe
KHv5SBQFM9jmBJDElT9Es16nkcjn+PPb6qH0KnK6qC/1avEiSxXv+j0h8xxk0XnSXyfECgxpO9Ju
W6l2s2uBh3ZP9Z0xLhaoUJt3qmGcOdbAohItMRxMmuGiTJMgDgliILRqQEIKSHHnUmqvg0H+K2Tr
Pcl9R3X6cZBL/s0/zN6xwh8iWGhhTxsQPJKSCOUrbs50ANm6oy+JDmODeFxlRNc2CDogDXBBETKL
NE++kXtYlU9HwcYBO7PP5MqkNzKhy3o0cHUBBCGeEoUMHS0w0TbFC3PprUF985y0e2DIJaU6O1Db
HDiS4KZhv4zCklpGEr0AkPQVAJ2Ca78FIQqOqSmtaKFJd6QTWtj9GnS8tgeVF64O97kh7d9p3OfR
BNvoa5JaKcm/x2hCGU1TL9ZVZKElRUtjsPHP0hA5UTXRnF2c2++AZDy5GXuymhEQ10FTW8e2TN/R
HiKufbUhvLTiKWrjL4CwN7llgaPLZ+rCR6nvO0Cuo+jusF8+lfHO0CdaamRoFo6uxXqV3F+5uCGy
upyDag9BCWzq299vnfLJJcxp4UqRaG7rF7CNGEN4DQCgWJFmduRzDLbi5jUgCc28KajySm5cWbsT
0F+OK1zck0Xfo/XJ0V26oSclKBFKAnBax/IY/Zie6HvhUCjssrt/sBeXYmKZpAwh61WJCl2T7qg8
B4y7mp6jkkiw3Pebcqe3gxXtyGYFR4apjvd3mxMkhI77yFsbZtOV67Ix/TZ+cIf/t1Yq8hqJxxj8
cg/28IB4GMrP1afpLQD4AmifG6eD+Sp7z68JJO9l3zjb3/ZyHX7t5xRBuqUw7PpWth9MeIxorPkn
WU0pts3S74ihNoyTIU1khYLWK53ASGPIIDuO0zhwKcqC2adl79Ai5/26gwMKscQL6vpZwpLhUo/z
eQG3yJiuNHFN0QTpVu3vNgjATEVUiJnlvQOmMtmcsDOY0jip+4mxioLzToGCjtrNPs0QNQNoLrgj
q1i+dq84WTIpVEzCraDSrWIn78q9S2dCtzFjnX2GZhKZaWB64XECht1ppFenKf3eL8ZuKqhwGq8d
tnywNwpBL5kkyuYoDaESNobz7y9N7SLK1ULFuyERMDPg2xTjJltNGtf+YDefkSHbtNHl/e7Vmzla
0OCeEbrjp0TtKRX/NsvMuhe3Pcb02N7jsq6tKI/RF2TfhAO6mNdBpj9oStZHKA6y8B/9h+OFkJJR
PsJmuPqDTPeL/DxBv4xMs4kEVcn8y28qkY2C9ICYmK5YTgt9CJqMVia6nwNNycJ3j7qc9TMa1GP1
QU0YxQ6m5Z9arC7jiMtFplpJCokoq6MiRhrvllqXzfMRrRRpeLODRigz+TpqLPsjOzJevdXwbtnl
2Z74p4IMo8OPcaeOYyOdMYI+pKrtBvPKORHpVlYfBtaAqbOxMecuOPTrjWy10jMh18d1IurqROr4
Y53n57cJ2ynnBvC0t3osp3hE7iVbZbcaGYuXsh7vnfNa23YBQNb9NHAaUqZIm4LIIElP5eljGPJ5
3eY4v7yKu734frK9k3r69dKf9Zq06NtpnI0CWv6IFw9TsS7XYWmsYPHojJP/OxgJuNoyAb3mv2qi
KVZzz69JUUuy49Mugbs6qJkTCQpLgrxM0GhdFi1ZDrKmRA6HqOzp1HqdjFp/SxD4TzeUOyb0GtPu
aIHP0wIBX4QFrgz8TRStAVxJoL8z8K62rmt8LG4fg/ryplh7ElJKtN2JA6cpKJ+jI/bOp0iVsRud
mdr68K0ire6N/S7KDgnWVS75gFiXfNs0vl07w4ga1GKWt1g9+r7Wu4Tc/rpWMoya9ICnf2JzRfNc
cUBh3qit5hxtPdEf9hHPBQXF9RQdCqwC9mZ3E+s34vcaLo8GeXaOHw4SbK80Yp8hn/i+RqP3eMOI
MzOiLITeOpa6cKaUT/rwFN56o8+DNvIMgGSHKc0Wv9byq5lR+y/2LWYREnvMZHpmCcf8jRVs7kDE
c9jOeu6C0yrvoWckzd79scYfTEym5Z1jvoqoMMYjr5nsmrkysqbJkJ8pnqUDBuKa5Yr5dVeByyat
3TvhSckUJLOZgVu0hzWLtE4nEYFRlMRNteZP4bokVK9Souq5/foOhCwstNH414JGzsxneLV+QeQX
3IHpu9yq2QtyVFQYDbLBmU1UkBJqMMTsmN1b2FCnMx+dHYlMbT9XJ5VtGYqWfksZJxSj0cTO5Bhx
xECytCOSTyZBL3ykLTN7zZrl/866eOXf2uhoxgG/AszN4rhXDUvRqCfrWmwcKtTXhlDwCRUrdrF2
Cimud8KPQ/+VEB75xmnYwL0K5zILZmYNsehNuP+vU3ukgFmTUS+TRcUSV5saGF6uGbaViZ+a5et9
IZ6++QSbWNj0pTPXjmn44/BH7HmsQl4S7FiezhUqJm97naGMOwSWQ6+H47p5c18R/QLbfbj3zQoi
VRokIOA2pXRaUukK3L6AnchBVANLGQjQ8Br3xtyHQpCPxDkC9+FGmHgpftagbRQrmtOftaUQuT/b
VSUPJkEOdCD7cph/v9JTFKHaayMTzwISVqrbGgbB/RHGKJP+6+v0/ssJdBQiAKcBeQAUKrQlzcxT
HH+aT700hQqFK7lGHtysD4YZupG4yrZUxhustE6XQVunxJBb1azL5DrY9ql2PyB7oZfRfSl7j9RR
AIUFm3v4cRqERzbsGo2XjooEFC899v1ghzNcS/m4I+Q+YWtOiT2H32+VICXRPyBbB7uIGl1hSRiZ
S5L35HiJyj3H7OXXglv/6wM8cjl3j/4QTC/rBegkKP7Xz04RAesFHKn/cHdnRBU0U1J7jrhozRXd
OSDQYWW75s1/KDagtOZaLysiWUBPX4BoD2mf82o4Iy0eZvYhO/MxoSdhv+g8f2O/RHaWubPzYloB
hU0eSflU6wzOo4Aki6epDK62ORcs6h7TZ3jr8yjnYMybJ+RsozVdJWrp2SucbFAIpE7dPg5CS2GB
MF0rCsPrHUB5PnrHLjefTEPW7gGVXv+cP0AYPZKnvUkHFO+743r4NWLlzaz1W8Zi100hKZzj5nTK
vZ7hL/URgszqFMFKIiWPTIr0ER0YlA6/BGyYZgtwpUfmiUuXuoNYOzC5buhkL1Co7HxX+L2uTHdL
+DSMSHfO0aiNMpQBYZ0Ni+/AOOjsOIGpUVtWMLpQO8LHb5B7cSq0S7aOlskayc86u+CR5MFPhHVV
pZMU3lZpw987YO6JR4xGaxHuCX0BxWy3tct5aQxdAoaf3epWivmGcHvQ0/cx8k7a8Yfs5PJlnXfW
cuditvuix1uVLQoB1+8RVLwCZZw0MjiXemx4Ip0alga6XsqQKcwk+5MMoNvmu5GunCWsvdyNdwkQ
E1BV/Gu8QRl0aKh4LDPbOwGu4PEF26Cgexnig/avrMc0rg6DLn/kXWbnjCmT6kaYoAVZHW43VRfD
5w+yDfwaVvjBKXtFS0IKuzFLDud5R43zhDqFTNyf8trDADnR70VirkkNTGaOuJASUrKyxteiZb+v
ByJxJPw6MvHx+9n/b64r174MCNbL/e3RJfp9dPv0ZFGlFkeb0afbD/iqH7/fLR+2x0lJ+gQeSCr6
71ZDU90ryYR+RH97+MuZ83W8vIoCEE1jt7oh+XfWU2lTkPjkxqt/DtR/LxvOrsBBE5Gl6E0IxjBw
QnLFdO1+qx1afM7aL5+3L01XXuwVSXzUDVTzcMjcRbjc8860vuCSJir9qFG9/RP+vwd4oCv6PWKS
bBjS6Cwqa9Kf2cRMscDDtTZzUdP00d/ZUZb/uEzJQ4HbA3cOZLlZB7mfrFlw8eZCHlIihcG2i1mB
5l8d+FTlbzc2PseJJtJaWcGN2rtDJJKNDSbopJDebg8+3+mHrp4HlQ67dueIAZBDDdlRogR3dGGB
g+fZ5QKpy9Nc16AzSoEJ7B173z1uhdAs6lHwYbcr7OUipRGcTtR7JFh4/7MQYGa2BfU8QIpoz3jn
ix//vHgA9SjKEY02paFoChQE2pkPbZwKEW9XMJy4o9w4KFYsb9IOZYCOuWWBw0NgdhWPFtYkYq1O
P1LCHemCo9KcdacBngUVqLYscffKZepNIdaOP88aHo2NGVM4snIcaDQDEOcPZFluRs+F1v9oEjr4
MkR1MyNo5KneCsAOJyI65Y0/jKOP9rQWDN4uASVCSEEgctOfi3hEloxW6H/eEi4fsG3KNH6ADFxq
RaIaislvlAHuD8EzTTb/FDJOosH+23FiHqm+CDMsSi/Pc3KjPstrVSMqZzmkdGBPmDxPIfA9aOwm
O4/ntCYrvhbUPRJALzEFvuwdh3pbP6ZziVRK0TQsMLCQda9AkyRjWSWzVnINx95jVz8/VGNtRpSm
/j9hGi5MXn+vXVJVZL9tPE6eqm0byNxSd1I1KxbXXAmQ2C3Ug7DgU0c2cV5KW1jrUgza2qYL1Aum
dmDO5G1ZCDCyycXbwGqtvX1L0y9c+/zGvSjUKR068RvAcMws0reJoo6Ypv6DswKGYSCC765/Ns0H
lq93v49ukO+mx/L3/gxaHgQlHlKlGKMMSRf8jKlGizLwaWKIrFRbjCFy4NOcoI3SMDqXttlSRT0a
PYo7OmjLjAdCo+i8x5qt7Ne3Jij7TuXd9YD8IxcDYse9m7vZWYPL2QxIIM6ptsumseFI2nGS5zn2
XRXUd28ZUDJQvRd9sUis7DRTxWyeDdT17vxEoi1cPO5Uy3kzxSxWnj5OwvBnk85UyWlEcHB9Kjxo
6ouDK+qE6YVmVlsKPfn8VPMHtQoSjIFwZQ+VnCBAZfr+cWxHQncGeVuG7uUnEpmBkCE4cZY7+7Qp
zlWXMcVeZIZ4qfrNL8Vacodw4kNaqGqaujL4SdLCFDBPro4LeTavGmzq2L5DPhHxCLLZgPVpy3FX
6r420Wc3AfDOJGbuxESi/q+mCXspUdlAdGppJDkr2HFDEDGx+yTW77KdKPCNLSHaONCxv+jrvK63
552oavZqR1haDJKav+p9640E/jY2MJLqEHHTqfR6CXDDefkp0+5r17fhWL7nK+zqXx7hVjAbSRg/
iFz+25uvdH8j0Y5z9KM616YXqZxNdYCNliBvBSmK36vgX8aHW0PXb0OFmbuQ3fcJzE3m1WbdLahg
5Lo6sNeL4ED1CafV7TBRchwFN6n7yeHW98n3/j3ihfBPZES/YHg9aMFwHaXv4NWzg3wlIPBgMt+Q
aEwMtpSlEh9eIDcRERFQaGm9KYsxrgKOKnAZyqDPpvmSQ+UxHvVzNkxc5v/Ege090ZsDy71Owreg
qGGPxXSwvKmWnnuCGGGjs29NDvM10ZULUfcPkZzO98XuPM4wleDc5vh/iC48hzQjCcJsG82TLgMR
r8g5wU2ukxcSnRcbgQZq9OBvUrXK4P3VeQMBVp1m9gcfBDrCiF/vwHVLpxgtRZJ/jvw2fbkRpoUo
vfxH+xke2Z/fCTzMxnNAScTZvooj51vK5lU5MQ5/mzMPIMMyd7fZAzqa+CLxMNgRuvxFX57WEoIX
ck4exPMZemYy21O+1Ueqf5NCoMVXGwaT6rBmeQ+5tQU+HPUQh6UK79kQuQvJsXu13HScCDjFDDUs
4YAXlHt4KDh2BkXCo6ve8FIJ7K/xavgcXDAi2/51juSGTbAzlIzrsQi88s1041F//4D9RJmGVNxp
xPv2Wbn5J2QZTRLdPyvQ6DAzzm7f/WF8izhW06vwC/TPyEiE4vq/K0crcrZNy+gZ+VsDnNFXFoFY
a/c7u2BllevHFqwkpuMQR5ioiPpV59zP3zg6rH/trb4YyiwvBwYu+3ZAdQ3fClzwZ5UYe3Jr/nfA
hxt28JaMEz9h3sY8uLt5a7bHbtkCDgAMdjkasgPwfZ0lHMVRHz3e/zwuwk/CwML9K6+z36rFu1pT
dPzYruxaCbIkJs3cAzfHpDwuHxVWPnl/8eII+o7E5H1V81FrqBPO/Z4vIO2WSEenm9OLEGFOHQpX
QwrS77QAzD6DbN6eprDHSTWtJuOTa2lyQG4eu4sRd35uHAYqiV0YL7+GcVKb3ZSQlob3O0R51urV
3RNnWFLi/GzES1wvq8zgccCkk0edZlsSNFVAQK9vYZaxKlbjuOK3YSEZZv7yGJdJDd4NBV+S2gcb
xTnw/mhGoCqXEJtMjsDYd+L/biPVze8GOdUrAsmKnET2wmzSc6eaTVy7WyXamvznTc0w7hlPvNOB
0TZyLRitMeAEG13EIoSibFKO7wIlCyEigJI10Qgjz4mUVaZpsp1/xJHVg0d08qv0i+2wuecZxZ18
Iw1bavOtOjX7r0BS+lBc3jWc/xXW2TusRwu+D9akqqHIVQK8cVSbQzMtrn4u7CJj0ujz9Pg29kIF
eQtVuqHN8EUW0Ejze8YbGB9TV42pYayN1WYjcaTjxmgyMFtjkEB8gSvGYQ9SSZHzZ8/KjlqNbzxD
ktvN12AScb14+UasNZLVVAM3FFtq6MnwLKdq02CI+raBNxqlSFW/BHZuA3U0pYQtNM0Obx4LLlRQ
EIcuyFxNcg0N9IZ6okNooQgPx7qwD5yZiFe/wwg1DpzssMQcwhsnF0GCQR67cxV4U/l+E44K17o5
7aRH4x2jUYNqw1k4NXBZpvg89q51VWGgx62z+8fv7aTrDUz8sW/3Y5RlMo8OFOtJ4GGOZbxxJcsC
RxU6BW9zRl3bgCFVOhY+Wia3HAkDuZizIIvj94u3SqT2KYkVvHK/DVocxp9hwxx2NZgakrTEs3WZ
9VaI7nQrl2toTRU4NUPK6unuqgmqEu5GbGRNP8fUNiV8m9HYQ6lZtotLPk/g3FHNBI4jWjvlxI8A
P2NyUXq+UvedL9+WUapbWJIegM34bbyFdM5WBJ17UAnKTXE0AQH70H75sAgnPWFesTBvgzrbDqDl
B3PvSe+UPsHE+1HnbJYdqdVCFj0tF7Ej3P5wypxkfKVHZ3IGxxFXj66x5otJWI3UxnhtEO0RbDR2
GaIesNQ8yGdEEcH84yy6xVOJUq7Gf2yVvYYEA/FD51zhfcpl2OWIuROOz9+Fl9GBXT5hy1fnTFeT
Hxma1BwQd4jR5GpDL4JBQxsE8CeD+IYoTOK8b3oLKi5E/4lZ9AhLSuSeuPxrS7fptTCskFxUms+O
rrnWZAFa448s6+lbichBChAbDfLIPlveG7xRdvV8SSvKTfuM8+v3NyP5NG8wgmKgG5p2f1WZAH/P
1wEyO4dTvrfHZfpnMN7EvmTBdSxpb/QcbSoQ0JwrvPMtMj/mpfNFWTiLV9rSxEq5BvTQtt3gl06l
o5Vj7nxgX5POnEy2iKdu1MN9QcD8oqTwgFZKPgaVpBSp/ibVjbXrSH34I1NAoSji+Q2Eb2EpI9d+
q2xNGQGqYDF8g9r84g/JNese+wwLmjrXlSc83++XtwaHSvD86hiC/x7+p+5pcbIQuADwiufEPVty
ke2c75iYbL9QduAqX5vLAUcHVS16KebN29lbDtjpvCVCp3Z8Z83QTHjlXjmFkHvZQHY9W7h04LqK
s300uuNbnfMtR//rJtt2YwapZNRoMH2mxWdNYKyditHZmDu4OpWx+4qtBgT/R93a/FAV/RuTTP3y
TsEqBQv+2IXtQfYERmagbxtUzMkGS7jwmdpT4XtWCuBikuxxP8hw9iTHC2GgEPGSJI4xizyLRai9
WkR+zjw/H7zHavWyLjCifHsVe9KX2F809Ny+9arGAwDXFaSecqtn3ahE4TiGRI8gSBRTbaDlT+1Y
Fv779J7D+dI+KQS9i42a2+9sQRRpp05zrLTCAl5veF02vTM3JQB+XGmWl7DicG3Nmq4EFeKAWOjX
yruLTdRejhkMLY+xBG66MKeGMei9ExeuXHMeT9S5hkXlZhOg46jSlL73UpBPJ2JzcLztFpUMgbcO
70j/QHQ1fpUxx2riX0ZLKMYfhEYmFfxIMyXWvC4dfqNluD9K5oe7cSjYfeDpl/bsj+o6NGjvRN9/
fV2bWqkifdEOn7lr6mZb4LHdnMfyWxvozDN+LlJTP0eg8MF8zVEzuI3Ljul+CUZod9Ir0PGaqwLP
odHPE00WV449wncy0tHLX5OgY651w5Yjakg5GARCD6S3zJnopw2ZrZqfQ8WhqyoDMEOdZeHOWcCg
k9yDIbjf3iBOIHkDQxxQ3Y6FJikqRsgJER3/mrIB3snDWY6dej6+2SJlEDdjw2ZAMA3pQzT6fZoQ
stMue7oRZxKqEs2AlPykYaKUlun4ql8tNnKod0yQiF++BZ1l2waGfrkspMJXs6DavvxwN4EwPabo
S8tjZQQvm7HmqSkQ4CnGYx13swipGNY5lBnqm0X3wc941dt0/UqIgox/zJK+VkVVOq5uEoeWSPrQ
jnuWm6r3AygzWrwKzJkChY5/D0ycxW6AIhzffO1S5gR+rFxnmanQJFwbz4+Qd223BGuQTK+Vk8pt
W43cmAAY4h1vS4bEmkKMK/jVDr048KQXmhxOP0xne9PIJJbV+eMfUGxy6onL472fGTUImTNNT2tX
oBZsDOJXZsP7D+YTC7H2Rc8b0pSGzdSMxDHNWAz3BUvpU2AZ2r8PppSFfFGoMSkzmD+LWVwtch7t
EhGp90BAVWV7sJyyDMmnrzql90UuHtSgxWbO7rH40U+PP98GZdBFzfhj1Q2v+ac4C//SCSYHhHxp
kR43dblnBht4Ib8ndXd5q4qHcaz+GsMLYzYdaXhy8wqywCW9APlzH+qZZAk62VUzgCguymSbJjRT
KIvtFriEiSgb8VeUBzQ8HiiXka5VnzUAbekIspXPjdHquGYuFdSUqZkYe6V9LYUyRmgtH5k6g3/s
a7xY3LyPRNaruERdzzs2KEj/DLXl8geY2zh0WFt0ian5DyaM+oONGRGiUKQRR8CPiQ+wrUzYSMLI
vipFSD04hJDDxXbXakl+mRZtpp5hsS448z0KlvJTCUFK5/xSrvVk2sGp0T8TfttudeKJ7sj347Gp
VhnwjQkjMCbEsJElIptX7iErErYud1FcSPwpXSNqqxobhCCDnQbpMYrlyG3uCdyLMc4hh8tZCbkT
4dUtqCCn5Uh7dEbYGeriGzaj6y0jgmCYPor1YC3I/nrJmElxaqvRAp2k0fzWCRfwI03oJmu8VFYG
pNS5Bq7xZxGi0FwRbBUeKdOA0N+3aD7/P2BoOD7ci6Ahgc3owBiXrsCYpMAitUay/UmVqQk2I4Zx
W/u3OKmZKOWSmNUADTNf9UqZHPOM+SYYe/OKGOZhLyLyHAZOv0qxuh5I+TLIvWIX48Gu4YCyrFC9
D/KevzN8VRfHCVuRJPnofHPkROb+YyGwKGEZA+TwuezkqUxCraADSrFrHLIZrYYMs9rnKpr83t7V
v45Kc9mskcSBScFMm34rm8UztyoymJ0tEUojmInfl4Oahqz+8/78pX2fJuo6EDp9vFKfiPKMEcZJ
hAm2yhnkG3fPmLxJsHPYni/BAY4mpRw8oxOvLbO/AeB5EK+piIOV205/T/cgcDtR+rVTrWV36yU4
UHMSOgeNCih/bSiXR3aOXpcyuw79Z5DtYcs/YR80y9ySO5bSpq8VCJHK8IEhmV++AnXW1jxXG6O8
oPFjXRK9kD4Y/rkOFy5QuZTjzB6uw/vbglQcmPCYRoBWwyJWyzRsxIOZYDgxFZ3l+2MAp6q2Z8Cs
xdLFWtzPJMCwb1R8imwyq/5uPdxZmW7sG87dNCecnQm4dESuPDe+e5WUUiqEgeAhE294ARZPSdAR
H818dBrMyY+A5oVCMtNT5HnYYY6MV5Ia3G4NwfLeW4kb+dIx49hmgD/7uC3VXxcWyROuzgCqr02u
o0QUocCEcNbLa6uMCT7emiG7WBQpksLn4eiUYNLPeKEXLYc+XawRlfxBC5sHUnDOCCnOUnluB0cV
IjXe79gaezh26X2ZF5Uyn8cN/72sdi3uw+p5CuGc58nBqEC67ALA2fPaHdB8KhOatqVTuBlDVxcb
WS4Lt4uGZMkCo+zGATDFYuWAOUha3ohu4DHFMeA2NXLXRiMcfhNHMxDp6LMLgT8reVdcMxWTZRU4
LglyiI/RqJoy1PWNLUaTnKeOVrPmKPnRTjl+FVSZSi1Q341D4cmASJWBAXOJKFQzeCwvrPFiGi1S
gqS5O0kkrjJd7e9NZxGG/x88R36CVnw9BmSrYsVLDBzRgiSQKwg8G1t2NfKrAQs3GWWjFVqcleph
HszZqkVRMwgKQtuVqf9HkyxxZL0jI5xnHUSK/CehP7F6GQc//s6AkYR148qn5TeP+HP8vVg1t5kq
JtT7o0/1rgWWZvVCqp27MO+6ezh7a8kXEd8fBqWNdYW9nO6tUjnINivpXE0X0otb6g3Cl1lbd8qp
X6VhXsNANiMRC7WZZt3FEsDp5fdIQKJJdmZvm7OzYttCXkYwLkV3A/6Z6Vlr0ott0inpcbbvPWxx
2HlRs1mhO8zUcAk8P8uX9jHLGQdgt5Hgcskh53PikGXFOomMRFikvJ21G7tvAF2blPI54A3pnTOb
ZFHmrhqI1fj7RxWEeXUqh0MYlHTJ5y012C57QiWONwsSzb2fN1UQrksaR+SvUWImiliA8+u64bQQ
OsmxRM2E30l7Q+53gM7ez/oWHReIRViTvyFaUy2mRflCb6y8rdYBViR8iTQxx6OJ3WWdItxUYW19
5Qj69lBIbSH3SQuVJtrx6IR5Rl933Tdlf7CdbS9rY9V8wHT5M0dWIlylQ6wGR6Do3iiajad97I8g
pkAzRDlYU34RN1hKugbZIHltV0t2XCt+UJCk1RmUBvQRlZYv+RXSqbqqqDez7WsMcjppBxWF9zOT
Qtm6poe63zsXaKgBTmWnFE0Nc4D4QuuNlO0F8LGrnN1XJqKw/cXWAyRZqA82vC5k11PO03DXaprI
emmXD5uoxwqFLU++80SI+cMHl3d7WyaLgHsFDLTTt/sW7h/GcU+rqHGDf1bySLSpK1H9hJucuTfr
bI4pVoOLBKyjaAm920ZpoXfEz3Q68SAJOzRRF+R5XNIZWvTQeMffYawCVLlWVIHLZRTQAuGbYezO
Vxl6iRhwnaAD8EDlir0Rv8ili+9cGpQnqK2BPqnzs/nUdateTMChQma9pMCXWG93oS6o8OaTsjgI
HMr1UxQeMazp4WarPMfkaLV3RhvRcXyFqsetTtQbViHErY4ONYEqzqVVcG79gSRQAKYoJVYdxXwc
dMU7ha406EQLpBiAySOBjz4u1uKBE9D433yZa5ClsL1C0+/4KPG46aLUFKdJhSjtan68Azvt1u1V
w9uVx/3GXybl6AiTr/XVVcNqRgSBudrweR8iHIsLpILYblsp7YCCubW4ed8MwXorHFC7vSgaVgPw
+XcY4jeIffmS8SHW/noA/fgyYLICtAkozw9FlaLKgSABoDDOZhl0tO7jrW08oiECO0OaFHLHtJnK
4fV9ZA0o7wPh6QCx5zpu8ecITwixgtYRq7fhQKOrfGvy9w2zWWzGIwQwElli4sTgVojRaRvdce4B
h7IVcKwXpyLx7KQ2e7rulv3ask0xl6BUvu8eK3DqJrJeZ+CDOu45ropkGBRJM2tXpGMt8FdZ4osq
e11TeE8GBL/ofMjdPXW3heVdG1aQBCT1KXFcV/5KaR063x5PCXU2+gpOuCD66zFS/5iP892CGO0V
7bqJp3/vmK5Bjv1zptydnrAU3vIuvxM9jXy8+w2AOlK/9taS/asTNFrytTv2K5QyJdgAtfBKiTjH
f6gysX+I7eWCaHZw7VsSCegsxP3ISVDabg2ESYmtKTMpFQofFuyGS5CEPChXxV7xdLoyLiFbsjIR
2kAKMKbhFMBZImZJdjRm54e9Oh+6iJotMTdJJoXos1jr0jgPJuQjp24OZxL2xtwJQXeLdAe4XrTJ
K+59vzGlTMtzZHf3UY0bZL0ueVHgD1s+KLXIiwqn2sB0g4goqvtReaHLv9jmY8dTX5mYOw8PeFsy
8cwYjKFH5vzg1fAjd8/SIpUJSTF7wstglpciR5QuIHR1oBzz5kFVn1U+aS4bdvjBmli4x15FuhM7
HF3ur6FL1jrBEVgMJ8QZhm349FGMBEqZZBFfgDZpYlAPPtLzzb1HBC0YygUw1cDek4bD7fXs9gIQ
EtMlye+DVlpFDZfIJESVt3Jz4kWNspkrR2ldBnQOQG1PWUmBPIi5lJVP77tfa9kDLVm3KjGM4HtG
QzgVAK4LvzoxXNa4AeiTOiQTfxx5/9Tlk1gtXeh8RzbPoqt3m4pLeTvtgXH5EtCFbSqqR0ZPbsCU
J89c5aKgvyUs3GrEzQZT5wE5210JElOVPsl3vPrbIRLHD9OL5mrCXiOEIWfh+aZ1IFHPT2PrgKXu
271n0Sn/gM69FubHCLcRJuc4EWzuLXFoPB9kUEwL/7yiTQduPqSYSO6mMx1/dSSgCBVmrWue8XjJ
L4faZbrKdYDnGWTD51XOnKLINeC3TBpSo5ymZwWBTioNignh+D1eVCE0cp37aTi1nNpTeIXP1VGG
6AUcLNUO7fLQ31gUcGBwyXOju2gAaOxtR423LJ634DS20Q6f3pYwoaDVz/20zQRHWyUQIeetFfvI
vePW85mfKXzYnLcD0bccFQG+DFePNGqdGe1loDspACQw088B1ibx/OZdlMh1HuQvHy1nG/4RkXXC
Cw+jJkQinRb2V/hgTUdzhqqNDjcvX0Egtl8nuelzGA8M7UTJD4d8bc0YqZ77K0aEsxOH/uLH41mf
y0wcjtldfuCYpQ08iqW8Y5JTCPVcW6X5W4gss+fE/eYGgWZmCGJeMFLpCdfQz/VSIbLY8/NG1xQn
dWR0kliOY1bCc5gAE1UxGaWo/Tmsi8VdHxJXtdrfjs6i9n2sDsuwkI+mpQhAzss+Mb/QVT3WM8cc
3eeEVGYsTPiREZtw1LMFIhUGGGswkcj9nuA4c949LI51/RhCnb+ZjJkWV6o2616/FQVyyN93vn+q
djVXinVudho33hTtpAr1J1rkG+RK9aKxW8TNzhARrHGDxbM2r34pTpEl6VUgp8Xg/NCD3W2xA3hY
vWCf3DCca4nywtB/KqSFEr6XelMD4qVHzPkCF+HfffQOx4b8yQbaVy3Gmzhyu4vsQGDsDyzbmCph
jaokwUeX0ksXGcCL1lJ9Ok6YLAyjAtTBEtMF+qPm1pIRL9/7iV7MHREsLy3BKdgeo28VdUY+/8g0
HlaXCeoNUcyzV87Bj9CSKSlAlnITd99R6vJ/Q64rmwr+NuO6N7sV/fou8C9c7za8KEenEsHZiVwZ
Mi6eKeF/Om7HdwTVhdkXRllU8DbDuvGcAlXf0l43GbUEkT7XaS/Tp05dZM6ZtRYtS5qwheueq1aJ
/DaRs2X22yevJjHkNF0N07QOR6q2TpGDgyk+i3xw/xCpYtSRC9DIQHUKVLtpP2Qu+ThgM0QbufuN
fWi/b0vFMy15LucM+C62qErnTipnTijprgQAr4QyxF7NiixX9UV9P9/4o9ZiVa4RCy7OY5539IrE
LJXCoOr8y498NAdQL0ofWogi16ifp8VWq7V9FgI73YYGCtYZFub57AToo+n3Nj47WTQj8V3zh/8F
Xl4lZUKv8W2Xj4UjSzRXUgsWIOWr5xI6HPdVS2+8z48QTvfzuy3i6PSq1SA98n0PyC2hw2twhVI2
OkFXlMWC/sI++OGnL8fYyRBECEQJ9+cvZv81pMzMjq1DMGV9d01t5ufvGoRjUebKGDEIJ+o3oCj9
U/YcfIYwIp9qZJY1nsEYoNrEemutzbOnue7cjaPMSb+QllELxQtdyGNHMaTx5dsq42aWopGQV+wB
6Y8uc5/8XbWDBN42a5PDCLAWZ+c/Atw0qnyT/wM7HMMXBlkgBt/B7nCZCHAQiSrXJuGjCsU+DlcK
IaOzffcLLa/DduYU5a7k5u4IhwQlKUUlJQNKUcL2LWzmCFzauTp68wnV8TVkNP98PPqkXrGHSZ6E
GEppFUfjZMN75N1+1O/64k58eD2O5igWPTrOemrrnsSO2SP4DVfA5Z7b+fDaSiixkxsoSGDlBDVv
edGEeSvLAXxMhvQGHtD3Laqd+NKghzbmPQi+E2Hstn9z7KCG1noRE7AWm7ZFuiwT1dAiZMsNhtpF
wP/3arLuJdUO8AyTmMerwThgFqmmQbZwhCpBTrSaW0XibP7O6YdHjl62VpTYgwh/gtZ+m7NhwTHz
KYPoVi8TLNvUeszyWoEFk9JVcxtAhplxqbA9w+PDUuJa1Bp17wV2FO/9ULslSjRYM9FjV06f/s3D
gMZEYzAdf8ZKLdCF94MPJ38RpvJy8AiBN4p73KYdmzIiPvfpG+Bfl4O2YQfYYNVfIKC1P34yaSuE
hv+ROSSyixO1EwZivZ8Xd7IbIMebIPkUGP8o6sWiTLN0JczWkKwHKUBsFYuHwXXK++xZu3brSfCq
a6CZXQEapAGN+83EwAVf8/9z9AwmOjlK0KiHSDuolVATK0ON0H/3goev/UMNMBtiCRMl398ZUm3S
ikJ/Xf0XAG6gUmiGZV8ExekxTVU9pfH3ovhSh541eKeH9Fukvz54O4EaxYz3pRGw+iN5IC/Cum84
eSZeUkYO7vwOtrkR2Z+3g1BqZKaToDY5ACP4P0JOJ/jHcCqHSdwb1Q9gkd7YFVqGVhamGtmzFBxG
BNhNBuCvWI1k9qRI7cOTwcIdeZpK3WAUqzl6TyPY/ULBJv9nFQHwTAPOBjmKjUm1/9kXjORGJP0a
Xdl6LMH6YAQew2UbOI8o8RyBVuOGBoj/tRWU59tA3G/InzRbKJYAx/PTGXnxXN1n42/UKI3fNpMx
LYkR8n1yXbBGrL0Na4jmAwXEk6oXUG3HMiMN3cucKNB9d/nl6TJpfmZ4O6Bz77z09oFbV7sU47YB
a59DHlc8lj9i/KOgos84ZRmG96wRtEBF1CwZe9SL7AwzYNmAS+huNApw24BTYAvtdMOBeKDpFfgB
ckIf3zCB8QPrASalajAXrSRS3KgED62aFGVUu28P/RT+qdJ3zXdBsHzgZGmHYDZjM79SCHSgr4s1
jpJD2YLcS7UH+G7DNWtYnk4oNAFVNwUhvaF4ODCFex9PXbulb21WceNp5eFx5jn7ihAClkTULtH3
LmkYVAX8cL9p5WgaqoI0VPJ/59fDuyyxkBk7OQrZHAjcGN0V5K+9FRomu1OLrIZSLLyVpbJAzJT9
Yk6scOGr11RkGQGzxK7JjWFSlS3m2hHj+br5mqZ7DaWQddpK+T2I7a+Gf6sQFLbSCMpB7fQYt8pi
Nn3CV+4yWShcBu8vwV3GPI0G3t8GtbZ/2Ot2KJ8ojFG/5Ef7HIUrSYi56mO62YUiVjqYpBP8x3dE
zvuZ0AxK2OEKOT4BypzTQAlCeqyvRqoynwv3z0agsV04M76lXssYmaEBERHRgOAyoj3EkDx5omm9
oIcoqF1Z4BESW6jSGX0S1U6tMwkb3L+WPN0HE/nl5QqmWOuA8iTk0Fb5SPw7dJER5PofOqy3GBIw
f0tVV3HIH6znACnKJLc/QBcANRjmf0W2HP2LmO8/9pw4Sz/tBa0tfa6J90c7LkcJ3+O2CjSb4W7m
js1fDL6L4yaqtaa1BEwejfdQ3kTC5EO0hgY+nqqgEs5NAczdLlbsrKQKU4yt8TU/+/lPWEb1Grcm
ZM208V/QC7rJOWYCtA1OCGWZVhQzd4YgKQeVFz7J7Z2zfZOM/tA6xZJwIS2X/xilB+CtI+lNjgRc
gHjNDy64YHbahvVZDfMnyqQveff05La0c4M9T51joHoySqmKnQ+3/uG2u2i3V6Zv/mVPFWXTFya7
bz+XUg+cLpBRqx7Owc+LHHnVYPWsJPn+hZyEb1pBHwwr3TtljsRAs8m8FgE8ovOlf2RqCf0cJAk6
qRiKMK6G65ee8pmbPU/iv5Y56RB2l24GW4o6zyGoXZVXbsJsAY6bc0RRze1/AjtFSGbnUSmpDWYy
EENYUbje4GbN0YVBEJ4w44ipfVtaHcO3PhUtir5pnytOvJcLPMHpCd2pztg2QSSvzWTKRMiytKYF
/Jh/vkouQ+DLdX9BO5KDKSPSkiEiCoROAIRv5pW/s1DPTSjZJP2EP8DRmJfM44U15M98tYp5m2NQ
Rl04y68okezElZp6ud/eO04XdlQdieBjZG/5HkSuxEnTao7yIEWFGrVgWKxEuEzrBYMpJu80TA9X
Qr0swXqEl4wIXSC8J5UFx0DR7enUQSSZubVWd0VPygUJGh81wn1Pd7r33OAkCR4M6skZD+lScFNg
KN3H3QOHPZ/IRmNZ5KlrmBWxKo/T5IAdUsexf1UKi+gCAWMbdM4xWchb6O/PbiSYwXRGVeZ4Fcds
OUVG9rHSaTCHy3NoMifzyEfgAU//XoclC6amVtMlR6kWAr4P4gWHsYoJSj8fCRTR+fmJboPKwtbV
bYc86depX1V1jGbOvm0unN2LX3PFdK2QJkTmw+1EviZCc0laRHJPl8DxwTP4fKIfGhX9NexCXnd7
p5XuLm8+yjBtpbndfTzBNS/06qWAqg41422Sh5KRhg+tejGzkgX2SbUIo8/bSMLZtTnfeG0NwOY5
YTEPeZsTH4PS8gu/JqItfovTZ4dShKnmJnn1KvB9GjGoUfTN+zpTXZpEVoXQyOm7D+K5gyUAQW1r
7mg2v7QL4+ZTNhPPddajPmXpOVOjpaPunqlGNgNrZwSvkp3BrgwT6et/dfblHxTca5uwTmnekcgX
2UAUEHPePiONkuejycKVuyfbVjXqq2WAsUG/hJyj2OK6pePvUEasDoYRgaUTkBf75+ZlLMDfGpo8
yynmJnHjDe1ieO4d5F7Ro/qPQyUefPAXSHVEO/qTqfVUcjsk8j6EBX2TVxVr6Myv9WUZ1YCXvBbv
ZIPLkPjGuNnr5DL6mvBV8E2MaapS9zMJG/Wb/NMCHoPugwER7jb0rjV7dmYvMaI3KYqJ8frRCXFb
Y2UaFOP+Y/cfRS1lOUyLE5z2+h2JG7uc4+HL5jEtB4CF5AG2gIX39P4XozUj7vkWjiLaYsa58nFp
tzITV9p5+o90w87YhcVAIqoijdKA8TjuoSLCXcbi3gVOsmui0b4eFMbImN3UCXJYDIeXegRIs6f3
BD3+PXKnHTBhR9GdHUAzVfCF5HE8+X4XcNWwiaSMkUDXu0ibV6yiLzT2NwKjpL7zdnj8Ps6b7UzG
lXkPKkCaXgycbD3p96hpB5HirnNGDAkxrx+Xtfo+eGZRM76EhmvhJqPC+qrNoSsHhViUQuXrfLIi
9Xwg/wadybJaFFx6bx3NBbdjcrwtPjMnH6PYhFG2IuKDFOy7TRqIqsHLr5eJ7F8AgnuJD1kLNig/
lJJiOd00OECmTlCX2/UpFoIm7x1bBzh/XXOfoqw8veWJFbLyRRIgkr0QWx+DiNDN65solSplzSiL
9wRv1tIZkWoYZzSYUn5sJ40qc6dLfi+LO9Z/ld8ToU0BUMUfNruprMIoAlz/1VO2pRC7G9pyERy7
JkblMlF5sVuca9Mu6A9JQ9iH77+dXUhgaBDGTYNaltemdFB8WJMolFngRx1s5MhmOPNrv3JVWPaN
+kXZU52/iT/dWtSMAAn2+BinO98nZUXE77WdmF9pmx6BxRCqkfQN9cNRDgw0R/c/3quJ7KOfy6lG
lpddQcFLgpObUa9VLr1tEswhDq+FldrwjUJK1eoy8TOv2XQfFudo9ktz866AMnkvyVF1QE4J23Jy
CtdOkeR3mWguU2Q5RLWn5mhf+cU1JI0f6+8sJJpuXu65bpVU92MbJFF2oz1CIGykYeuYCHLz0TGD
7bV93VosXI658aAqvgNqMwNxa5vXu97zOUD/hYj7sj3Qz+LfM4KftzEiLm3kwb/al0e2QVYUuljd
nez34CCLy4LocKYz1ZN34WaV2UgPS2m5h8PqZnt1d8qnF+3CkZP7c1xaXtt4Y1Cir3KUrA2gVzq5
L5LIgpni339YQpOGFWSu1T31TL+twxMvgWOlulDBaX1+MNfwZMW1Ak/ZELkYUvtaHkoXPcsocgWk
KAsmYxR05/TI6u+WkhzVC3cbiD5IRXw7vq0Nz4r06YYxLsqDmdP0soD2F4sAVcqE+qvKDJmU/LEj
xyLmBEW0Kef/xPJgZ49L3PKIivI2Cn09++UA7TYePfPRpaiHR1n2KLGKtHmdSdVdp1HLy/ifef58
kEjPomPamxeYoa2MxMcwpRCf61yihD0yv2xI3mI4fFHOoHeyL7X+Zmffur0NtRKsR5Z98Izn1IS9
OSrdivJBZ3tqv0nsHmN5DVQ8tKn4HaTi0tRKT8AsEeFcqtbRbkqbItlO602Hu6BoC0cy8wQ38NP5
uo2amLNmegPGVdI3OAfYkdA+yls6SPmdNx3VW0L2XtT4ObZPsx2NcSXyEz+XEeojhyxg6iJdXiiC
areauEiwWNipe8GDkYtftjdBs7120OiUnnR/ClQ/CVbe5nxX+4wj2VIYCOIe9exPKUgVyII9EgPp
IOKSD1ZmDBa40ika6t9qzfvdkyW8ySljhuI5k2R9nwZeCRy5PITcipI42EWbLW6kEpLu83UX71KT
phojbzasq2OXSYovZkeIU92vhofM6VM/mhUr2x+/PyQ21omPr9r8l31QSGN/B992gbRMawqQEzf5
vrmYisxn9BGoIbXupsND8Z8jGqpzzo8cZqML7BIC0GxAkZHt7OmIjaSTGmZjoVaSRqV3yBxL6DiU
BXglMvTiEwxIiOSvBY9MJ/d8TxloKm+ZyCiAhWV8XV/CAoQrhyXBzKYTQp4w7beU4vOS3OU194cd
NhGqM/t2aSL/RC47n/z60AgBVMOvtIgNN2zbkoFb9aoR7olL9G2S1HA9eieIeFw6hx64Rli1/qYz
vJI7nuffkA64kXllu6DMR0LQKvPUBApxkr8KZcJeJBl8aktidnbw6TcVNG3DTBU/hTsrDIMQCwg+
oQa2BHdpXk8FO7H3Pqbthde619gtkUayz5AMwz4VXE/9BYa1UQOVtLYF/IidqJx57IjH9zVqpY8F
6oi+4t+EIunAYNo1Mdoc8Y95XZvZjjgowtXJ+KRDEW94aSRrs3XlVXHMJ/AQGtvNAoniNckQ5MFG
v4Pube10qneA5nNPGjYutJ6+QNVxOZ7Lsh+mwdRw3AN/Y6NkUlu86UY59STHsrQReepJNvcx8Yuw
B0vJB8FWrn/hs4NS5zeXICgNW4ndsziWfD53yugltJE7VyhB9OAihE777Jnz1MHwaOq398xsnI5t
eLm+0gGMtwwImI+yu034esJ6VSSXC2xf5BjZm8X+jHunGmwYgA1wGnQXMKSNej2JzeDsRZA1le9Y
SI13MneiqfTHUyz/YCh5BI8sT/cNcTxN2I0H1zj/Z/4yr9EBn+tfPA6lz1kyAA59sGktdUakjROA
NiyN16wwc27YndNXOADjoXufjRzNmW5rsRtTADoTUveKORQrVMG2m/wVA/f6PqIIKhNAKQT1hQQZ
gZ4DMhjukOtNv0ZopoCI1wT+EFs6rJKy0kLv4Q2rzDq2Lr2vL9WwTM8k9trdpkn22YR5MwdUB+XQ
ocYcZjEARHqDLeLTOglMM1aONdGTzcKc2nlDXFlfS58iKByQ01lfRgxVkkpspDvwYVhM5xHnpv3l
mtr7hb0mq+N5GswLMilH38VHRq+3tx4g2pIL1vf9tSS+1tvUIxNbWjcyV1Q9noRzM3JomguxDyAC
pxF43/zISE5WQCfO/1YXm2pJy/wlBH9zvGdGY/Uk8yfUZR+thdKcnUo4oJtu6hCqs5aiwBSaPt34
KlD27ZVW7Tvy4j2bglYB6HrDvfrrPyKIe1r4ULsprOBxpnMqDxKb/teTc2sa+n/ZG05LakNkYGmE
IlzZ+8lWyWw7IsTZUaaFLeDJzNW6JutQig0m890etbxyhgEZLyYh/GQa0uxAaprh3Q1Nhv1HfX/t
JqIZUHSQPmVw/AP4zbDPdELokvHdwXOnrL7SPXW7qL0wPQLvMdf9lmowdma+YaOmCN5sDXgzogui
RyGngdUawNwSRdb3NQGn5HSEvBxyYIPhnUPvcKjrIt2ijcrahmdINx7z5c1tyfKtvmF8YNpNU8Pt
7AqUzgA9PhiXUx5TQBVlYTJkqqJ1kjTVxFV307i053WKOiqDMAxH5PQyGN9Pc7pY0+yIrkvH7VbX
rYRYa/lx2ApyX5J8ZBq+dI5tlcsiB920ox6WzWrOjeJ79jLwCqY1ka3NzOmXGY3VxhDauZvaAhYN
B+7B3qq6Wyu3wcUjUZaneIG57XyxvV+r0m2gYGYvNB+gyIo/ns8tsk05vbaZ0sFmHCIpgiO8jIyy
t/Ef4oH72FqrLMLAnEhyWXmzYXhj6FKRT8ncwIeubYmzbwmjhYyT3zv1VKW52DXeHuvS5LBSsyh8
c6f80AnfSn+a5qeGKwrjKcXBvAZTm09kq7sasrI59qCNWDJQ34nJReAFhqvIlivSo+lNBMw9e/YX
wjvAkMfxOYV+/mPgksL76YQUw18z3YmiBULjHIr1RBYEkCa13RH/MPwcPe9nLuypZB1Dleeamt74
3la2gjQLN1p6NgaH2jnGkVZRIkuY7/Glrut4GIMwE4Xp8dFdAKwpjFYM13NUolfRZxHH1KruI73c
EWXz/qUlwRlQdTFBi5rRqQoIHrF4EPyoFVY2VVCwB5mWnzgybYlRkiUxKsUEAPFQz4/uO8cNmEjT
Q1HihSUGc/3M0xTr9tE5g2/mgYY/zzTRR669AYtke78LnRjh+BPhIpx2DHJgUEVkgEU6UnMu8hqc
TA81qvDB/zsREGn/GVP6H0Wsh6DtRgFs967mpBnAmw46/BivuxKmqY7KwrnEc+7FZgU4TV6Y+8Te
GQdZQ5TylhQgDZCsnIA9W9I43HRB1n/RakYXVKqGqkaieUzLBOXH3D+BU7o8Cv4txbDzSAT+zBLm
CqEMDE8oHDSc09J8H2qA9nOC0K+aoXzkYwj0RnfXXFISsbKSgCEp3Nsqo1UpcdeO1oZezpkl+e3v
1fTfgNrf7N0s85d3uBsBLNfEbhKbMtQ8KGT+50Bi27gXERwQSLrmQJNxfAwU1v6bD2cvbdeMLQnP
QP+JaSxghu/KfmFoek1RNBkecSrcYx1jU1vshXvARkc59I8ei8KT854FZxZlt45Usy1tSAHGy3Wb
BGbVRwQva+byoVxgjqUFrQJ7q+lvSgQlRYmELPoKwp/hv/wZeiz5QDpN0sXYnK8ylzmFpCFsS/tu
WOD5Ghr1D5rHvLVGXPgjNXNQk2k+SiDg5mdhc1nXDEbgvbTEQyODul41TqWlkA78ZeVGppI7TxTX
19mgRHHae+P/TAlSTxfEO7QSfssrKmW3I2UeZ+zXN9twisfH0q+jzRb02OIFXMkapQsWei0F+jYD
jVfY3DIh7aVG8duLGetUwguO3Y6YUpX920LHcEG9kKjadZmpFAYY/AL+3PvcVN6GXJjSi317FutJ
BW6RPJ/VmhDozKhrTReal95e4TohSOjtgOEk48e8PbTky1BxbawUVDdEmBDoALMG/rhQirmW2rph
EszqETyehAxzNFd8Lp+X9V3lti2v9AvAy271yUYA2hznEkmFq300MkWaM2nQZgkuRslmqJibjsCy
1ehOqC4LVL7MnmZZ8aJ37Tk0CRGQ5VMDLB02jIiPy51YHQ/Xe5H6/rwKQ/77SS2Umw7dES6xML9u
zQSOVtQhQ20u2n6e3xW3GNQSmIJvn1gFKnMjNg1E403WPrUs//kdUmzP2VUWhKmGK7ilvwCeJgjN
YfA4AwBQbCuWebeALYxKmtv9gQX3UB0HJp0/0rc7HbXNvplDZwLWtg6Ld3VjGy5bqjEB0RtLHLhZ
wzwdgaFxO3ML8VfJv2DUVGt06MpflDXbFZ1ryH3ff1caB8doUl0hg+37AU0K7RwQCRnvhNdWmJw6
W537E3ZYjdm7sEGOe5D6fWx4I0CBcKTNylm5JoUYzkS+JGxkMNHw5URYdijH6RfE48QjcOQwHEq/
Uix5x+fBXgm4GFOXRB9zXRYPLPT3wDKb9K24w54IM8fc+bhPM8hBLcNmeQPh9njg1WlVRcBiq2W1
DyOry3pl2CEe+Is4GL/pn7D6tsROjioxRlAmrappKryK8K9ffy1Rwhmw/R6dqwx5JzyCuwNhnjyn
ysuMqGYSRwTCBPZKvlIFpiIXoAnNvkkz5BWiWFZZmpxtweltYYqLC5P7IBoZgIaH8FCmGdTt+/L+
6G1RqdwyPlg3/sKOhKQlZgS2OiwgTsqel/dpHJ8kFyiZz01g6jlbnfq/mC3g+EJFsEwv8Ai3CfPX
DUMZ48AZwcMWpZ2kEEGr56pOcruNUEZf8qfMKIzXkjASJDnAZRSgbulRqi8ZicL7/pYBkzHXd8eh
pbjCUAtVrSPBtBH0Dbx0Vl3jWjKDo5hVGBvugQfVIrSY2ER2L5qiSdD1xbxSf4Re/1UXygxps64U
r3kenu8IpBoz0IckSvBRaJS/Jtu1hteeKoHuvZv4zC09BG9crqkUYdFM3sGdyd5ci5aiPQfogpLx
DVrTP4pM6hNDJUOB1mgdam1BQzDDzOR20ma+6ZC4nKlQQ4WQTMWB3EGtTciWz62sJRdL6d2uzn7/
HSGmkL1iEiwXtdCVeDOSjoHwHWKd0S3sqVROtBcTzgAGFs5Jpt2ONzvHGJZJz4690WPE09ib+WoL
akoQSeEPQ37YSMjlcjkVx0AWvQSjj4J+V5FJiuodz3gQNMjUJk8AaFdISfH93ml+8nIxC0GGp6TO
pnbf9mzzTLO4KZoAUC10L7XWqK18qNeN35fFDa/g3W7/YLsqd7OB4wKjFed8MLjpo0TqxWy+n47G
unuSv5ZgN7mSz7ETsQFDi4QFeM251jbPAFDS2jw1lNDf/5sbr2+Pk9nPN3FXWm86Uc/ZW7uK++u2
hpGUPxy5ugpWDqOagnENDbgL2tAaKtBVJ8PEJHkMx7vbKbvwzTGu2e6WR6IDDL6eHw6TYPQMu6sG
zupmtYXCJX3A6VZjnL9AAPboaFfQuzE3XgHD04HFioctBVE2o7vvSPPNgEmqqahAvT/u8XfbIvWA
6m1jA91YH37QDFSXDoBKREMdXP2X6LsMCTWd9m+iYiaA3JYZMpiS9QERlFMQWZoAC4GDnjb61UmA
jO2SxsFu7OVZN+tykKGJXpCNwEqvMu63ArP6gArCf4yFEEfAL4b66/YbVdKJJ+SfSJSK7O8vkISe
dEMLgEG6eHxKPdWoTYdLVeVbgVFFJOmDzV/D/bo/SbapCEaFG2OhbyT9QWKyX1dxNNwIkRC3bAti
6G2CXMp9ftt8x1DFpVNIOfkoraWdeJoOJGz3uKoelLyqCjyodtFfJcLb5K/Ua5ph/xhWR9Cj6fer
NcmQI12M8tMbkhdTj2AUl+P5/fyXxg3eKlBSf6XpMm+Lk1Ofoxiz9cPAk/KtJ7wC0tbg1FVh8X7w
BMr0dLnyVH0+zFiA1snV5qfcxF6/OX6SItS8hI1WqsWR1bTeH8au5Z38TWuohp+5q1amoefATdri
JSVJRUsmLTO2OqiT1F7G6NH4xv+B1ibQkftn7iPsXZF4YMy7mX/rc+XA9pja+woG4P8pjA+cRZzc
cHHs9sdKP7FjF3/PsKn+gKUtATQwo+nwkZhFfp3xZJ064QzUxZty8I1wn+dOdv4P1D428svOyziY
Cq31DPKxX/Ekj2p+GrHLORNDUwAEDwSttVmf1YffxYsZrhTeYp42mAoZ4KSKVOQ01F3UI0lsklxU
aVp+VOZXd6Qg6YebIT6Ak6lPVMNAoS4d4mlrkEw9hU2Vf801pXSq11oQI4UKCu9v2Zo62OzvEunT
6liwOtS2IK5wIX1QJLmYcvpnovn3XFQCSG05f1sXmcbCLr6g/V93ZK657WzSFsxuti+RZuWKQzl8
h1AqsWAo36Kr17yMvHpkgJEUVTgiMLfhyIAHwkgzCmW39kDaVEkHE6lvWrg3sxqU836kd46SfGh7
VCuPOA+fhO+K8djVGMTtNYKvKIVRg7ef+JOs49wXPSQCGKs8W+74t7P/PGsiFK/rlzXLwHRkB69Z
zT5IJQF9nDp+yFHPa7I4gmX90cZn73dmVcuDoRbWrQsm9v2C5XGjSBlUsTfacbLlpJNghB3lUkmr
q6gjtlBpr1K1jkBClKwrSSS3prkbm1/DngN7q5IuQJfxALZryL1KDu9ko0pHtNJs9dcvg/aq7gy7
b9YLj8pG8CA574iidWwcSxHSjApyFWQ140XnTc6+FTXsWgxD2iMkzkjAG2mWmH6Lo3JH7sFPzRNW
ZpwqQEdjfRJgn8Ovvrj1PrQVVK+nJtcfElhOSyScEWZ/cbCdqDtDDeRWOZIhba1F8tBNF7o54Qch
IWB5MQXwmMOVZ+VwLO/lLKMwhgyuQ2d00X0Ea5ak4LZ/NyzAezbOVxkXXu42r4md1MSbE0JbpeSS
qYMIxaLGqVMqAk+hQinmxelAr32GBdG3wcwK6euf/b9nZccmXOhtjjR1ookAzu72iT0BQGJTg67H
RjF4fi1U90gwxiYqseuwX0MWseYeVvUJPNTslyYlAnPRvqq1YhVOfczYiP5IKOudBwUcHtWgt3vm
ndtLvV3mDjKQ4qbnCvfUw2lqf9nLFlfGEdmH3RGRal+1Ip3+1cI0nGMs39czh/ZcgwpHImq5mBuu
z9l739uDeiRHqz+k+6K1ilux2MpBAcnXVtSid37EjracGHI/EXw8leK0V7bQe8AWo5hh11ARUDpz
Jtf9Nxiaz/8ewJ/Mb8ibi50JOJgGbBMkSHSLtGfVpJsQXFDlPLYtpf7YxBWjw+oT5lyFq3YeII/C
cplU7vbU+rg5y9GZoTsr4hV2A5tdEBud7pf/CDaJPhkfPuUNtFn5WMccJ9qg0ziAgvN2EDVQiKjj
adYVyYpArDQXQsD2GwIuWJPdCMy5yzdDKwa8b30oyd0iPgDF9tim2WU4JVQiwqzFY3npGJNVRH1Z
asawNTO0tBjMzkuSOCCSqBibEI06CIEtNJtgPDVwvq7iRV0kRmoOhFOwI8m3FbcRyFknQPd1gAYC
jGstOA9l6G04ASCrZbIPs4ck6rHmp0eqXLsJUZodbkDEWxaBkg5gcwQ9kPj76o3aCrtnwHTAmRDU
HEvKBnezqKgCVoigwgszhPblNMrWX2/9mZjgEj5LG5Q68Qd5loN9AXN82rKyyu0c0EYN7mGKl56V
mCI3bblJ9dSWbhdVo3fgFe2pfmCQw8oQbAPYTF0ZolBs+IqZt7v6pNRtQTN+KzHpw/sV+EdJM+9J
CgJ2AJfI/eIAAwh0EX5oPKBc6Fm36nzNH2VbjBK0cgPJxme6bAikW0sTGV7J62MYf/uy+qdkQbsZ
MchMELxxRVyRv7l5X6cC1Q12zvl3DfZ5jZf0yR4mmAZ40w47WUTvZUR4KYjaidfbtZydK22DgLeo
1hoIGay0PbOJcmgbHC5//bzDgjTjhq7MZvo6fnAvqF5inEMf2yL5GSQ0gracidxrl+mYErLxUZri
rWEzJpzosD1y7052q6ytd2NrdQhqBwm7ixUl+NnKpSroUYgoj8ussjOx+inzg64P1M4y87w8B2FE
haYQ6vl8YlG35lj0Ns3wM8kEY6tRIdXqKPbs1b36gXH/WiJ43EOYi+ExZ/KENA35rVjnAY9VZ4qo
mqIM/VudATUK4T3C02AW4dteidBLAcfwLyhAIv4AhGANf8zY1QXjB3k+elioi4nOoaEumNsg87Er
Qt4F4bgVi/w0bv1X/VePug1GcIr31YNYhBZErzbU2kmVx6iL0eITgi2Q6b/I+GWiZ8iVQoSf8WF8
gajCQ6TZEP4b3rR/imXlEe9p6hJ4eb7xvipwokUW3gUc3T/uHayoy+PtH60Yip91HO9V4gC9tZTO
d0DXKS7t25lEQ6eQlBIeLAhGYZrdr1Yr53SaSTdOf0MN5RHTU9o/9X0I/tTMejNX7Gw3Dho6nVui
pHfMIhZr8qG36Ph4pHakI17QIh3pkExv3kv9+WMHI1l28iQhCMgkAjSs+M02zzVdZb/WrEirhzv5
sJxcgcx7ZiiQtfAXUS/grGnARMImwj3z5ZgVD5alkzDuZnSore2nhbBT0vBGJbYHGASi6l3yLVCB
xFa+l+C75v9B6185inXNSSRbpG5354pN1B2MJVCrc2APCrcs/3/Sivx4XiUq4neefnDVABF5WDw5
A4tOkmb5IOMWTogsFIq99qnV1jkjaeMfzTTUFSxziOH/DUDLKY9h4Aus6hjO0KMJHUkJiTmGPRJm
SYPqN1lzbmym2+ZaSNWy1n1gbXntFcNrA+P7Gsv4PiJjMUPD0oHNqUp8E5ZMh/GiAvKDr+s3A02G
hPDsQMgbHDa2tmqjq2QAKYJW01CfL1cMlx6Zqr0b4ngt4htHfl0KZDddSrsittW2XCS58Gvd+Wb5
AJImOrTqaLhyIF9oSfaamgs+pwYBMVGUEIFvhMk7cQZUJfVAHojYNiF8HXocNRvEO3v3MXnMDbJN
F3YD6n4vJuYkm56BO6FyazgC1al93TWpx7PLAjmyfiwHmm+sF+OmmxWREtwisL+81kWwmVia4VOO
DcSOSCS6B/97OjO9WFJHoG75usRfb40BKrm3EWbKWnJf0TCnYBRTPytt6KvMHYjl1p5fdUmuHsM5
SAMmUqj+ixiQe0N023fOfbPR1PqutDFxxlMJucjYoRZIA178tQWPLRLVgCQzB6xNZ8t8MrOrkitR
kYmwYw6REq72bB93Ear4pULqIqo/TfwNfuenvQiKunNw4MznKgLQTrgxveiLQUumyky26wLKyA/t
pqak9cxj/aV7lQjnWiIWY5mIhwgA3Ha3FGQn8fxXp3IDT317eoSZe1zpsdUyB8iTx9N9agRrPzhO
QewpbiqD/xg8xR2Gjlm5Nc5UoD0XXtQAwDx/3iReNJL3pnt1lOc4PniE9P/7WEYonFjM5YiH9poj
BZ5VHEwYX8sxP86C2Nz9dY5BRVW1qIhY3KXhDUpWZEBeo/mi0EYbDNT0E+55FBGUquljiXAiKvIq
Mv66WgWq4h5B1eHdoaQ9KIKgqRwCtrL0khD2cc5XappoKoywe5PpWEYjmTOEKDunvyheZ9GANADD
FoUueYSgMZ7eYb7JGQLRbz+JTlYh/0HVEmx2e3wmw1o9n94WdnF7cvygRVqeXboe0iNY9FMAjJ7s
e4uB0C+al1cAppp65TeFm9GEcpXXsX/hpu9Yj0zTlkkj44P9EsQDVzSzVWrBFBUMuPiq9skMPPQX
OXW5Mk/cIfIWD7GcZecqHMb4nuRuMRwZCCnVwneNxNmRW2v4iSv/i1LXKPJ7SGHyAC4J9npkdieH
6/FrTlSn5atI8xXnz4N0arH92GkNuc+65z1F4l4rlxVS6zxxEkw2GBnxLTFrhh118Dtfoy+PdV7h
IoUy+y1VkABLYh790gz1PeTruB8BqIESbj+RmVJRyHF956L/9GZtD97qUL3F0XUS17feOMqruxPg
XZN7s7mqc+cSLzmFbcl7GyuZG0x8TLBGZuN4Z1x3mbi7QxiYcgEc771GR7zc26F/hWdYrf2AiKF5
Cl/nNs0jEoPf2BfsesMakVUwX8UtXEIOv90LtU55wiEJ2LCTWDntT8Qso37k+9FpkTnAJtgGnFMj
I76DrEi/3UFxKlR5JDPznkO2vfc4jgssnB4uPB8aeB/m0OCHH5QatAJFosAlxnnf9BHZ1TtZdqQZ
3YyUxCv0NDMKf43sGHaeCDrHu6l+rQqdmoVARHLFDTY91D8dC1MdEWBeB133WzDeGo3vLqX0eLn3
KCJC0QryeAYDA2RjfxEDVykKosqh+Siu+2ysSYBJHshO/FkcI1k30VG1ksq9ZTXkoBxlMlLiF9MK
UZcM9B7nnL0AJPXLMeHuqIG+NI3ZgVV1VYtwTcQKaZvbYOHsawExMb0SH/UkeNHJmYGc6Nb8Z+eH
QlqzB0D3pXE/QrouYmwp2PHP5+5MHl9pzYwWiyXBSY6pM4/ZWtWPI8kJaehDswZYaIJoe4fixtKZ
zaF22JNxF15KkGIY8pkcLVIhHFqlmBwU+TnxBHXfznSjXb1D3ZJax5YkUwZbDnVNyWRvgzK2Wofs
Exv5Fd4I7W2JDh5HyieO0n9EL3d3GyV4dC/Judym4AMqzFonR74fpmgj4MAMWWMLj4KR85xRKybJ
jXoiLcNKwIko3LR7XcbJ+RM+8AMD2JvNlfjwB+Ok2wlPjNODWx9dWYYaS8v8ZN2/opj1c7pEMXeh
MwEYEQzyx6g45DjPldRmVHpeBxu9NdWcYPevW9ux3u6fLXFnWOC46ukGHyOIO57kyjyKb5L8BWen
P0CgBDkQRWWr6fJvRymYjJdDHASUyuvVYwN1Rwx53VIHMOWhhI0A4ifXEBW19cVcfMrVF3jSDoTN
Y2OakpmbnCmPncWwbMr4AWw4lqz91UMMrZrPDA+ZQRatnEeQ9pYzBSJ/YzXUeTvRhuZRsY+cTlHo
FtiHvbmRckLiZwDuBVkNZxaUHuirPLV2xQabCs9kVvy/QCr4TvypyPUInKxQoW1ovZ8kgXvhikn8
35TKZvhOnFfo/BeB6KrZJodmdsJDStVvgtUp1BaOdgQ4blXg/5zt/6fx7vnwPuVXR/cH00i8WTY8
VUo3rHr313UH1Fl5BPEYRJgOowpzZFGJujkJYjaPi1+bLkaiA6Rgd3LswAu4pnLUvACKM1QV0Ma5
2CgTx+UvcSAfiDNcbr2hpSdHptWvxD0vTnJudr4UNK+5N5ycFUoAlwXYplz4GpmflFWsLSEGZ239
AjedhibxfFfiM2KcgbDLcDyGKXfUdrLoj1r+Rtf1bMhGhmtKS01nKy3XbcldIe+HZxB2Vf0r4m59
/cXGWx059aTOgDJyikXR54oSdKKIMJcUP6w2OxvR3q1U2Yv/ad/fu5K8PilKir9UruDKK6T2VqhK
ov7tVdwpbemtyxP7rxMmpAEQGIQjhIfHhUculRuQuKPoqDA/kOhXghbKnonQyZb2/ezY8XEjjKAu
+NEvC6D5l9p6eD/x22ldHxr7vOeQtYESX8y5ZRoGiqiWuIn1kQLwho0seHAEUPvNQksxBv55iNn7
RZytVv5i349XdsnItYX5B+OFtnIPmX39VztPSic8j2GeQB52SMMO5KZyu7jswGSlwkfA0Nu06nO/
nqbk85lOxXzYoWGCfFjjB3OBmFrCHllYxxSjzn6NpYfrrBo5jv1vQLrZdVfjP9KN7wg4QqmpnW9G
CA5i8Zy5V2q3TKpZ9eRiGUuYsn6wvRqae4r447NziK/NkmR6xGf1jQ7X67VDcIpm0+TjF7CXGJTa
RxBXUnqwzd9ppd1XRdLvwBKUdmR2UKxhtF4w1gDerhAOnfAQyoqkmPMrg3L59KzqxpRKTSsXjwRD
lgWs9YUpyhr/eOhkCL4tLHMMEDinUzPs2YzK7uFmz3uPJMNUIg1RAZKPE8jERW8dt+rvYqdokCMJ
Sy7CU4PUOeNyUbL3umrc+o5DskVROJCxwtMsXLlycnQkhHX3IdPYTRRMTn8yHFGQxHJHMfj73vdz
5ZtJ2v5SSX7qNBzBKQdzn+mTmiV7/na/NbR21X5r6GMjcrwtzNQN8mh3sZIrW7Ok7Nj4wwplUNtv
eH83hOt/l5Zu93QhsMBSuXfyJe+jw2Uy5mPR37gEzrsL2/pXUbgbMjAIOSEtYQ1IWLGiHPJcAD32
b+MdHrHjIo5G19NLFTnxGoUIZcO2sRWQfPWKedw//L5igcQ9/samGNNDWfd4ucygMdkWd6cauNTM
NQEDsF8sFY534Y86ml6L9+axpFoUtm8f+rlm8BR92Jg7esMzTdUQufqJ0nEM93VUGe8k0tvFTEIJ
V3p1zHdfUnl/4HcypyliQxjGFnoJPcfIoCYraHnXVJYbRr/VC4l3YMTwYSosMS1dLdbE/CTJ8F1K
VifoO2y1vJsdMo2WeFNA9y9+iJyr93lPZmRT2TZFMQivmjxOZqFbHzC5EW8SemBdEVZ+IacaYQc+
RaxrMIrcyzMIkFuye7+F8ZQuIQjzOvNtuk97shOtzJIxV0RIjjLcU2zI0koVdpzd4vhsf56YHocJ
xVTlpHhimh9J0eHOV146E/hru13zAMlucUOHu8nOzXaIQoRUKZDsf0ZTLDuY7bTsRUSfohUiCwOl
VI6rMQOgyH9vkxckxdyVqZb3ku2m70DECMj/hvq+VTJj/0GCuX1rS+QwuLwTzSpSOkFCWSb8NfU0
CJR6QqalpdNpZA+2K5+48U6p/wtWwsomcxEmvY7xdKoE2HvY6KyM/OfTuaOgP+6tC1o9SPNp+zXp
7no4ar4WAMKZvuvToP0ITmTFQM+gdFQEq4B2axqU1XNyRTcWlmd6J0ond9ASfi1EmP/CKYZ3PckX
RXxzMbiwrT1b9XSHtLYUfoAAzQZz/4lkPVLol8taN95WrjzSWoTWPpqrEPbUWwJFw9I9O+C5lsY2
avqCE1L1Ytncf8Xse5/+JDKKI/926CW3cWKPdF3KrUxAXmaa6XGkj+r01JAtldN1uN/WELcX+5il
IDG8HgX0wz0zWRi3ioCB985FkF0xD+EZlbw0IYStDixd0dDtI+Nsunakr1eLI5DI4RQC48duKH7S
Eh8xg+i8RWvUtRgfLdRWAPrFv3ZYeAYk585JTTE+Sp0gftdo1FtCaEn0r0qAo27oC+sfvk3urQhv
96Q3llDRmmycyQiNiXRAltQ2dO71fmkOgWONqZkrp1oN9n/6Qzqs1vvfp6sWggSCaAZUWV1nrN+C
7Rz1bydk+sCVJ6mJPhKnXp6i8qMOFmKXJGEJzVGHbHUTSsSePpWgywlnZbuXf8VspYnwCskMkpOl
QdJgN6QOe9dKuJGQ96x5VtPALCfStf3+jpUlDAw8cs+nsVKJ3jxwoTCLKOBw6erHPUFLrNZa+qTG
Ux+cxKj05gjYZO5UPHxrwJh0cyVwZKmcW1LYJCOhLGiEJC0E6itL+wlJpnCGkcljLYRcS3RbYdVD
1W+BaUqB8WFZs0sz1Gl0i+GO8kLE1FZh8BI3IMKQZZmEyh8ecqVBjubZeqp3MAiom726+qok+i2Z
b7HC1CMGMgCBg8jiRk5LjCGieb+4mRWiHsnSkq6jcGH19miOdbKBjpi1/OmdqdgGdiwslUlfJ3dw
deemhxATc4B7LbFLz60CJByl1kWN3ep7u84taA2tRH4+hczR/XNPZL51NBsLNSQDGPvBdwd246LN
SMG8y4XypV+ivI/sZIWHWBSer4QdN3RYmmED6hdM1d2R1Z8NbSZZe9Q5uKbz0QHVwnBzlwATpS/o
jI0IgZvK1YZkbZNLGB4DyLQYn+EfEk80ryRXyYAwUtZKrWLB8QZ5YLthY8k8KFAmRjmMsHzc95Um
NASBIDr6deZQSXfJ3Et1mfoUVM+CVfJ+gs6yoN7Wc+gzwOaj3YsTH9BMO6mBGblonCYRVDcC0knK
MF7rgR92E/ApxtqvftOzX3grBljvUdbFiHw0vU/bPSh4R02PTGnCj3GzTB9STR8qCxm3AiAnPSVO
t6FAbtWcgOif3H0D1q7yeUacfcB7LOifDm8lZ+ip8/HSt15bphHiJKolvmrBJvz75YzYxzkLcip1
Uy6mTUMx5U4i91MmqXXuO/Jje/ymwvs0Q5X39xUnKa5SdmcAZREn+nRXwlZnYdrnYerKGtRk6tA9
ps6n5pU87mH+THfTSr7//98MQVRXsEjAlt6eI5JyMCImiEWG3XPDmnm/nZd8hSw3ZpRedfrcU1rS
GIBJ2FT92rtcocphO/JKW+LXtcI8Hji77+l42VgaKPEltAOpwWa4r3rKGkbWSh4mCcVXX3qu1mJp
q4biXsWLAjw2vAsoXOPUf2Rys76Ec/Tb3CcZKfTJKeqq3bRaakwCFT7tHI57Dsz/bwue9DcJA0p5
IpVvnobTwTCigZ/Id4p+3RSh1lwRhafRFWlloBoaDr3XAhv8yC41aCx8HmYQ1NUjab4KkHU9JRIv
7KgJqvvAu9xx9mVB9pj3tJ2NFtE67wZGkD1Hut1hQpOABOrF4gr55OTTsOs3hdwcK+8kuNHQsL4k
g6QqT3GqTCxYzBNBIZEX8qvMmNB2DCM7txxwbGiEFeRqywF3zpF5nFBG4rfy7C8NhxM8tOUA0us9
t9QJvFH/vqw/UxOLyxFCZpbQ2ChjNvTOKpsKIjVbxYS/fL5oPACZnECTf5brkfVikHMxvDDd6LRc
aPJcGapPjOblHhJ+aSDaX8aLMYmvv7AokidxXZaynjKID4U1zt88cppc6x0csfs+rF3nlwcS3Opk
MJ4upYTP7t4U+1KJA/GHF50BDyRVqVAIoIH438aeeuEGJMj8mLNP+65qTt9y+cJwHJ2dbsrPecww
rD6aAl+4O8+S/jd57kbpuKFD77rLZfVuwd3ycjCZKhinkFdO2aGX2ooRXsXiAVomOAGUY4cQ6WOA
h3HJGm9u3OFsaYRi9Ilf3Hbc8dnd3DFn1Blj4qacW9C+mNVPU1FMh3Me/PGObyyKskAdFF6zrqiM
Eo2slrjrLOgTobuIXKVAhiX7G6/H77J76UIQvdNNDlklyvlCDouwkGzuxCj5+Y9QeOhJrIPTjaVL
OFfF9oqfuq4nmps9D1pXsT1XheD/6TpU8C+kdiSWxHLuCfztAwns49wQxIh64BvFD1qjkaMmuUCx
AV8EL9Y0JyFbSopR75CnqecJHRSJLDk0rerp2oA+FjNjVRGGj5P/gma0tLW/zYiTNVIyBZdiy272
9OW3yJD6KNnm5Cu0cXxp1AtxsGxG/GanlwI+V42vkZVHqFw3ir3D8LfCJFmPuFBkCrjZYXfEaCkD
kzblO+DWoP7BWNFro59/NUVYtkymIiRIvpZVqDd6k9cUVddw0W7fm7MtO934HtNf7mTfdGhhwN8G
R9C0Roq4PYS46RvykBGsYZIyFuVZ19xS8vWO3D6w8Pb8j0Rkp87PGLLXPFbIOK65Io2kikW2/9xq
vOs3HqwFunudck0bVBl2qLANwHoqLDMNkYR7MjtgZPWKvms34bIkaqBJ7egKHwuU14vTvrGcCvgp
oNIxzxduKqT/MGDVgEPQAKruDbZxp2i67hHRmqnr6ompJ4w/775sKqE6v/Geh91wxrv0nskIDxZz
jnEJuQfr4Cy5ZQb+H9VLXoR9+E9AF1kR0nQXI5FVtZ407ylSufzHg+1oc2n/F8CwqZb8qcmJ1pT1
4sJSgaVD4OjrER4Hno1fIP23GxIa6SsXNcC47gSzJ69TUwZWSJBjUMNECD3mSoN3Rz1hNhChp40c
w5efRY4OIOCtXPVA2/8uIBwHJeaj5OY17RixSzNyraLuOdud3vFR1kIygKaYRldyqbZuQ40Nnhwt
miOq/mkpAXSjekldbcK44pMLcd5Xop9pVdZh26gU2mkW8BiJ3qtUCcaSaMmXjdqI9mv47zLLc+cP
VaSamk2EvgG01llbFsneOito9Ks/YCqCG1e0C8ebAMzNfwZ3PEeJQQ/wimlIl4fY5A9lw7YBOnQL
EifX2aLJH3O6wcJfvnnD+UaPQm+menp2hLpyaJ3xGau50d3fq69p+r0PZIKNzs5x3JPWDchUTQ2S
KQUiXFG3QNfTPePAB63Rk9YOme5ojuI0Ol+eMBtZnpngaK4wx5C9sl71Ug0R29qo6DFg5s+q/gGe
DGiJ5HRPLb3ljRFyRnZkGbvvSEJIsd+tiHbwf1Pe1eYxla5HVMLzOnV+HMsfajrUrjp7DwiVcVma
nuxhUdSi5kjzWiPrECYyIoM+NJG9U8bEMrfmHrBZf7L864sMwu5Y8HlfQOEnVBkmA/oeFiToN38T
oo/Af0Sa7wtsGtT1675OMi2hmhYHPTjLkt8/tfHelUIpqK+EBR6gG0/0gkYPVwkeqJL/Wv/wiXQL
4DNU89wONlUwZ+EaQQdxO6cf7xFnFXVskD66ZUBqnM+vEycnLEI7ZSCkL9hVNArQo2DhI7zH/k0d
5MwqQoKA2NPG1YR0Xq/T3rprQGyAO1Qtkt7EG4EzPaLTZXQKt+LUnLY+Rb7agJmBWIsrKygBsbaY
qROsZAtfhvq67i5m2TmF464LdMTKZSQWM1mnflX44vuI3a3fa16GrEmYqMOOlM4gf7r+xtRLepZB
+F58QMk5h6LpI1K+Bp7wYS+vDosDRP/Y1f+wqAg/7AYgTw3OHhQjwpX2ePV3Zeb54LyXAFXIEUcG
dtAdYg5oxoc9/lDo6arMP1/TdV5e4FT2b05KgiBQur0PH7sD7GPxCOeq7taqUMk8Ad/1ePQ4tCBO
+mZe3ZI2R1tnBE1oBeHVAvMmRKSdFKlBL1YwzgTBWtA3txBNh9kCNS48w/0aHSSLlaNRpArvawmO
VtKlguvhkWfX2jjz2VfRoGh7PnS1bOCnmrdv86AClex2rbqqlIFv/inuoTstMcSo/FjOoea2GSTm
7OzuxFx5QmIZwz8rJQeCNBbB+qhYbGqcNfmUVib7ipZcvgMcWKCZFhaTp3Hte/4x7dS9v/0EBmQt
H+LKIaxQw2FF9JfIIA51p35+Bg2OCPOKQIZGk+PHDGKKeX4p05t8JbGFc5yebmsfIh3Op8+Pw0pN
rRBl21ERpmZ3tUmem4CwwlfoHn8AVFFMCwOobqzTB6yyGxAWDLko7L16godeVDBb93nGJPtCs93V
yzDwiL1ZhfGIf0CZRKqtT0yWcKSROwZuNSFiCaUwhrbn2Phv/kCJnVjNrhlsIvP8xPvB6CNpaRXM
jg92OIlraYddJZVhggl9J/ZeTQFg2QwIEnRBSBPQyKjCOprOD65s4YCZlo24dKtD1Vz7w024DvU1
bq4bq81apH03pib169ae33yWXYdk88sSFqnGfItEfYeuFqD0DdZpg7UWkzJW2ruPeQB2G/oBvF26
fL1c+cLLewb/TjhzW5Bx/F1rzAzT9mUNieNpySXRg8HkXfQ2p725RGFo5hN7Pim/7Uc1cWyVVWC4
DbbMJM5CJkm0sDCSMqRdnwt1xZkhUPTxC2IIHCJNJmUMD4E5e9KxcXvxktpSx9s3uPz5J00wi0P3
HBtbzxAya1pfDOVC1qUzqj9H2662sI18mYfWwmmE92mEks9jDdHVcB6daF6RVIMiOlhsWxhbm818
LUjIZW95bD9vrLfnmvc6OxlJ6v4zERSy/XmnHsjqR0HY9nPVGgY5/uYQX0sh7T0tETgPiaOcVjP1
iaNo7/3l/4UoWNPuUYNaFsDhmo091E8S/mZs4F3CL7OYC3FkjJEHXKI/7FbFjoE95kb1znJINNep
ZYfaTrrSmhA7adHrP4OJ/uDY26gHMznKVMAWly+uIPwxsSJUWDX7RrE9vIO9YXv7sHQW8ITRvxXS
PZaKaC8Vm/02RMYqdmuMz5nzWQ1W4YtwHat9qEhuHJX4dzpim0uKlXX/FbdJtHi1NP0mBFlyjIk3
iz7dQU5Edv19M4jNXr4al1+ALfMXaPfCTvkiT2RUYemy6HQqCBfCqauEE5O9xH41riLvPjDOwV6N
cJUjkFuD6gfl604QRvbhVIynxwoh2/bY+im3C6WkX6VY6h9ATPqAxKx+DPUt3FNug/FjwljXzJ5Z
gJsYsi20eAV465X3/IfGUTimcHA0EOB6RJWbe2fn12xd76ecsiRyVGsgo75wemNnISN6OJtjHbW/
2kIPUc0E2xN/Yzjk0BOX2ZyodHRIoAgbG/SWSn4S4mZiHC1ZPiKkcP/lMAv2lJ3a/hSQ2C5vnCu1
FDIEq3ZZM8L3RDjiDMtcMKuD/ZtwLYkrzgnbRTCfJGXewMWl+f01IR/4CTGRkvkJ1kHmpUrOroNG
uB3WSelxnEgBwlcIcVqAx/JpemSsJ/ObejYN2Rt6ssEMiAG8TovqdF1Gd+8+NfIo0tTCspqN/3Gw
iyX5tUBmSOBUoxw74Os89isgH7UiJJoVtXUiSa7zOuJskE13mBuFd8Av53DsyHMmn1UMO+oBZrya
YW9SdezLb1bAgLc4NvJ7rcnrjeCCNakQabZEVVzVXUhRp5mfT6hR9H/l1wmh7BeYLFZC+oLaqgs/
bJv6P5Oi48/itrnKLj5F7aft5Nq1QEcy7yD9ZDzXM8pXzzwZZgss0X1Ct7kKqYXEInvkE1LkYAuF
k8uB7aAGkd+3YF1DT9gsoqKY9tEL4OKyx3KIlFR4xuuhsfeZfG1OW0esTILXezBfPLkTUlpRANJH
nIQ5f2b8blH9gD9dugYUCzNcW36OrjdC5oTW9Q5ED6fQICMsLEU7T+PqQZsiVx7vQj7iY5joURGZ
qVBoubVdOgDad2xYvHRXs8GlulgOnQevofxgbukUY3rlMCB8TmTgB0GVOwG1KMu053nVS6NgV91Z
AMDppGYcxldDxvr5wjikgxdjoqo5qhEFtZXSpACZUkcNEzZkZgEfGsIcP0UxwC37joAYXQQ6Gtov
YbwHAWihaJCEio7+ZbdQz6CnTur170ARtodQ0tmzZKS27sQcMDjcFCTMp6T1kBAk++nz7lg3TdvN
oDpTWKmFkPYkvqO5+wDyqmUxdTPuH7bcIaj2E7zHrYSKtKPyJrJJ+K7h/OF+8SZ85UbnHaSAvaxs
eUrspn1M6PZAPfRK4DuENp1Z26KcFturfOrPXp+o6OzAhz64xR3VPwEEVX++81yiQRGLWI4LtpCf
DIK0LtwXj9R3w5hF+HstRHJ0VsqHitnV+WiX99oeuoD36YqnQMAnY/CLV8xbBU00xK823nrPV03Y
Ts14ZQnDolnjHd+ASwC5s45fVF6dRPQHq2KoUCZOFFzey8qAvMvg20Q7bfRaSug4uh5d+cJKWqe3
N3ZrXIbcWl1sae31vHi+p1RuAL4I3pVS0rmsh8ipUiX+4fIB5W6NKh+tASgDUc5TWBEtgoyG45Yc
evvtxU4Lr93b2TI9IuZ4HHn0/Oo8iboFEkXYAvWj5ePhtN64Vw30mJQ7QNK5h5iVt4hNoQMg+TSx
WXpjGkb/3I1BX96w9KSegv0q8lVCuA6LlBxLd7AIy6K8UVbVSwCbeXJ3b7XnMnqNI3tW4phvETEI
BYkPVQd1/UREPytePsVBpeWebWJ99aU53ZFR5Z/grCc9ZG0vypFNjXJNLjY+NGqqlPlf/zRaTMPH
/GuInm1C1Gi3SFuy45tEimjn9z9zGVmDHkunwxx8FpvCvvTnz+SVgZT/HPrNO/Gx/g5/xyp2dgBB
s9YcxR708zhKskbitk3IVn7RrhBWx0uImPAV4ahc8iJlohLWGzDn3c+fiEVzT7i3PTxjVKDBNcoS
asXqt9tdj3qGXTzD1YfYKHU11pbDC3fqaUiIH3JOxFJ0tLPtxU72aDoWE+u0z5jO/urV0n5rWR3g
dhrNjCsjFTVcduCHggeUCA/yY9E2wzQqnoAnAM/Yc88tWDE7pB2y/TH0bIquLiT6zOQ1kr7ffKgi
iIIYfAjpiIdTeZl+z7tByIbtC53gFYHQlzNtYPXTI4bAffizd5NeFfJymnznCLtNWg5Dyr4BW+Bi
iZ7zkeafbvXSuiRTPudnCWEiuFLQGdOpAN6wCLg0Ql/+UyYz/bohUkC4BCDbxneb+HlvckVKuPH7
F3N+u7DAMojD4jvPcqzqn6JrRJTniE//5hqlkPi1jnvWjFKkJFlOmKXreKQDTE5ZRd+qOgi/W+GC
xGuiR0odMt5LrlcrGgl1UbjV4kjNHTT+H0LvpZhoIqKDBSTy2LOvLpezORjLRRlHMtH4AkdA4sCv
ZltKjb41TSyuOIrcJuq66MUuBM5iydw+zz1/MKlBh68vrPZs2NfupDSpan9cbGabWB6mqq2VtdDK
1VnGsorO7OXMe3jV6klOBz7zjeqorfLkDRgnTZe0Ud+eHGBv3jSQpmfg24eXqBtzMLjeYd9Q/WXx
sTg3v04DGUrlEXBGo+iTpF9GUjZp7SP9QYuu239O7DgIB8phP6ZolZAy2fgSf2QnEbcQL6pbDsE/
cazlRSKBMbCXckvsiNFI59b8PFtQkuo+97vf8CvLoKJN3IAwPqynpyDRBtMH0mYsnY5uJGto6AmV
ftfp/HcXLS7UZ9xv+J/YtWZljDdvkiZkc8/li9oOcLRBT5o0yErMoWnAt8jQ4prdhRM+ZIbFoD6Y
fP64zve5LXU3Mp9/ZvMmVWZWRIpsnHvQNZzvksIMzz8p7P/WE15Y1Z95DLZa+H6nEPccv1IOmqOD
srApkKeqCE69hFrf5ibFkR+2G0tLKQWE0GS3kWc0OBbRVHHjbRgbw/0pJyyHUIzklJyki5BPlZKW
SjNdlMelZ3Kq+X7he0Yse/f/krgtU860CRBuKrJQisEGXigj3VSIweYTIJUl9xXl2Enw8k4qaR7x
U3jHNXF3Uc5bA7/0fCQ35ZfXRpneFoT0O74qL8vR49DyWuSerI9o7t0CJ4+gwkMRCfwNX0xgagQc
sZdB2U6tA77cqKW1dcm0TUGrexMhcxG/awygHzzEJ5gNRWwXRf6piubcfI3M73W2NNLcD3XorEmt
QqiDlWKblym20MmywOxZqKZamWcRTgnGIeS7zEAzXFt7fFYzlxon8B5jPi+zQyrG2V5rNhydaKLp
fQGbjHYpjgzbcqiMPKxDwx7xCk7Csj0enw6hi089xNJi/IYGNBuq4r+HSeYBnHQW/VeRMwX6TRQs
d67bVadd0tAGbh0V9pA7yx/0eoLqNkygSTcEs4UytGXjACIn3e4PhCGxSqnsuYB2fLGuCkQaPBBv
CQrGih/F4EHdz06bgPwEgPUJZXDIvsvTnPB5/KLP6LSdGBUfGnmATXmQ8ZQEZN//zRkmoTPaOzaF
8pvnRLd79U0JhBV1/2aMLJnpSJlqeIBlVstYQYBa/kHhXNVzTesj/p3guO2/5u13ta1ozEl+QCpv
JzHQy4G2zQ5mqD7BKM9heNttYQjBbI9rOeGHqxvT8laa5JJUNmy4FnP9PmGnuF4C/uHylvUJWL7R
ptAssKUBiLs0I7WPuLSL2ofQZc6VzPPl7oEdWKJnYUKKxIjGgx2G3GGCFS5EMOKcQQBOcsd7Kl4P
pHSNICDQc48MQ3bQUbnqd+ZzizlLVsQvxYp8Bz63Yrb+uEDhqZH6WV6zywxSWjsPiwoRbP2p2PRG
ORktgEsdBoG5C+Y1HZE6hC5866gCDaz6mYyz7Imt6DwrMEsRU2b5dZYgbH1iuYVnY7EEIDhd5FL2
Joc53c1E0yrLkYBOpHL9AwCmU5YGb2ZGY1GbwvBrunc91SH5iw/7y9Hzs4KmmZBdsSs0Y2mFm4ov
U/idWr6TQccGU2ysue1rhn81jJjoM1WaEmXYreuof8k1WejRpUK8as3uDkzRXPGZEJagtrjTKZTA
7iUfeQhH8iqU8D1f62f7Rob0ZVP265v58ZasDcxr1xXXk8Re31l2xYuYxBAUAFKQHxgdqm1v+sK6
DtJmk8KIbbW3JsC3EZAoKXv7huJOABF87Rgr7pZhnRm0+Z1yPjXHKjqkmnJAjh/LKONv/9rg8i2N
BzoZeKQn3O3ceYtjCDiXYNIb7VU+ve5dQwIS/1DGpohS6cNpGNZ4seisf5QmJovcXeiOUOo42VE0
Zur6DJaAgZNn5EnDfnYWEz5KIHOEzeZf641kN5TqpPz0eUHJoHDsvguEm7IOAP6Bc2XWwbGE1xg1
xkaEEKEQERalHEiFSQl02wCJSAhHptJIAdymd69oAXXoHOC88BEWwnO88lVzyajdVIZZU7HjYlEE
7bj0Tyjf6Bga96nOP2pFxD8etcNVtkHVa9xj7bXQA4P+8QXDzuE3nzphph+MyThVnhEd5Ct6bxWt
7H1b4UaDoAuB6bR4nHTkSz1oExgpwMKKMLJeXnJTl7x/yESo2uMcs8+vcl53+mQnqv5GOK9iv2z5
/NMxsiuItAnlAfUcXevMuh7V3u8B4b9BLanlaWpEZ6jiT+yJYvB/PT7qimC+TOgtC98o6HoSV1oR
PtCYdf/wdK3E/Ud5kf7vOsrkvXYa1wZg+JzogTJ5ieTryTRLRGyOpkmkFz1s5+pMgKbHSYdJtanZ
3+lJM3C3rmKOugyS1ZygV4dUk/bDB0F+8iTCk14CkVDNyN+ZtyeCAeuQ234p6Ku1X+FuKbV8FEcS
DCySzC3BMJvSmo4NOByhIamc66Lf3OxwSDzPo3saFR8IEpwaztavbgLBmv5BL/7bkaWKmoPfsqhJ
NHv3RBnumkk4rnXsJNvL8NU5L/eMKCqkoV8Fjxe8F5bKwv8ljVn8ayh8bNzOeSkoRbe36vkzLDaE
IMMux69dVRAyP3AXfyiLkyFenmquekiFNiPQ/FKnV69Ze4PgtlEYjghK6eR7xZawMnc2LATjG9XC
V8DEbD0+TJqhIvUoXwE55X4RfvlE4Mv/PBLBkXzAkG8zab8oi5JFLLFzlL3qBLhaUyQKKgm1Ksjh
fHkBYMxW28EAwT+r/nCdvkencolaLmx44B6C/AokhHOFAJ4CxqcALZwzWXq5J9AqM/20AK9cci9N
f0ZiYMZrZoxg5WfTZgY5PIB63qqTW2nYHEVwerLSm0UYeE8qWWNPv9lqm6o0QyqGB2uTT+4fcOFr
R7Q74+tkMchpfMbk5xCe9RzAIxdXtTjyeR7HGVQq47hskl0juSnz+s0T60q/lEaNT08OqX62I23F
LrGvNguBIsPAtW142G/4jui9kRwqkfcjJhYyQl9VZ53p9n3ucXNb44tJJHBxgYBy1PkFArx7y3Uu
wG1MZo4P2KvhKILiiXKCFi5Ead/qS9pIVIXNXhH2EGPfImitRmtGuCpur9Z6ubcU/XHlsIs+SkoW
F7QjGMUwzg+G1mbb92Q9Ku/KZq32iRjrLHFVp05a9xYUrhoQxSDydMfLvQK+ICk3osGEQwN4+MIS
/IgppuXFnp08Jd7r4TqQteU92hHW/eebY/ZUlQplh8Y8B4VluQ94b5xUJiCuQhy0XhrF1nvaS4fq
7FdxubI6jfWr8dPVZ6MTXC+E56vDHrOm55lxv13eQT9a3g+s+n2CTvS8Zs/QcUj1fllWBITYlcY7
0akJkML2czdH4Z+n4HkECcfe30RaYJjBlbL4gyQUEDaKo0N5AgJanRgTe1qS+vOMW5vbnQuVT22r
yQgh36CU/Kl7FYC/C/djkBvisaN7DM3bBveaIB9Nt8kptGSioj/hdZ+LP0I8pUcyLKjEcOsZITe/
FGnbw/ccQLJXzPZqVf+EUmwtQADOU1HVHec41EwS4hLJXrT3nUOz1q06Zo3iy6Mqv3W5LiIQhZKK
uJOd2WxiuDPwvufHsMHiQtRgOscDkRu1OuLXI8ToWYchEruQ+tW2tROdHasOvPgrUF3s743AJK2w
69hyBEDs6jdnNJLQ0QbY8NV3Jobp2GS8el8jkYnmQPcz5cR+sQ5kw0nLxwdfe15EYm9NALYdcswK
pB4FfXv93AHIUHZzb7kkMrpTAGtxJUCaUSx/ZL98EzdwDJmjmDde8jCUcjHGhUdAYf1Hnz3mcAMF
QmdCfeALN9EJUfVJGtmn3mn4Z2zm7EaPfvU13hhIL7dns1on/YAA+D5QOlq9JMcpCxYvKKudNlSG
ZSexVk1a5gCzgTxtJRfhug0LWvfD7cFJQk79SIlJKG1at/GwmIQ0guLKU3VMylkbxua9Yrf+5l0r
2Kr5t0/KJtwKsGxvAcoNiBYRIiXBjOfpqCtGQbp3AsiDoc+nm1kgJX/qdfqK1++mGSO+/1a/DGJu
Kqfc1kwG3sLNpxJrKtzYIWO/X25tHxffsB9b5Z7bLoHDQz4F8/AiTgjf02DStbMERyJ0KmpBjiCE
f8CW074w47VALg10Og8aPpujmjYjKET533lYKXYqB7V5Yjlq35fsEog9+6Bwhw87cHwFcu+MjCIJ
KsKABrs5uuarM4UJsf4Pdqg5cmYnHjzITaB5HjbjRrd3SRfuA1cXLSu6pRHyRF8l5IH+vgx7e8a2
lPaAopq9pimoRKr6rUGSvpSdanPUzIbmDBuBYjWFfnud8VX+25VKgfj5I9OvLbit+epJQUsE091g
Fx9312g6KTMTxZST7jFuHAMsNjTkfk2vI2b+TD8Z9+D8ufoHrCUD8Kyf4RHi8V7Mg+76FitnklME
3BXMAogFmY63JK+bARacrQQjXUBMQlregNFs1wxDDbLI49/0/itv9nXcrgwGP8klABZu6zz7wXXF
B60We87c3rTHtkyAujqJ1mE84DjchL/RKFCwQreT9NJLiGBCXTgmiRjaRD8YIzLpfnHS1Tu3YQJG
UirrkI9WZhaGDKhNEUfa1ZLrN+U/aOSjH5SdT2fe5CnhPYVm/p2rtVdT//aetQukJpIBw42Ha1ly
3+MQW3+oQkqYbVCCc8su9dROo/DxrjJI8aBlrnpArD0CpfvSWoXdLOQkPluRLnMbfMBrLFYV6gXF
YsO1YoNGly43Hd24Shd9igrBls5EGk+XFP3vDuCfHnwS1KV4I58T+ty6LkGnf6VKRZAIrDeB/rfW
/miz4JsLuHFqk1eqfvoqcp/cJ8mV9AQDRtfLFtLwjX+/PIsQD03fhNN6hhA46ZZvaSRPE0g4spDx
U/6nyPJwWx4cpi0K5599bbljw9gi5ylo4wYviksytSHg6jRlKvlPsf7lSp/IGEpLa8ataT98jj+I
RDyrqN9vmftHjTaiURlasp7jnGm5SNZm1LHeNJrw+++I7Y7wiUyMF8sxMFRVQexXEOQcnwoNNVJo
4AiYXFRgzvkwtQAQ8heJqu4KqV8W3+FDsG2DHKlSIyEKjM0ECt3+bHOgBCl7RYmjWxYRkX+OrWHv
Uu0DqCAZVHO6y0b5kPvX0iq9mTBGBjIPinatXjPHbF+X05fhY/GzK6JSIt7NyPpJVCwJGoIUeDjZ
zyWKuH9bGqevWHFsoa0qTQfB1XsTeSNOrwStUoikVAdI7aeOsLg0MartAo8wU6meRYbVjYpd4DV/
mCV2APhc+jFv7ues/Yp0RMesSAk4g4eZS/5Ed/RleeUSu/VuUWAoGJBUIm+w4kuqQ3lp1cRTwARC
hZIBfrwumE5PL8kHSEl0Y2Km1KA3wcurTMWR4yUjXbPEn/UdtwFGjNps8/6nRGgWx0Ypu52O1yTn
jp0DN9vEkdGF3ypOE1nN/iuSOA2vl0r5BOXAZxt1NB8l4U8OOaYuSH8ByAt3jDJqkKy5l/paM4+2
7hmtatoxVSkmivJkGwpPyqv5j/+NITAWyiHvaZeGXj2GxxJJZ4DCOKFdjgCTgtOCnTfIQiuIYevv
zc9pyCovBqCFMhAGyxaOmNaN9CrNY1YFtgcZEGFkaUPWUMzs7iZGztn2AmT9L2+u/xkrgQfhUYBK
lgqrC3MPaBoI63lAZPevl1yBu1psy7lq5jUvajj5WBWBIVeEYgXbOFQB9qzdd7sTxdG7neBfBm2+
SMe7/R4oGGkiq6ErtTmp7GbD50XTW9SH9pPmXKz+HOVh/pUd7cMgdV/lqzRt8pWuQm5t4UgG7Brf
Gmqqcv4tuek7MiFB+xzeJl00LT2Y9+uE0P5N+K3RGjbQ1hvq2As4RTz0ou61mD0eaq/qTElBqizh
TU59OjG0mfvt/R3c8z6LpwabGQclfWBO+T6ZdT7s+GOS9t8snjd8zuAw4WclPd+3zFpHzqnQ4BWX
YKDKLL65E1bYLFo2xn8JgnMmewLMIoDe+o04v1XZfTdoTzKOtnSJr5H6meqDA4vhLIMtyg+Dvpvc
IdoZIqlpB7YBTdR1UuuKKVlLpPOKT5Kq6xzDVThYWS5FYqnHjEiYBSCMM08FCEG5qYxYZqTVkZ54
C1BVyPsr22W/oQ7GZRJJuJLpK1QO6D1jiUfiyyLjivp6rWja5euwtvA1/0Mk+jBbV6O7wNmvA9zo
QDAJ4Mt1/ZpJMGT+UkFIlyldzLDGSF03KooLAYQZ7AWG7wjgqxJmF3ANKT8WitB3LlDrc97JrYEn
XSN6Q9KnoGch35JW5Pa8q5hn4tq3a5dcv2sGYxLfx8IWIvgAN186H7Fb2jduVt78ZmN8OIhIvpr1
59Z91gUmv5YziASCo/K89TVwlUGiz+iGv6OYpsUKW+3o8xkAYhsC3s1tqn/QHAbXVVfVYYOCmwYL
Oy7F/qIXj8y60NydhzIMWz/+Yp6AYkw/MAmDi7w13T8FxUeqPYDu+VQckckpserm6wHTFj2By+Wg
0UWzrudJFqV5+C79dVi1W6XWmO+JDh0BHI7q4FTp3dNtI5I5EDDK8R3A6p4/ZW2Zdi2CewX8OI0N
PYbflCpKczUkOSTFvn+GZfJ2XoExjaTZ1Jlvf9neWy8b69tfZMqz9o8O1Rlv/Z60mWPIw/bW0hI6
sTx9qBzWNPc44UlpkqYINYE7Je/q6voJSKwciMGWa7Bn6stLf/WIH9sD+J1uGrt06mTxgKY4ksjt
F5GCL0r7ewy+KdBgjqHx2vgPlYs2K4ozLCJtH51Df4PJIEj8aC46MY3ug2rdFRFPmER5sgh9tqNr
w1lXbkPNW5U6e30GCcgnCgrTWaUfZxK4fs4wviVovOxQ3sgkMhC7Tw2QGGH6+PrKwqbt/WXfAhjb
qtuNZmMy0YWlHeiRbnAINJ9t0GUWe8LVxT2lKGSi7PLXwSJYoItYH/SNW6PvqTTwRESlu+WbhXBH
YH6JWhmxZ8uhqtY2kjLqXUP+DkmWxV0ezN+HbXXgikoH/P5V8EgBn3vuKdvxUuyUC4e5+07D03Cd
rohsSM8yJps0vEMrVVVrJepuQK0CdriT2lOi8WMmWTzqSSqOU544jqtmxXbnKUV88GbTfoWlZvsX
xxB4zZuymkzrJrntEgdgl9QVP0Wh4md/hmRnBaFkm4RVrsK6/oqIPKtct1q+RXFFy0JQ9zw7B/04
Lg83OyupGmScIBJjHO0i/PjmyFnv+NGuKUJoOzF72R8/+z+uTxBw30zVlUvczhJEwqvDGWX3UG7e
TKBoozMQBm5/p8ledUdxOWN9b1JeX3K1h/PmhPp4De3DLzC0cwnQ9V49VoR/chdQ3pGOlxX9fedU
W96UuUlmbXlvQcY8wR7sjFxQeHzfG+Ozd/MVAfEoBCp0R0BBiPnO2blY6bJFQMw1eu/iiiG6nfw+
CvALJe+aTDxlxDeUPkZourilRt2GlnKwWiikLMkAcoEiyWZUg2bs7xAAEo5X+JZX15fOZvMizXqD
EzgVzJ4jjcpR9tVeA4eTubm6CgtTa+3kCKbKDRpFTKQeliLSzwQ+d+jhZprb7S7BGc9Hdh3HL2/w
7S1BNbLJeYJaUwB7IfZcY6Hx5WkkBww3MAHOsQqx31SheDU1JI3wFr+ZXEvBiFZU/W9oqafqVSGf
V6SAT1LaTQyEKG0Vp9ca8NNANJQGo8NBUPj7c/ICPGbnzDkn58vj0IPs2WwBbNNE4b1NfNHf12NQ
phgke6slrtDkK/Tm1m25jgHxq/P8FAV6n9+uHeH7xl3th3sudoCBejPJoAeYLvuMTfniXbm+NeFd
Wbe2d8YZIIPFTEw30Zzs0Xl/uG8NWYsykv7MxotCHdsnMnzO0N3LHUEp2qP56zOk/kqQ9fvpIc8I
w/nOEevfTXQD0C7qK+ST5OGp9lQDTYKyLHKTFa1oaReGTO0+z1O8RI1FE8Gdgx+5vWGmPrcdC62y
qp7nz4wRFP5vuPqhQKsc3F3B8fmd+ttEJl5HUc6qSCeJgLbHzNlOejDrXU0apXGP7rVVVCI7cfN4
NiT5N0j0ck5xvE0efh6PmlgPWZf90Z1lJSlQqvs/gbKj/sPxQ2xTRgD16IPBlt8nuZbQ4BRWJFu8
WNZMQNtqrxjSAvrCmMTphrv7+Sa8K/6myyrWMbweT4oqvfup1YEedNVRf8wJTJAX9bMt9oFaTaW5
ONOQZDnCNpGCCdmosQHTwKyGKHC+KG0gA5N6TITT2sIVUPjCxUDV+cm7pDGeoRQ9pNtGPdWM29Ye
/2wYm1ETcdBFBkPqhSBC2WpV7G5nNcJyjMoCdGSHjHZcDCpf6zsspXzuBIAVqoUxXZGmB0Tyv/Cd
uc3w7uV5BSF1kU4m/midOWdDeNXeZ1ucR97ljXlBe+fb2tbbt5Q17vV5Lc/BBf92qiv8937sAdTE
BLJomr/WcP8i6aJuamuJ+5tGQ/qvMmjwKdDsvbxHIH+9daspwskA5mJXNdYBoyzhfljR6WT/1DYh
ptflKuHjeYYZS36/eG/VmvJciPMKH6YRTWQANn0yAv+nqKVDlrnomy3keRIKDy2l4mNchre7eMfn
sj1eExyT9Qma119UvoF4LGcAJ3U7m9z2o56JHgAGyrkztG0ezPWluoSVHtb7vHHa/JUEaHGVKQCn
XwAmkLmGjdVVWfPvxCaEx0Qc+1qun8e1V5+g0mMtzKb96nLU1wXPCSaI4tjELltLK2pQk8kyeMKA
pOgp8mBINKyvdoz8NLJwnZSMdzoH50eAbzSJuniccn3Z23kHO7MsDmUrZ389Dl7K2Nq2x2fmHB1E
AT6XZOjE+cXdZu37xBDNKtk1ZeUx8/vysh3lhiSiby6Byb4rFg38RIU6dryUr6xxkSrirMyzKw4Y
xb5YO88ctDPk0n7ANXbm/T6KPCQJqalQA3FZXVD8DPajXMs/TqvNFRLR3lL8y3Pg9aCfFvMirSin
NdOO8bhSzhMfvHeqP8k7gxzMrRgLy/6DvEWgzp8ACny01qF3v7LXMLXMq/k0wjF/Z107QUP359Wx
a9LlktmTTmrLl7oyXuUKTAcaEDFkqyonLDdxEGlEUzlNwN4BgVG5v2RqF7jCItpcgl6gHcZHxLtj
6lxjix1GxLRYTENeHQfakJU7Zqz0jkad4+iI1wr69MW8QCvkyEk8YXiN/ER12QwayjnT+pz50QWx
M4SkGm8DtRzQ1rjXqaqbpMai16eD3NgfmJ8P6x/+2w1QsRTQtOtSRS7e7P+0nHEyMhGDcukmy0I5
6iZry+g66ObOy+0RcnrI8SP07zR5UIqoF8qECLjjbKnA+iImpmZrz7bGD9XnwEDCg3p9J2K7pNlu
tTTg5hLww/xr8P18ZqyOrkJrqpD04lZxTPtBdkqzqLHFGsOI8mwIkKsg6afvsCHOL4HX3SwaXNk5
pohfI75Ndt64eNbod+FEIypxqDMY93MxYA+FyMvscCPUioZyea12gnE4BXyO+lcnmeTKJRjMvy2F
zGJaE58EMwV3RqTtFdOhAnyYgLX9hUViur6FtRGgygd2JO4ZMmP49D0IvssD3DWqhiOciwz3+mqw
xFwjhOJ/lF12llu67ZbQ4qhWdGkz+afCkLwRNSgnUmIjn82jlGoDWLHDhJZ8xMt8OqfNmEAZaclR
+p5K6pygSisNC16I2RxMRecTpAnIIRw5FWpJ7XHuqt+ScldmzP09mhdTW3i0Ti87DFVEk4oIIY3S
6zn29gS8u/Ete7ddJVDcFfzLAL9O6JI0L+myFbRmW7hmppiAuOO4gkfNBuKrsg/wmGq+qnGZ+gI2
eXmKAMbH1+epmiWLaXibkn9nbNXmLGq8o66xYEwDQBUw9zmPgyvQvvC+o6O7sUuef9Xl8OK3gF23
QY2ZdybAXbhHNDlXTwuRO0lktizj5oYJ3/+Sz1QEpwKioUadP5oy4S5I9GMyLFPZUyFgdhGSLmlW
WAO9WScXk/YbaT4FTMQwUfJU1B0FhdWhjEk3Mz1vn9OljrubdJUtsUj0DpAwgTORGyhKxIKBNYF2
LePU3zg31Xu1jeAA9qHcGNBElyozKNYckvXhdMpD5CjUqDfKKlyTMdFarfRfj4cPPY9wjJ1JgH5f
diZe2nhBwKHi6ob7ZYFz+FRNLq5lKIGhzsq1Q53pjQiND0gw04Xq1Jqexut919kgXqYTYtVNMA2B
1OB3HukJEeHDPxQZ+2AhYBHz/VT5hl/l+q+BuaoK4hBSW3kFOUSRX/78OFHKoWsSphMcaN/+UavZ
5zMiutZ2rR0zzQndbsLgCslZIeQM+sLXrxp/tp1LoHTzFCeWDqebd1l1Jmf1fDYaoS2J4nYA0c0+
NmUZmEFkSytjacpB5ibn67tJqH55aoRBryKjCtw0IDvh9+Zz1S+oriTT/BYVbQ6SEvQgvL76ZT1u
YMEwy6xEhJYI39XZSVP43ZYyViz8LaZcf4U6TUT4tA4kFkaS3aCRK8qsJ5v/8+WcuGJkwphGcHBr
6TeSA70/DwiiR5DGo2l657sGybgAHEsaCBUhcBW3LjDIr0S5NKPfGviG6K6BNVB78KSxmd4BmyP2
LSVpaLWGTG/2mjG0umiV0hUzl9EL8n0mi152tlhSazu+OOCgWjTNmdFzL0U/ar60GbDPJ+2kouVt
n5YWrGAOic+CXJKa78ID/9xSLk/WFLjJau3iJZBa6v1kYD7Ef+J7inv9sSC7v39NwUW92r+HQ9w6
Mu/AbRMwmGWaAROA64Vofrk2t8Y64ICG3JGAFg29EztwNJdlH2qHHOqX6pYAQM52EqZcqUtrWyt+
uEVuIRKv0pqFbPslYu6E2uv6Aw1HHAkx6nrXltoxtPGwtYEUDWARY8DINb83Z4eHXQYnwUetnCyF
0Pt6DcGaPJ07jtnpT5GjC7RtfFQ3Bet8Nk6V9PlkEXF/5pXVtsFHpizBVnDFUYQVjrECDEZAAoHX
+Y0Mv6IRPe2rJ0y2CP8T7f/4mSnkEYC7O67d2J+oiLDqA0cgrkrM4uLZgR3KGrGB7isGHkwgm+Vr
rbJ+RnLMGS3fr0+hDujEtYadFopsJS1IsKVYWWw66ziPmChfzZrlZP6G4TA2/wOBjY576b0Bd+1k
kyWuFCpqyg36kUhCUfgGlTDaB4lOq1wm/lLkupxVYgs20GdI+7JjXH6Ck9LibtCWSeQuMPcpiMA9
3dOLZccCQSk75bd4pqknb7RaX/FDCrtR32dWSRk7RBokraHZ3JRhKUbYHEGz6tg2OPeM0J2mhJ1V
vJPvoQU7TK9RCZHSHrLDn8cuzrMf33Nf2L5xSwd7p3O24EWtQr24AITRGRjFEtQaECmbAI6Qa2PZ
/vJsn8H0RPQdC8ZQnJvMNqYagx0jURIkfN7HEZ7QikmrA/6VzDBG6rcHdRyBA9D/e2RlUvd8S+RY
/XL6cTwxpf/wi9W2AmCukxol66g6wgmIR/5t3u/S3bNksHnlnZARZdzZ785QQ7gMK/hss6One3ot
2PCoR4ge3Tu5On13NNxeU+IQkfJthR0O3je9k9/ycqtocRgCXJsuLHQ9HLBNw34+hTJvDnlS+xMR
Bb1t/D7kjPVGr/1iiarfO3xxu37Rq4WwaG2UQpHIW6CRegUUtubADGMQsYb6ufHex+Wd3JzCVkg6
1O/YYeR32rf6DjfUfZooAoP/o2zE61IdU+N2jNjahMPgWD7EV97LC8SfQB9yABi2SDPgDR6QYzU0
AXQC2JiHmgK8t1A4qTH10J15KejtYNIdZvakQzpa1iQZEQqgOUy/GXwHrnWyzg4uLQTpCh4kZm7J
au3YgToFMalQ3M5OUuYzcEJc6cz6pjv9nlAVyxmkN2RSHoAf/uJCud7Ax8r8HlmA7h1RDorJjq8l
sMkIbtJYnctfYjk7JbX62x1aUaogUpZAruKJl5KH6NEy7q/ZLqDLH6NRnX7pkFTdAGVeKhMULPeN
DyHKykIIS5hHvm27hvVyXXlvpP0Jzn0VBApUaWeNYAOSjCgwtzXpYDEFoNPv0Nvh79VLGuOJh7NM
JbPeQtHq36IafRdK3QZ1/sSBGo1bSYcOwqGUKsG9TUffGCXsKQlpTRYVeexQ2cYNKW612N8kXTqA
PWt1XnhtCw0YAVV5uPgL5BqFVDLApDjkWTJCzO+hTIBu+b8dFbgAbPBGE++yT47/86YAmFhR/7Hz
Tvymc7e7fxih/lVAV2xdgTeoaxF9MVrWeEc1v949Zajp7qKjb1MKnuR4kflqna0ujDTUkFliLDg9
qddb22ny/qOSFxsSd8z7gub0B/S5KBRVkc3g/ngaY+Tlt6qqmfJ8odgfGGAhUuW/SRZUF0a4ui4j
O21qawQw7mGakAc4VGNTQDNuXOcs8Pihvoihva8yCKkRPEeLLMxREXgv/le9ywp2+H8+jdXDFFLA
iwUT7dh8l8+QbavOqpDoheIeHvdfon5bjWCBuNA/9sye+2pCHQJ7+2BD9ZM2Zmu4m6MW+cnZR/m6
bX4s1met8kzt4NjARWqQ7vTdaF/PQIxgU4tECPodd4GLTLrtCpcpQ3EBWotAuo5pA2s/HWaM7seN
uaU5WhEE//pqtnCdQDlHClxOSnvnM8IxWtpnzSBl+shhZzMa+5qrYeQ2jsQSpwaEqYusDVRdH4ga
m3kwlZOl2AQ1BPU6LVr1Hza9fjuDNQyvF2KW+p0y6VKu7nnSP1PDxAAkOtyNEAyU0AfBlYoZiYsp
YSBNrndUE0nnYxL04niSjudDV8yU6BxMEWm7Xu2a+ypFYAETYiPhyorOBBVHi8yEgYhFfk5uMmJu
GLfcQMTcLDKEtZTw8mINd/M+Okjmk8MWlq4k/HpwlbCyyEfj/qhB2aF8kEJWGnHcp20C+uXNQZLv
TYBTVoLBMXNiES020awgmyRbeOlv8wsBYxv8tYbh+5oTWFyohF8SjtIk9wO6TgJt2vPjastsULxk
RQj6AlEaFitRtk/20OAIyuQ7f521NarGME5p2ySNDr1pdx+o6C4m9/MKvvjBd8cJCBSfqSzRz8Gt
geqSc748+FhXJmJdp28lRRQkdFi/8Y8cbsgX7sq+dWdyuTR7IKsx0VCwP4zYC8oTP5AK/vFG8Yay
5lUQh4p4lWrWF2rAJD5so4DpufZypeNWx3VRer3sT5v0Cp2EUDHvHSyfVPQMFWeO/rMuk5m+8ZOl
K4IX++ze29G22DWEOoeqLVOtCLeJ4N5JhRWxeTxTCq1Ykm6ZJl49r70HWsgG63NSnfrbfwtTjgQl
C2cx262E5ASrzVywOVzolp+8oGdlQGbpmX8rJHynvoYXovXHOeQmPSouYU5hgdStuKO5IJIUh6nM
sp0BhmwdCu4YR2Go8LfRzmtOsApA132amQDEtfgv1q+XqbeEI9hOirkzZh/TGAJTLZq0O/3MMmEV
tL295GwoqJ1BCntwv8al3u8SLBi3X05dar1nNcMuUMZ2jLO/X3oni1yriQ5u41Oz6zJz8Xc8XcBM
ASzHKgSbR3CBLkvMJvKMun+2WWGM3hUMJI8Em0WEBpnuBbidLI+NjyI6Zw4rRAq4OsQI59upFNLu
B6/LzIB3ECT9CsHdLKYJrloYQ2aS4At2wvVsomB41kPajLRNTSZut5OWH4IAByw/T2592QLHSO2T
yka1a6b6odbzktPTii7IOwSNoatsr8VUpgZ+Sc9mpoU0/jLhWetySzBLLRitjEvBjfaMQDo76C5j
/UKMqFesKWXO7eQSp1XMdQeHUTCDkZRIZTSQQ9FsweHTGN4byE31WRvVE8HVg+ZrYEAq7sT5TESE
AsfpAh30fuFW+DW1Q44wU7C8DhqnJNAo41brdC5YbSNFfn8jCy+yx+3CLdEBlXgv18fD1K1Ib8Fm
ZKx/TMCmt7Mhu6v97NosDHbthv001Jn1mMK6Q3pVmq2jQGrxl1Z8j9BeYBEyOVGEjUgdGGxYP3ss
YjbjsyjDc/6XrXwA4LaqnBKbuJUdY5OtydAxpO83BYJFm9/sEVYHePmMHgaEYB2G1yDZIZPUPeme
de4d6oovhOikVhwwKR/2IqQlNgGOXWX+pTjlj+eNsEu6EfgP+nyB/iZ9be3/sp8t+ZxCjAzPKdXg
ITOEBY5NzUv1qEd+v4nXP6UVK3lSoaGnFQiHqFKjaHT3oTnMi8zNJ+3kk/jX2AuiBKd2c/xJoe1Q
VjIPWidKkfYncS5swj7NzYm/1xhTEg1cd8KVoOAaNoEjesgy4pi2GgFl/iO6ciciH342uo1zXzVF
5iBuUVOtXTZJLMvExaOdrQDGCm6NsJgjjYnjXSHrqg6/sbg0qyW0CKf8vIp0YONMs37oMtMIV8/m
YoLT8ISvcw4ydSeBbe4A273GjMh6+gJLNUyEXx4vWXZiXLTiPvt2lrEhPq28H5YpPsgK43vFuUAV
o8vzLNhl9GsFmPuMOXL/sEA5/8fA0PLfspXytP1po2bc9A3t5TjsmwDr6iW0hSpwEtr49SWO3DDz
17Ifm16QyHb4ToCnfsufs5NIfqLEUqdeN6I5Xs/QFMUhvaknwOetYS9HpmDbaJri+nJxuaov1YRs
NQzyOeMKWNVTQPJj693+rD+zRSb130IcwJc/0zk9WVb/GVeiiKJf55/n8UpiHMgBzaxoa5iglFqO
HQ4ZxBzJsVkS4VpDcqtep+p1TOWrki5LJQa8lQPgofH2opax2Mdb+S1olELCNhHiw5PIZ1LYvFT4
EAuo8ge1+oFmeLPexfAgPl/DloDfbDPqPrg3eSovwEvHV/eIWLm4br6aJNRkbdSWE8PgWj+p8mjm
OrqqAQTppGf/5hQL6QXKtxHocVf1GQ80iKAQPJt1nRfeEbVJmoSzn4ejVEI5nzHfGkE7uzBUJSD6
u1O1Bp48iCXMoOL11Uz6P+c4YBysgdDcsN6uIDXnLWe65TCfjLrPj/jO9GENyvpDmF21xSrmDlwI
AeHBya3aHc9Dp/iui/G+0qed6TVFdaxu9E569LqrXGMVR9245zYdyJp6
`protect end_protected
