`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hTCDc+asW/tBEkbiwaBbFmNMVZoDIFcAY1Xtjw2/5qvTHrHxfjowMxaSTdMaDg3UjW0H+j7OosIR
k1LvNj9d5A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZSTMgs/LbjErzH9NHtGXsu+wUOxrtBka2Dwwd5+WgqsTn1nwo6yr+5bBE7IgRrYr9r5UzZiofPTu
pNnDSTkt404JAQVxGBoHEF6wlWpLvowa74xYZg+Aac4SZ30LpgToFmDkXAlaLhkvrXT/Ejux+Uim
szhrZbEWaHtwX6/BzNk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Tprp6nw1jVDd54Xf1Dm1u9TK24DNFYXUErYdnmETt+ODG6rrBqZk6L33n7nmdLiOSsU2uMnKrHtG
joqyTXSqgeFMATzx6W2AI5Uol4k2/GIqWRK339RCGceybJ4Nq8JdzJsK0L5a8iOsiFHk29kBCepF
PCo3g0yINyGAy03PCilnYVJFMEZWDxgxrnUuSQ64wmq8jRAuthxUURNqwx6xdEosiIPgiabRofgK
LH4tc1Adh56PSs9upj48JIWjNF5Bk5tsfp8DGAwIqQEz3R/iO8k/tQ7cAsYfbt+4aIqgZU7E+GQu
E3YLwJloH/jKtLyTF03aYk6JmWjYU6DT2/FLDQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aVks7Fu7AE0DZAqytEkKo7vhq38Uaqwk7TMz/9bGeHNTxS9GZkC3gQE5QEivi1OXs5k8JsD14Oum
j1NGXYl3eQ9RwoBEycLNilyYp6lyHeW+bns+ZeHrwvcveQzXkTmqo/kVhql8Kyw6n5uYCTWgaYBr
n+m83SY+ly/2O++pg88=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VLxvk+kn2ZK43mWV4Imivw0/sYDs1FIHNvrYlglwOzUif/l9R+KRCReEHG8fltOjMOE8xtSqXFJL
smZzKwJWUy2h6c7gLO+7W8OVkjkTe+7EAhCkxBTYsjVa3Fa5SL0JMMjUil8XGYUoeK/H9jbh5E4d
+PGLXdiabEaV+H6/qMNC7jM1H4D+iYuVMxONX7w6QOw5uf1Mitfjc1hc9S64QksviBT2MsmCMlBZ
zckw1G2XkWMrmlFxZenhfZUr84nfcafcoQtc4m0qaqpzCJ2JtE5ZBIGVcoLqmCSekmwpb9oY/w/y
mZyQlu4brgvGVq9F7e/u7mI1J6o4eQTw3g7RTA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7744)
`protect data_block
Yr8mTeds+09OY8u3sv8e2Xt+0+O9lefpRyYfbfkcvnmDvFKPWz/eAuHxX8MfCUIXUfXWKcQVptSL
MIik4x8SZCbWgaE3LlI0uB9V8D6oqhCEa4U8P3DBN6UbidtHOhRz3lupWQN1P0GOwMCfNq1sWmDW
2wzFQsyUiQ3ffhd62d6ewRCZTFiY+e8Q108K+NQMXK2I5bGrtbObddvIIBAYwO3q5az0fgRbsnTx
jszBGSdHi0GwKoQMrdyPSAgr/hdV8nGCp6AzZzeeNtaOeaiBmhsRbrY6Isi4LriC30DxgOiCKHEM
DqJ0bSt5N8OcwfmfzcfEvibsilF9v55Kk5tv6IwLaTXPwwDJnzjYzhZyBtvOwSJyRYp9XREKeehz
CSLUMddVg3TGoO12P5WxCBCAQrEGi87Phi6ZoLvpd9Eb9S/fpxwjbG7/PzXhoOplskaakWiOfl4g
igjX3UhU0Olbes9C18GUpHL5WL6t5jIDvb+PGYFb7OY2msTHdMK4zsSkKzJID1RflNYUgAmF2aVh
IwNkVJIUCh+yW++4IBilJfHp5sJ0g3WLOqjX4ueRwtaVAWSMEQUSlv4dMTEGVcx4IC7x21MVtX47
zu2U+1jjVkwTObT+XRUEAK/knLy0KRrW8l86cL0LcIDwHqoYXxxhDSIF51LHL4JBN3tTxw4PgT33
GEc35cVoBpH9TUAbXwL4KBZKFOHrr9EieMtT9mcQ1lYPzZWSIwjjItTLNaso7WrrkeAMjdYYZZHe
p0Wk26+TCC8zdSHJbylvDrlvEmDuoRmBX8YZwTASNuA6U7jgbpgaLwn/m+AjnqK1RwkFPVqzoR8j
2Xk+aCOGZr3aVJlDyaiSoAUHb3Pg2FnLCayDqNn01U2IXuNCZW+ABiwa9qRTSbQm6gtCYNa3yySQ
IOs4NbMaB/3dZPheOti/fBkU5Kqy7qsA8dDtGXystSJ0ScF83ctT8C1gezgejGpdr/Db1N1D9Kuz
Xfly0LmkJDy4+y8/1CqN2SJ4vkoXrKMLO+zy8Qtal7vFxMlWSl17dFcgjOVyIpwgjNRRBk2E5wtK
wu546ugI8PFI4W++au+u3udu4JQ9AXVYKpC01Ld2cAD32f7k2opfAHMjL7d7ydL4Gxx+s1geTmHQ
xgUV+qP6QA8pRMB7upsqcjm3eFAdjC+05zQHivDD7wiwLDNFP/w4tBOqSr9nfN73xt5NwK1dN012
W0emCXWna0KMtL5FKMeBAql5Uo8M2ayejKdgVON6Rg7Px5PdwQXCzR5LjqkajfAz25CiDm2pdYiD
wQFCMaaAIS/vYg90o0kWzUE/hAvunlgpMnaSiHsmCXNRyZ/TkP2ryLuld9ucQQTq1mxUAnBGZmvN
YeypaIO7y8DUMZc2nqfLKWE/n6qBF9M0MWizhMgDro9PqbNkXXeA+3B8/9+4yfC10JvZnRjl7eJT
A0QiT1UJXL1yJ9Pf+9E4tpliZRsDJiGGM1aMPM0ssDdDUGspxZ6rNTEw1AL++EhssihBUMxHUaZ3
IGilDuLarK8/dM+fGty4e48aBJe/6qB7m28k0YyirL2BtVz1w4oWDrmFRoc5jyik4idNNuZMA7vW
Qs+OuXypgFN/FYNQMD1MgRwqoXlTd7ZvMRg3vjaF9shp7VLvz+huPjMzki69I70w2gSXwbOI231b
A7qlD3hTN2k03qa3IVvFdbTDAcwJ/XSa4tvF7tM87m9NhMR99WmpRSp8q5UrqEqV95SChNuQg7jk
cwivcYKVH7po+qlzIOm/sJ032OraZeFFIsNnoBwmSCg9QLObIHgBG2saOFXG7h1JeRVvmIvKE0Fd
lHEFoupQ3whJLUeJjtZY5t+qA/Cq2DUpEGLKvT+/m3E6qDE7BKhH5ARtH3fOFUxq9I6+zJh2+WKs
7cneAJp2GJfq28O4dhIt65gQ5CWR4qZYGEQrqPF5uKEsCMLpNn6eoGsr4ge89r1qpzxbHWVAAXDh
F70PkjaM6FMtHypMAvZIVjotAHLcDsVgw7Eh2//EXb5UV+GYQaVAcxPlJNQJ72aACPnfDEMsDcL7
IhBTPJVNKeyRKr+0L8YSecgcu0047Eu+lcfFhAygBae0v9haKGJAl6yCo0/dWCFH0SNjmchrokpp
/LVvjnP9F2E5J0pM2vRZHvPa31p+CyMLauFHBM4tl1mHxEcvTDEcQF+hZQqVMWXZkLjTocCKNLsP
wS+aCABjEUWbc2yUAaFMpkLlQVo71Z/HZhSgxvSn33fyugrs31DmQEGte1vh1h5GMoMD+6EeQlhi
m3TtYfErMw6wbJL/1a4M5KEDUnI8/WID64rzQeE10OnnxHOUiJ8WWa+cjrjWBjUK6efFsuOWyisg
WVmVauETNdXu+fGu3kFUM1E+exJciYgnvTwLjyUiIKnCM3yCF7Yb8iRDn1LKizUNtNmiON7xbqsv
mlHLzyp8tJQzppoBNzbP6J5uP8OyGryvEI6REIpw82bCPXqHBC/IOALiUxiKwbuEgG7FVZ2YXHBU
U49jQl/KgV5Ny6Vuyk4zwsSH69dlWMvg2gnVQZjJmJmyguDQxU9i5epi+p1ni/hsmy8w7lRQ4sTi
n7M4uFYOkq1WoWJ/t6r/2s73nZ+GGh3Ml4RCDIrcWT6vH+KDZPLZqWLVIweeqaXDNTr7ywf8JE5h
LyZzjGzH5mWBbfGSuOOxyfoU9H594+L0DW0dJxhEX86kjPYpFZz+vEF0mZBizLmM6RqWmJgNGxP6
edhOg+Saf5DzYtMcYpYQ+ULwLh5BM1alpNut8ClK1ICREXGqnRnj9MzZe5jMknuBPGiwdq8hgpDe
E6SzHl95KSC7lV/BNqzmkSKTb4vE2pt5CxegiM53nYnFUOy8pyO2sm9Yj03wSnG5LxTsVIGJc5m6
Yi7+lYvXWfW/f9xA4nCbT8DAmfy9ghbtkXs7W7pFo7rNBiO5cwwlsOr6w3WyYuF3PUjm1tseCVU2
MJaCNDoRd+CDVsSW55yJ81lNT9MXrngj5iaHuJGPgB4WU8uUK/YBb5RDeKEvR7p+U6ZDD6uoVIQE
QbdjGQAHjhmsL1WBiJ/sKQGhbkXnEXYgzO53XwLTIsodVaFFQmaY72KEQYs8gVCEgczxEKJ2hT9d
FUEEEv+zV0RAB2jBpD1Z0hzgzafQHEVvCNwszyoKEj+EbZ0ey27YXexeYiX/F7LYDKCIS4wZHa16
gOfaCJa4VW4rFqmwXb+UYbRc2hvRYPrwxr61B4H+USIG1vcsdLB50wNjY4fd4Zc7WHsYqAD1UkVF
fljiT0sqIVnwke5ACkc5kVy3D+sux4bBMwnWGAn1xnX0iZL6Z3iAz1ZgTzNoLrfr7upi+5EqgICW
hD+XJR57AqumVoD2wLoHGmowNW7rk3aYUnPUCi1krviAY78RtZsXe9RPIq9MW2zXEeEwnlf7Akzw
AnqIpREduke+/fmtSsY/FXLvFTV6tN0NqEYBjSIwEJ6B9Cjh6jtDlY6RQJkQTyD9V3g9ErHmR6Kr
p+t7u2JBabz8GDAOYfGxJsWTTJtMmp5/0dCKEsM936dYPSjbrpaymQG3hAggYX1bw5QyCCh26g90
tJsBinHJ5UIo1eAs6GrLdaW5KurlwFxE84JX//RVy9RjGgrUg+fjGM+cUwJnMjBpppOWbdkeypRz
ASwqM8ct2IOX+mPovhcLUj07QogOLvxFpL+gWk1j3TIErK0Zux1UPYZQoAMCUGiB8bTd6xaG7V6Q
IPqtff0xW3+GnYf7Q3klZmm6fQ0KjD6CWmPEZP3KZBDb8aQbqkBvbRAZ821uePByJ8o9QWO7y7Iq
4FQqE66FjqjXFeyhPUxOF3uY92dkGI5+moWpolYpY9ChRH3ETtQJI4797aSAXh7VvX2tU0lEHOvq
SURRTIAcZJ8EUeNLtpJWc8P/n82kABROg3zq4DFqxniOnvqsJv2lIdE5wR/u7On8BXkpx8ARZk1h
cL0Ke+PKVJix/CbiENWRFUb0Ac3XohxmcxRd8kDylSyQi626v13qYY4yYL14S83h1N6rMKvrHZFZ
MX6jXcCLRqG7E7gs4aWA3aNvj8UekR32tWGjTobnTC0mkd7msUGcXms3ycecAbbWxDB9HUu6SfTa
j8OS1Iy7pkR+eqLeT8PC77CYVWrw6fLw5waIYIe82fA4/AyHyMrHWeTyPn/+ZWqGHsTAqsPQvo1q
2701RFgTvPxR2eH7m0uBrFHOuJdbQyRKA1gxia5dAdFGNzjruF2rK9AcPhyaIS1cVX5ctI56ljLx
wPfxtNJOyrzjWACtQGRfdMAPcK/JFslFIgfPxHn4Dr5Iu3NIM9lbQjYUe0QRIdwmYeG08OAMJNS4
rkDvAgf9gNLlp+yBPJiuH71uiopWODTjF0UnS3cAtpA9qLGbRa8MZQNkxLWbwO4/6FLuXS5l3lty
pf/WNHvrFBGgtVWL/na8TuP6p5q9h7CcI+GnQTLEap/kRBLKOIcqA1nm5aF8tkihJkEYO56hIYWD
sj9/acJL/0kUop38LKGR8vdUdkvU4exXhOUJ6FMcZL0LX2xfGn2H6hQR96k7LnfbL6La8eLt2o7r
kwOEXx6uw2l/KZFh8DYAbowAGcuQMSctw/mtk0AEPpf4FtID525dzDMaeHnejdX+v45n3nWrDHCx
CXh7OKsVHT7vp4uKRWNjquVofyLTZ9DApxsiIcH5Qzv8y1FkPHNjY4IE5A/X5OHCz/wrQRBaqdBT
+tEp50bo4Hykqtn5t0wkaskYevYG/sYjPtdxj31+0GFd7hDxXloSVMps9Mc1Jr7W/NwyMRa9mniR
7hUXftesa3qZNabB5wulMImRd00PJptf74F7FELCRoZbUxfNrpd20qxH0iSG18oupcMsOy/fuVbi
azUMdZCH5h3FyluuVfBsHwGmJQQQxBSmkNx1AvRoeLmR6xNBPj+MTswz0PkokNGrJUaEv4rWHR6k
37ZHnv+GzYR0QaVp5wt5oj+rYGBjRqcYfirbKSeqdRaLD3vDBIZGqs+H2He35TD6Tfb3z1+mkNj4
GmXNHXFC7NuIeschux+z5kCRzeqI102FVEKYPVbhWyWxbNl1/BE9/dWOA9WCKea4rdWU5PWZdlTo
17QVrM6MW5bJu+HwznQ8sRF5ET7JHSm85Blm9CHRetziQ8IfQZai1Mhf3Ia3+dyQAib9a+Zm3lgH
z4EnZCo5RptowMO8kgrBlOtPwQ6zjEmbR4rKPSm3niGX388X50LVPgiHCL8f25NtpwOeRfKnQ+pu
Tr0zB2TxvpKQcCz6+EG+ZYG/cNTEwx4BGoUlQIpKU2mQNf2P5kNGu4f0B2w+AvkUhXM0gkgx1Nsv
PyiWCDh0MiTg1FX+TZdnbfzlsVshMrcAMlXAM67/7htaMofjSgqG3notwiCUrMUJawE94arqF4bN
Du2Z17qIEeKNB8z+WLxZHHxHNC60LOgKBTXAuPPgnDfwcJ9nE8G6U1YjT2U7ckNhGQeZqsiSurp+
ck2X5Y8K+ilWqjGFH7aOxyp772Nf92L7Kw1SVxV8wMyi2j1f7v+wU7fvdGYqbGe3KrAXk+cP2rqq
CfDasJtl2t2vHJZ2fnZFhB6fOrjlLz9BB03HXlt27hqN3QdL3ZcE+F4nJMlGfrrw7iZDsBlFsrJC
VjxFg+SoiVMW2i2TUyDe1S6UN/hKlxCxMMHKQ+kkB+vYyTLD24ft3Hmqj7FG7z0ltSd+qPS+j2BB
2u5g9Q80W1Xzxzm+qbro2FHq8NTh0iTwWOE8iWC4YDblOmy1j0egXNk3fEnPKwVk9oRv7Siy4KqB
NPBkD+WZ7GzqU6our8y/d8Oaw3qEhPfhnIYo3AjwfXOn9WP/e3QGpVJ6Sjp9pRySP7AESwUTZbOy
M+aURguqUd+WrGzMSIOyV4Q7HeD+44kNWSLv/bjXRkiBI1jDQ3+5reVOWWZOSjlqZJz3s0WVAAph
/6WECc29w7/M/SAGYk4krPwIRQ1ec7DNRnABaa8lby2W2ECjPk9HXK7YpLokw8pTqs24JScPpt4y
9L68u2B+NHbhVWyWbldCGoIRMxfZIJWaq/lnDHF/bw9u9Ur897lUQlDKodWVQ1gMKTAsJJ0Dd+G9
1uhDB5Lh79S2HSmrqaYDeqplH3XLuH2v4GjyxCnUvVXuJgWux0RsDAekSu61wqqAXV8XpQ0rxTDZ
okh7FfE4CjlLw1D6Wi5/vJUUYCGwb1n2BBwMSw6s9rrxNSVWnTVvPTt4gXE8xCSe2NGNMDvtGGZ/
yGEtRxZ8SiL5t43NUlTDkVlzGUcD5yNSRzeTYKuKcgJ7UxVy0a1gyJi/Kg4lcwVoFitGB7xPt1Sn
q0yQnmndxgxLTvfHRZzLrcDsGN8yZWGTTkfcUOksgT9nhCJrHW11HsWNedG2ICt+IXb9ZLPKeGm7
tObs3Q9dNZRfrufhHySf+8fekeB9hoPTvW/8mx/iOnESwTzpJoX8NsmNcR9+IMkx56gFc0SLX7FJ
XF5Qi3NQlVvMt0bopkPlovG88UKR2jRKxuKyVCOQ0RC4Z+SI4SSuH1s48EXCJ0BYPdvggIGmXjsE
ZZNIfOw4pJJ+gsTENdA9a6YQYIKt+TIjDrgzGUUZ4/Nif/Km5g1vMr4JqUSADHzt5lBVhuVkvLQk
c2zUu8JuL1QPEkyY2Sspe58DNmL/mD0sPHjz0ysI/g9qUmsIHfRkr22HtS95kM+DEpczPYEoiMF3
2yxIP2/I7fPdy9OiJZN0v3etO63PSjhUFKekFMBxInFc/nq8Hpyru+KCrULkkBkOzZwiPjfCEHFG
plqL0JYAlyq9lNH0UNeJOzPVNcYD7VhMARVllRMtnaP8WUKW/UQ2H0zBIDpd2c6WsofE9wvEzg0C
MqN5Z/g1UxyTl+ZKOnh56TvXDncSoZgQlKVBVFeYwwk6j4i6cujGS/TxSpYoFDXMCQpGHNLh7t/k
yZQSRaphKMdGzbIiuc2NAMY1DK6sgYId3txyMo/wCOhaSmE/8yyhqxgpMlTAfXLw1kLg3ucPW2u8
rTtAyyAAzWF80q9fhdQ3J0RgLI4gwV8BnoH3+gJJ4qJJmEqXBu74F/LTwd1CUa1SLuUKxcO874PP
lIVVY+JwFcucbCRInBPZaewtCdUNxctJulVFLnk4SzPXlbti7R4ZNzj93tfgOBaslgqzMMMm5Z0Y
AHKqzh8Xd2gQzZmrttcNgV758OgSxZJHZhHJ68wPyHMDRr05OD+ItdWFyhWN548LYJX3gZu0rJiR
BYfPyNe1SPGs5C8EpDOKhXeJ++y5KHHierjczzVaGy2iW2eTWomcVW4xARw3/ycXbq5wH2mZWYwn
8N/WWw58EyHcBizzSd7ySlvGTxo5W/mk4I361fpWfErTwZPeEN4v50VbJWzMPAwCvhMamII/tUhI
M5M8G/5IDoLrIynOAv/mlwe1snhluE8mRjMF+GC0r6dT+wP9c/YqHjIy+WANFqGQfq2Y3rNAQvM3
PM1RzFsno/+Z+1tIsjYHI8lFEN4mEO5pB5DsE+27XKbdc5Rm+YYTtd3jDL0FDMvJQ55m0pCPf7Ui
1aGiKihOC6QHLF74/HCsVnYXuVVKznJ6sYzPHWwUsilASY7yv5xvu7E6iRyyP9Xptj9DV5mp6SFR
TUIcO43qOQleRoWDii2NHKrpoO7zzrMtpoxkvWh+1prrjqgJkx7nltWcd3msbNRqR9KnYpmrb/0h
+kqzBYGBhCXnRS7uUVOitHyWlK7aNorRBRdAbu7U+hMCvjmc8J64yJepH3tZsSOelisHMCU66bR9
YdpWGBoyiUUQ0W42ngxsK2QQfzcE3ZoCROFTVwys1Pu5ygGaVsQiiBrlNOMg+tvr9Noc7HeYFkEt
Y9fM7zWcxjR5gxqcKhxkt4DNu2m4I73fLLIx3XFcVLndNghzTvrukV9qywmhDy9KAVF03wFmXFsU
1+HKEW48WB6/31P0vRSLujpNE5EbPSm6BMNNy46Dh7v+FMOz5GqDysRm5gI/kfiyOB81T3WvEEbr
Bt6UrJsgieeb+BVBmxqLcNhHxQvkpTMMIuQiH3rkfs7Koe3F+/Cgt956BATaU92rzkSY1ufsS4lP
u7KwgBgm9UzGiZ2WNLp1o5Eze35AO8b6CcFD8RwcM6w4xMmIjFxU293Bj3JWxcULyzGg1ifOhH4T
q9vBxTpf1bfNQF+/L/wKaOd4/HmtF+3CHthZ59I27i7NCs3GnQetDcnVGFyb4TCUsrvssxN49fBz
S4hbisHyvxTPRP4NrLod0QsJUPL+LCxTc+HgjvADC7BB4INcQCt33gEiNp5IT/1SIXI5uzR/IPgv
buFVuhKwRJdffTgfIkN5+Qf2ZJiAqdVZK7tmh0Hr/p1W/Ft7Cc3xWqdbpj2umLta37I4iXLqPQk8
cODVY9UDrarxwvUVrG5hk8Bgdv4vTbIvqKlaf0nqRiSsk6xRW0/wyxt90/KNMwvCMzaA3daA2qwJ
WHQhVBxfarXNtdtFFC06uXIdQFRZeWWTWrgpMMn920O3i0nLZmMq7OUTuhSAEiXymd+0kTth+C/o
FQhasnCB+1Z/xBz657G8FGgmGX1ImZnX1wr8xlKSDQrj/2SeX+Ko8avXANp4g/E/lCQq9VhqvCfA
Fdt+feFWb/6pQUNsC7valbVZyDQ245Q7lGDjjdYuzlC/ES4ey0/SFeXDmodeuKTOcFyUyjDQ38WS
U6wDR1M7sCjlf0igopogco9zeO/5aCJSm+561xAoDGKUw7EXcuLTsKLd7O8XgFihtqjQVADtvXlu
b/Gk+XDTbDDVjaVUoFXIsK5ldKmdVt81N5vIv3tvHIMckazfD9skVA296om22EGIMrfcqoASuywN
K0x4ZyFYNpNp41Rr8CQ/h/B0g47QLZUjtNCITdMqkC4r+1G0oJOhUU0cj+l+tjAlnH3/6DVRsKUA
jbs8qQfhPkDq01cSaR6uuZUEwIUKUAejqC5ORIRojP64ARh6WL4ZjaDMjMgC40nGFk7g0+GRmei3
XLswHlHuj4G/CvdngT++ky32kySYo1t4LZ6DTfhW6D5KpmDpISMbvPnnVcBGg5cgCdK+YPD65cZT
uX1/aPqylcJybIxc4WntwmPifMlYkmFBeGmch6bl2NLQbOy4SRTv8JsBGpZbHPz3O2w1Lf4d7Cik
65MxpU2S24kb45TDGUQeZNjLYDdDAe0iigOjz6s+hRzPex72OuMDd5h/WjYQwnpmlmkiPB1jGoRY
9GSh30VjzdgZam3cplTCRVKei8ZgFCUoluSiXKltRNlgPcd6rzICb/hUTmJc2G8fpGKAH+UVyIpC
opCUsXw0poZdCWxQ9qq2c+iosQm0uN5cPGHnvmSsvY89DV1AyzVCJoGC2IDzh/813GQn1nEJB72v
2r5VVngejFvTt2mtSoJ+na5whipi393JiwRaOa2Kxj/1b53isp3IW8aYot+c7TFFmac/lhghNP3b
nfqvWRkVpXtvGfpjQrhoZlQwd4ixPXGIzzai5AE9HMRD2+frog4sF+1/q/2itf4r5cNkbkkLj3dJ
gtnt1p1ComZK1FUP05zDOMIl85wrlzyFrctsOQ27lK+WH2VkpsZLFWbvuf/NwuKXCwi04hZVGtsa
AX+GFB8Sxz+PWJExpa6rOCMyWo5YYPBF3W02hvurmnhh5zSymDvf+JQ4VlncUvmLKGqWtV6xzdUo
frCDVo+kfShjKdgq6fp41n7++4fcYh/aZa/VgUHGP0kiz4nVxvywnUJ2JCSBH3g6eikbC2iIcO83
0PIWiQW6O4Zk3R2iDBYdq62G8ou1kY+udiQxmJIUiCD5uJ76AFs5OqPge5eGnQCsu3wbFa/Fl8tK
g5mgdp3Njcs+b9rfOYF9A87v5wxe31NseQWbZz+zDBxGV7+vGZOE4gCBKrIIUYpM2vBGDvqEfyk3
WXz9qBjjos70fmH6hr2bWk+bOZRZyobORhZVcICF2+QD5VNaXFDvy++e21jsRyLICFX1ruwMObhW
e9Xeenx6dpgNl8h7pHHOtOggaA2AZbQyHdt1Z6KVDACNVDCUcKm8ifK4Wn0iUeLbLDQBWbK0QARA
5qX0q7ASKa4ahihJncMyIP1B4KitTT9uEXYfcL9CTfRT6XnsnMAIaelXuP3fUzEAcrAVGA5cvzZy
CV6xuLgLsEfKg0kZbpvQffFk4Ym8uFA5JNIi7Xwq3S+tJiwJ/SCG0gMyjgIVotbjEZHNVntTu52D
zrqLFJZRQnzXnLFhOQ+UVyEj/oXzSYQjMUUKv+mq6CZERCyo3PLl4AhK9AF+maqnM/U4KQlEtVYu
FPezK+bBjU63qDOIcFJ9vsThwgPRVuNnuCH1cQ1CWVzBkQs3mb+7MZTzKN3XrP5u5g==
`protect end_protected
