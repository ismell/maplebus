`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VZz3gA1OEAo0GderLFN1vAy9VjW6GHfNIvzuIsiYL4pObhfFuD92v4JXddeUi8Mb9uiE9mWeniAP
6axurY4i4Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V/FHqGcuHkuQA/mXo5Z6hby0fYqv5HdbLwzSf6RRkitLROmzZ7kuem6lbOkkdKPEq7el37wV7LLB
lS7Z0SpN6+NFFxvpJwmAXsxAlmNILJUkYM2qy3RGTd18wZzOLOD3LW/CxHw6U/8KDCIE0QPR7gPZ
MonMc1sdRumiZxCH6p8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MhNvJyoQvuBNKA9BY4qs8iuN6gsubuCwSLP9+9HALR7b3OaTr2NNpcJWL5Z2I5y4M70GpNsDLMPN
9x6xxl6dDjiJRZECV9SwEWPnMOiCoaB+AsXeT7vUUtbJNztLP+IJM8m4GxoaXa82G7GmovIGBV/w
4I8s3WETrKiD+AzsZGw7+K2Rv9qW0odg0raG3Nf3cg0Jj3QVcFHpKgJBjvYUZ5EulGHRyU9ez7w6
y6RJfN1K1RY6s4t66rCqdUJUgL6zuBnooS8J3bfZMDJBU02FgqcqfaGv3VkgxhqebXTwUHH6dt05
XvK5nC5Fa8ivOVaKTCai6uvlheV1U35wjc4UaA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rQ7j2Mp14x4heUZNN1sxi590D3svKV0yVp+Er26zbuDVzZY2es4L4i8KGLZDZgWNlJ8KygSbSSmu
AMrgF/9J6L45adeffFOhMlUSE3dKMc9uVglmHX8+NJzpjX5dYFIRPf6r2tIEsYL669q5VkCA/E1w
OYrkIhxgyBWc5KA4bdA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XSzu0gCO60UCezzrasTnl1P56lBSmB5WoyDnA9GcGthkxKlRJzbd5G8JQBmzgeQ/X31AQOI/hSSR
0KBXcFTa4p7F8sfh56g8EO9ICdlNGlmK5lwucB30KgGIDn+D16gBT1WrdmuBInOK9hVfZpKxtH1C
vNGY4AZdGokYQo2eE7iEU2Odq01QNto1qz8mklUCahoHRhjnyHMerh56TbVU4kjgnoVqlDhf67S9
1gulUL5I72iVvZt4D9d+OrnhSSYIHIsZQNCxGgLPpQh16jelRUvUb8ApjVQqxWWD45oYQxzToKeP
cjW5Qj2B5xwGT/QE3ivcnwGi9iOvHlavt386EQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
+SfTMUYhoEZEGaPCN6exMh8+5eINx+9h8XenvZKnYT7lUL+SKIud5B7JP92jml/r022nFvj8ljEq
tNdfF9RCQGGTHNZFMjYkXDv3AR66TL+QZKuZLZWXeNcUYnnD9SKG2ktEPEeV+OTH+i17D0dQ4dc8
bTXU52lZhc8JkWmQWsu8ynkKhqD6BWq3HkGOlzar6pn+tCzd5YncrCeF+VThPMaAk5jH3m3g/w2q
shWfF6W50/ZK6pWfVJaEKW7U7W0hPjwY7YHIv6wk/4Jcp8Pwd541tlwVviXKwQjgLbi/+ya/aw5Q
vYOzlQORcZtlqJ/CeO1zAkrkbAcuC9SpMsBws6kEA4yPxooi1EGUbBxQmv2usaJqoZPrUC4AM3s7
XVmpRjfyfU+u6hiNSKCJAtNK8Pf/ZVdOKrTF0UJegfeiZipCFWYlhEa6Vw0cve18V7/celtgL6Qi
02dFMt1MnlCIdiKBeINSQhseONklNm1inHBg2lrRZ5XuOdwt6AR8DLy5LFbzz/XotZjUj9vBDLZ2
8k58WFKvW/AWi0Ljwb27U+NmazCXYCgQH8iPRWybUx6am7q/HFbgCTWVa86R3uAGU8Kz7w/SiIGA
ClEqs+5bCxCY9YpO3yTjQn7JNsxMI9G7lnyf0fwoAYJYILxPy3de4EuZX4H4j/F1DKCkUZvShPC3
ng9lu/LnCGNXEdDmP+kqccxCtS/ya/YdcnB0JXG2jEDT/XhPYof02HdktePZVeGgc/+4TxPYBBOS
YkYFkpf2HK4bAOWcjQ0/YMGV1WSGkuheG0ZOAxxJ6QnZ/2u0i7FYir6C8ndwT/WNLifbO8aZentK
2R/AcYVghfUw5wkqdhl1payu2drwWUDm0YaYwdQOT+E9YK0srOSEVIU2Wb3/33y+ERafmZ2VMT+9
Vp8XPrDUnJbmDnK3TfxLCXjyh5gUpgnPk0dSInFh0h9gT4dXxO1nRA5535HNxGNq+JOxZJlgrrFm
Tac2CUXoyV7aP0Xe14PldjKnkWjCTIYLtrPgf/QCpSatYDczQQxPhoopicnFvRoIe+HazUC21kVL
EsQ2TL6enQduIEXH+eKlEG2Yj/9m3X2d0GaRre5K/fYk26T18/HQ5cYn947zFNAZVa72+QEm9fwg
qFuCAfWCy5UFtyUTLsRnSceaWF4fQa4hyE9sJNbj3RCLR1MO1OU+NyP8LCX2SVST+Hh9dIzXWfjR
LtI09v52T55kfbdxy+5YPssCOJwB9+KoUhRmBbVb2oHvE7FnYkW15aa8Uw6F6uBpSBL07NwsYwZR
bbuccv80jiutzHh0KsRxI+JHSj24nUfZ0ofM17xOeacEqnEsACqKoKty2SkeTb34Dng4ApYlG/rH
upureRjAqyOtsFzYq1SxsowaOOcXj1+Iw66GWrs7Bb+dwR+uYhvStKhJjrqigEFeCDZcx687OEkw
SLnCBUM1Jw2POetGI8/b3N1Gz0viUR1dgCOMo09NLXUm6aQkYgW9B3jjqS6HRjG4VV9DS3kohLuS
HP3TlD4vytI3+uaMPHfLi14oWOeYfem79e2HuqoUbR6FoUWetnbGJGZe2iWCWg2SINTGFxm00Onc
xLtWRCGasWYBw7j+ZkrHQWiX0k3XIneS+9jUPuq/TegyrbMwzCzwJmvEO/XdXsyuawoTLet7rqhv
/S9YDuQgDFQ1A17sWax1RHLy5o1ssg9RBw58LVCBgqGDJLzq+jrakMiPc25EngaDubDWZhU+6Dks
HRYt2tfBq+3rqdiyd6RSllBQWMo+ErHVfNpHe6/rf90TNWE8zSSGOvzHn3ssl5SEbdvknDMaWszR
9xJ/EhqWDbBRaW9OnSNBnUHHeXCWCr0Q7tbGAW3DFJO9/pM7rw46r+HuxDXQ83YPI/6jRkJWklvg
cOt9/PfrplkSXryD4Mk0mz7XD6ZkRd3UR3gkGBV6TbMrQJjaokzGJidNzBtozgcKBUv2ZyO2UYvY
r1Z3KwyfTVjRo8yC7EtVi5bR2pVuQnxpawgCUqsdXHJEXSNUTyIBJuidg8A9rmRZmbPFCbBvflrp
vR06UPQuzhkPM0MP6OMUdb4bWtCl0CoF+7gCfST89acZ4J8l/jyxZgqmozk2/rY8eMyQZoxmuZI9
EKfARwISgTIblcj2A9a35MlCnCuE6EGHGYxj7g+2qiVm43pDl4LUhie/uY0haizTya7qhEWCMpbM
DHKKeYgAzo5eHPSz/3E35PBqKqhsDxF+2jQvD8TOQudka5xIsbFyYiKIGuEVKPDfwvFr4Wb6geuZ
vh6sK/gef736VMq+NMwhttBZWWblU++N59/kn9QhHjqtXemIPmNjFLTY1551+K2Vp/ReLf/ItugD
2yyELVibvL48exJDhzxlGQSEUL4OrEUzZhZNVijIh2POY841oo4oDbdTpTeO9rqnaPuBNwG0SGjY
aG+x/OVSuvkoMOP7ltEJ8L6frcxhcIFBaCb1mstlTxHxJGV7EuUW6EHMgHs8WUdUCqTygpZ5HETx
XmRM2w8Hp1RJoNUvVoCU8BlmCLxwxgPQyLusCTMf9QU2vQrehhr168+TWKAFvBbOfeWJsXTmKmPd
KoTb3eMQdOAHIKtMXDB+lcQ5/gtr1KrVw2GEaSX1azNWcm15lKlGXwwGK0xpNXwuUwr3B+RXuHB9
khcHu6t89MuCv12y8ScdMdVjcGIP2wGYBpU7ZWZPZN4HL4vOA0Arly72YngI6ncA8pK2i9F6Hddi
LQaYzWJXVq0pCd8Vxi2UtRE3/2cp9IftpROGb3tOkkBSyQlZhMEiHYro8Uhr9Xq3FiseLszdQQMx
2HttMaRSo6X2Xw5Byh/obUeCOHvOFjvd77tWi2ZjxWxO3lIfrd5uHJRkQeeayCbkDt3niDXDmfBn
9wZsGelQgnYjd8TgHTqeqt+18C//bJ+C2ZNzhSgmDKCHbQU5r7j8QkW4bJqTcLidcfmejGwYX6TG
sHT1PdUQtV44faSaQYQBlYYpnWgB18nla+F7L5wt/HLXp7dfNXSTnKK70S7wYKbOuK71BJXnVV6R
tBNKmwBh/wS5EMWfkK8kcfkK0twlzP9xmf0UHVAhJ//gTDmzuk71xXD/7xTl+ds8DHw+f7Y9+kiv
OwoN1kfP1FF8kwNujzwRj7ZFYf7TUTTZLq43tPN49qCNr9OxzwqjmS/4mapkprrsJbq+eoYz2vuK
NlWb/WJdKAsGcI/+BxCWDPxrCu6eiSWQ4eu6/k9rAGnOBWqVn8vBt/UyHtHh+dyKzAGsG3QvqMY4
2gd4ie9rgzN7oJRIs1XVMBJh95UPMozuPPPN0XS91t69HvIzFHpP5LPK+T+qS6awiHi7PZFmOPmT
r1nrrX8rIeDquQEJg/K8iO4dpJCK7X1uGpKQAG+iSKuJH2hAEZr7aZlNvLEvqu7Pe9RCwJ5PGSs+
+Ldp1BHxGiyVGAaeMiiaTERsKaevqvg1XtjUQEJ07q86FoXcaMjRoSEUv1fUBd31llzZkaXN2/7A
+p8s4dCyQ4mwmcW9I53d2fsouI8Q1RvkO9o/HShVUI5h4sulFO1TxLgXTqe66YnjBF0I8H2JmYif
/N76hJvjvGMn+cDElOAFvcc1fLbEaggQiuZS6oyypmCvg2yhE7CpnBEJhtQTYnxnOCaQQSZGh71f
CUTVQRtWcLgR3jlrIDzSn/CdMP16P2mezdKg+lp3/vMMKF9yUh2s4uoqA5IAREnqFWlwrI2JTvzS
VHpXZThIuSAMzypQZbeG3p5aHq15TRkIggF+Nvy4YK5RLmDTbWobuN6WgwbW4ytxgah2+/MP7Jty
pI25N0+99wprjGu7Nzh3uZJBhEYp9f7jipEtcKcxLFIPbHOYufDc0u6p1OBO8stdPDn7UUGwnJfc
wHL/+gnyGp514f8SrKYJyouXmd2CtKYb56ZudV+J5JqHkDY/+CijaVbmv9gN/NjKJ4t3BxddUigf
WqQ9bKf06UIRucEnFBlNEfFn3kRUapB3g86RcQlvdXCrN4tNDMejKm95iXokAoO4g271B9rFA3+q
IYJ2cnizKxWi2G8uQ3TDGDVUDgM9MrVnF6cT/O/dpLWjFr0cUT7aKXAfI5uC+lgUowLo359tcU0V
KM3Gh3dpRUQJB5b92zJtGDqClPKZcUu2uernXtRtUmNIOeX3+h/kvKjgpA6wbtwvOmoeUzcqCxs8
FVx7vgSYbvEY68IBQqau0V2eKhHscAuzqwUFc8iGVXA7vzOEcdBXCfPrw53XniGVkL1Lh6VKpRvR
yzlYGlDA0ndpqw2McDDAuK1xdbowGLb5RQ4+XNhZ0SkgHzti+H6wMsE256lsCXoA8nBP0Bc22ZjS
fNKrL5pe5pYJsKZdTk/3ujRwb10y2uEt3tv5batUtTXVfaG8fX0Sjc7eXzU57VrikRYFqX3CXP2p
zBRqqskl/YqJYD27C8MSPyPSSiQYvRkDbD4tU38VQBBQTfx+nB1ouonn3DQg5jTh4RweKZ9OEX1u
E5J4jh5+8cRbPJ8DwKyS2WkNrAqVcmdQ5QYqiEakTSvQxDzjoI3Y9a5C3bFzLDjjhH7ycWb2VySI
9MLZdMYWZSfPhiTXOoyrhv0eRXJC4NHAmr2mIKsoTPX8+f7GcvxjgPJUv3Y5QmgSpsXNKAd9zEGg
ZCuVhVChqRvv18/jgKUHQs0hAJyE/Lg70Bh5O5A1UHYA+ITLPzFZKcu1wK+gR6GRDcFDjgaEClL2
lIAMUzPe2gbdSLhFkPMj7wYHDpso7dPLRUt64Qb3YT7VzRkWE4Y+Wv9i5JNtYACI32MaNa0yXTlv
NlQuk4e9zz6sIjdZIY46jNQe3/R1FU1XmtcvaDdUt0tphLpV96QNS3htw57DFiiIgg735LnAtRod
nNkRfjjSrcTTlRdnGE8xNv7qDnI6ZdA3CW5PMmsVko3EVqpfSbRHqCJsyXjXFQynMeItm73A2Y/Y
fmBl1p7k5Pb1kaGTZkGyLDqQGW4kfsDpL2mXaEqnBdIQnxk6GvX5BUPe7CVRQGDzaFKnNc0iNEra
6by6yKqqlRBZqHJfcmZY41k8iRu7/9W1+5LdbopU6m7NaGRsnezmZL3YTfdGlmvGLNWC/0/XApnn
OuUDFX4KhVIlun2a7R501pK9EE5mrpxe2Q7OHv+tOVEuQQ887/EL1r9wVOmbZEHR12zZ07gj4r/v
eFmv215yxNd01mNILTPN6nBP/sNcAWqFRO8JTiwp+sj/j/tPY05YOgQbqMZdf1pPLLiLpXpfLUQ1
73HhbhYKzduzZQQne2AYwldUj5U+oHVUbXuzKDr29FP2X5htlcaRm3IEIXL9jIdi/MbeCajX/VPP
+4K1FuKdaVQdj2Y6PcteSibd5+k6bCUKHVIm0ga+XhspuTi2f0/qCnLmDpzfwoaFYBPl2mUTniWK
ILDX6xcgrNMqjbCWF2qS9aMwIxIRo1Pi8TPLBxQEgM4gvXxTuvHvwluRksS4ddrZWHvRYWT7o4wF
TN3dAHhOBaG5rRdYKVQfGsGx3sr5ZG8S0+fzRv+lbf1i9L1yE6fs3vjkIllRwgicIMr/Re+7D+uD
FA10ipj2SuLYGNI9QrOsoROZnYTXdUathKj0wpei7Gj6I5VO4Nzm3Gx0KVeXTIGM+Kb4o327txo4
g2wRANNCj94bBdBdS+JaPuAxieq7gXbMBcGO5FJ4/waUt3Ln4LwGH4M1sM8INl+fvXegoryAIGI1
fdtzL+PdaxNrKA16ERfQ/udFQu9gAnxA5eWNJQRgAnVPJqRetxex1SC68lsNkzw8o5ihh4+07BTi
mad3siJogE9rZmlpUZ61cNHUBq9TJ3dX0IRcsHY1lCr6dEnWvIAYmBOH3PU4hPTZsA0rBJRDslc2
NS3LK5cTeQ5cY70mnZoqbiooWIQfkSxbkUVz8X5GSnhkbcggF8oeYZn5e8qhxDFsgubhg08hID4F
XtwO7TgGFjUIByVg8WDhOY9tk82WHZTORexsnDru/hUnSFh9/KYLS/RjT5n4noJkOX+Q9wVORzYN
/1rQ5lMHUCiUqNSS514hLGyaRMCuVEKqd7QfuGuiXXWrbgEdg09sI7WHKf5jQ1Ei1NFE2ALzdQjW
1+AGnHIkzviFMltb+IpCYTPNtxgO6RXwDht2UOVSFgoy4e64qRYvo4cBOtceHkLn0v2av8svQwVK
Bb3FZbdWQeEvaOmoKMcIp+fDiHkTKyxMMI2CZRMLaaQytHiOGlY3hfQwXjaEk7x7gF2jKeYxiUrA
Ul924JabF5zfdtH1qQSuyL4If1X2RJ1FHK1SkWMQWHfGJZfiOr1cAXZchBua1Kn4KjbmI7BlJ5UR
cRyU4q7gikDw693gskJ93s5DDfo+Tq6zqXtFHZWaPTTsdKJW2APoajp34C+D1ZBlhI8XfIQhVyj7
NR9eowDvgpiPKPWNvPo4c3xCKLiXRIJQI2DN82whv/QzwVUD9woQdio43jMa+Sv1wA8Hz79iH7lv
29ccEzFuieyekQ/nMBSH2+bXhxTm4tbgculG1nNxz8rGg+Nd4fDQsRqt1+b/SQhPXnmQqwdYwO/Y
AbK9zCUSJVnoKOIgxI2DJqvBmUQAHRTK8muMvvgIAfuWRmol9YGRuHZbyl/9Cy+CgF646eD6ln/f
43TLV/kunqWljkgfTvL3Ud0F4p2s0PNoX76EXfQ/dl9Uc3T4+jDyqSHNQofgKgvO60YTnlf5Ggf1
OKfuh7jOSz4Krr5nSYIZYvAmxzA20qCJ/9H2k/MJenIsoRC5STXb2sk1Hn6pN6Xjz5URPa5V911q
lh9njqsDzMQh/anNR7tA2zG+AucPwAo5qd7DKM2CIwQGTB3f7T5ZbxkL6NQcLIl1H4NsEGZhjhUv
jqzhNVDIDWDyNXr0ukyX0nNKDn9JutrdybRKqtEDvVbQDj20/Lbpuh0nF3y5KReCzOdG+HVB3msm
/tgOB4Jk/DvrMCFkkYG+PEfhZgOrYkQvvcRl6uBuM+MVA8mDwd73cq85R4VepT4ds8R18EKdeXnX
8QcoKNnzJjiflWfUZqu+I8ykhrQ/DPq9Mc/WG+NDqx5Ui6z3MooW6+BOce/t4QEpM+fH6NPYRg6Z
NIHeHSddoV6QlfoB8dA7m6QLzE1oI+/Rf/69mUNmUQIyA2sbGJJ1/foQGczdJt8V2bgkNjfcr6Cs
F8rbMeJB+HzI3fTqpwqUhwTm/WDn5pFVaoa2IeX5/U/J9TIHVDVPngW30bO8387rwBkwxBN3D7sR
wX+016uKcwRFwHpTpe//fG4RDrG44FgqH/QELydCv+EN2TNUHWOjk9tqZIIt8tB0w0t1Lw3ZePhI
Ue9IqarulW0A6hKKSraVXOZ0iYlA/bhnbooE/kQaY4Dul67QWfbMhQlavsxOds7uRvVp8I7LUD4i
ShAWIoFKQVBDYR/adyNIfrHvFv3zdJCWwaJNfpsdfwaOrnlekyf6JA9DyaOrsYCK4xIYLPmRdTP5
BcR6EX8fi99PHlOMtOgMJ76knKrzK7nEDkvMg/duI0UsoUXcTk9MvBWpo9jQUBoi0+uVuHauWWad
Gpq1CvpMxYB2esJSxl6wJb41ewuYdtR4YvkC8FbJK6pTJYgG8+/SzjcpMFoJr1dewSQVuRA5EnO6
wwdlVTVLeJGSdARyGHsN0G7sikRzCqul6Fp2s044HRoyNKY4eL15r2AQTx+iyiiqBSvTwoDNVME5
iMNQJBqkxfcGZb5ecoKPVnm3rfe36t4DMX9oZLoJtdMbariM+cNyXlkw0EX/vy9xY4AB0tE5i7kC
WK3crQwur4Cp8xIzJwzDJEKU6O3Lm5ROVYdSRDWy1ZByW/TB8GsXYIXcRcRPBsJxA9uncV0FwlNI
VooB7rctavoEGqC6/EwVSyPB1jz3NBZIAp6eBtpPXRkML2nYVHA0/fUqgg8a4xmYD636ZI9rHtBI
UOfqUztlPvGEsKbMXSyrYZFjlvgxbdfLL8kTEdATE3EsH27Uy5Ua3V54epUxSV3kFqCRjLIxY/7r
Ds9MEs6tMyvnk9hrid7jFmsvOg5BpHKAYDNrb3gnC7SJLQINXaEBo88RTmULBBNwTV5rc1TQmIMi
5/7NadTE7Mv5U+pK8id+t2o/BDchQPTBtHp8XljVw5k6I3mfhUxrZGQEuYAMBEv0R6OSfUSVmLzo
yLUsaIwxgBCKyqUhdH6s+gXrwMgPd6vE5gVMl71N//I7wuT+XSMSdwRtXED8+HxCTdGygAjXa7rQ
tJOJvJNZ//oLAgRaZb1DUg2nqcmaigz7nA5hqplF8AlJeRaQkPdm1ZZrPUFyVzBvfMNs9qhIzAsj
7/7nLsbq6buFZmG4yye6i8L83V8i9jWtbczWFdnriz2yOpRlmbOzWc/+b5UKNWsWqWNUwhETz73G
YVARytV4JIphmtE9D6Gn1lCW6jqKaZ31T00IOOhRtp1z6N+jZ6Gr3787WV3n/YL6ZzuPjfB+XXs3
0rEuXppcHUG1itQTqKBveI1r42udPmGLY4Gx2zz5uZhvT7EHpQDL8iEUKyWRvvzQmeU6WA/uoftA
VsYTq2xeDNJjA9eqJQSU5oMiAfsRaotuEdQXgmAprTIQTtCkLvpTbkFnysQIisZ4+Curd/tkrqr0
eVtGMUA4DUNpixZVnfzrqdM+s1ANo+jAEbtkaaQkvl2O8xR8chwRrxx90DThXOEDZLz1pgH1RC4m
ymyLawgqxyNgeLXy/wlSd6NcwmEJdcYH7T8MrsEvnmPLzYeT4/a+NQ2c9DodDC7VsbrNnYFsPKKA
nEWt454H/VqxOwCb3yhXqL6vRJKkzj/SLVI9Dh+FSBTIcAd2WH1VWSksk/542EjMHcU1MpXqK0ex
mGTsfi3PRizcvCNmQTmFyWrrfVtDr/JGRVupbZerrFiT4hXyzcsA+yyNf5xrhAcFMQtnQV19S/8H
XoOstvDMoz+F+iD7bUwunXptsc7x0MZfiWtahNR88QsEW2MVU5RUiGa4/u9eRacPACSc+Pj+FvSO
9o4q57PhE0T5WtSP9F3M/LzHTN2QB3UsfumR1I/U00tkZTBqbXNrVxpWush0LJJ7MX6CBsafPxw3
0mj7+DL9IrS0OGDzUoQLM8N4OQWX/9guPrmRIBEoiiuxIoUr0B0sOWbeIM2GUK0uythRMbcC8Lqi
JCqsA91Enoh83GLyviRVIDfehmx8ZMyfANnAvJPCBRE2O5H16pkHMA04JSXQsG5+6hrBNR3pW/zF
ALrDM0PsSFeVekGE+FVyOfjtA+Pq5jThuOWBJOOSLWew07UTUIsFFbT6ZqAYogQumuHzryVCl7vZ
/mjrCFM91Zd2/kp7IrwJMWnRUfyF7bXdzSIRIy4CMaR9IuR1dLnSfvlDuLoMoBkgyZXdJTrz2o2q
dfTmSVBbYZZKhLG2u5J5kyCYckc2Q2FhO7zpvn8UjO9WcjQQ2X3Bnylp0yGmg67QfqvYifMsW3au
q0NqrBkfwPCq1VtloU8lzTrkI6owbbwpNqpJjADfZ/NFvvtEDWSQUeF6tSe8r2/6kXpC6UX5Pxmd
vyakYoc4uQXOXN9rJpLYijethYwN9q/x9D+IztrUrQtTsg7vYYK1TpEIKVQKsyPt5fCHliJI3lls
aRLTHcYc2gkiIqIICxs7VUPgoogf+OegwJPYgiBUXWjo62+ub3d84rvEbrieUNjGK6TkmFSy5ctU
IkDv7WozXPVmR70HIJ65kA2tdmuaaf8XIDH+PeT4C63aZcU3ksnQFDPclP64gBnEkI1NJRMjlbE2
FNZZq4tSQQMYEhIqmrac5R5f9W4pf/MQb2qd7s+YYSEGm7xNtCA8azTn218y9mWkvylnfH07VRlL
3DfrXpLhyA6oQt7UHqJRav+wAXi2tFpRTrUsjohgICxf7xVaIhSYsDz2lzEXgNDlaujFZFT8eA9J
wwqWGin8TItJMXhzSQBl71et2GuoWiKcGieKBxKPGuAwZuJHAhsvw04nUWiNajUGoant9n/fTGMN
BSj4YURU1FfG+FN/TFC+c2PIh9xNIbCmYS1wyE3w//1XePrCcOUH5YtLy03RtZwjde+bBcwc495D
DXxgY9z9ydoS/0IFmWi576cpUgK5CyVCi5ala8crnn4thGB44xU9EfludbiCu4KU5pubYuakxggd
TreK0+e1BrNeJBWrSMpJ4PBz7BTRxN/O4so98b5+Zm3gx4X6iEVV0EB0qOIyJOcpnL0rGKDRp2c7
oAZjXKrIoSv1csopCplY+jwgTgCQ9lGyRPmZMgFch4PhtAJdX4nfmUnsmE6xzmEmx283N5zJm6jc
4Ov96DWp+R8y06wiw54USBXRnGF8tZWJ9vHvU16vYs2ih7kdY3TFBSMFYKtUFqmb8v4u0NKklF6q
1zOw748DDISz3RTs2iTbjQbD75cC31WqelRDG7jpJygJvf+vd78tk7dPxfewYsjNYE4uSMM4g/JB
iYHDTUwY3eMktBrHJsMdbs2/bgMslwhhWhGkk2Sok1NhxFLiRJuQB0QWTGM7IumSlmtV91ACVBPA
4b9DJSHSkGBj64l1JGbLmsTeXnvW84RTssRXilNuL4dCDw7A6K1+gQK4xiZ1u1lbOqrj90BF1tmI
Nvf6ar4oTdDduyOoIXrslGvW0IAyZUgrC9EFAHOXXlW0ag2u1O62cIZIEqyvr3yKs48oLqB85UbO
WxwKNKX2uLbwinaVnoDSh21nKzMhrODL6VcenNOQLUy5LxTsN2R/UVZU/sxWG+FGuvPdmKCAOU83
DG6GQ7q1omOmRgoKvLjXWkuZW6p+lvZiF6vGVYjZQS4TZDH2RsEU/SoaVeB8hsNMJ0L0IxDmOuzf
o4JovKjpJ25o2G3cvFnuqzk9BRcE/UhYcGaBOrU2S3ew+mb2gL5m2jGq1oFhUwsJXMKZWLo1KcM4
CjGlseUQmcsP2oE1haL+41ig8gNsw0lrWm133OD8k/EzV4AcgfUbyAcX4S8qWYGeg6PobBEx0Nrk
xxRm2fV6S8gb0UXYemB1nEzbTbMKYkstgu03kBDZxk2z4WUVYy4baMp8+09tzj6BlD+Ob0Twdeo8
5JYYRS7cxOrupdqeQCPpiYu3IMrVW1KsUX49tNvCOSjG6WmkSE3lzOLYA7qPi9cVgeEH3d7MiCiH
66VdtAViA3NLTVygmpMIZl+qtgCs6TTPhPVLRmLCED/N+nMOTDJXiM0oUxD9c4sKfmHK1peuIkur
sqcxGlpYytRFugwDBsy5jvltvV7fWuA+J74yGJk4vjVfgdDb7ktwCwDY9A6jCiTC/FEjEccZ48T+
nvTSQ9x4YYzav7wcrsuIRk75bo0Sh0SiUNdvsev5uJn7X7vCmtPSpTe9i0GoK6BgZNx6XTAS+yQr
ayccGX4K6+900Ux3ID+leXQ/VJsdF5E4DOYZDf4DSZrLKsDpqkvQCAd/Ks69tB3KJ8W2SdfapI3n
LFfckG1DpqlVsR78cwMNdv9BDcFwkVC0mpMcavuExPVPB+NpPJgkFnNWemfxd29Ue16pef/TL06K
zVH4k9F2ay0XNAmcCzIIrgiPW9qZSmFu6f8eZaDHIQlf/08MbIL9F5kT+juNgOCvRbk/7l886hLv
CHogYxuEy94yzWAJs3Oz+qdqj2VWRtq1yqJu3+v88OqG1C/u3xYfhP/cH3aXA5E7Voy2QBxixe//
p8KHq0PWXr8UNcize1yirxhr9Tr/5eL9dZYU9Kz1kv5c12ySsdsGx1Dz/PSqoNr1sN3MgcMdFQ/T
M+fssi2+DDhaObEzsstZlNzCAUrTuztUdC0tjSu+14IewBjozbTqvETVQi8DMiaK65qxbXrPGrE7
OFPveT8DT+rmYoxzGX/IMrfP96YJutQyi3NCrxwKiXWgQ1dBU8gCJ/gF5+ldJalHzKx/gkK9MuXw
9hg4ObEOFynQ4k1G02W5zJR3HcAlij0nLzt+mieMU05RWfSn6gDagVD1VHd6YfmhSWX9brWlgL9S
IHydcbuTGp1Mk1+TUl13GO/tozr4W7hfE+QRd5V2yZFKpZTxYbNWIrFmzIu76SYtg2vuHSYjl17B
CwEARSDmmVkuiAA2h2zxQ/TWMj+cfqbCxoadN1XA9CwI2whI0MueW0jQDu+V/nz7bp+hhNmsNQyC
8jetgpMgDQDUqm/OwmUp/iqgKJWjNFo9Bte7ML4YQGbyl4E2uxQM7rEhuxH4ftr5oYko2afW436J
2foFRQZiJtRSfjT6ASfhK1+bnPXfGZJtRCOL2zy/y+lhjRM2m+N7WN08E2yCM+yNahdqvBUh5Fuj
D1O8LwVdV6B1QNJhqrrpS+9LVgKtmifQAn9fSoWhoXXdSWOQSTmtQOg/b+5GubJLaHUsrME2Dh6R
zI8V3GCAACho/MqGY//bilVG1a2aI1qIxr0WFg3XydOIQwg4WPfCaF5cWv6Y4lMH3TVYrORABO2k
oJsg3W18MFrDS9yzt1o6RiddEBszhGLeliPko0mJPyijiCg9cU8yZU7/ddBtW8WzH0oYsMmSWpbM
i/TkZfAAiDCYbVZ+hmRqV2R7SYJ2VFxLkFnQ38GM9KutbfrbbJf8dge25NAvw/sW6lGxjT5RT615
ftiyYzDG7p/XcYgHV7QQaqHVNYTdzgceExskkh3cKUUYjOmAqXIOj7H8DxxvqiGzd+lB0AXedIBN
jxy4CHy1lR11gh4YK5Qnt2/GPaWcspK1JYYA7eP7vcX4VeOG0qLrn9MRENvoLClAcr+9KXGGAXc9
OEipNUmFajlRL9+WdDMm/L5IdJ2/ozTmUtjcaDs8CqYFw4RHVk+dUVq3RC/kCSad55qdvsQpv/QU
VTyJgSfzFeDUAIoDSntt+X2ZzMJEoU2Lzqsk5+ey6h7C/pqyoLRrHwHirvPdIH9+HLUa3wgU/8Oo
IbskvNIYVFTDF47MU0m8kh253QW4OvTYk5WSqZplaKORHHaikFRgHb7uEODxGNwfH+JH4cWI+rhJ
WiiF0Y6idFKGG0+QusdlcQB30BU0xSZZISIaI7MDjv87nnDkuQCjMX/0+nteG9Yg8N0BojqSxnZc
UQN8tMsQ7hNY5P9UNGCcgRnDt3tgaPaONQIira2/mTl7HFqD6grzOz1lKhr8qu+wFO+7QMkkiNiX
EES/TANNhodvgMvt/hm9FWax1Mw14i10Sxh9x8fYKebHXVIeeVrtqYoOXaDnvrE1VFVZt8kyAeo0
DUoCK7kdxIo9UHkTAJWuhEFTN6XCmsOXiWerHDcaQFJI8sgv+i/m8aQDgX1xAAthuunapvM8JpGM
jUDJy9Es/lLcna6BquQ2u6EOar61+fVKiEn2ixBIspSzCz5zIdNDBms7YkpLzw/QZ7H2Fx3Eg9Sl
6PWjmmzxyfA7hhcFe39wjOKqQxJdsL5kKGNeSUkmlmAZ3DOM03ZNF/OSytW8sBFYvrx7MlG61DMf
DZNnWIQdtj7qK8hNkkDW2T++afFP6Jmikq+Y7CO3lx+CmwA6UXOGwvOHbFE8itWteXqO8cItFXQC
h4GR6NlQNWsrnQH5Eb7Z8BRlqaeiBkotNzLW1AJspZdU7M7qH/FsmfiPncKuIxVOaMuOiKTdy0Jb
2H/2BvRJ82Yz2D3DfWy4FVr4NE5rNVR4lL+dp1SBlBW4JtZA4WOML8putvakPG0e3Jh5OCpUJPEZ
itWRR8geAMrce5GVrtYBbTF9KtwOmkNeLmwyrqFAjl/OymQa3gT0Z5+a1q90YELKJ59SLrhJe6+L
l9HYZx+g8Yy10fdwSHZkfLuGV1niqCUrv+z1gWr4lkdkru3gf9XZLhZioOCSb7ySrtoLz60HAdkv
P6j6CLjgqWQmZer1Ov9U+iSBrOxZgb//rQkpZDDyTbnY9cv0qIBgtmKqE1a+q9x2pei5KKrKuIno
y4ARYXw2jLD75DZ1qXieHT5Bx0HcXFhfnlQggDWDOGau5jzpt4qj4L9UB0VaZsWLk2iQkJ5huNKN
czoaAHaN1QeOYaPVqlyHmnZ6tU948sCBYMOSMbQZt94yvtJXdYjGLZTkQnIGYDnRhwGXMhi1WIJr
Otap66+BzQf9N6mw/UeRbZ8lGGOBiRKStUTPJ/jsYErawnF05XGLVx1BPMKw2qLCl3TFq7MgtMlI
YqTT1u3iUCVd9vct12mTrDuA+yNCzTN+dkBSVeoceWaTKEa5kLAJHiLX4oKG7jgJ3DhAx2AYO9FR
NS7odjQZ0zxQittc75XO5pflC/hgk7o1D0XhXpB3nFvhhgkxPR9zoj3dw1x/iih45rsNEGhl3Ejr
WMJ/OXZ1hdQcwPsBKOlKiB9kE0iMiBiDk0WYay4UjpQH1ziXtlV8GelKKHD5B9i31hUkogsFczLn
KInbpJZPVwiy/B8jO+9YKJDABaXN8KWiAQe2uSpzvEO+9WOx60mOj7ucVdRuaAdto9p9hqppjgkZ
oOkFDr5g557KyB/86Zt/nsHsLuY6F67VoNL5Xzpyw4uT9NjfimXC7YlGilDIfqQkYrBgo0+EsVO3
DtwV5r0UpWStzS6cCMb8INGb+HWrQdHJRgfJ2EUd45Cg/KeZtaU1MFYFBd5U1PWlh/6KOGN5mPkP
ou1VPx8fKLIvFr7dACTT+A5JYMO00PiespXqokx/JhDMbrSu0lHsnzwIL2cA6dAbgT2sJHNpCHOp
oSfDDA/mB+A1pWI51kVw1gOfytdW4aRSs94/wlHIlIgKyFpm2G5O/P/FE1fOH7TGYwyX7Fhxr3/O
hDLCMpn4PUuxv9zbD/r1SFb0eIel0RSJGjF8k7yL5I1+0MqCO4cTmhwJzA4n1nLTRiE3tzCUZSWB
thM2agQSRJTUjVrGsmtePJ3k/QEE27b+QFAkz43YuXu+NsWecSNx8GKrMtyaF1iXLhoyZdGechrp
Nsx8LOfprQhDK9buSl2oLs7P0c9J+d/hpxJrI8azi+TPzGZi1vbFAH8xYvKQT9gD5zLkD+svWeFW
Xsljwwus+rloOjwJvcOMKTnlGnXm9rVJoH7962bAwPC3A5HsIr/KEYric6d6wjiDzZmMMTJmCUcM
v1H7eRWKEGyT1fFtm1RrgL7MiX6EPGpMqXnqVIgL/TXUY/aVvkrmlYAgOUYVFzsvHlYEOODYHyTk
k4OHkU9shJ9LXqNzgerkUN+CI+QoLv1lZg95rWSzfWoao8Wgal4uviuH51KqWAQaM5Of5NmXjETm
dBN4ai7ZvAWmv8A0aofCtYgaKaM8YYc9cRpqp8BuJXi5uQDM1gSTakqBd1JpGBseKBLO/54nqDNG
b7sOFkN/o+Js4FwArJ22IN+NPkXcN2qOigFapL2pU+UkuKewvtJJTpKdpbRiVRolmfG4EunMO/hW
RZIlgEDCZMkk/jtZi5VoJN0kFaasL8YWAYhRUZVgz6KwA3Gg+5pAV/HeEmUWxIzEkQ45RjpdaHGb
YttXVi7VKUyD9dfxsnxXILBRlq/lsh4yDQG32eAHy9I7p8vEhGZUxaNlxiHOHf2jY76kKKRHQ/0p
aogJgVhXn0Z5+9DpazQlarrnMROV1K3fCM8dizr4wNMd7oImHk5aO8jbTeKXw3ufGHLQ23RbtnzU
AbQdILdh3D+X7/hAAP9tDjyLl2I4FkqQVOt0c+zqlx3Yfq3T0ySYEP0jKP88SX1bY+euWrgzltiy
zA913hWsMoA/F63k6BZ7esASEKJ3/8F938MIJgZrjKezhzTkfKzahbV80oxOXbqSw/TycEPmdLpD
f9biSu4BqLXrerjIYjWyRMpr2LehhR5OZ4JGivhyBuk/IyawHCpnNbogv6hos0+oi987F614qeuw
3V9zmL89txwLs/ac3cpjWFLcVptAhbFq2VYaFrnh2lNkTUFP4IaL4pY713GtEzB0BJjRG3JUJ5A7
8Pp7Xw1MvQisH700mNN9hq/kZTCa68v2ENRqkbO8ruz3bR3P7xTahirP2PHdTYNLH5RyIsPSxxso
ilZCZW0UJXRD2aNVsmuc52/myo0n93SM9kOr2Ehe7zWcb6gNmaU/manV69kzuaTbQDfk6mAq7Ad+
mWeWbZEt9AOdLCqcSuj3V7x8RlohPgIHOGNLhSSJYQPEUEyOTq6dfCZ1Vz4QVQ+Ugwvk+qYU59IN
C8Z3bB6Ya1kwuPeimh89UEerLAzmwzmRkmoS+BO3DxVoN6XUyVWB/6kJ0M7WIEbw6V7xAU0fhz/m
v0ALCwT9xnpoL+pbPy4GrnW+81Rmq10vsD035b93o8oSsEfpanmNuOrKU0RDoAAi493p2KpTy1Jg
EIEc+YoeEH3HEY0CrLJ59YtBejDXg7mkaQqW1KDmUdQ7HICMnnuLmdwB6Xn2u59dEM++FIl8w2zL
bzanOyOV9PsQqxrYLiyvcQg3WX0vxX3lSyAqFnNAStEUDP7Cx0+g1dRMJYDEx7VGDHmWUrgl3uDU
duZyprbnlwn5+ENzd0TR2btOZlJ70JA+uMJh0eueU1kimAp2jMzTVu90RqM786HVyY4ZhNrWgYfA
vxkjPsV7skVjOEE4c4/ZtCMQXb4TpRKDTEuIEfpAeUSzXEDO1Tq22/90BNQY5YpPrP5fFd8vgDIC
LbQvXTUcW/w35CVqGSzhXIbxCIQAAub565CwqLQUZ/4/QSZ8g47ypH7sC8rVKP5aRoWV2I64flQC
p6hGReVzj9x4oA5XEGC+Gv2/tW4+wfd87rmvf+DEwXjDFg4YXn2zBpjacHlcRQ75QlTsmAAN344A
v0dWVEjJDs8FfsmDCVd8+lUTPbS5BKnPaHTCH0sUv5gUNiYys3jY8DPGPIpAEywM8AcL2ojtKrwg
1EGU2SvcRqJZi14l6xPwd5auJFrPHBRZhP13mJMEUj4TjIn6oVhpUIVepyyCXCsumi2sWr+tNYf9
a5umfJoTWpAxeGgv4e517jiZcUixh98qYK+xTM8XCB9vNcWKD5olhsMiY17EPtlgd/7VJYq4qFsl
qsyKrl4ciGXgFj3PekDp3/RjpfGwA1rrmzNkVqp3FuLty1g4sXAsCkJRqRK+vS0VVpp4/TVR1dh7
3qIHkI9GQEAhe1ztGxerCXajygi09ktzjG/TIOfLlIgPHDZ3Zh0HGuaztfBMjlnf0FOdALVMg26+
Lg5OVcfczFQU1sCFKxGcpX+Y4XSERZuMTNVgtR3KPqfV445baKATG5fG9LnV/1mK+OZb2ldc2PbA
vQ0MmNdPFS/bKhdB6yEcZsxMe0S9qkDGZ/4M0G8p5KX3vWnOum4NSVhuX7RwdlRbXnsxjvjgfsMw
jzuZZ3t2NFacrxgkn8TS3xq6BDOVZj6ZpP7D6w488Qc0xCf3/43exr+vs5LAd7j6hzzgCA22NyY8
eENVIe4dzYWA8SBsNJx4Sc2Ae77O8QbzJMVBUfKRijyvFkJEeZlzGtWy+CWsgx9vs59TbXe7Omay
dS/7IQ6w+BBBs3x/cp2ZAQMoPJkrryJn5JorUGZFA31fxOmXB5tDKe7y4ZZUsx4CkjF8MWaL0+K8
kDZT1GMBsTA2pIPh/ELaB/mEZxOk2TwGdLfR7ZAws4lE6dzNuTX6S2l8isFCGRFrR70JQwGfMLd8
b+rq3dG1yGqFnu1AufOZvHws/+XFJFyHc5Z9ZRF062ajpVVOgbb7Al4YidRc7805TqsmN2NI0YKb
Piq7uXR/d94MNHpLQioTs3h/NOg8lfooMzuyuc5MVoMgvyaxETBRAyZ9QJJpJkZWUMqlBr+i5kBb
JpTvxcKCDIeDo/nUTbmpFiOtCNE+DQOO71l4dc9A2UVLlgWSLm6qDlC5zecpLiqh2j8o8m4eeNpi
uNa6Cjk0ISWrWVEQ5IZPZwBADLRGKmae3Fv8tjSGrb2lFFTEZXhyelhtxBonkdvU4vkpTu7iDll8
eLgsnm++FsM2Q+I1oBqyJ4uaoxvP/YFUQ3YbJjlxODKIGz/SwSm98JRJKS4857W9LdMP6/r3brpY
rngV3eR0Yxx56SPoYFgLNH1CLeLyoSmFMPRl7xch2jvFbXX2LwkQTMLhKRB/7TA/Ef57N1ls2mZf
l4SloNmtuX6RH9IItMvKEYtqB7E2MAEYhVc2XdC7iZjf6V+ydloTlDHyhcOXhY7WVFjzHCri23iB
HJvuAwBAGqhG+/Dnq7n1kjEON7V38cAOJzTtQrlOCEHBIulKBsZJr8i9dOB8yZmZLWW0K8lCkfrl
5CGy67dQUAsrcvzrYuYX2To9cKhaynesumlERnoLPPQCUSQ6qzK2vUaeEDOSIMaztJB7OfRdgsYT
P22OiLK5QZcgcWuzzwiLz7/8HI+Ywn9Q+tquiAQgDbZ2TbgrJ0kpusdq0N1mVgiyM/HSobBLUkuI
VAZIe8vSGV1VUGWc3PykNXrtgl5p2xoeGWPa0s8CcHu7Swnj+Ai1b13mqKTIXEmT26xP39ifSydW
wZennhy48GJoWWq/gXTCDkTL8GajUUp9KhL/byUldo/IDE9DoBdzswCxRaBf90X9hqLFSy3QD9AQ
BMERKQIdN7JofkdKAOtkcAdExiWMG1LunHpO4IigGtKk9vbJ6rCWc9riXQ6pP8YSPo4cNynFYv9+
qaLiwiMKozhYyM1YbWXHsWbLYKwskW8OSiYO6nNbf+RccXFwGFPaBtvVCFM6S74fK5QNmjayQ10j
D1PWOo4PDu6h35YkNpCeGiC23pXWgln3v1IMOej4ojKplQ1zQSv2Uzh9+RtTFPlW4g/piikyjzAW
6Lb8Ys4ntJA+H0tlibf0C5JzhJYv4d9M1Vr6bB+aiXYgaszhQPAp/ImC4tCIGVxWc/6SKscg6tY8
p9HMZe20jju4dplCrsO5Ul4xX455sx5six+sliF49J1kO+qfZyUgzgpWwuK3Is6vfQa7tSz8vasb
mgj2qeMOABcP8QWniJgijs7w6nb2k/NI5XXHdYO1jsVQxBe0Esd1czIrUAcWhk0l2SeITRcJuNmA
DdXSu7t/I01j+Yg6N2sSo5OAXxCVg727N0gxfP1dInivA9Gw32KASiph2XEJlA6q8w0ZT7a1fAd4
OJVgty9szrGY2xvhc7An60QoL9rQrNt1YEz/fbwgFZJR2oSSNAljv5fRVY9/JCoKb7NQKBnn7VFK
VWVJ5Lqr8f2aufomhesTAbaVfg/G7PIW52LcCAtha73nUXq8gX0NN7pQgMxGg/HqZUtZRrToud40
cBzfpyt/IYzuCppvP/wNnRn07H79+jp6KOqczr6OLu5p+ikP3xoN9jF8hkCWNN9RH6bXytpARCqS
UxlqpkvavNq5zjNxvqbXZjxjv43CYyINWvcyBIQTJZKB83TZP5keEn1tvRuTpwnqWXMcKRQ6eGmO
pHwByxVSXThUISQqTnbHaD74C/5F7r1ldx7s5xLwR1JCueO7qQtEk8hT4x41BmFSdC6JFl3+ArFt
yI5l+7yKMO7d7Blry07TdtMLWnhIV8CnT5vtWdJK1OEihKUMP78MUdBzhW9gWeD1yOGXhopv86a9
tRn51VIu7RjdfI0t0k53WT9le9cBiqRNDBuWy/+P2g5TF/CYRG1oywtfGKWA529lK3mbgGBmAUdo
lYKwtVSGK/tz9Om4rwRtjae7X0spUqaKX/wAUht0oWhgOmLYHfALlwlctHVjbkPyVenESZiNjvW6
34h66pTMlcRGJsGDQu3m8yn5GgnvdjWo2qEAEATWvyzXgIqmR7hiMCs1qmdcSvF/M623LcezPcq1
cYZzxF+I3A8czuLirLrVBpNYR4lX0C/e2ECUc6WEoo2XaYsN1By0ph0ll6YEGWNaHm15CKWnUF2X
xN06vbi8FsxnZDO0bQXB+qKD40o867+nRYEQ2tuCIZM6fZi7rLL06IDphjFtMeSugdZuI+w/eREL
UbTbYngl2VUF1Lbxdn4CFFrhoUoO49u1d1Mwo7uo1UZCDfxlJCvZ7M3OwUd5HJeewPuPnXoIkDKB
ENjBNzG6SkcymKtPQURqbmNcidOMK83lWr9zCBi3qW6cAnTpRBTlmPs69tJuwneb6KGdUBkeSSMh
mBWoLpjSAfZDmVbEcaQxxjkkyEHJmb13wWSLoRmyM6vBkB4kE90vWGe1AKKDigI3310YO1E537ig
w0DiFYXCxN/0cQc7qXYFf6Phel/dbSf3flTIgK61DPjirVUgDPIIyJB3SCgI2mAA6HsMnCyMLJTf
PUDi9g4OAMd/3urvNoSaVLWnq2St4HWOTY8BGygavyvB7Y8BsyWpiOFnQjMQmkm9UwtnRTQ+cEQg
7j+iDyb9BndQzgexViyx37tiNBdMu/TLi0NMeQMomPTqc981zz7R/mlfsXEdMu0noLZoZtjvWz4i
q3RZaX9ONzNUVkIFDWsl7M2gwJqvieBR/8j5gjdYGeLXKiWjDBN/ACUuRxy/4tDKsxQEsSlVNziM
Awc6GKk8Cr+FMDmDDqZ/GN/YmHj6ckffpvoh6BMGfAqGwZKxS2/oGUeKqNMHaOeQARmHPcSGXS1p
wvAZWWppNPid6xOLDrvDAPvDip4OsmY64+epyNH52O55lxfmGQRf7MC9fj2gDIpQtzvZaSvHBYh9
DjC1F6SUPYpgMYSaAZYTkRgAg5XzatohXYCsKCQPOgJ68ikOagHlo/wTM5qMOemEC2v4DpEpeunn
HCGExC+STP4bGKkGf9zw5UujOj20w3hfpkBbETVMF1NQ9m1dEAlmX91CmTAbS8CH08rEM1teeZqE
24CRmIpVJPfe9r9rTVJaQKC29EEutYrsGSsIUEx9ms8VXP8+RAptUyCd5ZxIiCEfRvL9s47haq6F
FYCQerx/uwzJi5+yKNADK8HLY/2AT5UqZ9qo5dkgF+55bZyk1XbiWYXFgpgwdmLqv/e7wWBzHcE1
k5gRBGX/RmFx8cuDrcXyIfLDYmn0axWURLa49BsRuZHjJ3ozmvTSQYwRCURJCHKVgjU7pzNmTtWk
rPrm3Jq6BOrMA3L1/1Ji3X9/lHRiV8uTwS9xHvGXETlg24q95zs8oWbFQcKFNuVpZcw6sjsWxmWZ
yu1OQmgxMAzQ0VAK3bQUIuhOfGrTkgUKZgT2vUkMs+1NdCiuBTfsXfAZwh6DTCF3jPcah3tchJt/
g5hfIcYXyb/gIk9rOt4PerKMsoEajXewrGlAktWsFrSu3p45lVhhrCYSqJpv/HBtcpOj6KekOBId
Z7upubQGUG/3r3/q1S3ruWwrIk4APCofYA3siIwV8IlzqpCK602tF4VB9chIvtNLuNRuW/vSt5lJ
uM433QvoB8PRhkjdOCQq5QJxH5CIajXLc9+BgHpwMUmvVAXFKbFNKPP6Wv9erKyGiqSH74kUAvHl
/tfxgcyE4aTEB7bq9WjUJlptebUF55iqCB5wU8Yfwy73/FLWXTN1H4Z4wu2tZ2EzMohedFR4KgUA
uFiB/ZhFaK1hxu48Fr/AzHe5temy1f8EKhRelN+N6C886kYyTygnRzBaqNyc1/TVTwXvECsYgCjj
co3Qx3VFa+xR4XgLXIrth2BdqxQ4V0OxXY2UYXIBOELjFofStAV3X2MkF5mVwb3dCEUQhQ5OTvDu
clUllaEMUex14gJzZjYIAratNmYvEeKwSYirmcYPLZ9sqco+2dbm9M8iKJaMYPjfhmbax03GnUeT
yuV7jCQUaYJVyvGz6Hc87rphmFnwSO0xN3wiUALulIkSGxIQJm3OFwTHOQgFUqY8e1YXxL8AI804
sGhgUcLmfrFofmoSb0Hd0Dgq3u/lk6LUSMIDs0Gh3hVd0Y9xix+MgWFBQrsLqtBbkYGLRCFBLfw+
MFKloYd0Pm6YKIsv69bjjBN93zR5A5DEvYMxkKYlqNjEzcoBh9tHti3zYGuOEANPQBMbbJzN5cCv
IzpII1TqGNMxOHhblaivw8uTrJXV8sQlVej9sK/X/onCvAEJp74edTxZN6C3muumEMfAG0/JASUh
/dTq0QIUYao2EJ8w93NCpHacifUw1qnnXqQSI96EwwEw4oc01V9j2gfGyUYYuLvjQI+vatNW79cB
MxdF/TFDCPb5xSskrX1Zl3SYHYy4xlfZYpH70gRwRje9BAJWZJyAo9vtY+r1fDXE2uByIW8m1icz
XHILK+CU5omzplR3bcmUxOSyY4Q4pJ2rAZR0lt4bC/AD1lnFq5fnpMDs+kqtbZtXcIiusne1B1PU
n3PPypQaVNS2vN7N9/qVaIjH4K90ZVzUWSlsJ1/rHcv2fiJgrwEmpaWBRxAqOm1AbjkNRlBdFtuG
i4okcxU8BFBW9QNGVM+ijkXb/Lvy2QiTepdKuX/bheiOMwdF2A9tV7H7PWTOFRaxgfolELWzxr8Q
RNHFWjN4HUCKBvaLFfR5na+LDtcZHCxsYBW0u83yRROm2nWfFAKbNbUFUhE8ZDHr+/HJECLurRmK
55wZwcVy86aFDcyJoM24J5DtDddMkhSnnriWUQWUDTjhap6Yio+wNjnU8/uhusborrkELYRsHREZ
qGNL1TIGrhYWF1zZCWg8l7uOnypW5B+TQjVLtPnSmoXM1CKas42KtyZNKbPOSaU4+oLX+6UglRVX
KP1VNRDYFjFZNSopXsZ6VDLn3/4DFGS9SvM+DAAs7MNq8xrGfc0mClvAEJUi+/qQ25Ndb52b2wLM
4R0WUKpHJ5TLutxMmTOPOWxgj9BN9QbGbnSqDKTFLQYxdNVg2e1iOewe/ErFaFobdVQl8ktGDOnq
qwv2+KTjRBETgsnES7HWcliyLJd9XalZk+XpPvDWiczxRgEbXyxx1CVLrQp6kXl2QRXAdzV3NgW7
wJ1lP/eyymHDDtO44g0zYcFYtlKnWeRIh10wgXJ4C48STZydBijfbfAzTQ3yva5TOROSRYLKaCEC
mCqAEOsQ0pt8757s28lc3LYZVIek2givKNuO/TuWlqjykJcAvgRcZaWFdiuUbkr0lHkOPqMr/5dV
XAhjUdxH9l3IZ4LLgkiY0XH5rQ4mBXyjqIY97Ifbeo7Msbq47PahFl+xCSMGmYZUOXgZ8SLaaPgj
T0SAxxyhj+4zh8/NH1te++/3txD6UpulwTyPLu9k8GbxonyqXHwFZm0tWtF5wqbgOPuztpw/fCZV
HHVeOLROMiSfzjdmQA5A/8LfwnQo+c4s8mAbLvj8bnXayv9lgXaVFVs39AABZNWphAVVTi1Ssxtv
tzyXRKY2a6wFqk5Gq8bqithhw6bh8RcSbUEiFIxIwjVAEEoWVO+7IN4qXtENvnREUyKp5hK2IgJT
SbOe7kpErBHsmEzb0R2Jfpd2RfBDqg/YuTERHrLVClQhHMUhX/catIg9OrJVPXhN9S9TjrnUTcWL
OK/9sNsByd+kBCyK3y3J0YC+8f5vaPmUK3uPXrsHJZA816NLQUgSjmEqfU0lmtcB1p+sZ2xzRLu5
0MzqULTe1HVtH77FyHhGIeQIQPOca+0bYftc1k+0dj4fMC4mLdTV0rBoY3is4dgVvo+N1YihNjgI
UiRif7e5ASXsingMPGhPSJoaLvetZ2i0BPQ4d4pRA9ArL/XmTi9E0Zhll35YOAYKbc6JEpUDDvQJ
G/EEg8IYZfNmMTPborojspILJQEajTMSIipK02y58TBPv0vU4ww9gZvcccZ7nbhprTrjJ39JrZ/K
WOZNaA7qhpNsQtWgJOgQcS7xF7rhUcApBcm2bWStcOpkrrbTeU9y1QXp7JU//bGPV0OV2SQaPz4v
5NyIEMymFe4S9VM0yGLZXgmLz2/hIJu9gC1jjBsOP/EKuuXhjyEVXzqPKxG/2y6C64kC1ib3DUxq
zFWR4U4Av5Qpn/uHoroyMHHQLYbNBQZ530aHvQnevHriSwPThIb+f3p0X4J6X4zR+1Ii3U//ag7x
+L26RLg1CKYzm3V/Q1SMlar9ZCBOw6+9UDik3mL+jtLMLj6nxNWI5jBLrvALCVhkExdDYvuzvbyc
MuMejZl1xU0cRw6uvqY/dUS75AW/pU1uaQX+K35z1qf9iq/SXLqMmy+ObOyTS+9zW3ry5u17ekRq
bYpTWUZiVA2J0NPRJ9P27/qpSdUnZl4Ubn3fW2wg510x5QVJWjK+aNsl+uVg8id+4E1HtFzbumqV
xGFqlVSoJ4WiYqPcpulp+aMGJkzcxNPXKbMiqw5+TKrgO9O3/FC1ToLN95ztwHHrOQ7xaQJOotdk
Mg0eXdXPpymFBN5fSPrvAE+DmNbjnSDuttdOcxDcLTYUeX/ICqE8Ze+uRbrs7+ElHYdoAsgDgCXH
nmrhoz74bAc29AMsuN1ExUFzuddc88ePGgyNe9N4bXT8Ao2/0lKP2hWjwnS22kcPS+WEJheFpbMG
MnkMlwdozd47DSA7oEhWCcI/Ju/qBkfHOyYvzSiswl0ImWxwVs762UT7HSsjOvInsMGMfaKJ4x5d
v12jVkdFPjdQ94D8JkY58cQOh0JbSlH1uxJ61oI3aEVbld1lCMnfSPsVnqUSBRja9GXezX3q7v33
MO79D5e3neeyoq3XhgpkDohUCem5/b3H7IHUWruhAHSbein98Lv2RZG7BmcEnjVyXaZ8Zz+a7fl8
3PwIDzD+26XYToBhEIwvcJPyq+WUafx1O6WE4AA9HeCa5TVaBt6ytt4ojcBTnZDmx5VpC9CNCQa3
0PJi27HQpJ8NnDMEV5LTy9RUYVUCMT1dvxGqFkHd2cXtJ27hPeKtlGiPA2fFbJXCES7oKPNIUOw8
kp/0xWOEw++MHpsBxQX/KtEPzHFKUyee4G9HoFQJZlc/WGv/6ZPntGba7qEADwggmpogk7+193bM
nqg7rBdWOTEfC7TADPf65GJUfgVX/omVtiTZbFtWYv8AhgNjM/U0iLdE2786vrkU0vKHe9STjPun
xOwsTHtbnBbPOMSp/anho1eUVz1aKRL81gLLyd7sFMirbDcS2G1hhmuIgVazueWkQHjy+/r0c4Op
Qz2nP3aBXTMzZvklf3Oa7YUKvZeYzyInfucxWsUGNk/egnlJEIes3lze4fSGmCOPGcNFiJ8h/K8a
3dmmgzmjSvFB98zbrH+X5RsQ27HCVn1AvFxM39pOJu7bkeZcgvtKoj4iRs+qSGO+Fj+k5K++Kycn
Wk69T1SWqT9O55SfQT9TIjZINa6HNW/+6WW2FALfYI849I5ywdP9WsFuwSmS6q17XKUgOTIhybAn
Jjw3uOIkOrnjvbQoWMBAwIak64wUJk+SqiuZzOIjWSwU470uIG4wssnOuMUmM1WdqKNfxWVMgPjM
ytznqX5xvXrM7aoaWnFuwpAMfmxY3KsJqX5k2UoUyF7yrTpUEsOOd83/cZvb0ErKzBD5d3UeqCdn
evKLaiL3VME8V9RHONTELzwPm87oI64gFSggQPPjBwTlR+0sWaTK8DrUeJm21kAC4DMjw/hkeJmz
vQw6j1eyFiBBMTigWY8V9zAkQp/nUzpToJGE456v2yBdT8t+Afpm6h3/sQjELf6o3Rwn5Sd2ms7w
0g21Lt6QTRWkebQuP9Y8kO4DH3yjY70sJefIIATKPabCkL1KSTMQdxvEax/J/Ft5aYyNWg34DuUK
N9RMdfOI8e1iayTzpqasHQ3MYMouaRIsotWzL0oVb1bd7foxSAUu0QrdQ8lJJ9FJdoR+bNxvThvo
foVoLmB1w5s5lEBGD2MihmHUKIpjEBN8qsxeAo6ZMEwTZeV+7+oiT3qyiMeTaWz0sL247V9KaPzu
ld32gyCeGEhuY4ilL8o4ScTo39/kbc+SJJG63D1P+lUW//t6x8HurSKTIOzepk3pI86C8mPf8P0p
/LQlWtlVbm0Kp1tLfNlYAfywIjOdVvakwaUX6y/rSwxgB8qnMp6bQMIzDkRvYLZy+cCFdMVap5B3
vJ82kmFe+3f/3x4a3BH+Qf9SlyfhNtS1xMM0DStzRgO2MmZ5l0XVYl/7VEPy7slGUFFeqSV90755
PjMroodFTnE2zgBZDeut2ODguQXs+vcyi2xVtA3m0uwqGuSNfg1oHgW1p61peOXsc3AF3YRkDhf6
WDtguJ66ykQ60SAm5LLDAM7bsauDiSaGsLHPhBcmLv21bcvymrekCSfY71NI6/OWQWaFgQ1S4H3h
+3r7U6EyuGXC3OqYUmvTQjGSA/aNIk2uyksKmPlEWvpuf6ey8wbU7X4M37/mVvwwr1XyIeLNLX1o
jy6uzZaR1kxZ2vcMAp6q01wtFHrk9QS9dsA1X9IUT9Po5f+L0a6OFSgODgXO15dkNkqdHDfmbuIn
26r38jJuzxzN4LWHqG1UEzNNDOAKmLXPJQcTlp0k9ol6XhGcdpCIIT199HPJ1Ydt+VP8oZdvM3iZ
d5EpBqMLj4VGcu/wZQOM788/s7Ve5zxWQl3tCoiwsUfIupuvS7xHj7AZKQ2PZ0doZjl39sHQLAdw
auFzMoG+cbkgYAr97RlOl3oWL9E7TndnJWnWp6SsM4gQvzCtg+sGDyfl3JUPdAFRVUgunu6A/1pA
19iwxpgS4UB9F8UWCLt99P7p11La6kkCuStymhN/kZLJLwhGrePWghaGhCqzQmjUtDyt4qTU/Lcj
aakRx2Cwr4A3lVcqhXFwroquiWa1ifGlvkrRB2A2v+iDylxBMUE9OELUEBP1/Q0EsbW3Sl5nqgW5
HdNlUxNHSY/xYCfXrILv3NgMwphqPIHxLOqSylg8fzcHGP9j0Y0otnGyC0EPFhyjHztODa5iwupc
13aqfTttfxN7ogTLClmO32SkcdmdqFi5Xgf9kA8w6yZex+27Q4bmR1z/5ZCqvq4YcHwRqr3aSrJu
n1JZmNv4zr6vSEk+vaI69fJfFfCweRdmaV7FLvNke29e4GNYmoem2Uefu1Fr8otwRELYFNm0+gRZ
A758p5JlCQKnv9o8u1z/05WfiHw4G7IsTSqM7ojKuGRBt9/xS4eaeeSfOOQBGS2UK8eZD9L0sPHX
JegLqLnTlL0NifQdiHf1gS1hWYIGAwPiduIST5TYaSRwGAkgrq7sDj0T5jhvejHh4NdSikLm0O6U
X5MH4rQMQxBPVyQxLhreEFPq4zE3cvQ0zyYOLKzuPjJWPiSnt29YGRwM9yXtMu3A/Wgi/xgDRuNT
wTTtloLcZVa54l4YfrYaY77YgcnZKaTrjffBt6G1S+q1RyB+/n6S5ef/ZYQ+ylH3HRPwt8XG65Ih
Gv/vZvtJqzBZs4Sg/+Fh3yR33J+jyshZIsRvVjPPGa9+/1QTPX6+/5Ncxniod5B6yd+4hPw56L05
hrmCv6LiCcx8frOwdswcHvYOh/65OvDNhQl1aS1WO35yTDNg7ImnWLwQn9fJ7k7eSyvVgcnZme5f
QppFyEHsyKj6lfzSgPsGthItAt2WEAZxjOoubDehAHhcaL+j90u4aVcxVdWt/V2ErQSZTeprxNF0
AWe/lgI6PqQ9SxGqhmerNSx7T1uWUfKVj2tbWkPgr0gRAwugGacR7WkHpSYZARmjhRc1JFA5v6Mf
GHidl7tQzPjlkJHW79TaVD47bkAvVO9Sften7Bt01hpR0XyonDg1ZSgtTawOzwKUHqUFZDZsznsh
cBcrTwWbyqGzYPQuvf24o2KuE+dQ+scmvlLieUXMyxskasINifTCm7SuCpIaGbb6IoZR0zxe2Ald
6ehn5Z9axToVUAXidOFBCQuAM6PIoR/Hr/8i0dIfJyUGBJRsyOelHUKj9zScYRDo298aTQQBcqmX
dvYSvVG1R33CenZsRL5VNl5VgLny6EOscBVbs2bsMATioox7ab/+UsrrQzk6Bq302G/ug0guZB4Z
KYVlhX0DjHuswbgC30lyT3NS9U38nPlJzFqXX5PsewN2GCn/G8ud5roMzBISnuiJ3+p8gtoIMFtn
m2MJWZL94VbceQ5oXgIvMa6AyQArsq9WKCaA//3nqXyxSqWtFE/XHuZzsZaHAIS4zu9kvUl65Gri
1mHdGPyYS9tCHd1AbrIv3tTyg7S/gX6Wjl07bi4KP71YrR0czmyDolI0MUQgIb1zwgDIOFx/6VJr
6taMoY0J+LDFzLi3Al9ZlbGiNNSft3nUrVbOu6MOXtdD0/Ms+GN0Yh4peP6/E/nPnFgo2QPGLZTk
qD7Stso7dUNWEJQJy5E3VLDTAYhpLrG+8vPm6d0pFi9zJ6IieNifsQ1ZmRlEy9Inil2oHv+XoEOZ
MjZwjIQns4HDqxMynQx3Tlm/N9JKAIqMN0+K+oJqUtpRGYIgbAEcdLnYTl5d1RW2hSDVJ/9KXbHQ
oC5IdYKZtuwrAKO+Fg4D+uTaGcxx2bk6i+do4GAAR7pV6+sQU0NDvwZkQApp256iNf0QDLOfGw53
g7LqEqBUcPjvC7h2GFZ9canZr46mdJa205VRuDaWsLxSmlSPGHYSJFpqwV4zm7YbVhe5qiSDSpnr
uMliprNSmrJ8Zl/IxIp+FKABdNpMrUKnWOhXwOTFrujmPoPzgf+Xlo6Dsku8iRRRllOG1y/rGl8i
cua38rSWDCPQ5PGBTOFjpXmq/HN+yGFGKjoMzElptpC2LOyuXO5rYNeI8i4e2Ev28RbJZYPH55Uh
b/gOzDZgezGfcpuPgPVwevAIO+RacZ2wXmwI4AcRfedreA8ElzYFadvTIwGiafKH8pXkDyrAIMpC
MW4x7gLnxD2WoOsDPv1ifEHLKErMMl0IqU3sZVhPHyoVsB8nOnL035W312SoyGvLwCAcG3ZtRs+b
BlWnznQjKrTJNka61cWl2KITXZI1bXVGYnJ6Ehe0lkc6UqI9tULwr05mmsLo4snwnXaz4TJbltsE
wo+sSfNcMRTU8CIrcpoYP/p2i9AikzOoUCWUgXBgOr8lSprybI6Br7/XaDmaf6wFfuYNaNiruTHn
MO1Z7XrrsWGPMu22Ega4leMKdq+/15HbhPb170v0lXxdMO0bReq6ENabMkul+JAphpgsxizZCdX9
OYzHvgcyvCFMqMWWr8lxRIfBem9rNH/XRiIR5wBXePdXPyCxe7rTIyK7Esanb7kgbzy4tznsGpFW
DPaWU8XCD/I5qyKFREEO/xgjyFYcciWuSa01MvuuNtAQmLnuJwHqJ4KSp2Tmkb1ip2WpDjc3RqFW
mCxjaLGHrgf4BJ8jURsZT4cTlRgwbV9Og+URKnHlDUT6oYC+88PCSvx6DoL8qpEEXQ4uRCYFFC1R
Hoo1kjQXfv/sF7olEDr27VxVVp0Xm6vau6awLdiNBlCeCBOb6RgTS/EHnUGm6Z0QPrBtgdpq6BMv
iS1Ok2lFPO2cy21v504nXSruWMJWP9o6ee5cSeCr5UWgFAXcok5MDmomf5xGFNbySdAAMPW9Xi5d
bI4i5a+ZNuYei8OA5VVKT7RN8n+yvQELCKfaKsdMoe/VetBw+Vc4tal6MIn52s/+cIY+BrFjpvg4
UgZe+6/m6JgvX+w0/zfbaHfrFIVfk5wE2RJngk2y+bPq9Qcx9m1K3GNi1q8YyTGx1b8deNti18ra
WeThQJJslik88D5p7YTtprPvg+jZUnU50Q8nLcFj52GNhUzVNWjNZ4RAwaePiGgFmp+T7v2KW75y
e8mhw9rB3qAAyEcL1rTEIgrj4t0bym9JQHOeZEdWl/yCMD00Xe2Dr3kOO56/8YNWf604JKqEhwug
qIptUqKqjZC/jFImNouIpC1qV4N5yfSwgB3zs9QtTM1EfZrduA0WjED/n8r9/QQ8lOUADlk3d7lO
lQsi9FTkQ8QjyOVacm3Yf+AgayndXjB5ntPevsbfpJYDnJZc49/Bc0zXgezimy/b4xezEHjf0iWn
Vub5e9/u1lMjy+HB+Ex4Re9RPj2I+smkrv5L9dqlrOUJt1IXkocraEFMtXcdtRbEbkwKuywNHwEa
bIpQ07Zb0Rb6t2Bu8cGd5jVwX+j+/noRlHbGVc8QHTv8fODQZB3eqOL7TqYs5vAQSseInO7yML3M
XagRn1JHUUjfftUHSyE612MPtmWjF/g3m8L9QwPpKJw3wMLw3nPwjU8XkOw4bRv3/JCEBRszx7BK
BfdslgqegdtRsAeMRzwxsoxg8VGdvUn5vQ+cLITkc3uKePC1NxtwArhzd4Hc8bvO9vFiWj3/gMcX
lYeVnd107MqIdWkBoKW+3R4TPxjWJm1oXsxE7hhxV9utkW93MJbXwIzIJl1Db5sElaHG6uJRVhmV
2riXDvHxsI4drsvWelR4zTsmwlmp5rxwe4uDjuYXN8vb6BBX4shqzzdRtDVJg0gjjEl4ntGpFyvy
TYWFk4RnYgaS5WPXxzQK7vN1aYKpwrGt8Mk8QH9FhkSBWJRkVkKlEeP8ylpNEi8QF5MwYrc9kpLh
TLrdFTvmi850PBFizIjCzIe8JTiQSFev2g35zXIhaOCc6J3pDJpcqkVgHbqgwS9GLCCaR5r42kD0
F0eRcT/8hX5HDzWMfF0029sD07HpNXCiW6xf6q4ymOSpvzmaHeKgdWLILhwWw9qot/v/DLw5B5Fg
pEcvlxFCVQU0BAWF77ngo7E6eqQJ/heIWwxFCtNv1XotMp0oEwRc8nWALsJT/NBtGuecBalDZqvd
U5jvxJZoJ0PSXFNUR1smkRiP+LDCuvpMspJRrOIIMy+vWdggxjSKTpRxNy0pzklIginNr4XKfVeQ
04pOl6W93AO7688nO77Ohce3B9v4XH+VgBs6cW2ef0hB9M0qFnkBrfZO3hkn1qf+iX8xN3IwFbDx
MP1OhK0as+cANbXV/W6gVgH5KpFZFtk0FH9Aknvtxe/HHFVi6a5jnr4kxCJRAsxecW5QyWRR1BjY
LzFWYXa+h7ZznyxaMjsiYtpiJy0T/xwOqgjDmnAOsM+vV22YetC+gEfu2ywQ5ra/zYWCB2vF39Q2
sLKW7IPbgf1vXe+dMB0aLgFUcqFVef6B/KOmC9VxyElX8i9+Wgz06cN1CI8Omvy2tXokKl7A6Aub
9OJ/6ZIPUwj4mNWYwNTzZEvhjc2a1Yz988iZf5Ev9orRLd9IIc4hZOFikRowu32Z5U/i9b7KtlVj
wyQ1UxZKVwSAPdu1DipdSzhmBNjXgu3s4MQ43jqXRuOSD31d069K4hcvFDAyQbP89asFG1WeM+cf
ZDOGDkDfGwPgaQ1zJzpy+g+U8ESATs4df+aEY5OEpVkVu4OKnbeJ2BL3q/W+Pohs5TRZc91v7sTu
fb6L+yXXvOOkxOeqSdPwAROZOVGc2c6A/sfDSfwxzky+vAJFtv7BtTLTULLOUz4sn8DKCl/i7wZZ
JaUuJAbN3pLzQctPeeNibGeQNslSJbvwRx/uSOAqtrC3HUyDQHOywjyDbCoUlxJ69aEqvrX3DVuO
w5dk8XtAEOkVAwZWv3njTWeFNS3+8ZTHacBD8I3p6CkFLT7E4/yhZGwdS3mtonXUqS0ItPh3BgdJ
sNE7KTfKLVCAM0Tagda35FMyTy3eGdlSWl8Q7uH1/RG2RwVgicVA1lh5A2sdE5LH8w2QnAmt5NIz
BvnJT8aW1ek7gXQlJxZJg6SYaTJBvMacVXsyLwKJP4frqhAdslxOt70I6qsjY0ngKWQrHbf3/Csm
Js1W72EzCOrsA/jejAqIYnxXIwYXQZnMv9e1OF0HnOdzvKuwM6H8a2SimJsz5+sYmC10vRGAKxI+
/PSGrue+aB0NJqUrC9c4ZzMIjUoFeZhCi3kH0aU5sshgPsDW66UtCJIy/J7DnjL0CdFMaaBsKrqL
5qXmBXp3Do1qcsD3BFwsV/fWH21yVUsdIxAFfRWuov7DF69I0tC9prx3RmsC6mnSX4PDKC09uwjx
zbQjE0gKbLClLVhOIAyhUOMveWFNPdoAglhYvsqNz5b7kVMYDzIHX/0D1yIEjwYiGdo9EZZWbBiv
P9IgfcuvBRxOdq51f6Ig16L99BPzjobIdc38KLJ9PA8dFHoY1WSfqWy3usCdXpGJ2OIgA1YeboFs
I/BuuesTuk9vs3VKzIO0kyrUQLKqpQ9cAj34zyeMrC0stnIjgfgSkizwbRLnPhj2rGJCcF9DQZd3
Dnbw7SGFDbotctj8nSVFnDOnMRHmy+R3m/txvGzJB//zokCIq4giUxIFWoiCDXE11Eg1q62T3KQz
N7W1Cyd136c864oiKtrACpQB+n6M6YGFlCSshhy3GmubemR5I5sGyf5dSmFyGmEQinLmsZFGg1zE
FNfDoyO+sK3tERV1XBeza6z/cqc+5VRqZ8BjfcMK+n9TXyi3ZMvESkmpyFo3+n6R6IM+iZKeAbNn
ZhRhlZin994YVJQHp5G+sC9sCZUxhOmj6K6BM21JzUzArDxmdDHuiUBAkVN0fdU2Ir/Y1ODyAGAq
rciJ3pb0DK1MW/xmuKRqpwCmjE486MSG05MWRmpDvDpa+yF9HZHQKOjk6xmAO3fhnBBDlgjlan+X
n+G/xTbYCiBILyLYtngPkMrR2dH3CHgBWySgk/Ue1hR5OHDU5ALVxtKacy6TEklldj3KAdQrCQk0
JwFwlMeze3OdmlmVt087rs//JtVDL5RxP0jQdndJzUenHACa8znx9EVsiNb76TbMc3GS/am+tayy
UiXpbTO56r1mz6tRJLjUSTuQHctlkksIJ8832ajvykiZ1Nxi+x7JFB/mDVJqlv3QpaYndAcpBGJ1
QrEXorjKlYnNYy2Eg95y+XhGcWn/r7aNEr7E5URStPvYoXeeHnLZszJ4wTb4+TGtMYg3nvXaDPPs
yBML5gKgIZZNuzjCErjEqDPGBTOW/kwoYroDd0ep+iUxbKdlbK/nDNGtEoYX4IvkSR7DVes2dKq1
7/zhTGW0DA7f1mZEQx7C4DgQOwqliDtJsbc6AQV+AxYqAfO5YTsZ1+UaR/V45KwUZ1iju7YG82bU
i4ex8rqFUrEVWoofVZm66LRkousde9wtTyqJEvKz69RYKdFyxn0aJ49H9aekfUQ6dtscZ5ZAJgJw
F2EhfSnJUmHba4MND1A1S1mxzG1S+1XX9GGlfri4fmGp4PubwTWNe5bAqfz2hr8meKmVROBbn5Q8
KkIibBkIOhgQWsabHl9v9lm763pz+v1tnfvoC2pdkLD8AhqYx7Dd45ZrtpHRzQQLxVUQ6ytbzjSB
0OiiO0tCN7aXpZJngek0SGWqMsbqRz2c8ya2LGooPw+Rk8RqSSsHuEsA5gMZdFGtEYbYrx/8QwVW
v51A9LPu9u3+JqfEFybZcKiKGf4FDo2R9MA+MCr1Kpnlo1nhCjh9A/LWDxeoLHHzA96fV+h7uFBe
FGboBbSa8O0IriXmi8seAOW+UqlRusMmJLwCfyhWyXP63XbuFqXJTgpX5da1VjWO1960eFF9rypQ
srIF/u/d/zNGXQWS9LrAcNlVROT8wwxLKXUTtR3oi5kXGasT576H8Kwi8+8wnkRm2CFjFdvd9p6R
cXMUHZlC7UXUtk9RBnkFVJeluP9OzRmOl4MtpTvomQjuhc8FE9EtEcAVtF0HtDicQDrwuR21W5nu
lDFLNKv5eH3MEllaVYGBM6udQ6zytMwGhhp5YRn24NHBBOAUaeKpCLvXOsyymQxUu0w8N7JXL8/6
fbJ4+fGy9Hse6tOA7PfuBizapn2MUcgmDaMKwnAuWP4mPpRpuaDxiJ19xhDghM5Xm26p0bXZFgg9
fKxK3mLg83RUE5PKYGgBPjELVsWSBAdMmNSOfycGROAnZO4cqGoo8Dhtiev5M1x+8vdd4xkpeLjF
4fp01gsTwlsJgLQLFdinH1R9FYSzsjVBJywNzqfY3ocodMexKvJFEUIRv5rW1RENvC/Bwt73l6Zd
vTdedyscP8xoTV6GLWb15h6Vpu9wWSir1bsMQpJyLTRCSUgplmZeKANcR598WCPcxGBQnHmS2zwQ
cg6A9DWUYnEF8m1NkPERbMUBNPAh88b+F1eA1ZSrWsEKVvVb6CPCbeGadCw4PI3fUbNmRolAjQl8
3Bmj9IuVBQKmty0Ylm/BeZK3v6O5A3MmTZPo7NbnsyPXxHUgRO7F2lxyWfkz8/WTQFHgDxq4nUKu
XG2BjxyX+JY+MOP0I3PqVM5G6hxapIo2xWJ9+ql1VOHMQJLEpBdx934McdtUy/eTB/6DqZOgzN3h
9KXTVWKEpALDbykGki85FKfsGFng4AO8nlu1sEvMqBxnl/z/5zh5w5TZnN+/sdcIcYPFaG3MRH2x
3cYYqZNczDovPUB6aZNDnmA3yNG8jzkCDLqNqAVtd8fpFEa2WnuVpcCiGW3LULtOw4ogDryda5la
YIwokkwLE/hGxe3uaJRPuDh6aT6pJbLiGiNkOf3Y9YnUY3zKfF9777y/9VSoNu5rurYf5oxVtEiF
hx2CqaJJCoyyTdgX/j04t5Ij22XGUwSAP6VATUAEJ7ZuQKi7xpMh3oOigKm72QDTX5GvxIRRc6Ju
P5LM4xmEmPTiPeC9w6wY12BhZwUAglWG5P/DxiL9ZyLVA/F2s/k7AuG0VDG1Zq+zQsUbGUSI3FmM
Q7YF+rpelSQ0ors8PM4dsa0YCuC8jun5YGEGo0eAS/dZzC1CCvMLAtOmSKnh0I230cA/zj7v7W8p
PE/HioXKb43sFq+3wXUDjtKdiNysHv5V7sI6b5uB0pIc0tr7B7ZPcLabsbRQTGzKdpSnfYaU9acW
fzsbt37tycvQ/WvHjFHryoL8C8XcexPvE0Fv4JLEt6Nlw71bO6/f2Udwhl2KVhZ69e7+2uOuGVZg
7aX6+5+PNMO6G4ctO/SwndxSvzJfm5b9b++ofhYrokN+BXvPeSyV6AFylbivmaqzZ0L7SlTovnkP
Qi0NTBtzV7OWSI4m23Lid9egHtqEp8Y7B7vGKG+xeIgVDOecPdqxH2AmgKNqhKi2buTOsdWNqqwR
RClBAM134mzc/YO9s278csqp/hkFp7Jr37xt8SFn86NB9LH/pehoTqkIBgEW+DCd9gkOSiQrA+Nf
i4DorQzpXGBMPJ7rJ8fjRC+47Ym4//kiH1a/i6TxEAO85I2VNCSbMr107x1W7GBvABt3hfpR4o4a
/FkMtpggLRPz4jydmUoP6Kuvs/BdTUwgGbS4erPhJR1WKjKJzZa7PrBf2rcnQCunrrZostk3N0bj
kOAXmmE4p37ZE2r2wpZsrl+kG0D/4/9aSbSwq2WbnKVbpnC5sS5pO0skeEhBzJ5hGMke6YkvWtRb
6OO0AioPZsv8t1gFWnyccFJpgyw+meUFoLz6IcY64h3wUVxX4LwQ10DSRbsoZN0OeZw+7o1Gi75I
gfK0hFzgEfHxt+tNUSO+9Eh9vuRbtFmnhJs5dlcY9FY5FNY0SlrKq08VI77JfzqCbEK6kin2ui2W
i8IuUBqPAY1ZwDYt/o39NIIP1sYjYk5LCpH5APPQzTobzoXBcvyRWDhanYXlJ6i5vRMXJUOqMDh/
DPgNpVJEtxYAvV+plfK7BWNMhY1M1zFsSoEBVkSpaVj6EpmWimaZqaIe7TxCDvB0Fdtsx635ZS/p
rWflsVtuAgtouJYB43MhzzGEZW9ce/ZW0xD57zqtNKvhB2aIo1pDgQZGKwmqwn8YHDtOD7WeZXXW
qC9YjVCPqumCFQxFN8NPVYzX5MvLnFuaY3rAD+vXz1VsjkwbWARJ6sQCZzIlQEYRtRbGAuCAMHFq
Fs078pNzn7JwfgGGqGUECNp8HzxE5zDkLg6UK7hOCOYhMlZm6EPurLmNr8tOOMGiQgvQHU0oe6Hn
end5w0IDB//GrGmz4yMECeoSRmwUUtCRXTe2fbnC5cqI4ZQBl7VXs/CiuKpaKf0Pc7Bf+BpJ8WVw
6CC2PTYylGSfVbjMzd45GO7TkTNJXZzXCh1LQEjcFZ/zAPDmxa4EsoK8lmh6URelseis13+5QWRy
mgCcaebcXtbND/5K1kdI7IZwWmA/27pb2xNugPLZVSl1EE+G+aaTuhEyxv9+P6e4HWZcm1VhufBp
ogLghFd5lFrBL0xNplwLVrus4uQiJe8AJBwNLpJLly3HN3yctZ8cPa5djwykNzR/B8B/2686eVbK
dwd2WoTRprHz083oFV/AqZstLN+QoOSA8WRRNSEMfcXTjqHNbbsquUhMkveP1KDafSWAOeUPx2HA
XHz/lntVjoHXw8ddXJMXXsKLaclH1rZkydqElwwrlKIwKAZSupJIBod2ngX6jGU583v6a8JPOCy6
8YXfaGosRbjCl+pfMfVjQJ3GJC6+L1dXVTkUFch7017GRC3V9UAmO1wyslowUaN82T4etJNjhFsb
NwLN+1jmuJjZxx5zDaeRVhBSkkyxtHcQyy8JMKysig/Q75HkGs1AnI8ktRE1K/lNzTYpaH7HlNkD
l94PlVWZCrUHOXO+rsu7vZgbmBsjmFeDaWBsrpLP6aPKQ3NK1z2fALBLbYx3vkQBjuFdyO7CbP0n
6zDi8zCBpJSyM3mD3Xg2kSSKHVuM4hqiSzRawl/vxR8kzOyvafizYjCM8r3iWCgFk7e17bjn38kw
wSiZP1nyH6mz3NEOi5dt9RYzz1cngciNfb51gfD2YAnr62cbH2nZ5yOsYQl4wAx34sxw2wSVjxW2
I9SueaM8yMtZtnJJwGs0nks68p8jF7navfnBfp4iHeq3GQk/HH7TyX9PfIYjvcsEnQPnNdInd4uN
zzV/XUY4QFNI5hyau/4xmHktOBZo4fd1B4f/7GgytQizdB0buE/NtACJU6bM31Yb7Wqip3E6WHOp
GUI3MaDq9WDryLX1f1nzd5uubnEx1Auu5iPk9lLXOhGs9xyqyBfgQND9uy/SYJ/jzcR7nEFPyeYU
BP/hiWiiJ/9nQBQOwR/lbaSKc8QhFCA5t/aowEqfZQW3DOSIPNJn7RxggXE9EXmeU+9F2HDD/1Sw
bEtKT7McQLfnV7HtarhPFzYCbffNjFevfkQg12MZkb2d/7MxuAi2ZMSvzjr53WFDRfwxMknqCaKm
0HCYzlsWg4xY0hcVNBfu3N47rlzJnv6zbioBTAkJ9XuJ3MajaOaKN41hpSPSvesbq7lO4JdsOMhb
xmSCAi4RIbHGoeqIhArbtGRjq5oZ0OTj0qqV3QdBIflnQyjWPFrAsX/fLR13RKGnHc2ocPsK92S7
FUoiK7wkx+8k+Y/epb2pqat3hHIu5jYBIXJNpg2NczxFFzSDLvf1FjVWg+MADYTK3Dv/2AAqvkjk
bn/uwNSAVsNTUBSJ3PZOTZgytfdg3CMzXFT6wXBfF31U5+TpD7kRGZWMFDMCcPc8usGenyAEUW1u
CWvpPOzQGU9KHXRDY8gX8+PCvoLVyq+LpPhfSiVsRQptvPG07v+mSbUTBgNUHihOzHjVatxF3USx
BC2ezOzqfGX/FLXN+qeHwu/q9oZSaoxoLg/7LUdIJ53xXpgA/SM83aQ8csG3+lVaaELHJRty5gGj
kBQenQKJfmOPT22YMj+PWshh8/Q6KpaQbOytFQnjK+/iAXzvW+NHD44u6Rzw4H4rhtoNuW++u5kH
amNoesZb+L6GNaLNGIl+cD7bC4kLO4xzgjIOBDlwIHNjq3NLzV1mz5QfBpiJI+jC8Ac02PO89fTK
RrwoJ/XhxNI8NM7YiN9PPTW7AjekKoTMm5B99EUdNEe1mBey+c25h0GnxPRdlXrlU/lJPQMra+pY
EWT1E2J7vBg46vRHL6aJ+94c7C6U1/sONx0ya26Nu12TJmkhW98m7twplHnlfJIgytgr5mrK1L+m
Ki9ffCNRyvR2MvBd6wnTtW7R/eJXgqjsXaESn+oSZn9sbsEBtuDPMNVgZzXYZWymD2/Sp/BQ2n51
VpDn0fW0/p4flOra+x3wX9QuXEsoJWQfh6hmcwK1pEkeqX1qAiwyDO8lbrvEJwLoazYyY+7TnMs0
gvtO+37vwjH1MBLUFHLNu/GzHS7Dom44rVhUm7NNmpi3g3AS5UVdmIc67X4bVn11xP1WxGXKhRR2
/D10LSUR6DnV6efOKofOXmwq0j9vDweoaM7C/xJCfDT8ZMlrAp1FGTSEezmfGPQuhMGcfSZp59ij
gQN/dN+gDLAv+M3DVtcOY9bEbIsfIhwBJV6++hlqPzI4F9xJPWHVqmXzLvlqrrXQ2ggP6aMz44f7
HfzHFFmWTErilXUVRYiCcIUh99k2YfemsTNXJ/YtUOFfJffiXBjDcM/1SJm2GrsZVV0px371hh7W
gwpqealq7Secqwce6rB5I+hQXY/Y8sVxG9OvhOk50/rjUR145VLNgVckBh702DW3rtbVDcVMrZNc
t/WkLU80Is+df0FpXvlP+ZlDOqkF46+ZcZ0WbObje2no0eLhsdwR6CTGRyBjR/uR28zE5JOVTQFA
Ghwa7/O8dy6ac4Q71vyjU0FgMLCqkYMJJeu9aEsjsgIoDqMi/7lM2aV1qO4Wm5NIEJjzq6iaLqRk
jHlHmva0y8GjkWrwnwDEeGps/eREjI8Qklu364A/g6cne3zGeQr176x/hXXu5keqx4YJ/N8O5YgC
o4zhZWfH2A0XHlmzgLL0LKGIKLV72sv/ptxnGIKs2GRLMPBF6imN8EPpv0NhaS7wXUoiYmL8iYXw
ii0zTikLrhVKZTLx+hAA7IfbrHEo+YuRQNKjLEp685CIMMYuIHHtX2boiW56Bx1HAaTWS2+75Oem
lO3tJYO1tDR8aVCXLS3lcWK2Zkn4EOa38BQpkiAGdGfcWZnFb1Ck7kz8QC3m6gRIQIw8aTDnmhay
7R5wgYFr+2wNhtFj/d7kUZ9d264TJ4SW8CJDRjv4PsviYFjZa63N8k0QBnIRvTjdy4IKtlshob5n
KL4T0nbwq2qmjHauQ0QOY90W2y6RUdWYDsLqLFAEfZPcVzz23RQcOaLkQP5awb1asiUOWdDYOLm+
Ssw5ICaUoJlLi0KLkX4y+/h8z4dFu7PDtOVQunZjyQLPnR2wPlhOVLV++G8TfxPFeAnRlgXZnHBG
haeXUuDy6yPzxiQq+Ufdds+RmaZvh6z7HvNS8S33qQQ6ageXS98UwRyswl8RbYZ+HZ6LkcCL0Omv
QbggxLU8VkyDYzOPadGoTqelj9EvIz89DufzlMcMjp7nM8hJRb0CcsUpu+p3ZNP6ex7mS8FRdPmB
46gjDvZD6EBVmJcp9yl56GwrwwAsgoDwwgjdByoguIj3g8ovUbIkKnGzWMUNBssFJg/3oTbOvpxS
mqS2QiKd3qsIKN6iJJxNTQcQp1QXrdSExQtrohplVBfPT3dKot8Pl276ypFT9lauAYm+O1Cdqvp0
+QdQCmmyVFZ2ni4/gG5NEqNKwdf7+TJi0ujDgSqusxFLlDXDoOEAdLOlzNIIU2Hmw44i62sNxpET
eE17zVPGoy/pBgEZOK7/hNciWZ5oC1DQAph+yvdzED8r/qiBhsIbjXSZR/VFGyAE84nqeA+WfMzO
W90ApPxNuWLZTGRdLNa/yfJi1VNh4r2w3oilw7kj2Q5Oa28L4Cdz4w/UxAdKqHI+HiYBLLi9inXO
PBemM+XcxM61jpqIlZdn4WXchMjAKhik4oFEU1IAD6Ds4aB/WZTZEtA6nKmr61RJO87ou2HR010f
0+T753IKrfSzU4zz4mN1PGfl6pTAgxJhqvnARONLCTwwyagDQ/DQ3n3iGDqlZtp7eJirYKupK8II
Mg6hVBMvA2OwK15wXd9llFfszX1zupBxxfPjUJXKFaPiip7rvineK1bgMZIt0OduXv19tmplnp3S
7fZe6axK/YP4SIimlic8+W4oGyW66h7E9HwAxApP+mSgbo5d6/Hhje/omi6h78pm7bbgpN11/Qao
y/klEtWXEJUyKCB3E/OqcrNqGBKEU57pQdrTMJaTKx/eU0ayrnXDuhIpkcW4VfQzd4kDoYXs6ymh
1hn3A5nSUG2YklVX3p59UNiPT+Ligs16RDeZV1doQKeWkV+7rU29ycAaTEBAUl4Dl0U+MVQ5+e7n
NvUiC4LKt5rry1DhLywAhRWRWxyy6h3AfK0ov0KMiq+PzIn1caWD1LwGJxTN/5T7aBDEftqfcQy2
KVhfXJDSGnTUwCl8XpYHpZOajruMSfoSOJjs0BDye/tZxzRmHz9h+c9/2U2YLcXZrTFNBzD03xRw
HSnBrVtPzcK/aQJuZ7T8gcKHmo565sua7OvEmG6Am/a2RkhFBLuD0cEj2y05OBsKAVBxfa280eqO
v8WNuGgRECUYprB7DfZwQzysSrpaVkzzPSqG4NjuFRBaQpwWkq7YhzkKp467Y1J11ExX/kefzk9C
qcdv2v8yfMbVsnqgVT6DAuh/xch5MgQHVx86hGC465QS91+o22w5hLdC5By8gZizclaW3S1xKxRb
eH8nwPpsaXo6l2Zl5owCQk81FKEm01KnJyIMHbfCxjHubX/8MOyEhqA7RB3+7ONCgET6P4UJsJqN
QjSuFgOSqwPuJr85DBK21mE7IBFs8BiPqw7xGrpf2m7GCVvBvjr1WMLyaCCHfiR5qtz0xSPvwmJK
FEXN5pDkXhIT504nN8c2bJpJ4wcUIBrFh0VNgeSp3MPYsSA1T6fPDscdDWIOJyGglJ7cE3GMis76
Pva7lvRQV38+cyUhDv4yGASTvywEF/1gm43o5aXSpyLtSa/j0CdJOzdUckfaPTv2zGQKrP6nQw4P
CHb4uPy4SygML8CsYVEl3RaGiKNGxXixv5FIdf1w6tv6KYjNe3vZpqCXROQ63SqNCJw0FeCsx/vY
n9fBH87BJJN/OdAxGIUOEMiu+s7PnGSCR14/kqN4uqXffoo6OBA1J6kDWs++gu6jnNca8geYmOiK
HbEZq2Su3rfPa5s3EQpAFypVMnAmOlIAHFaqOTCo/zCjm7jHSX/A9YZ7JMha4sPGN/xVmv4WzyIc
arX1ntDE1nYDbRqjeiwx4kXLHnPbzdKSINrRD5ilKk0FQnxiKBttCFvgq7DtCBCYm6QWQI4WW2oq
OfTyKsTtgYrAGJd/wqcRQshNIRp1UVClcfOkiY91gEIM1eBKBLuxPSm5mCYXfKdAxPz6icTzW7Hs
fqqhRBGksoJqHfUAuv73qIvtx+tqKByz6ZeKDJjlVQbnI18BLt5QQFz4Jw9bPRg6GlMO+m4hW15m
uRFxdLeWyBvhGccC5lIu9/3PKxLvahI8bYrihwVxw64sQgSfQBd1E5SMlsZjkNa3RwuzUh34G8NV
ZM35qjwz9siBNg9P2R7mLKj58VRIbBkOwIDDK7jClX9EqMT+OV86z3Nk5xB2dU5rmM/wgF+MmDnn
uKWKPERSlEY0c0jasJDD7Qzn4hT7KsyhXs3P5AlQXIc2FtIT586rILiQV7wpllJUtOeHC7Rz0aGN
VsjWpB5bgUZcC6S8TI0HwglhjBhb4p9aq1wngn12MhnTv/5iJnDNJluEdAWk7gv/gLDqe1oOSDHL
he/GrXlFdCa1NamkdhNYkHrk+j89HgfGO1W0SFNjleksQEBZStYMpFDTzpJSGLg9xNaIPWZt9Pm5
TvoaU2BsGmxK6KEN0ci3wBVc8Z8xdLz04lTqzaHLBIkMUB3Yl7UMQUIfeiHVjTqhbFFZJ4YoMF55
jk2lT30WIQ0jMIPerLbJHkME9SmuepfSboqN/sxajUjw4P4633PCsnIGMgJg6QqwpoedZ+GPakv6
jASqZ7NCKjzCvpXmul+jAoWsgtg90/61KJMy8c+ZP0R3hRcYKbJ8Xp5SM78eDMRB81WFGFnFsuNQ
mtr+cU3YUSrp5lyZvINP3ufYVtSmaNo74fS1RNT0GyM8rjmojt1MKUNKnH7yPynxrrX/gQK6O8Dl
UurWZErXuNVupGtZSlm3ihdkaWR2atFHvHEKSvfLoWPtX72bcCybefD0ESeZ5N7SHCuHDSaETjJ6
VY47xjnuOYb5YPVVq21suzsV7JrV1UuBtcXdHuHAmYDO91PAGYKcDWNNI3RsCE5F7VSOZCjRbjRH
38DrD5Prn0dpID8mM73T8mRDvpkEv3fxi39Q46stUSNQYikxFcg5EeCWS/rL7ckgrD3UxjEFYcxn
8YLN13+prH1Hj8bXUw0wmCyYvpwfr2JGQaJtHP0EC8vNMuazICWKuCU+q6DrVsrUh6oOe3RRBgqw
uZUgcxTfErFSdDzoT0yEQxGkNupGpKAda7nXozpBlc5Nm4ZI7wqpepaninP6b1V0scwwBbEZ5aQZ
dHV6XYSnK+VOvnYw+ALaJPfIiQn3W2/bDYWpoTVWq8bVc2ctmE7yjPmVVcWhYYdmTC6YY4DIiBIF
sT2BVlTEApVEA3BxHfhaTNzxccFPWEFEDxUrhbDomXrB68vzyDiWNIOos5dH1JWSyOi9cgYOBRIQ
/K/LITVZjVErBp88adyYYt+wqsYXC9HA7voXUrsMmM3fLIEOLCcnF7RV5TWi79jcORy5OfV4nkEM
IR5QcLiNGbY/YTUXV5JZ7IhHknsPB2eg0w3xXTgXXT5dnol0ZTQLoFXKrl0DjNd27f7qeq4afZuU
R+5HLBdesUf4TlDc9ayaK3eapZiqkXCqe6Etd8zJM2zeTLBQCK8ED5Nj2Xjc6nVUgTqmgnDYVWoQ
Uhh3M8217vWdjis2a7Oh+A1x+YwUcQHDM3tpcfaGEZTW9weigsld7DdKgVD8ZCTE/+5lqH9LDsUj
BMwGka1Zt/sJtOdQiUr7F76ycY5eMQDG5l8PARZQkWWc09HTYAxU8wW458SivQImPRo2VbldDywM
ufRcnLlsuX/kY+JmgRrEU/kRjMzHaT7R26kU28JcG0fA+J8s4sjnt0FEdfmP2rNoOILMFfcNXZ7q
l+RxGrtdL/3hZs9Nv3HwxFaegQfVk8xT9CNx8KsCQQ016Y0Jv9NpK1PzN9J3T3kStXweHu/rv+tt
jarHBQdY1Y3uSul+YY6VqxirHW93jCL2yDGafsgY51+KXJCkUYj2GHBxd3CaTYXTPZcW91lerQRw
GcVtg0ZbpmlQ+6xUzjFikJYKVh0eeLSHP/T3RWiLeMK9ZSsbfal7AY1/UFi31ni6Hytf2Hr5ucdP
iwMRlGZML9AE4VmrrbIkkkyF/fbyoqvpgJl8XJ6lOuq9ZQBqJvtK33/QBM6t+2JzAhXBp7hXPoK5
sieR/G4HkEzp3MmiBOYQyWd+mOO+Di4/Vtx1lEZzqdfD60utPNZ5ngmB+cdLt0CkELn16zcta3ds
791UuIlknQkI8Ia+7lgHE73xbP30ft+jcFTBwehNeYb5+JeEoet6+yrqxGQIcMxmrqXW3sMEVVxk
xZu/oDlQzf9+wgQnJcf8RB9SzLxiPrmGEe/EdTNiYlW9Yn/v3I/fH7ABHltSrW5OBl+aI1jOFasu
XXQdYfD1bck1sAnPsmN/UzbSDjtGjS0vdtQe5xSzq3FO5KuThtIrz7cfE6TzswwnDsK1+R+/yId7
0Wts+jRrKsvq6LTD6KxkWMTOOdz4U4gYQ7LZo8HF5UvZADkG5l2UJFsG9qeTHm1pfD67+gU+VIJ9
y1OKbNCbcnfSfJQZ6aW0e7RnwqCH1K8S5RVhq07rlNFpOcEsC7IFtjnchZvZqfOw99w9zxsJIcOY
IVSRd+0Y+nfz8cnuprsDjwslkvzKMbrLV4/srx5taAP31RdpUno/kJuIwEqqeuhTpAQcp7G0q6TZ
olalWpR156lfZ//GMpTLeMkut8bCD+CnDn5nCHenhXTjARlF5RXROoYrpY3lNSTGxo7OemTk99OR
lbBGL+AZDTreHRuImpYoZvDoUVJ4HGWlnxUWtzIo2k27+mwaokPX+crBCiDILEo9eAd52AvfNpkh
tSRChINfcpGW3mP2oYKUX1FTpcwWEdkYbbaV8TMEFahb9k02LAFAjM3J4FG4VsyzdWrOF7ZnSz7e
DnXZx2vBM0Xhe9/6HVa8mp5dcQ/qik9dgtJD67i+bKOUk+q/mzA8Bk1NfAD1I67/Y/GgcfSoS3no
/m8glCaM9WsolIoC5ib+clAXq3ookPDzZDprkRsrK0JhnjuIKvB4zJhlze0AdTF3On+Uq8OCEWCg
yeEtqMxEd0ffMntMhxzBckGVR+nnENnQPHkzNTNG3SZCWtgqg6Q7V/gLCkefgO3VLu575tgLvyGw
6Q/4HYdxqGONtWUcaUxI1EDACQzlLXnQoxnheAOPL0uxQ0HSdGloYceaRvGjtNQ3ZMid8BWgG6BV
jwbWcakULmoSMDiEL9LpPg6qhygFgPTAK18HpAud1kwgck4ROBNXWA66kE5GiKU5ZZejXG/LBoVD
eItZJKb6CPYmCnHntFV8FXYH8vpKLjdaum3iwp+Ix6hTrpENcKvnhzS8xxEWtjygo36Iy1NN9Uiw
XWJsugZy/JdVwQJwz8rrVuBe9k7jQtrYXwJzVx9v0a3PjmtoVARStLVHn6SGyPZ0teA5+mdKuRaO
Oz4KboOKwuWocr5A/IlCMdQAW4/PGEhXoGErpD/jNZrmo9p7fbZLTJ3IAw4JE0b0yuAkoDBLTDbr
AlEkWmau2bilfHbKZi1bKBujLGOa2KPeD8n0vEzyLfTfISYGZYIsnarzzy8WXFpxFY0y0nwKjZgm
oX2E6MJ/dmFlhBmK9sUF1D4NgodtO7Juwj1q1IIZ5TrRUlZYjm44XKW+vCKwHS5cv9gZ3WdunxI0
k49wkU9vRbNBSjrM27Z3Ecu73NLmLU4xR0FMODbOoPsLPH+vj+q0OpaO43I+oSwCmfsbVWDODf5W
GxL4d8UdCRhc7k4DveBAlEUKasRQc64hAfvZAB5IqqwixF6C0bq4sSje6O06lwnODDuwwlOfWY2T
9Tr+pS3TTRjNoO6FiRxmPWXGGFeyuiatiTgG4pvvuxL1N8ADw4UrS59I9/bOUrkPoJrkwtvnGb8P
N4VrAayvmUberZulYYMVfPbQ8ZH/7sLRg9jhuEVdzm0suAEBHIiCTKZxiHI92hxBTCDIm77HsueM
zhMnxJWhlSMx0WYa4yr2Q8e8n2rdKQucXDQb4Lp2jcpB2fQADvaSEYUsMnQIaWZ++lCfPCTjjhBz
vkkPLGymsN8+n8yzrZNdv3KR0bfHGKzoF/OtemS2PMtkdJhqIE/6Np8j5ylq7diRKi1BlDQa5N0h
cPWDxSZX4Dl+g2Ly07xEP7FEALgV/JZcXYQvkmobX6obNjCL1CdLioVpJTipTp/F4aZMTmBS6WXP
PCp8SpoGIh58t1KR8IFAHD28QbUsJnw3LtYyqK/zI9C7Lni0cMk0fntislxD58cH4ZcFVh38MNVs
0UOWMSO9mhRssMevgHWWNdQsYlYfquvvB3nKpD0iitjM39r4eyqhKL1ySENrK2wgUADRY16DW8Cj
Lv0B0vstAEb7GoDRcTL7/LoO4BDFBFVyzkM8ELezsphsXGyfGNh52C2f5O4Mgi5pjuu7XvL1fpGW
a1S15PzXX07ZAH0OIY4eXMAo+h5zIqudIAmTMtKF92co9mwxmM3i3QdASU+SqaotGSbZSmv3iv8J
YvcPU0lpKNYJsCFisrYQAkJojWYScpjx9JWKUSV9N5VaIsn26adqQ3dsDd4+2AB+RID7kANp28op
OUv4AWuEAlZzvnZa/IpfXY4nFgh4UCgSD9U3FHOfG5cmBlM1buksadr77F/dxF0hGxZiD2AwOeih
u2t4sm//x5qrHa6MQhGzizvXqVyG/hFyqfb4SE2Kv+lhDFTaEjxyeLBKCIiDpN/H/rOFqjpMqVN3
kGG0sTDpOEyN7zf876oB2JpCunJVfOw9A8VrVgwTd5G5YU46fN5AzzyFUmt7GaDlNOwUUSnx2ige
Oq73QzvfMPJFbUVKG9rJybNNwm+1m6ZKsAj7nCu9VHozL7Ew13VaEeAZUo8dRhk9rpJAQbui0zMm
npjbLQhmtDTqdKhxThWdNN9HmIy5En1VxSu3u5D/drMiFAHwBjoAF/l8sTCuV1C6HQ9Aipo13VKv
ZaIQ1QSMM9JddIg9fcZK/y7iRRQ9WpZ1Me2M3rLjbODbWvcY2uWT8Hjf5lbJKEKBTX2awIvdmWvz
4Tkv8m+1KYz/0vmF+0XtdTKL7Hg21H2CaXOGK+OcdF7KPCRpYtSaJJHb6PhbBFspJTozcVF6sRJ2
JBl308DD483iC04+74U+nCGn+bdXziBhVv3dQO/ilh2SxDF3xWYGZs1hPsWqYE8yYWWTr/8XQbQa
b1L8S8mCF6SgOW6mzKIH4FkrowoJ9vH2UaPZRGSZXXDjGftDz/7dtSn38DjEUl4t7/O2hMFYhCDf
QHKwFQd71CmWbC2Yi5wAOouixxQ61znLDPpQv2tLE75wSJexozm6Zf7056tW372tEn4fNb/gaSsu
h2xQUtVuI5rqUWV3NoFsj4SCEETBAunrKWz5urlPxhcVT5qD8CrxarUKAXQbeWm0pfpMtFEPp4Ft
D6Dhc3ILlxyxZg47j1ZskVljHnczCXgSKbmPKFgNKLDrUDy5fHLF8lQ2axBI3U5XN1fWEQX5k35y
ROkaVI4tOMByl+Y1XRpDN2KhqeIQe3KTlpM9pPlrUBQI3mnOz8KBGSwQ9vVnjs+d8a4IWqSDjZpQ
Iq7I7diVAv8nzoHAJXp0Dwd5ozS/FK4ahr/E9LJUv5Q+6L+xeUUBSsJEeCD7PxaEckLj2xC6Lmp/
2j3WYy8XoQFxNTw9kMotsT8fv2VIsZzTzyAqmDZPwxu23QaG26zs7qwUzHYcGrJIlUzrFKkR9hL3
0d3sHx67RbTWlQzAGd5uF7ynFKgbJKecv8ZKv0S/x2OWz+2TFzZww65VljbPtTVeREu5J5NQDVTO
mNEgZc8XumfR45HfJmVGjmCaavUJoq1tO77sPAu5JhHrxDHZFntysPt6mDpHacwld9yzOVt1MRoW
c7oWbwx8mxkEILOq7elneIixc2msXVfJeVAKMje6a7vm7skroaQBB3z0/Zyglc0ecw09eUNAAL1u
Yp2h/Asd4WOwJ6i7TrKpBuBEorEAi91ngGvaF0nV1GWua3F0PQe5pjPEgyS58mPpTY799LgNj7bk
UJG6a2de58NphE0AKRHzxWwHjC4rco0YxrwLuzDz/Xc7iVPJzf+ftp/ZeHMTj90oZJdYrymcSdH5
0wCHCsm6YP4k1s5xS2TZKsrwMD0Ibu0tD5g8mGYWGi5QtbfDkTJ1h2WsUYbJ1wkzKUs2tRBrrBu7
SdECPIW1ZABnFBDcMvFQwrgw5/4v3L/9Uwtd4zus8lfBHopfR0aItO1K94rFtCDJKS94AkXXzPVr
JBQ+yrukT704kl/tBO/bAPatgIjAIbs5+/+tXXDoE0hRj0xFX9NvnGeNY99AB/6T8ZImMORyw4qm
YtoIMwFNP1itJevqvAvh3Xn9R5h25SUZm0H9JHdQQH3TYvTlLbwLQ7mGGM/I1AD3WuW9jJOXEJD+
xaeaWZkpA7e32DtLAtjB0KKGxI1S6nhp5DbLHi07KDqjgPpa0vdOCehK10gEng4uA2k7FESWhlh4
tUp8Dv2QZvN6yMt2DdgctM2cFUgOUMr8tYPWPxCfYdXf8VExmQnS1T9RyLRJwEpX1Nus+epe2yqR
+Jqwvlj4m2cDZJqpXa3vGyCcbvD6mqe9dx0Sk+ZxTDqIs9CsR8GPqi+JwuCGusiebuOnm0nI38v0
Q3y/EIwSibNrwYrC6Cc2EIJ87RzU0NERM+ah7hOhdix/i/uKrMIkxMzJgYDx6kcCZKg3i68cWL3+
2o6okmdQQ5DFwhgKf4siRnhe5I/utflnrYat2rfIZXTq7+nSQgIfghc53h4s9MjvBa0TqKdE0Vbi
tMw7n8FPT1V/y1k6zlIVCk1pay8fRrLegxbwXAvqlYMD/5DRj5vCeTNtQGCV4+Wz17GOOBUJTzbb
qUJD5WCwvk/bs4IFX15/pWNfVnE671laTqgZRsnQYI99LyHNwM2o9DgFAdmRdCqctRjtk88NnnGm
7bzrNuMm1lRqNkYronU6hMx4NryKQ69roK6Vv28mnXPYDGbG2SgmN9Coog0k0vaekQ7DBnp5XxDS
AQE21DScPWwW8optGvEjspPArubOup/6lP0lHoB40HegSkk0Ylg0YJVfYeyyuQC87mafdOCOgQgg
VBfnkaExYo0zU03/r26vA78aZMFHkawoRmlywDrGVXFxBo8ETZ87rxMDCRwnEP4dUAxlvxRTS2W/
i7yVBicF/HDrsFoEhZnzuCdUWjC60lBNgato5Rpafc7WJdr6NJtX3KhMgA7saAEu70AHOxxCnYgE
TT+Ohrm1Td21/L2focjBgqdyoZBECITxoT61c//oKubx/XhdLR/JNA5CpJSd0Gyew6K8Z1P8aa0p
1S+fnsIKwxJlVaovxz7vQP2u7GBUs9EL0WOMRgjTNU6dx4j7j467AJmBupeWdjVW/LxzMb8iN/sw
c+4femc4gJMSoPwmlNHhFbCOosT0tlLBAhyZj8BsHmMmhqYPivU9bIh7/CjFuJrApteh9bFtX+U+
w4bC+VLnd93Tduizpy7iEMWnS2mGeZy9TM8cCM7sQHmU9yQdd+FhkR01Xe/GDdBfZLhcH21ifEQK
RqVvmxhun7qLvRf2KpBN6dCL53kueno07auIAwdOExCsSGrpG4RylqYQ3/WTnIiI4lftcI9BYNW3
csaZIiIp/1fbjwDgtOM6vpsRJr1NVCdrfgB+x5dsI1n2NZmUSHo9HnsqmrNI2nm5QmDw/dPwGXge
3UAiqEzQCENv1H+4YDt+tD4snio3boPncnfP2/w/bwoRScRK5KvKPf9F0OvfDyFJiAjmb/swKG4z
zg7bHxUXuy1vcFsvzGSTqxOZOzdeLUFBWr0SKHDlfA4YWbt05Th+ZInB966aVHHLd4Zax5ahwsyT
L4WbLqzVs1OZOpbsZ6iyg8TaCCxOND8DGDYM8M22voxASRI0C8PuZVDq2gPsTt51nXBdcS9XGP9C
LbCQiQjQT6o9krYXz9MGtFOS/HePtrGDL/IReMSxlKICSDi6JFZM5+Srwlnu0BbBmfirGun6Plp0
6KkqMDYta0DBX/m4QbEbyfseBvaKILrOd1ClqBBpB+HOESsNsFE/giroc16HmatvAHoe56QoBy7D
n7yH9tOGeJ7oQMrIMCQ0wZrgJegijQ/J4t5wHXGl1RMmjXJ0vEigNgZaKm+zp+Qd5+XmFEkl1u/4
34+kuMKlxitUkpKcGmtF9fdp4pwOwNx+80qPyP2q7cXcFgCRneTDsInFUry5rSkky+9z7qYlszk1
CdULeXLelS2WiSS/Bh4sEFINkTArHN+aTD0BIq9fr+NwTZ4FlH5sZ3X6o67+NxkgZPo87PrInjxj
tZO1pYs/dFtyZ168sflcuzmWFH5hyPMCuHk1PZqfwluvDe/fgU8ohvhQKU+GK7rLAMLxbSNdNcBj
IvrZI2MS8Q0tDNo985Vp1P4RPnVlce5yBEEt1SXBZfDXPmWxTZilFl94jMVxsRNUbJjcbpGasEmX
Hr7ZchZdq3bsbyG3NyWhyrMDQavlKN5fyhUW7NqXk3pZHq6G2YFxUajD8KEHrcgS+YxvxeqW6vgu
Vpp7qa9ZM9DBgAJWPc5EzSZd9/kbZ/JRxaQWAoG5TPjPqxM5Z2MVlfVprbxjN3BsKYhEszayTm51
qKp6CSIu0QCvhMN384+zzJ6ZcDzXmPXch9Pi+zaomfNXDafmUdUxlkXCGxkYaR5BdVMcahRdAp7i
MS04DYG3bgwn1iz4dJAFIuIicfuKI6jIHuh+o+jwyH03u8VDGMiICNpoD1hNAkZGf/n+L8DyDCqd
y5Qw+hL+T1Il/0gWqOhjogEXflVAfLc/O2J4oW3KuCO+oBjjV4rV7V16ezAFgkMZQRGGXcPQJVUJ
ub73T5kc9DTARpSH2PTIGJIhhZvQQhfpWJSVMf3U/bVpnamkx02bCKQ+e5acMjshEwVMQgY0DGqH
iRnCs28GA3IpeXrobbzuUYyThsj3QPNq9YimeDEZallk7fSM8gsv1PvRZ4kSYZ8DcOWHzBM/rzaE
fsjPMgBtlWzrs8JbGK+2QFEq24WhDUKLUXBtfekeeXPXbJsGlplKOZt3ZLXxJzflotSG+fx9yZ+q
6mXH3X71G5fhg9C3uWJvkaaJUiBAsdXZPh66Zfnr07mdpAkMAKeNc1KvK4kMwbPQwYwzPg1xvNUf
Cd5vvFZwI5d/y5ED25ayMJ3CuBdQ87cykgkk0a6FAJj38ATvJh9snrMGC8eE0njiamd/elLYV+BR
wT6webujvfKui7raoT0cj4JrOtLvyLDkaAuSwr+SgBxVSfJZHvBHI/yGxLg0lA/euCEmsibTwip0
Ty8HtrTpUKlRqCcKkocCn9/OfC+gNwXJ8DlLis2g3WvWu+fQYCLMqFDqhiY76DiOxtbb31u0QgET
2mUKQT58ToGsxW9FQB9MpM5p2uZeILKkNqZR/XtQkPUREM9Zsx7j26Hj1CIsvCK4Shu7aWL65kHR
12naGWaBTe0ZC1svSyJKcqsXB46zPU8RBueHtwHYkvWAlkB+hqCbQ7kdIOCitR2UQOvSv07oDoUn
t3iiNq3JD9YhJgrJfqLVvAr1Ib3zC4K2qq5nUyfVqwYVTe0aMngMwj4yuyX88SfsIpF3EGoiXVR1
PBsezaL9yjlrJhHt7zxr+EyLBZ6bm8DAqDoCkovShB5ZeaZ4kfygL/dCGbVmhM5aixVitFAKGv/L
0lDXSSU1H1Iv/DGNys4dHXppic4KEH8biMhbt7AGK45f+CYPBfxhJ0Whxj4nXh3zcshBXIXyt4NG
bp8qAMXBFHipcSpOHFf2wq5SSj3aOZQ0Ful7UUpUjf83B/Gt1elLqtdB9+tpAcS6CCOjklKxSni/
D2yw1SYOOa9xSFfma5QHq5e7G0DZ7vnLl0PWr9cE/SYSDhkDH4sT3QJ0dqj7DeRZgSE0t/c5kvE5
h5O6/S9Sd7Pfd0JiF7dFEy9fI60RYmVwQthWz9LO1t04cY2slb5fb0acSJYdIuXQ7NBz9XinGn3+
JQJokaO2EPtpodJiZiciho20RpSjEb1NfiOt2ZNHS5oBuN6T0CPNvr/uweZ9tjsQaUf51AvatUld
1Y+HFH3d8+IQ2Qun6h9bpvNWCre1svNiToMWjMSAqVPNU1x+CxFK0BFNBIwwzq1KnYzzA51YB7rP
uNeYW4xo1ESWooxi03mwD03yYyEIvYNm5mOnI/8uBe7yiPzG6sXWiNApJLhCKANeb+I2RNejunyb
iYw7wqHpON/RrqX2dUV0uQLfIaVUykqjA2x0CMR7Ty0qGbwilV774kkzjIRTq4nl2wq61r5QrNzX
A7LvZDAwuahfiGggR+ziKm2yiY/NDAcSZYbGABf0YbbIj5FiiDneADawO0yrXEPtLA6v2IvluFUx
sybHEGwp/eGItjVVemsNLKq9yG9ylsCanaVZWPjRvzd7pn+zVTBCSftcurtvhlcTDI8yOEqNc2i2
xNO3fyRI7D7J38ak7e+JpEZSOWckL3r2+01hjH02F7oD98Qr5DsfvN2H/r09epeLHVSdALyQo8dz
Yi2mxjoZE8ZdIayTmyI975zWu6lNuIQM/bYSeFGJ34Bk3Hfy8sblWXQGNgt5IPQbjFrz5Orod0Rn
cGEhlnFEnjbSgymQn7apO63t58u7FjjVH9lC/mJ62wIMeSJgevxCPNXZ5jfzVNQIJAONjSV/I05Z
lPGMaFcIqx+26sFK5Zdek+8XLb+pdJ/Wbqq/qtHtn+qogJ0+RHzIbQUjHUOQO/Bu1pGyRt58qSq8
s0Ej9fsPYERoJ2B7fPyDRichT6vdcYpI6yyU4N/Bll6QDgmxyvxeujluH6pth8chO6r51oX4Tw/S
m61cLGy+KBkTNu+x/UBin3yEuPp9kHALExmJj4Dc6rX6dii1QPk8OOW2LEFeEowGnG3rnsKkH0Jc
dYaTo4AkCczkA9o+o+IyT8Tj9HZuletnKVdllQXctTeXfV8POVBqa6iQEq41atFULztAMlHq50ST
u7dj9CwfYeHoPAEJJiAu9zoYSJ9ppCUzEE3X+OAUdh2vvt8EKoIzAQr1poi6ETn7K6pODEatWmcz
LVI2tQt3Q1ktZXUFQTcMR1CX2xQTfejsAHup02zOXUAYPaFHGUJW/fhE0GL/hhkCrVqecQ2UztaA
LEo6oGii6kPtSL2cq342MhV5SRVU1pBgT7jZcfSwJ4EM829nxiMA+mX4BnGwr4cAEk1wwykzdaS1
6LekpYROl3r84tlV1I4sQw3Gw+9vZMpfuh6008nglbAJkOtMCJvhbAmklQGW9k/5MfwYyZhGmYen
WYastCZoIM04F9oTFxCt+y4JosjpOLl3RTWyu/AygTa126CID74Y5pWzFKqviN2S8OsYM6r/Znqx
RuOk6nLIIkNY1QqdoA5cxaQzRoo28FlHKwT0i48K1JOm+SEkEFF7bsmB/qD+J/il6zp7Gc0fmltP
AUcAMW9MqR1hFaaaEVTee/7ec9ZsHkv+5H4edq8sy+nNr2LSfxeQn3vIRtv1A+scbLV2z0+tIh4e
oLFYG2+a7lwCHK1eiE9XRB3aaNgbOTiVQhIH3o/DZlASBR6EK4y5daeWyi8EH46e8dN908LJJWwZ
YgH7d97/KKkpe4mUvnq7AggN2p02ZBBiOatDuUMGyHN/jWe9GnPkHSNLqy3HlQnQ5RdK6XrBFe10
LdRdsyTMxnZ7e9MzCp+jeT395eDTBeyNMwnfRHmai2A1tZm29KTgrtY8y/U4y+t3cNsV4px5PHLd
uJsl/r/ylCRupYYP+zKYpaysImZdUS+92Fg2aNO55SYc5Ov1VzEcW9juW6SLaOctkCkFKcfwm8f2
uS8qvDWWfrnC2a8S7p4Ce3w8XcN6J2LfQOlecfQ6NQ3eo9vHic7AZ4KfzNYvriMBro+zGXvsRPYA
73HAtyr7x7uvavWT+XK/GTrtIXFxeEZT0HBpAzpA0d7dJyfBJ7WHavkythFVHBZcP9buHpYF6f01
80PDyAFoWzYO7YvKqibUOu7qVSyd9uOejd4E+pVIDjZrUrup2vFPGfDBjEarBilEz8yfKAx7R2+i
psmThh8vbRbGQmPsYqnHcZR1LhVW54QAAkSR5iVMZsPU4E2gkCMmZEeWU3gMbByOtP2Mv+0qxRMc
MoJwxSVL/Jqxha4YY/QrVMCXEMhh/9OjoYF1E1s4YVUAaafJWV1P0LVAXjz6NucVzR0k3SW+BgED
7fc18AMl+rBGD6pROVERABkEmaXO/umiQ0l0amNSYFww8yqT2k287kPBDzR0B7JL5TPaeOee/pf3
xYqjb2YUNGcZSU9pCX9r1VYEKR1qdU1iZCNd9Ct+7BkpxiRGo4bPSmfNDpFw6T/JQc8h9EOO+Dps
BqG4izeY1/rAV4DBYMMGDTYQg0n9Pe3WY/JZaJYitP1XfWnCZjzFrXl7QJxbuBKd864bXrhOhCPo
yyTKQtiox9KioPZ+GVQ9kQ4ajZbY/p4RJeB9SqIBOMEx2KP6cf0UEqdSM6jUyT/BvJObXaqpFpcH
Pi2GLokEaSX7XkXv/KPVo6mWcSBHdZ+YU+ykRgKI6szeRL8gm86TG8V281t3iq55R+yCHR7qNOyw
Z1iYJa49nThTs5/p/nFoSiqbmljKEiv1/sVu8GcEuhNaHxxJsNRYuS45mfnzdU6IHUARfwee67+e
4+gjK2zakd+L1GbjRtO7ttmGruQwfwcA5kh2sODugqIzWX/O1Nfp7Slp7ClMGOja21+mda6hkOC/
80k5WCd8RFsiZG7JOk0RlXoZJk7dtdr7EuRJZ0wc3sfs8BFGQtrZ0oN1Z45kzZsK7Cu8n9uePjt2
/SwlVA6swz9M1oBMMgylTgsCMTF8ZKplJ5vNQxQyDR1LBILAkV5ge8lSQ6jLLZr6s3+BFfnKbiyw
+c+llZkWjgXqTCRL8DTs/F34UP8fqAB4lzk9B5eUfmYjcUbPpQ7gt0QAqRr0Hcz6vHx/BZfr/66d
Shy3QEvlueBrdof5hxsSl9mwLROQLxPX2dE87UkIVjuGOILDO09BuW6ZiEIb4oW9JKHuO7JpG0NQ
Q3QDb4PpndInv2LlE6gNgnJM3BDfdFK9Ql6n9lHiM1uMHxXc1SQoI0H9v5uTUKzqBMrBuJKEXOMo
zc8WqD1bG5G4DQ2hY2JstEy5Qo5/hhzhPqFTXlPzJBEF7GJBu7goIr/1vhSBXCdQTNutH3sIhmnQ
mZ4z7iFhqSX7N/nltIH4vEKS7ElI5KHXUX7oZVYkrIcaiYesgPHkOfDGX8JsydlhD+lj81Txr9wy
CLhBn44QGNOoqJFG3GtccQU1sqkEvZWzTzl1D+mCQNeAp8ILbfOzzUl27LFPVAdJRsf2AqYQNGf7
hJGwNRVTs0dsPaNW8dudy5x1dI5/0GLN0jNHpJfTYKh/Y0AyMkAdCMt/WHrjH9tJA3ISwwASwyti
nOEE0FldlhZL7MuqqtpjpPiVZmWhJfKmtnLCqanYdmmQlOT5siu3wAxPIZbz5nYwknxUBOCrHjEd
YaNyISPag6f9Bdmz/lespuHIQHdIsPq/EVZyzC8issL3KUYDq30omU/ZH1H1zZUcHQM/TlqVlvoc
rI/9xhfxpR5JA5QlqMjVLuexhS+raLhjsPWeQvtbvIKbb3nzUsEezb/CssCcIXI8ALxvvF37AoYc
rasdWMmhMMKNc7lLagt3CONprfV2fmgREsXWCkXikfONR3ZW9sl2kmgPD4+Q8QQ0D6j2n5rn1Y7m
6McKli13Ys1otVvzD/ZyqjwKez+7q7FrcB9mQKnaop4As8Oz0A8NsXI0WtTjPOKUBJFCw6H7Lebz
GxDJYPYEFzHi+v5x8RRq1scdyAlS8pgB/6VAtTHwcYXulmV26WgbHO0+pOMyQZ1O81+0oxtMMe5w
+3dUuWhVdO5E6waGbaSTS+/Dte8ejid7DcSwB+dllohhmDlg8eoHWQenWlUPCQNohsLg7yLaCzaz
4+r2SMoL0NH4nq8EvebNiLcj8HcLZQ+ta0/CL2sokpxQfQzLWQR+EBt2rZRnb2YDupCtCRUy6EuP
KMIpuABGH5+Oigp3auQC5ImLkMAlXhyluDqVrRXc7jBHDXZCS25Ro3poTw9J4bzUirylmBg5ge/V
Esqv1mk7ux1Oraecvd92my/yvAnNtynMCIpkzf//fxOfngW5LPShLEoUNuE9Db4quPSFBhl4uGax
wVwuXnRcRvi9nyhtsgR5sFxmx1h34rkeZYFOCg1asioqyIbJdYfTtA7RFd4qVImdE2HG6sMvGhB/
U9QYXws41d36dN5FLOZfNbLsDJDameop9Jc3jJ8OpzXYlI0VlR6NeAYf0SO7Omy4Xk7jNG692xKu
9eTzGnozfq9SjzQlUgYH6jFzGv5cp8IOw8jJXG5k8oXejyi01+rKJ/fr5TBdIpoiOCIeMDLwzOFQ
oyxWlnoAub9yy1aJI4Hd8HvZvMO7axTq03e3SfWk55PyjluUS/p6vufxdpEXih6ubH93YGUMs+dc
GqkS7w7FAGjBZlIL2uyeurLq089JKGaRhHbmGmUwLc2pjFilkQrrnLP5ojnnI2U2e79QT6a77L1x
Uuy58k0CkiVtrfLSxgSogKXHRVWkrOmtHe4W8v20WgVo8IICWPuNAV+i/uPa9wzXAVwfGSzxxV9T
Upn9a/eZFrh967h8pkjkqVahd6imRBs8lmee2u4Tpslslut8rjC+XKKYMrLScUuUPcYREn5iaUPN
aN5X2/vIFwaYQx5qoEI1wBnnQH2qolg62/8xZfzouzx5N9cjFrh4UVUFaXtALNaOhc7rT1Sd6uhI
7j7Wi1zb/RZzIjYocS9da90ZKFx5A5mr3/7N0999c6Ac9DWIJy+ws9otUx46BAq+O1O6c6mExMkL
iDLgyCEtZN/Enlxdft+MjwCl4RGhnMgE5lOy0gBVuxVQapTrX4w+6Z6VSmQYVpXMy8+wSlzBAoPH
3AwuU2robSzQ/Fvw5QbNTuugFOCbXCQNtEPaxFSQYMJdgvyLX/ioE9DAmuX/75ioUOYniUoPTJUy
9f675OIYicuWrx/axTLysS8E6gpispWwbf3kacRtf3pk1E7PV8MvQq3OBFv6tkP/FK9DRbJc9glI
ufx6R39r1S5x2hwv+JzdhnP2UKS7li5qSSFfpg4S0Ao6ggrVYpVY+CNCmTqLZ74c/kqFUN4ck8f5
GLbcQBNyuoslAAByvoesstP0orgRiYnXjMM3PGWsDaBKGMlLePK92G5l/T5KOdwJFCEsME+txOn2
8oLM/TdUI+cBTQIR65DSHphHUYYYP+2G+s4uuThbzoZo01ZsYG/+wSemU8ooRrPBLoR7KZvx5s0Q
O9hf9NsDqzNuygL3mT2JSLiuOqUMKSXJBKRn2gcW1bkU1ENg7uFbDFPW92oayjzXXhNrfNWwbI5G
YNtFaXf9y5YdmuyzW4zlfpYHXcIV8NTHEojjlZ/L42/vF1XtMdj4heOQHq06LIHBssu14wwRwHuK
Pt8u1MOD0F5OHmhVqDBm6r1llBn63J88zI6O3dJiVa25aH8l+vINc/CURksT6K84fA7qdlupTsPc
YPkcEsbuovYC7qwCHUKiU0egGcJ9IZru7Ic9bA2XtM2j0wvB3Z5jkCgI0RYpsUhKNzi93Sc3wZAZ
St9IbGoV0pXR9CBLRlcYzTHd9dKoKo4wLs0FPyjR5trdo+lcCuAZdF0fFaHhsGApCkEfy787Wo7J
un3fjJ/vqCj/yNIyfzxjZILC6ihVGmbMzzkOQnWtNAopAxKTlKIMrBAsMvGOJMH4lD/Qk1Wi8XPB
9v7dfSfrJlgRt7unZg98YsYXEjj1P4GsmMDgdGqXVmts/jDWKtg8fYswfacFIC1+ZCH9fia1iJc1
I9q26LUCG1l8aw369E6+bft1drRVozkU8FcIT4O30yfnUoY72b+IbilJLBpl0xtJBxAxUcyQHLAb
WsIP+vsUq1Z7aenFEvYOLMk8DsCcIpD8EU5rYmzO80OnA3BRR3t9p1b34my5aYZYhYzNTlSgkhgr
6ekc4ic8IStB5MvNqkHgDY1qe9c/HskkVdltl+s7Xz3kak1YUmbyl8ukLLlVrPeQnNehy1Fhs8LM
f7Jxj+9v0IkU5b+OJSAMGqRZoTUFAX/MIUwxuOeFgYdWp1NeSwua8w8qgH2laU9LoHV7UGcD83ZF
X4+CQZhyQAhp6VgSLcHIYkfhh940I3pfSzgj7Obar8YGu8GFMMQucUm5zw0plJFdSHcs0RN1WCod
8DZu6oKA6MkW5E4ks03rjUSNFHKpBCutHW4wYMcIhLPt3BHKn0zn8E8+L94c8z/snA/xWKQZQjJ3
VTY7H07NUWMc38zqEv2HSfHo/GaHSUzPYBMGiKIBWsjmniTvak1nMLji908DghqD8x0ccIo6TA8R
b79EbmvwE7rqlGcHHG38KCpsprbboOXbThSBnGjoxw9NdEJ0r/jzmIAPCjC+iH1zfbZa3zCgdXNi
AKGiWrDXoNz27RWdwBr8HsSH1S5ZLGZBTS9UE6ZcrucelKibp6U/vKqADNHKUIAlTgzmXdJrkW9J
O+Y8OkIKScI0LujiGrty23qqp9LqTKjQdFf7bodr7BETsr3J31DYVrj/cIXLyVhmdKqsXS5kow6G
qa/b/XRJy26FhaJ4eR+W5tfCV58Oz3zsrgKkvwhB3AwGYk7xujCY2ceQlmwAT86+dT2+az8LmqxJ
BrVa3Chl/i7BTh/GXFKMeK6CUXSbEbhKtdcYRrbuLlnbKFSfnqt/DfiBSxN6t0mpCzs/RS0+mjd5
GYh73mwdIIbn2AKSprJI6EN1WZiDBVxmcZBEHYJ/JAAZvwZg5hYQbDbfBJ+MeuYWj18v903Y9/zR
pueRSanxHlQwVQzXNLfOfLMb7m/nYU8Eyke4ishr5MUyVXptYRdTwssiUrQImUiSAQiB3mcQDdX8
cTpo+FCSlAhKmjGKI3Km9XIX7XJFpNL/gtLwLx24QX14EnVVrX4PlR74kEJK4g01Wa7ECXLB6Bov
dxSJy6nCl/Cq7qejdGLTcVEi/ZTRickfVx8ng5IQ/f31axzfwL/qetaBiFosqfCBc8kdNPrNXRT7
Y3GVfW8X7ArUx6VnBynH/BRxrDMpBDZljVwR9eMJAjpbtuaWD5X3FxPUBKudTo3H74na/nOaeUYd
c6sWpxtbqrg93hQmPEiUI4g/caTnp+ssElldf+BNThlf+KJaNEw82W+dxD+aLW1bDiSRffhGFzWw
n1JfDJuLlXg6XQu71fCgYgPfLcJ/n4hcWRDsaZcBKT3ccGjMhSeBhAI7B38pbmUBzIv2eQxoNeQX
1ntuthW3AFLFYUWvjSdet4zByWtdpH/NltyWqddWd91j8Cr3BIS3UiM9p9h57/aGOshTBkcW8tAY
aKrSI4U8L9PQnVRTT/B23LVw5NO/nJ3l4x9LKFp1IUz004R9wS3G/PqbLJ+p5JKbzbZl5DBK0RmY
o2+38WJC135tRAZvCxWS1DyrhUz9Do89EqzOC7TctnKa9tQ+bkDR9OONJuiYH//vQ2lij2a7T1xq
qo18gj3adOpXL+cliamI5TjAHcrw7XzPfZSZlXi6WRNT5a7XREx7RjoTKD7W/gVJDqZRPA/wE9/6
nDHuLxcEqyFc96plM7Nx3j2jLDePWLxao5lUo8Fx3LfX3uKglKkx4lNfsamdChCQjfNY+zf5rt/Y
WgToUc0ZClCz6HNXkT7QrZtdj1AMhAG6bXxQp8hWfFcazvPdJB6IXUzpjKdt/ByvsS43R+nmb46L
Tci3sT3MOfkCBmbV+Tm3KeRnnfWWxaZ5WYd0W/vRivsIFTDwgsLIS5V+aFSwh2EZD6KzXtxW3EZK
3kYtCOF0k2m0fjNzPO+s0kEHm6ZslA//bwx2N4JvZvtAh0akrRqK2Sq/r/BGilqXr3pCJeECB/kQ
TxnHX6V3tapPqMyaiS/FioQrZ9+tsgVvJLNSfQKBvQGnPrp7oS7c5L0cmeUYWQBeTlPvSzISkcBE
SlTpuRDAwJR3JgAjHExFzYNuMsT6L4Ys7IuZgTCF50kK3LIkLTwfGybY7y+WU9pwhO/hg/vEA8hk
xHas7Leu4fO7Rddohgt8UDF2qi2CXsCLCp/QiobKNVrWa/5DN1dGVYL3EEvEkfrZA4Ipv22duzHC
zWH7w02m6lcnHRUtIC4CH4fhD8JH6CEjHIN42YxtPrvMkv5aurpT5U016vCOlt+k8PIIN52cNaCL
D8o16JoBK8XmZzPXanOqEJEoGx4N22ybUf3PZy6bT+JfdR8yaNMD+5KLCb0diPqevgXfWpVvhylv
Vomvvc0k8Y12btjZH83uxecsvloX0aGrHICEh/HfD6yHbbBaXoWmakz6I962HgtLAMlr3oIKOQeB
Ust03vRfIPgH86uPewWKUD2s/+fQ0ZNbuuKtUzQEGQMe+ukmWy1H5PLcl3A2MBWyjDpQwJjIuo3j
QaXscS0zAYtqn3gU9Jm+CALitKK5FZ3VOAy7xMKFeAjPLEgJrD/Yv4vSkJF1iz6nCXvSBYsi0R/F
za+LAldj6mrEQU47br6hMcO06pruhhzsYXw/TmxUBkjZWIZ2qyoeZtgDVaiY+g4ultW70LwGx2i5
R0Ow6FFeno/aJlYyQ3Gh2l0ELwrxs2X748pPxM6xwsqHfaeOlewrA3Y52RcmGVohLHObTOlesZWv
7kHwjYLvKDYHwF7NEdIwRraxbKEQBqffGj3eeAYWzkoCJ1PWTlJ3OnGMDGZR92RrXDd8Rk5VJ5GF
/qNfc3IslGZlfoVP7NXO5Z8p1EgcFhBuBG+0NSWuxsV4oORck75MRnvNWhH/S9C2n5cRh3TIulQi
JtZDbd/1n56RkASwINKLUSOPt0xFUhgLImc0G0UCpHNhVr0khzjIY0TUcd9Mb2yblsMbIZrgzoo/
wt1RJzyDRvldNHUKYD8yklT62aV+w0prYfeyU0Xn6ZvHKbyxQGIZ4YoXNZzLS7bo5Um4PnJAth/+
5GkdqznoED+PGuP26ffcjs69p8PzbcU7fEllAwRKfJfYi9o3GMBpGYhJ8SSTVmSjOtH/QdpPgIKA
YgLAMggqEIZV376FLjSdytxuRyYRzHKKiFoBizKysiS946PzuLw1+G3t32J8643A10IbrNpR21yM
//8HNbYMkU+tfggMHz2oGQALL1iywtKizjQxqsNMrSNjUeu3gtWGmPTY/sByGLt/+7TQu++/Sc6B
Gk7B4/nOECeswC/YN8oaLLKIuasv4gBT2uBHXED/ocffW6n0bjBjBo5zy6eEiPIKMxpOA6S/m1zA
UinI2zpE/EEluPPqf7qyzR9xFEcMRp+MN/C7T4GnV8+ii/MDz1BVutKzJS3PiNIrhzFJ3J4BczSe
XGcT5ykecqnji7iDkMN0rqVuYlGP/vbMAddioe280b30i+/beXGazS/XGQtk6iVJx/3dmqV5d+Ns
tjdbU5Sy3KpkBJ5laxyU+cY2zXu21ir86QKmNIzBOiF2IqSTQWmhGsI6j+TJ2gVCT+syjy23IN7a
o79j6I/C2l2mRj/X1I91QdaYdhPvM+fdXN6zPprUm0Z8ISFKWl3pell20tKWqTabgGBge9nqeDga
c16IzmclIWBY1SMKtzBB+l5XMprJ2KBX8lKd/aJzVZiLP01vUEvlpxNQyG6I9qAe/aYJ/DZyKKeV
G89Hb8XVjdadGhPwmuD6bEXvp777NRJ3JHaX9o40/nLNY8pCFIhFg8CWgWQJRnpViqGUU8IE+dt9
0CzkV3zStnHMefbI1ZiMddUfjwRJI7tVruZ1uy+Vyt4rVb0XT+7iASr8eIdj4abqHTsDCc7bglNE
rq44H2VKBXa1TQ0jFQlIH9dGloZSUDv2ABjWz3U+6m3mPg6wc3lR3RQC0TN/QjFvur/NXYwypg5y
+2pmDAvBRDLvoeSro7SPK2kbq6mDtExgMSPCrp0II1Qr5Oqf0CormD74mQWHLWSaHQJd6PwAwk10
h5r5sTIN0FMerM9PB8/NN4bgh19hK+N/OZ6EdiBGIJW6XutpM9+Bv5md7o7zssnYssjH4Xavooke
oA1+AZTnYNBALEbjx1JgZgfrJvFNM9noCMzdyGkfm9Oc5PSxwqx2ylwAluHKFn3zx/ERU7JaHpTG
LRKAiT+jxPl28fzD//hYwgmIrpQDwcLTCGP2Vh4sX1bwaj4nCB7rar/pnVZv/TD7V7SxjwPfkyM9
E5tq6ZVbR+Oj8GiYjs0KiBn5gUw9jnNPA7b4lUiOc99xivj3NqWw/Iv3/rtIo11BWGlBRbMlbM5o
/p402YatcVHwDVC/JBJnZcTzhkEeq20OdhG57T48rx7hhonCNsAlqG/zPSxtkrWqfUyJlPzlFHkS
oqJirPd72Ho3AenN6hYxpIp401YKqFrfTQefMWtZEVa+eAtR2HM11gJKa2V7jihV9jE3BZzgIThR
cP5jyGR+NLRBBJZnDSQ9vh9M81Q9xrDjea8y4Fb0vcovcE04oAlLCEu1mZYBzfENJEjtLT9Oyk3V
Af5xAmst4tsvNAfHSoEGIRmuaCgL7UPqozNhng+B14A8L0XwYd0a2wn3fwjMFzfiw6b4Z2UAhklh
IPBOtBoKnU9zheIbvYHXfyyqS9IWRPJ7tcYaM2yJCTdOCCARlSBZSDAMLOqOYrMOzJfrI6QfQM0d
gXK1HUn5LSptq1o80KBgG6VLOqaNyIFWTZ6MCR00XYG4P4iIltDofzWF5i3nntJOUfsyYtsOQAmp
cRbuwILRqTPLxtxXDnSyBwyMwv+YVGjMiEff2PcSg5zhAAAsCVmCNMSAdMHITNs/vtWYKVBBotDv
WO8vwM7741RHqu5Yux9k1CURPIuJoPxv1wY+i7gVBIifGN+8LQNN0rZxBaiRuWhxTu5Xsi7yveWZ
N/ngxFasIdiJgpQ22hINZqWD6PPpi7H8IhfGmEPclpfbBr+iex7a2+ATTeZi0anAgg3rHxATbQJF
1iq+oCPnIS4ZQXAOW6xPEc4ECxU9m2jQZ4fkRi18EV7JkchQ04YHmPL59mSEZF+rXT6eE/vkpSG/
hleIjtSzjM25hLVi7Meil9W7X8E+atN07c2DTc6079p/LP3tzTxkZZRiieQmXsk6KtnqEIS3VFCs
buC+XExg+rjZjlOu9Cg2LmLy8p6LH8BkFBUnqx06alsuz8LZfsA21bhUOCIVqRgAW8hQB21DAHCO
0yg9kPwZlNcigwZfmYp0LVVfpjfqNLDNjYrjz16skHskC3gtmiG3rePY+zQ763q1SZF/ZC6uYHLR
cYCirkNjXBXPv/5wO4p0vnFuIn55CsMYWMv9SGHNQ7IRu0GQnOEYII2xd9skBrNCmWExC5kC9K6w
ymhWo5/0okmqqep8zi/+R2HivgjiuaLRhTsEzUE0q4nrthYivROXgC1Jd915DmkUQrC4+lsmbUU+
qEWUK0tVOBQVnpSTmL7KCPXqmOJZ9aw/AXBLVnLBYJkjNmuUMpadMW4FmvG9A6rBuIPlI0M9G6BI
xE/eUqUG/kNM7p3eN7U6WocSY05pHdPk1cBX8PWzSX7F0Qzyr42hyQjqUtxtIsz8UWF6vdB50mJl
Oksaqf+mbdHLUNCBpTDYa6aM1kVq+wyvNKO5TmeBd8kNJYrAToEI0S6Cp1VI4nkZFIxV17wqGcFo
Zs+/dUk340QgpjFBGngmJls9pM0m8y4jgoTTcpyrFZTOjro5QnqrhUptLaK3VgRcSKxrMayGLWbz
iDd8rTiJ0OCZBgwG+nw7cHEFNj/jo/oVTuJIyvmNgTQU2WMx8U4X//iWCv+GoP0mVAV/IDV0NCw9
gb54Iy5wWmdJFROEHMWGBClPbEdBnNZp9b5ll2Oys/66bakHk7lufs2I2JZymABP0tMq+YOhjfR/
O0lzZUBN2g6lIGgwvmZISxQchkvErzUUm1Al0+ir7pnxwmoZx7pKXYW7sx/uuNFZ2a+QaPR7clf+
XK8wY/0nfoO9iinNEw5LbJu/IjDMt7oMJ7gYM3QC0LVPqGzzQWO9rvCuTJmULaLwz05J9iGHYxeX
9V+asnmcoyXhtJnJBKg8A2d3opfr4fbF5m+yGMi6XCDhBIaUM2AAfeMgWIM+pAYUNFrTwtXeQJ7S
dqhOdbxBVth/AloTWLMA5103UjIkichaVG8T/lAsrXYpn/vk1GDbTq2x8Q1KKiUtDedVEchqU2MX
tI3qF/XzhPVT1VO9qR9DDHMTg+GQL1lswdGB5ay2X6o8UCQCq4ZG+CVy7DowkbdVoy/yOG3Kf1iY
/U/ORyaxt4kWQB01XiEICJX8eUSba+8pHVoUOvS1BzuBHXARJImZ1CVnNAheNrESwOCh9XpT5QHw
pqgjAkVsLYsDaPsED3gCp2OkQaG999nKXdcj1k+FqJJMMZhxtiDgXegC7iV13YFC82hV/ZqPYG+A
Mrw9E76/3+GduzXMlQTDUfrlArzwl0O9xdseQFk5tVNQ2PY+EkjARp9stGC8p8+HIFJlG/8nNkLS
lRAg8eRewnJX4kxU16x77nsHpbYAaSS3YuzaTVxl2XVTRX/ocxCiUf5v0b5aPkrcJfSSherhopGw
/fQiCNai1L6iGCtQ5SG7Vbx4vny1dfQdGZSLoqXayPElelBmrRa5qJY7+OlSyqtxYNwBex2d1PXB
8fh6XU/IzE0w5/yahcLDPcrSDWrQnwcgaPA0DjRIgJI7rTehR/7QWNdDRDb01rnzgIO1mwoVVElQ
rPMTs28Vs9lplIYeM+9E7WuRmi00x8Uc223HeobfdksrNPt8W+QZ8jy+D2oX1M3SUOpOg3tn2JEo
3Tp+jtcWY4PMN5V9mpLdM7YDQC/cRaIgVHuVgpXWUiGck03jRl5PpchmJXPtkrdRNUCWK2jmQ3LK
BpxCJVx3mCCIddo/w/o1YPV/Nt15rpUu9R4HubLBsRN/SRUXsOQcvlNSgb6cjIJRwVXXQxta0ZHM
sOw2q+xFddYEgYssX915/fV2ZHdh9or3shhKQMMgf8V699GPja335bA3CHaObRd47TrC4xG4zuVt
mGhBTmtA9M+lsAXsAQGPnGNR/N8I2QjHVhouc0WT4T2koIbOtzDC7ARPEbkLZBIuPa9mBonKO8zq
5V30rTpIQtv0kAMrq4fGilx0BPS0KdZKxKGePlFsJK7N9L94q/4h1yaiJMhtkxsZWGXCoRPPi8d5
9U8zxCVZiOyMBAorPizAv/UFZU8+eHsRwBNL6jR9tLA2nUxfuephRJnIjtroei81CHongNXOk7CS
2VQiwHJ1S2RlgoDYETkXfe2B9soTem6ZmcIz9KBzcGr3KHU6eLCPPmx47kkBdhe7VJQ701Ppiii/
PB8prwPMaoAgpaZ7f3siIiCkdyHU7+oPpqP2BmZjakLwvSmoQP461sMW+wmLofCSVxOny4dcOZla
MW41ksSueAi6cWQs31+OzFc77oBshVPaqbygJCYTevsN/1WAifYKxf1S7c6fOzuO/zYVvt1DXObq
8Th0E+7fI27Y0wJEbdkf7Y0K0oY2ikhuK2AaC2lLhLSr9tiz+uDhH8lKM4b7ZKGrAh3JVDJ/eAL4
WB18J84sLUK7UxTVipoyXiwhyhEMbkp92zMMc7vZecY2V4Qmsmy2WMZ6rNmCfGzeizha56F6GQUP
1GecG8gK0J4SjJGc5RMWdAhicWeNJGwAAcNbHoqhUrahjunFawL4MCb2B5WKjnvzXXEFAAdanZ71
C1Mg/w/nMMoJ5H90aSg0S3c3TDvVOhdg2cCq1/78oThxdl6wGIzu5fqInXH7sTvMiQhL3rdZnbmM
2s3VxZWpVh1LZ/y2rIFC2diCbykdTf3c5z7OigVne39qnMeVxQJIYQqEYJpn2Hg/BIIVJfEIPSPg
zfSvVxwhsYS5DLZzgZCd4piMGUEhhTWLp2oqMbVGuX97Y0S4OarWmlyIzPpxUG3wsE3GcRXk5DAB
OJf9Lvp3kOGvBZ5Tu/8/psBImFgocxgPaItGXUlmkJ1wiJdVBLzmm9MexkA4QeteUUdDxSsh752e
eMUJXPtjI37bE+3MZ/qZm5jqlxJl9QWLWM4jicQj96MCZu6QygJXB2HHWiucIrUGfPqXVdsY8ZiN
oA+n8yuTwZ78fMRTZ3cUjQhKHlNHa784SH6NnIBr87/YUk7Prllq7uCd8oQOXrAOrPHH18+9kjp7
dcSmGUTtPiuGWQhmkF20/qa4BmI2Gv1JO1d1+l+6pxaBvianz17ZR2owjK4jXSVM/D3cdJucTAFF
6f+XCPF8RniROPZbsrVkEs3BtYRP6bv0IOf4gzMae2zs4fKpQh1C2du4zQNb54JoW4SEsa56P/IL
rYMoy46EkOhqQthhjQZpYVylSTDrU4mI1EFLz8KEsYqPoRqmXxqYjqYLkbVn67uJ/BqIbgG17i+j
9DxPABVyy0yPKklnH5K91jlmFIw0gyOXQHDMLHbAOf2Z6ggOzeRqSzJXxOsUlLRlOnRGW4FaESSL
8tZSTYx2eOaSMkjyKmOXCsou3D3dBUhul4SmO7YB5Dpp9tcBnFsQMcL3RhbnTUHnvudtoO1iKEW+
AvcD7h/TOidFRhget1RwQH60uOvAFxrBOf0Uk9+liOl2UltKqevxPsW9Tz6JmmtUMqxOajDNEoED
MLgOzS5W8XIrBZXh4CtD2Kkm9LRAWiVHUSwbdTlWM2j/zaobE/nhUCh5a5nflHNKbAcxJV1RnsRw
dRbYA2ICGiLisDnwgr8gA75JPodHO3s0fouKgpeaQolaW3fkz5yXzPaLUW+nuThJW9SxC+1Tnfz9
lWwGLN6U5AfpYtkLzQhhEehGmWtbaaTl/0B1WXGGTY9ALe3LJarZUsurRBnffetiagJaMR1t5m67
cbm9Adh+JfXEaLy2Kp8OeERW0tRy3whNbgH3SmlgYOJKKqQ+8zYoSxHdGLAvnmxhNlgPtXrBh4b8
TnvbZWVlEdiBNHahoIDXk1qztrdXb0t8TipMOCNQR7FOjyHq8ekgUyCFFoSi42dKFKp7CkN6c/cw
cAoJu55Te/0j83c4vc1dimdQ7vIqWMDnmg8gg/+br2OY7+7z7eBZNtPqZ+j4kmGYewN0MaMacpiH
ow3tbhzNvllnCwgdLAWr2VPHtBePrlXJlHSZqlsw4BVAZ2mZloTle+8rdwutrFDQUIOzZ0SI7xTD
sgvg+BjIw9HqfPDvvxbD17kAMY3trv7f12w5NBzApzaWac9aGbm5aYVKeIsUSedEq5PA9sDqaNxF
+qv6CGVOhNX3zHvDZsYCsvn9zoa1eZs7hykstckXJynwo7xoMpiUq31xCjNA+7YM6OJBebjSEr4H
1HG1yLPHi1vTNqpFNRqlywx7l69yZ5PLqgpSGNvmU9BVOVlORXcqpJYExuGY8znzPxBJtThd1G53
hucDbDRgxvEuaMEQ/GrtV+LXXeN6fdHY685kFYfoyrR3hXxr5pE3m7RRY3FigXOavC22Zxj81GSf
tlCjZ02pBoxnXOhsjkuq5kCARLKDknkI7MRjv7Iwy9gbZrT4lp4X5hk0IBFGRihE+GDGJNLdH+XU
F3Yr/hVdAC2vUDpteMEQk1z7ETVYQ77fjV8oZe7TNseqD/MESvGPCL6gyjis1byGhYVp8kCNJPxV
33Xv2p3ydCDBC70Cr0bIlT1lzvscGjfoEQZJ0PTA1ucgj05wyW7891Ve7ppnS5nPTPlQlusVY7Uq
6S0kr54hudmD007GSMki4xZH0zvshGFU3zqVZiKrNC9HYNkG4ZE+7QUcGfvDaVq4gbkjltFZwu5n
9d2uQRBlBPn6y9k8OXPcM2JCK/7ejT/61ZzAhc9806IE9U4y7AAE8hRHYmEbBCC/GWZWhZlFplsW
OxZOl0fdJIN/zTtHx17l3QRi6K12zqfTyjfUZ8FHbdrhaPSg/PkTaqrszHkqTD237nBTo6xCIZV7
LeISJdwlOBPfhOZJ/QLZ5d5Zw6uPIQv0mjch4miQNIath0JuWHs6m50UQYys0Vxjx6Dsvcka9jL8
WvfQuGozlF4R8vkVn1jz6I8ph2Qin7srsUXOUCRNUlD0TbGNL4pdUv5n58Fs/459ktr6cpbREyE3
otdZ/LKfkbUlpuxN6d3pGnf1Ol6iIq292TrDkX/tUeZHd7GLN5afKcDBciYfryWD9FNXRtZQ+NjG
s4qNMt1LoM/VvGI/yR4/gnanbqkAt2jkKxp6AJCe0g2LOTSJd7QT75kpPMJjaAdlYnYALKsqRktf
Ae6xdBMJLJUME0s/psBTcNsrV0p6ozYHllS3gkw4LKGQiNolUrdzGwicoP91k099seevVcfpyIIC
R2c8kkD8XpOKwCiwFdwVwBdvtv6sm7APYQBhZ6xzM7s1+IRZOgper2ho4KrJENf/trjOURCcjSBD
HqsPYikGsndTd3GCxiblcjCabnVVatsxsSqEwk38bCe7i3lmGzZK+pdjNVsdn+Bc/RqZtNBCNxkI
qjqd6gB1Mz0UHrVdoBA1hqBKOogtLmjSmG5s3ctgQAPPL1AhNKb0CIPgOLSllqTTOZ7LQv1u6DSW
+nhSCPO6clgAdwrlpf3h1KAP7nG0OTKifb9yXDJ1YnGl0CCTC/kd+UQ4hA2LWTSwFAuKa5+EZjHV
21ERBv8Up1tq5ScElF3NQfqbMjV+LeSIkloTcrNvTpumZYp6q/fsu1KFmuwV3LXqf6UpQjpuCMur
yKSpkYmSyBbCLS/0ouVhFSRdSsLyySsBEUx8y809l3OAIi7jocY/iuyKQme5rZsLhGT0903AfyKh
mGwmK8R2324S7yEBDC4GrAHXMwquQP05LkyuQq3QtSI6VhiJd2WRb7EpIdvDoz6rYn5/A9jEQpP8
9fhWW57tFEd/nvnbdOxIoCLZMZyzPupI6BsTy8HQDLgC9azs3QhHRudhS+4IKAToLuhsdB2a297W
f6uDa5EI6Ke7NUFcq5tMQ0Jl84KiiNQj2fI9tycvdxl/9mcgw+khoeCoML1+xdm32DKfQQeGLLF/
P32KWHvXvXPk2wA6ICvv3Yy/Oj6pNO+71VppiGr+hnzRoqY4XMhbb+vQdqosUkjRLPYQljqDEuis
UJnM0H9IPCnO3nr7i45Ux7aZhyk3idGorUC2kwMmWTrUKvEFTT3amx8DzkKk/JzG/Lhwjb8cDjsa
WrLsOLzrUyiRLd2Dny14ujsZUvS/OOnezbiYaJKd3Z7/WCr/hOThUl5D14lczvzWjlurP7HYNXOw
gM5TzJ1ilwpXkSrSFMiWaXNXZ1v0xwJzGNlO9wM7lxakTH2pbSELHC4ICngsmUx8h44wv92dZhfs
9BjZf+G3InvvaCXkSa9mLxHEApOaSf68PlD5QEpxzMC2wcOF+hyOpgNtBGuZZ2r3C2GErbPBfuIZ
1YjfwNEnKM3yLq6At4MiORc8mZsq7hga+5Rqm8hck1RTJ/ilIRhwhR+EuEhlLNHqffo8GP82vnDJ
GfgjI7eDlofere3tHoOHWnmoATcXhFGt3D+M6uB4iQ3R0Nne2Rf3+w2Cu8Em5SE7YkTd+ArlqDBv
vu8iN6dRJpfAjsjASzhekRImps8G398k58MhSIcnTN+igxQ9VXxYLgep/6rn+xejimjUwLW+YUSg
Ewfal+u4FSFmd8XD492lXbf3wN2c2TruTK32Xv1WiJAnWEf3PlZbx1Uf6wwd1YYjtnxexlWZjmWQ
y0vWG4CRmGYrW3+wPzDCiyNOlCcKkXGQmoHaZUFMsMvky09NxKhU185JceJ2ABiIlK17fmZM6gfa
jsUyOESNjMaqkUEfCkgHEe+Lti+2mJZhAebxR9CHDIRp0sQ1H3l5IXzBXkcYqPg6Gj6YSCn4r+bM
a+/fvr1DgPX9kHf50RU0A5/TbApp2RkXFQU26L/uUhXTnfvxK3prokwDOegCDXtXc+UTBwcT8LeM
ijRc6qeEOpdgnqxGG7HZM0Muih50XM6RZ4b7tRh7trRjozD0xsI+k9WgFddkEeRNIFtAYglP15DZ
uxL0lmjDI9LqQm9TfqlGnbHxubkAHq6lzUkx9QuKZ+PLiaB1u4ek0PDg9Kv0nQUjmoa2k5T+oHnn
6o7rrZvCAXIPaEqA6AkuQL7aOw2mtxS+kAayD4DsSBbU4A3y3dvPDvUOQuwAdWqZTj+x4zl4L1Tg
zyMavE1mV1p+eQ6/1OOKTKbHlypJ9nfrJrhHqlyyG+z/P6ZqkGkctRNJrgJcy9skhI2QZsH3P9RY
D7Bvarz9ph59DDoJB8/7k2fXKVHpeTt8OXKCFPkFc+A9jsdVMJzcYzJkvmA59leLb/pkt1OkLmn7
0M+gkwHn4PmpSL8+gLxuQepk4SUe4v4gFJWQXST0aRRrdZm0COAyRwHVBpCAXqQZ7wk31mdaBli3
MERkf/vdjh4NQ7/3cN7u1m4yZn/vaEwIIpap8JSI9PmN4KKDT586qlAR2R5tLFiUaMRZGNMhrAo7
7ktOXFH/crlx4NPSrKI7w+3Q3W/t9DGawrpGdHaXgrE/IsGH76TgDPtmYOCSVireF63oCZfOfAYo
XlssUDCaYXXmc7eQPYCBcAtZcPrie13vQe9ohDvmTyqVZwcHNmDqZcIbBxtQyEj9TKxKM6CGGgBt
eSVsUtLDQxsZqddjqcjGARq8wdS2fhLoYpFkp2/Fv5X4AWVL+lkjn1W9qqRz0hiMCCYYJe6It+6W
eRT4Rr/zfpfvyNqQa/3F1gjEPIgOcZOvMeW4dXhd6/IkNeFrVRlURCjJ32WhiAhtCVrC61ZJGBF6
aYmNqZ6hMc0x818mQV4BJLkPRFQOL8gzIUPpiD7QQaCnb1dPft1/h9OH9DGD+tQ2iNUIjzccZ87w
KL1tamTUbuLAhHyLbjsS6ilV0xw8YpQVQf3b3v/HIhREhOw/6hYUa8AACRM4FyQ09JyftDVJ+rHW
48pATvl6GY3Xq2JhlR/pu+eSnIc1cqcLU6fMUgy37wUREwiNsANIHyCl/9c8juw+6khD15+m3FoQ
JdErY8Av+RZ1jqGujdMGqOw5gyKdGlx+iXxbx9lpHHOMh9agqBAUzolMGARqIWmODmTcqcgztV1Q
5f4oGjN6a2a+C4WOZgDDiATe13JpmmTXHWLW9UsvICT0Ub6H03GoqBsx4DPMuHdg5yjPJCfRpwyY
J2IEppeEvllZAg35RNF/ztNVylbl+bC114WDCtxPskr1/oCnYVZIvqzZ0lpk/3Il3eB47GAs3RJI
4uUGV5Ayo2DghY+1+Cay3HePGq1BXlmMv9Saz3z653eJdFo0/aehNEzlJl1QSqiiM3zoQKyMAB88
99iguh4/MRQvIXzcATb3lDmda8kpZ2L3/hXB/uKTfwGj7UKNAa+Tw8NZBwYFo5ceLXccl/3u5YOo
qPdbx7Y2EXHCFQJRSBd+UgZ0xnzCYyd80dA6Z5cpf5fJpIJUAKHwxpN8I5/RvEdcOi8kSHV9RZwR
wX5EvSSow8odOxB84kK7cXMOYwxc9tq/TJ2iQrWAQgx5uxc4pN5uhqf4aY3fyh4KMaFE/nnugROk
AimWkr6ipZFDgZ1/pq6A8PFLOUnib2zoSkLTUu363IcEBXMV0MQhBNEGF90Ue89gc2kBc2rNj9P3
lDEvKqg+G4inph5M7T3H5xApfe4tVmmE/3D970XR+xfKtq3F09sA8wtuUajSHBSF6rM1c+Nl/zKE
l9g82S9dEH+cyYXvY0jmzMogsXXZuwKzx2EM4Zc6RSWjiIQ3hiNXxAtwf/pv+SWcCwKui4dEGk9h
ZxKtZ8HBL/PK2kzNLF6PLQNqev3Q5ZBPhdGapwsVmsIXBioAAEUROpYHrFogt7AlfpzZBFzXWccu
eTAZVp1iO7XyMkaoTgBPjZlyGdGwnz6uA9PhHBirfAf/L6VMTaSBSAqQniR2JRg2KMHaJTqB4Imu
J4DhqgssbVfhLmMaRthV9bgt+rdH4qG/ZxKJWkLsUbNP6Fo3gHlbOQ7hsFsARpCkQIzaouWKCJlN
U/49lh0eC0BafCZMdcoXhj7ARAjmRRJHQCFfN23DeMN2QQkwA3fT3ZBLYVm/iO2IZus8UYPg8V6F
/I3mvG61WtBvFGbuo4HKSV7ZPOlTd++FS7U6KWq8v/phLdLBAEpoUEoxCC2F8qJ3yzs/yfGt9d9t
ZpEjCwPdrCbd/E2vNWCDUrOKB42zubTnXjGRf/ns+44lohpmSAOI94YD47ozmusrPT5b0QhzK1zO
wFTBR65I7WKx+ddsMpgIrUH/KEVGwDNCFXz0cl3+mGyUjGUOx9F1WeqiDtT0MGVzk4BmRWf6WB14
w5HUqx7bURYQc1NUHzkrPOjLMXhQsAPiygdIJZVg2Us92U8g3hBpIR01kNkWc8CQgUaDnFjWlXqW
Y5FjgQa0OfMAAT6T2jIFhBmsY2qDgvv7+U9QlmGkQhbaCWo6FDC3H/fcEA0Axjck6CYx1E+jrO0O
KPe8Q8JhpDn7LFftpuB+Up531whbpWFmsk+vGEmg0wUFMY6z1GvH1YOLFVtqWDjzkYZTD6ciH+Kh
JzI3tzZL66JiamXz9flaHevHrJtq4WCgwYNkOj57vrR6dH8AJh+p37CaJU2KWmA/0D6oCnhkKczO
87asLuVU6TIp0xJRZqmHlRPqJ7lCvkHI1mJuhaoYSZDq3185ZAJzPzjcA/3v/c6mXklK4eysjtF9
7zIqFcdn9x8byBYjMGoOf7bZ6Ia0QwnQpdmLwLcXbCy0XrDzyRyAQ9+gAuxUYntJyvlKLcxD/rqa
+7PKkwQNjNlmQHrPEBy2ZLzklyYl0DA5C3c2izttTJazt6KrB4g9N3oxwC4q9GobgaCwdTUFLTM5
o83Oio4CHf9tl5CQj+SVyIL5Vh3TnVAMdjBnQ+1mJmbjFYpCm6esvwQQkXpH1JabmraC5D+aCYcP
s2EYxCImnB/WVLQ64fDvF1VBrpICBz6cAxHmwjDngZs0/h+AfRmQeuW1o/JKYS7dVCW0estSr3GY
m8IpGUNC8KnVIxZe07fK/TlEHJv8c1U2jGa0B4PsR3sf2lhpd9z4QB9r/GIvIARUU0syYFxtyX6q
tQ7JcMwbvMEjIm8ySIw4LfIHsU7ey9+bCh+gKnvlfVUHGgvUh/E5oJ3k07qos/5u3AAoSXsg9s2e
gRBy/j5/S5WpQW9FKcVMfUYj20ewcFndeFkDE0stcZvkJR1MgZJaFOz6u/HOk4tNEI5WlXCm8VyQ
ZS8CnfIC2J4TK5RZtspYSTiNItvIOpyPPhTIgtW+4JXjEBRWXxsrPgOEXeEmhVdhZnhIqetZ44ut
US1des+4lntkmp2Q7vLVI6mBL02D9V2k9XiA9/w5lJyanaNypf21Abu5JkV3BYeDyHNdLMI0HEx3
s4SEMvHgtHYBzfIeNqjO5Gl5rbv3SHofHd1vRTZlDA0mqHV/KDxSnzuVh+8xm534+CGtrLNz1luf
HYShRplg3zVo5MHsitN25UDmHmDctZHTnq/8elq9FYfv0Cao0nejcFkVHW4qoVMAX2ZPV/3MlVyo
ookBRMuKO5915qvLp2ycMgxzaGWok1eN+oduzRMXxEODLctFVrSTrwLXHZ2zP+g1QkGq2pGwE9Db
6WsvQFyzZUZgh1cVbThVRNyET96aGbgbGi7ybFsIY+7FqYDpHZbFbc5dE/o0y4fCtjxqgISqPtrw
nuFD9Fbe//Q11w4d40LoxQsDelSlijzUGk+m6hh7DzK9+wZuM+yZUlUpWZnpzGMYqbWXjJX0wSRx
AdYv6J/19s3bLgFXBaVMcV1DGA5hUmWulEuejRPgspXuGhOPOF/Y6pOQF10f1s+NLGhzJb6ENPv7
/aitP5Mo56wluQqW7FD4wcf3b4NzRkJ+DxEeLBrIPVEYuyTtK7lIMqd9Bna0sFdCvx3T66+H8bpT
3f83JkyqpU1DZ96cPx3PIZDMkNa2F6hC9c1S+mG07OURm2Vn+Wx1SxuTHLi4DnzVAhSfdis4CiBA
zZi8WBfCGpYZt/MlRicKvn2r13EdctQi7OSXI4yypOrKYFUWlu4wFOYLEn9osjNkaZRYJxjOs1Jl
tk8N2OA9VrQ9pXAFgfYBLVfTUNOF/hjDFE2LyzJAsdxDBSQGJIR0pdpPgGaTdmp/hnADdXjrlUgq
4Eeevp8hNZ8QHhzhg2j+pKK4WXxddIapqQalepwx7RjcfQNWlNT56wlQDgsnOgWDMGJVV1DsyOEM
JiKLEArzI+oCvoKiDzVDDAgnVkLwuF+oEJNd1rhjdr2GzkoYb9S+pqqRI44nbV1l3OPa0jsEQYrv
arl94evNmok8J7H5ZxOyi+PB9UAsqdmggD5mHEjCDh8MtSJYFx5iuuXLGixvXUk+a9ExI4UgmBdL
CnMCVeTY62Wm5WNcLEEDwtT+BW3VCdVaOAKTBoZuu1/fD+U0zFRg6/7Nd8VQ2lZU7xITkQKmoMA6
xyeoQiJ8JNO/s4tyxu8dWKEBYdtRhwWp2kdnZlTIIARjnWkP/Cc0iptNY/cjhTg+aX06gDEooObA
YdZ+1Nfoq3uOWvRFkaPQ6qbtNq/824zqkVwB+gQYvttm+X+TuWyaVtGCy3m3P+zUGplvQi8RiM7m
Vs+MNZejeGO97/ft9WaiVgSJCOiw0gYXSerm76Q1uoxBM5LGYvCbO3bVbkhm5rRQB9HjMRkoulGO
1dGf0YvwUdZAl3ZbRz4LZ3eIqqRVe6R7nobRFQt7pUzXmwhUzLfjcMMHnqHURcd4upDAktscftW3
EFjzWltIfQMtr0JhDQcCs3rQcBA6H57mwnCgbW82jwC62gRm6IIA9FIFx80ggFPmirJ+fyE4uppp
St7vNvdqcxqP5fFynFG1Cjk63roI1nJpeArJkPytpK02HtpPsJRIaPZIUwe5KO9RnIC6Kf3wG+U3
Tr7nq0i31ibv7jpvKiXy52MA+ZO15GCFxT3lcmpOtySGwRRQ/vDyqm8gXUhEZgdkvCTrtgl4QIjw
jmfKNIMXYMhLpNrFSHmVEZPs10Zy+kdqvtgxyhx/eP6r00yMfsgVXDoaOdcC2aaIo0Ee/pLfsp9R
qUSjRmPnsKM0ggFZ86FIkX0rCd0SfzA/JWqBSVem1VVW1hC62E3XIZB8kC5Ry1IWDgHh9j/gFmHd
vzBQb85bRyoq5TVWv2rt1pz45rt0OK2+z2OIg2eZilKDfSu8//ons8RjFU1fztcEZ3A8P3SSAmnf
WdxqYrbD1HoiIBYX3+izwCrMfRG1ipsPcjyIHTlkGboKibyHuaOSQVddak4Idsl3yjW4LHWJpm9y
0KPNJq5XrNVf9JY+Xzbb8nQtWMCgXaXE/eqfowzDWVE/Tqg7x/qRaPekPcV5jzz45y6kJE6De++w
FIWitUB4hO9CWeOy61rFHymjRmeeFRWwNu0H9puAO+vnqi+wBkw9pInizn4X+kxvnTQlgp/mSbkR
6ZItVdxaFHjDeYWoTJDrlzq5zEfUEgZEw7T0BUgFs1d+US85XyWVk3XYDwbUDM6kRmFl9tCKGWhN
cLTQKLQ6Bs2rxTxoRgyulzqLE5He2RDVLa+FmuVdrAxyCZRt3YZpjkmd/SHMSjjjj85yGIZjGv75
yyC8/0xwiKrcPvndunz65bdxJ4a+fE3TIeFcUDvJEGL6MKEL2RnyWuSr0INMvDULnLNb02+Mp3tg
nC8ffkZslXoXE7Ab3JWlYSS+jCdV2K+ph4/M0iHH/wmpj2W0RzVuuJNXtRKe++IhSzs++21xa54W
cLoLp9BM/WFlFPWwyEKNDMw7UMj1/jTyz38bGfbs5r1CXfvqjI6HZF91ahDINOFYWxNzDx+odoQ2
Jq9RmgCRlttr5F1pQozgNboRjpu3UX/navvgsdrsk59BfiRhiDwe1ahuA4xR4HVhT1hmfSILyYED
eqBy7XwdtSbZuV3wyBMK/xXNQ9kHh+MMcfqiwUn19g69AesFJD1rM2jdrrREXdWse2/tWqIlcnm2
zYFpsNS5N7tBG0e5to31Ae8Tma9qZmkM+cVYpsDrb5WVPWHUZ0R4NABOSX5XuGBF0GO4Sndu3ffz
jXYueMg+yijCthJKlofLaktPR9jhTsbC72F7B2YyqowDr6f5vSeyVR4b9RRkcUs4fMJzAPUbwTO5
viepHivvRh8cYVAWmJcRGVsLSMfvI716oRx2YD0J8Hm9HPZspOyKszYB7+3UDVAKD4OMvgHVQAj+
MRylyglqntxHvhsLVfyV7OIa8YLAcavbA8BZnWiCRn7rlxccE4hFWWtRQC9EV0wE5//bZfEnzQM9
hBeRy52kT0FklEUY1tYolBE4/TnR7hh078vm1Y3IdW5+HsBy4x3osfZAD4C4RWwyYc8V82qjKBBu
OlVuRu6g0s35FNQFNiXjcMqlxqZVHgKJp7otGi9tEWn9la+1U/NiVcMzGSC1Oe2BbUS6BWUAa25k
o+ubxgobx4WY7zAi53wyRGY6+yH5h0ClSrHcjrDjCbD24Nczt0oh/wun8zRqiMhrz9L5JmvtSKAr
Bz/BwUslFqudPJ2LWP3qoBujv0TiLKTloQRZV97bT+bQxNmr4/DLs7gLx82WIkdzZlVakwjf6f35
vgzrR92hVrXcif602FYiC6cqldvBC5bTGo4d+pKcGZxJ/SRG1YVNele8zMVLj+H1Pjy9oJpVZ80i
0qnEPmzGF7i9vAvrcjrRK5Nvxpt9Vc2Mc2Mu6wPFHyWhZLch6RRbkWolpUXh9754QZMuKrGpYBfe
e1huOzD62QokRI+lyqOV9zKZuQqblwlxB0/U1zaE42eUSfrDn+meRX0cHgHHw6zHo+y6/0Peyd5Q
wTPgrwic6IgnyC3h42X0s0z6V2qSnvd3pWkdcEhBOQIBgpF9XcD7cXDfmm+F4UqcXVcd9Jw0dzMy
iKBCjID0RU3YtiAmIM+dzN13vSjSUI5sNWKqtKOEHrnd3B7EPIFCbTyI7eWmIzR+d0OqJq3YmMJL
tIP+ieRtAVQpyQCVgkcr4t/MypX1rtGVx9p7cICjTGWk5Ie+G1ihaeS7pr7kNAMdR+Hd0aMxpczT
nt6vl3zJI+TcjDukl+E68O6O065rjfayr47VJYQ891AzWr15XaiJDgvIAmAwNiBwIzcYzgwVc8Nc
ZhAtTo7ATuEkrsWAp1pSEe0IhcKz7ABwyLqRBzsfxRKumdnKgYeoVEIWwg2S0lWS9mDnCemisG4O
EtdCmAt7ztK7nvK/sFvXbkeSi/RnSMCVdAaF+60ppISV1S91xIa7PGE3E8PmATqUt/5jXCvNoxcO
3yRkm58+jS5RMKYXuiyAdHqWVupEEVGybj3IPL8qriBIqbkxF002eFWQz8LHeSqIzwbhKvY0o7Ak
TA/W12AfmFEHiAOnG/8AxJLed1oYMKoMIOVxIw2svp5pesQROLNFXG3oAiKF+iW8LHkUMVqagDcb
4TM2vsbvgT2fxnIAQS1c+q7hRW0wYoTDz4rTyqanxAxJw84jrSFwRZB2+sgIyF0arWDNix1Gnoho
91DTYbxu8BpywMATCpEGt+AEZ5CAEtxtHj2oHG8l0NbFlfHwAg6s2q3lmcQNs1UrihrWMaNxPedL
3A8qd7Fpxiyh18JZ3QI82kFZ0/V4W6GeGfsdmkZyWTkV5EW7+FPU/oAn4gDSj9jRFYJUMJaUAfWa
jh/6upAGb4OM8jAfmH8eCfQndvZ5CjRchQG16DGd5XOnQR2M6pvkDXQSMFyW6iHzJ24LAYkvFOzR
TgpXIcNWouVGIgJMMtaBwnT4KcSCl4NCdRuPiwjSygpBWIb1FmTlkLVZV2GCWaR3GLJ2JXZaKYoZ
ow1gCLDLhWubAA3132e/Kg4eKVqf1uboDMhdsnOA1VlpfSPfbf4IHh7WP4OuX2xmkjqHNYvx08x1
eFYrlVfbFRnRPAFq7riqfKx3lD6BsARVlpUcxPYcksyZ+LyXTNtDQgYtwPdP9433L4YeyKFrNnwK
JuzCy08HstbRTl1qYTr6VezT+iiFFaxPtDb2BzBMOifkdpmJVttbEad+DiSk65SB3TYK8z2+GeEI
ZokKNHjbwMXA+/r0kITCdk4ZM6eDnQ+M0L1sKVIMXdq03DgCrthyXgMCnnq0Tr3D6tJmSfKCnIwR
gH2OPhbyuK/AgAKoJ4uaymUchGU7Rk0Fc6lHGVbpcMHsra/guKmf/yWPIksl3H798WeTsQJjHuOX
mwzWlLz1zuO5k3an3yE0dOyiXOZWZObdpnINWcPzaE5sX2iX8VpEcb4JLyMBwm07EMGHiXMmBsza
WRw9HkPY6aG4hL6F98rmrKoDEZOfSrcnfPGTdUBFJHkJy9kNmcJuvCKHJ5+O+usoPvSwqAPyvM5v
wJmduvhd4sA7WGLGIqAlkUmfvHDBzIMs45sOZovY7EoVci1DAX/qdqfzc8kJh7MZQVBSB5zSbekD
vFI8d3DLWHW4vd0FWmVnkETSDFd2UKk7Xk2aeJA0FiQKPSpAY/6kQEjE38xkvL9ikVRKWYxh+N/B
x/pRA38k2eFIkHW3+TRpnNVWBuHjEKqkT8x7jHYuVbSCrz3HeA/9uyL6riEX8iQfn8QbW49b/dn+
6BM3GyVddt0Fypt9GltvHCxHblQ429d9/FiBhF+cRXF461UXeLfuBX5icgG25SFvC7jHMaq0xWxr
PBF1RNEcHggS719dWQkrw7HZgMXsgSpQDBp0VMSPJON6eBtaIq9f7j4FKSxAP/N3uZ3XATDStrvK
gL/pcD7iUDi50wWiILgZ1rIyNvSlManHh/mpCmMPAFaoUgBpCiZ7lNKy5jmA8I14R+ylr8CsiG1H
a7qHfdDeNm58qPUHODe09U2FPVxmPNpBZQoKGpac5UuL7fjWYAnEt5c8dc6cXK2vOHTEyCQCs/Py
4G3oMghEvgb+fg+n4QMwrJ1el6NS/Lf4s+vyswaQQes8HZzYmNbRYyHtM3m2npwSoa+8zJWdB246
6jHx1Yq6rTm9bTtfyp/6iU8VI844rCCD5j89/iOIQen73QM5uawSiwZwF7974Ae/rJXjxiXQCeqw
XCSxnb+8SGmmnNM5IY5aVVY4Zn8/8s7XpakJfaWZ5JIU/sqoV03mQbKryGn9ZNNCVGeyOKT2UO0j
x6RDQAXvPRWUYhO7wFzzQekdRXJJAnvlvEeQTDUCYjatqx00hHreNVs4zPdGuChxxqa8s14M/gQz
rrBmbr5AQLdAXyKXj98y5aHYS1wVTos+EQD2vARq0TwMAYh2mAG/ht0llAJv824KQFTHceTbaEVY
MBvjEp+yM1cQ6HVBDa1H63VLAkRHHl27i7mn+uUqN3TGwed0K6YK0kRw+wJJfQ3FgIwU69QuE8Wg
eK+7NwfwZ0oqtRbTqqaw8Eret2eYJWIDvI54iHIhkSTcXanqlLJopB/9Nztl7oXq5MvEiWBpDdA6
wIAXjrie9dWoQC0pFAaUb0UMb21G2YTuxnNH446DHIoYHC2X7KiJm8J3bRsuDjNrBEiEb1c3JL6G
3rwyUseK8Sb1GSMmc+88U+BZiBY/fP5bOMbfZFAnriUyi/nL7CQNN8iC7bMskXheGPrDVrLfxgRD
3BSub1UwUBe8QlXqYCNeaG6TS0T35EpWEHctluRF+hhS1P0UVmTMhBqbOWwO5a3k8bzW842LiTxF
TBoKDJHIvkkAi2ULhjhqLiYJ1Pe9TAMkvGTpK4CEwCs4kL/hLvVMuAh5t1z5WkmxbSPvSOtZEMr8
k/qrysIfrRHLdCPt5Rt4rknS9+FteQec6JeOdhOgbbRWXgOZp9x+k3GZFudG568UIHtwRhf+aYxB
NjWQyDI/T2+Z3X6TPvwCbgwdqFdbnd9bq4tMIWwYzpjYbdbJ7jEbsIGr23roLvHG0L5hLzDzFTp1
NN1ClV6PTFbq1hkhYqw7/KQia+R0P0ByAQRrAEMlTYsx0I4CGPRHIEJZW1frVbs5YkPScjgWSQJx
mKDUDSU71CeIBa6m1e2VmjYOdoddGus9yxvt3Y/OE1VuLvtabin917BWp/4/cF47mCU0oBcr4RHC
Siin6D1hYmyWoEi+iyFmJBX4XtcJgjovyq6eWOff1+3qvlV9HTSTee7zHE58TvoKx5YUfKrtzdMN
sydWrgNaZrknV0T+ibj9LGK/HU8Wh2CfeDlR4dbw/bU9oy4FITUSA32ePUBUV0GZ+dSMQKr0rzy/
OryEkmVbzgV5qJhZFa/pkCWVs1qpLj/5fLjNk74kGMW8OClPgmaSgNie1DrSItLN2+pb6oeCiWir
ebaa82XsgsiVaCtxyw+nXoTBScoaVwdJuvvMn3XP3AMrZWioToeBcqgA1gvgUsvac6UXy9P9yXz8
AJKbvDhn6eYI391vK16H06N5NBMC/lj00sjpfLEcP9tr12O4WswrLcWgAeuX22INwo+dUQL44fYR
v2MPBgWzW7xOsGAtb6Emi58iprbJoVLPNIue3d0kdS4tHOjlTJ6Lk5VN2yTWhvEQI6hgR9vseVml
Irb1elKzps5rJKrz7c47eLCTdns73AdrwqssRzkhwP4knr1ewPdp1RhLB1o6KpJEPyTQgvdPrhAD
swRWZigqzz+QvmOFy1CfYEEif9B1f5UR4aui5b5uKMy4e1qREJrVlmtQKRCCgw3zQ3984eY1PtJL
y7Bj6zB08zD/R0OeXBToGO2seHoH51Wwr8sWHhfM+g03VpPGqD4oLd5PBIuW2VNFEiNWaBPWXp9k
G6Oa7MPJtsWbJ7jH8kplrrxPukkfy/Wl6OIvbhmtOpfLisU+m0Y7pxZg85VYHnVs2+7D2PFO1D7O
7OvmPKthJKfuAmaWhH/26PFykjVIGE3CRCyJ8QauM+Rtqg24y5vBHvKGOvKMdXtktyn8/UdWsPFn
4DrMVVhbLChaIjAToLJXKnquLBtIN4ISOUEPbwgcnqcLHymwO2aDDTkJeFkf+0YJGGYeEB6dwH2s
Y+F61QJKKQx3hfNmXvC07JEX/Sph9mg7IC0lO/KFZEzmIdmyXjDJhTd7uCDHYEABuLbn/79hCCoX
cQFQ4rCg/osqf4qPvUs4JSbqBULqkljadjl9/EpL/VWeH9k6O3STHu4FQWDvPx/w2mU09Q5NWZ28
nSuDIbB1gUJjbppDDXWa17sTZFBZIz4L71KNVw/Lseqx+BbaiC8rPpR+c+3wtByCRpxdBPTkYB2v
WcueLySmytKPialzQ15qB+9nKxFhiAs+IQP0BkcE5yGm27X5WyGa76Ia5ZuYpRtTtJVApvOpQcmd
RoiYjtlEnmZmlJpjhKdjZmBxhTQwI8k9diul7NqgUehE0IHzIMHEH1BfOdzmsxpMNczKpqLrX3w7
29m1TWUi17ligXVv8RcFM80h9nd3aNvJ1E/I/a81wnFRFcajg+DAOvOe3IFZN5I7bFZzNWk6YgdH
4AU325sM1bIj6Agnf0dhsg0DZmTeG+KcwD5iWsrZaUhUQB4C7V2MJFm8i7C5O02/U4dTCh/Obb+Q
4s/d2nummpNx3sMaBEhHNACjjgBzND9VLy9EKtfBSZxfgI1m+X6ZaDGzJIR8OMvnCK3AerNNPbOd
d1X6LvsF5gmxD7l1A7lmcaMDYgOS8d19xzEptiVGycMBZI/InJTQ9RTkss5iJ2NrZLHSFdYeeAAd
FDaIE4X11Ryaw8GNYAdKcaobQFEeYITtVaLJq0fDiUmf0h4eTnvKljPnWWpamVUG4msUHPthEAwO
loiZ31/VTgubl/nKAmWC9ajY+yqaP5oHObvx0u3qiYYzriU1YsDPVJJs7VBVK52NpxblSJiSXr9U
qLOW0tKgv5QvhiX9nhP7KIsBQKSL4xXcqSnuq/kx701jIVD1DUsc73AFf6W3V3hYHy8a0XK25i2w
DY6lBPeUWbfNK6l+DJRkkHUv5piORnKcpv4itXvAGgvRWOumdzK3mVL9/dex0VO1vfEuogNt+vOO
FwPNKOjuVmDJn6P9gqc7frtHPGcJl0TMi7QAZOfYm3VjshJMOAG8RrYfYS2eqq6GV3I15c/uqH0Y
GlIK730+A88rreNWvOUTNlDn/0TVRkUn5Ip96Fx3oFcJiU2/eCK+m4LkNfb4aum6Wv7FdXSOCBO8
WfhgWwRXAqhAPV0IiRTgi2MwM+wYDohlr2odc63KWZU5id2VOGXcLapGMS0suw4tfVwlRdXpiGEN
usTavrs3cNbIj/Xq9buua2OaWH4gdMGUiLK00k7wKO2qfQMPz2QNJLYHgfxwMcsFv2bwWc57fygG
vxjeuRCfOmF+TER2hkgUCEH8C9m+ix+Tbg20m8E3B35PnioBc6hA1FZItOvcPTRaISQRKSfm71co
BdzfjFVJxc6FomvtNLmVaiIgKiWNt+Eh4SIQtzGZf8h0KGqizzqJlzlfUtJ7DirBSyZ5NX0286Oe
OmQaq/KCWk8Lr1UPlAhkT0p9KoFgG96rsGc5UAhn76H4SgNcnYoX2o7QWnnZn1us3F0HCQD1dOve
2WRqFGmya4KTqcfipcXrc2BBvtieYwKgZMOKaBXYhpZByVcQobhJa0Iv3OKbD2TBSyQ+o2EF645+
ubnVNuYxP3uD9FdX57xUGI4ShxW2PvttySyYtdCwOdQsGjUpcnq3nnGh6VuP3b2chOt5XaW8pNZU
quxacPM6K4uj3PgEvUG6X+RIKrx6wEsJFQTmEgHDU/tZ+9/0kjnKAZx1O9T/6YinLGrb1Apo80Om
vpUHvCgW39k/ThkH9UKrcBCG99OjF1GDqHKnsOyl4OHz6dEN6b/5dJa043hftXMJSe/1zufZNDyB
qeohaTCoYBiCEHS7W86SxK1TfFlM719AKqLuStQqwEApgY6F6r0zJvntNX/KJ0WiD3OupIgFmUZX
xPAF6Lnb66+GOPxxAToHXAX4kzEi/BceM/7WBKDGYgVgMLUTeGqrieZm34dwPyx8fJGQ+oE+8wkH
2Y1pgkOuZNl469voPtDjFGH4QPVuDCdKeicfsw2VcoRNgHAjvbViWiJqcL173JU8zjZ+drOywwrL
VOAEqUIpHFM7KeETfVJA8QD0zqCCEj0P+XVByTdS0QQFKUyvePG1/MutFStJu6oh0Wo0rOIw8HQP
nJogZA95xTqqAFE6J3OP05F8VVC6B47JH5o2g2fdKanRVF+IZXU6oytjdCPZEOS9wDQB2YjiBd6S
RAwW42Ac7H8WmCTgywAEiQHGQMnZqjNFoYMLY9XYqj7HHuz2Vc80LgZADlyzBM0z5lrKUI/oL1bq
7llYHzUaEU5uj0g7luL4Zj//WA+T3/DiuSygIb28XHD1bL1UtiXctRqLGbaRqVO3d4yKFaZEAZhH
GUEM+/jk2Cw8OcPZHttMhwskWptLaMQIFmXwdWsCUGE4w6UVSCFpP4bblWzK2eRO05eH4oxCtimQ
l5clynU9LIfc65OKYJj2Y4fNS4PNwPpmQ5eNuR9NyuLTm5I67PobMvsjbOvOLCzZiXrEUTMinYKH
QUjA7LJuq2stU77msP+TmDRcu8Wosm591Ysmr1DKqJQ9Hn/e3vptvtBvA5c3ES/eBYHoVKTFRX4a
s71MakPQvEUjW4szoKFFMEvZ/csB7x5Ty5OhYFI07PkTLTU9GB4L/HCy0JACXUyj8p8ibwCUNEQq
9DBYoZFp/DD/UViITcfRoGn+xsXCGzn3vCHoSRJ7rTCRrRW/x8cC73BnOlwNmEf0P5EwwcbZ2k2w
Ugkk/XdAzJyd1r13OeF8gCdV6ZO0x1KipgSja2Zbtt+7geaFEydRgJOcvrxdP2IhQMpbvlviGjl+
REvOV0MzoPEdrv44eBApAVVUWmMamAOyKd/HRChf1bMayFtgfcgzuss3kktFDbqR41VbK4C9TFFv
xroeN9wWNWxl5vSgm4Yn0tXhCzE/zltHPqpECivHdHhU956RQfeaZG/tDOcQI4lPPAFlQhWZxnRu
jHBvJLTt+Ygko/cFhu9cLpyuF48ie2k7ZtgTyaP0Nz0oi0wEAvUe1A1xeXazvDgarGPu2duPt5ud
79DswDcz8oE0EbIDNnaRa94KBNGCTrGV5PVc9Iq+Ub1A+RC2jEld2RzsWnQAhD0jkW4jfsICierh
Eq851lO5EnMcTsQV4sDFqdYGooeMMsFZgqzSEoLSrd/2ZUvAmSkbZ200aTIVEg23ft7Zy43Yrcnc
1QxRFL5NdITBEJwxjW2+NFLGDkRvAHrNzKp2+QswBw4NTX5xp7guk+ZbFo164XMyo796+bRyaTyW
LG00hLM7EJKRYk9h3WairfIQfIpEPo1Cx1hlDEyJBxiKY5lJOpHWWhODsY4UN4cXiUuqCqdbvnRf
Aoq4RmU2KLKo+2+qokO6xij1rQ4xldUGPLY+C9O0KT0OYyHXkJmqV4vomq1ZUAZG025wiZ02irpQ
WqiT3nagM6geoE2Cv44HgDk8fFYm6MSRP/4S3NY3V3rM1DJXG4/Vj/1Ixgv4jwXsSGO14YsKLm5u
i7VZbmfN9/rwqO9QPuxgNlx4Rz7aiXo/h7UJ4IAKkYNQwYaBE3NFw6KRtr4nWd3es+GFZLGMq7Z1
dhNX7AAhSMlqg8swKNH3s5MOgh12muNqLUT5L792oy9mETTMCsNHavSZVVLcItx2yYqmlJfc7ABW
WbdtQNKozVwhDThkQJYWPbajbEApLQvkOP2vjr5o7hFspfEtyaz8rk+VEsULDbiBUZ7wgqI2BjTE
eesq2mgVa18CRvBick72UL5BhptnePndo2h0ManxRw6AUX4gAVx+505KNQ8R/D1LYQFNZr5hWdMU
gEGTlieG4jjnyoBF3mWFjj66QdRzfwRn3zu/Ul7eVLQhX/xG+3Gr9mAardcE5G/kDPl9oOFNL7BN
LdwKEk2sAfnNGJHqIA8yp96kz8XFc+UD5nKep4i3Z08oyqFo63QXC5wkEfTlgUJEERgiUeMVyH7P
/yo/gFBPYg/HkowItJWPODGJUshbLwvkknt/nk6ziu5SaXTGetJrHOsxYtwyjd5biQoZdNuwAOKh
Y6KXGRovKV+vZ1bZQh6Tq/8iWl3tUu+NkWmHbzT2q32aJOX98pgC3V5z9BxCmjREv1S25IE6E15U
DdTtygLlM50yTeoJBrp/lrROVkh5O5sCb4eja+e/V5tXwcWiAwn5cHKdPaTn/dzPYS/df9i/ADXw
LU12K4Bk5vC6hHDI35NI47Dte+DXxN8Wksw+aaPcaHOBJ5tKfKhv7xp7zmtzraUng52R879zUj/z
DtyVgLI8EsTVYDAaALLTrIJBG5RVfC8ZXi7Sp/Xf32p5YlnZ3grnBomSwI3wSQ2gUtVM6Qhrl6yM
aHghNoNjQFcz6G6o1I+RWCqjt6Xp1hDAj4Uvu1AHa/8tXDec2dZhpitpQsMYmArV4xWKkQ8INZuG
XY9kqF5zl6nmqsZpeB8DLfoPLrqWZlpbcpmh+7kdobFjR1WRqreVOquPB5WOyMVzfa/zm1MXuj0e
9i8mXiltDHP3LEOjIvK72PUs2k4eAZS+TZDgFRxOaFXO9Vq+oxOT+qNr2Ke2uQQ9432NS9WF7Pn0
1LtmIqNVChoWMzPQtG8cFjGGDaJXgt1oxWeMqPKF89iWhO+Q1oaknZ5fVYRiZINZ2ksTbOBsfJmh
ufNGxBYSiNmacduCnpzx6/2leubB/1Z5vONhG4GpllqEgx4PaZY3TPd5psQROfb0cyFxx8AUH1wr
lN56I9j/qzYiHrvNoRMrkCtBKhB4pxGsdS4/Z4tPMg2+xFUIIxSXZodD+HxRGU5OWuxya8pNy/G0
geGsXxk7pnWVEnxnDxRt4WGrkI2bf1ccDDW0RQkAJW1Sp4U3yh6Ki1zUKqzlgQY2jobT4KJDvy48
32zcu6S/8NvLV5fXp+8UGWKE7gzpeWo6CyAH8hYXdy3PFtEwv2GOVQhYxwAiso+3kxwReiYpCgjI
NLl0F2CFKmGvoaK2uGFod/HLm1Vv3cT7Pp57F39mRUOxzdKSwoF9COgFdpWzKi26dWQL4wf/hk9t
eEaVrYWBbthO6AoRWqQIUmrBcNPxG8LDILkY6dQKu4p6kITDXV+Ug0QEzXY8totdh0WZnm4ocw1X
YORDHMK8up0rStTgj5gaLAtzh2LZuYmhnwXhJau7TpbcHBQUMncxPgQoXiEtTLN6P2r8uET0kTHc
fRII1XkfC1xzAgo5X8Z/CU41MGaXo567i1LzAxlE9v6OuhyN95+RPjHztUXPkDe5oFL3psLGiWfM
8zVpBDzak2B4uk7u2lGSBpbVXS+L4favlqCP+K+jDIbT+tXzMO4JKIFuH51aq8y9srwubZYAeOSa
nASBrNQDyc5kXCcVwAwpkY3rOPIekIWwA0rPvIDhkCFb7CjbCTz9TO7iBwWRdYYatHWfY98EhPez
RBiNL9u/lcJtW4s2RLwTAjywwF8k6JRL+qa8g8K8Din22twfVHitboGQRiSEff1oFzljg/rZUuT+
tpwbz8CHr3jnftAGy9Uabzi0YfBjsJo/fkf/k8N4DI0M4A6rhJodJTa1VrUcRp+fPaW+Sg1s32kl
G9mG+KZ9EgXEz6H1vrB7Db4tLU0mCgM+8gV5XDSHKHFgAzUcAnbnPwWLEnfV0MCqZKTsaE+vWn/n
WFTJvgGQ40BrwDK58s2QvHbyPj4txG/LrpU/ySnnTsobpQissGr7E3T5+8yyOgw6ylvRtL4ldpiw
nBcRDtRzcSciY/aGbV2Tt0Hmf8OYKJRQhm8YH3N/mtLDSKkJPwsVHYhz10kSVl8kwKFpnKgaCw+2
Hffm5/xJV77XExP2zEkp0ChC3ILPNuLeD86XbrIf0YAMaL+SxflrOQTzGskZpA2B2Sm+QVnvA4Vq
zQfYQdcKOJEsaqW0/wX1FX0uCSKzyPgHR40xXqu6twQCEUiSd99IymBCU+eB83H6Q3CBmswqFCvL
A3JHAdD9qNpLzTVqIpG105gtz/Ch0dw6ixp1loq62oMC36oXOUcU2OOr12abdHq45+9B0DIf8BSH
yjvQbbyLyrCKeUQKweD4lVjNtYj/DswuZkv+6J6/tcC+N+BWNWCQlxmZgp2J3uj0kPK2wwHQXHQs
q/2dohbnK5Vdb4KUaCibiGFekBateJXGUbngqiPqTeqH+CWoq/+2MkzdvxqY2jf/nTB/059d/0hG
JhoZwrlu/2at065LcrY6HPLemV9Gsfq+xlc1MujaxgFtdFV44GHkGvp+tHs2dBYiWIk9Le2NGIF/
Ut6UPsg3Ydz5TXtq7amEW8qcNTjVLy8CqFRzbGzdPU2JTDzFTbkdheQ37kil077CQIoI8Vk3pyRr
3V40NTDoFFwJif57m82WQS6rhpfrHvq1VJz343wMnnmJPKKbHxs+lWS0G+st0wTm+u/GC44GZfjz
hdt7LF0zKLpnDgS6SdtRSRP6u7qid8QVnUM/7HNrKpwXATRQJKRMMRX2q8YY0cP5k7qe/aBMzWLL
PVjgTCXuBRHOaRWK2Lpapdx1t1dWiQc3wLXYJ6YU1WUH0XqDgQXXldl5Si4wR84rfGe+s9HZhQ3c
XEdfmDuz6rSgn/4xcQFoLHPB7xT5aOTVXboyHoiKqkr/VpD/ZrMXcFjB/Me/9eLtN+maVsy+XFTY
pe6Wnqno9CmrdXpGFhK+5G7sBEoSBUA6b0DyTTiMDGWOhhV8rki9gByADFYyX1X4iz+XtXt3+Eb9
AGplTO3LFa58kbmUP5Owr6p8fXfKhBABxqouUgJ3Ub7J75tHC9XBflp1DkwbVg4omhFQwtEy7/+e
uw3r6e3GvWqfHqfg5bYHtstMc8uAGVIairHYVvRw/Cf3KD20yB7b7LkJoI9JzquFKn14xAAqPjOq
QzsVmMApetnpWcvCC2NqBnBvLgpa2RvG9RTo04eKP86sXmQPwqwa9rcmBFZLiUpPM8qo+gdvZZgt
eWHNhr5U5mFmg8lD0iH2UwVM4KHHOGVkdmCX7a2u1rEUs74VFnKgbHieVH0zpbwb/ECbCw+uSupX
YrLeiKJM0XGpxM5hv/tWj7rV5t/wWZfnAmPbtFry5vdPxWwK2Ij91kfBwWgw7wxDZaj0Iz+zN6oe
bRs9qCQru2RLN2LEyb5+XdfmB6epwzW53EqqTe6b1RrvnUIDdE+c8NPpJq6suMLo5H6ogEV7oXkq
p6uUO/jhSuqy5Rgz47xReu3U4+yDgSRhvF4tP6p3WjMpE9dysMMSEhiOYWlRbymxuCT1LnO5fr0Y
5KaWGAxZnBDUm861Asd7FvcGcnlZZNsmGkKMTZUBaWKjX3qSL+PhPhUAPodDBDlSCNinHBDGJSsq
0us73gW8MTcrQGaxkfTrFXr9YDmDWCaQ1MOENDvgbApla3gXGzeehpApE4i4SC/skMjFBJRj50p7
cDYvgeYfhXn0WgY1FeSQAWCSAiajyfPWngNKPiXdi/qEzeO4I/KhPWCvph3SyclCZXUZqGRzyArp
WW3GomBwgU8oywj8UBZjENLolF1FKaPyBi6wVFuehQCn36QhpWVCBGMAj/9LoUY+rkOhB/tu739T
Su05RqhzXtbUx11BhjFQ8BN7nO/0zoL6JwbNNe9uuIp4G5RJp3J9vFljr6YM9dyvKpEBJeNOp4jh
cS39GpCnCfjt133jCMrqOqhBiBDuBuwYkjCSzPmjdiJPknV4fuqhSNBr5UwAYyEyk39QUjLnl/MC
hnKRhZADx56PIFxhhnVDT2UjxrA02xYwDKf4sxcWXsa70BXhHlpu7JzgYvZmMxq1ckL1VmCAwSHe
/f5xzuZdvrMWki/ZlTP9DURuGBHwZxMdhqGjCKI0q0VARqm7n7N47xfkkETW+97ZVZQYr9cYUlza
QYhbbsHzQmPXUA5lGycM8l7SIuF1Q4zRggkT5of0ipwKjlqXDiJ839HRR6kUuptxiCuNaHHLU92s
ijqgyH196qJJlU6Go3yhLk+tcr1HqUdUMqKazutWXodttv4GDOYFpjY9tqJw+TMv1v8puQ8pZNbq
ssmSBt6FA9dTGB0aweI1I9gdp8qoCDQ8GmQTKANyVwtJkBHWeDD/3xYpgixtyd4Bq/3s9aMZZKlg
TVlRYfKMnlDXX9U3EozjBrp/IxBZhDOnlXiRNDLzItgfbNbAxsu9ghbOSDiWfGSEN0aYfoZMzj5g
yja6mxdWo4YnmdiFV9pPrDUDMnCTGbBFO2rNTnwG0K70BaIEsGDh/YkxQZlISPkVh0JLFYCFd0A9
UBheCE9xbgR4HYN4IFyjhvnh1JeNNyC3YM7MN4+OI19Cy6CeSetQxAAWL0cl17r6+lcWe4hPLrFz
tizTSg0Vs8Y44HvZnTrCn8WM5JziEPjhz9JOBEi/bHoPpbB9mn3b0S9hs5+0BmhHk5Cos0U6FlrA
GjrSnIVMVd7cFOeVgPZdjWxyK+c7vuLEoJWg3hm+MJY3+MFEdGEEnQggVxLh8GaeWb6E37uvqqoN
4KrrF+q3b2AX52fMzvqOoCfmofyUXpiRSoiE9+cNLfQfaXm+g2loC2LB0UfRbkq/dQVko5I6Rr/t
gWIvXYtRQ1bERR9CMzG4Sw6ikOjeeNUESfucZJjEIj91amEH9CUSy1z/HuZpMtafvXuPtWhBkRMy
1+UD+nV5apZb+y3U21LZqLfi8Bh+B1EQM0yNyjlxAvVptItmsNcp01CoUuoVUNyrmciR4cjfAENq
Qr8uUPCSDP++SQuL3Z0N6bbtnhRNvWQjDm11c+IvpTbdw73714WwNGSnQ5H1G+em3tg1OxZOR0eo
RZW5aKarKFmD1hD/NhXnZop0Bpe2djyn3IW894J7MByIcWz+/+4WxFtoyT7SQD0JIEfV/k+tfSpE
fQv8wnhsJB1tm2WljbszDALJm59mZq3vHu+/lqGTMv1VCl5AtEAeOuJa78drfI71tm+9azHGPefN
mLicwj/GXD+x3hCN2DRXSn7o+/u+AvvKyJjttWm2gZvbkg2Gt/RsXjvXoWP64luP5HB7KmACP/li
i5loJ20hUm9d/ppUkrS0DcJVw2PVVXZL/5XXssRinKPlmJMhDpqnK0WPVs8FvndLpnCIf4cv1rN4
zBi2rL2jZC3m4917GqsoIu/RPfe8b6hmUjTxjP4o4fyiXVxLo1NnaFpe9yhvb6dPRRctehK3uo/1
tKDsoQckAkFJQcxqLmAUm+aOfsXQc6sFrFLF0E7c+THtMNP9owjTB6TmpsJJYk7ytuaNLYl50P4p
bRmFDmtGDCNkqRphrrExIGhA+1QuPHT3SETccsxb5h8UhQDZ9mW9VJlc+n9vKOoyxOwMwO+bTstV
Kp6q1aPkd2xvqoGYWcY9O81ILDyB7ryLkCwQhkiUoQShb0CzVkMuVb42+M3qtgLfTU9wU3Y7bpBb
Mfiss8A2gyRTHOd+Cdjg6mQwvs93kS+AhvNiSb7RmzmFSKakO5/GG+1URqxiJCs/U1F4wY2S/8gv
yLEU3u/SzbYCn+AGa/t+CEijivHErr4STdzyU/onFZ/G+T7CxrO0eoOdvYYmk1jkegExk/DhA+Z1
rf+zvGkN/JT+9Z3jyQwS84WXaqGOpYfEs8gTJHu/31SNOyGIkg5JOuRP2CyGy1euzJyW+SvfM1YT
JGJS3dK9f962DBSxhdl1roibG8ESF5upoRgT487MBo1Rn5ZPYjwD0irlZRzVMNawftFFn4HtYcME
6axeZFtJ5MmQb8WBMGFcfOI2znoWYydAcdahiUmgVlXhPalr/xx9p44yQd+KBqRKf74iPyDBom+P
vUnI3/JNVTTnD8/CaNnC7T91Q3K/TiqaKGalUZ62rNUMD1qoxDgJOj74MoLQSCAax+z1tXMbWt2R
PX8l9ZR8CYaYYPkukFJmGzp/C/YDQU/O+qIXVedgFy3pFKdf5kYpo166f1yMuiZNuR+ACWKr3/qX
KvovPmLJP29mtqD94UFpfYy6w1i1GZ4VRiBTlqCwQrKHpbgMHXWRT0+q8XnI6eemCr3l0OalDu4r
8BWQOjvnoIV7Ab0gNNnjo1IFeAJQTOPTcfDWhM2p8oHpWIFUzQqzhkkNfteaWkPxL2FsbomcpwND
/xphPEWcKroVw3oLxdQ3jr5luyGqBByPbB3XjalPz9yGh5ehIu59Do9Pw3MJa+tSXUHjK59lyuKP
ZgaXA2J2+JZ4xxu90c2qIow9/jJidHc6gz2/ie7rY+TzSKQ8bvUZTsFZm9sNJFVQoB7pvkds4Z2Z
lOqlN85MfDhJYo2Qh3QDRp0MgDstFtSWRD/zfEkbuCNLALeQXRVQ/4OwJjhIPw0qNXlsjlqj35Ao
Wr7dwZlwoX315Hdzb5ZVPaeHw13GkiseB3J4WnfyFCWQVDVv//yZzwDJfMfOpt0/8m7AxwQnyJUk
r2VD0pn3LvhG0PsXSHDhT2rdMxaBzfF7sAKImxpBDEhHSwyRx5j8n+fVM11Z3hwQLOzMFmcd+xDe
20Aa30D3se9JFSAivLn15731o5umkA39hM2Glhk+P23cb3AiY/ncbOJm+LfsrZis4818oysiHPTy
Qo0T2r4Is4ux97URDnJ8rB2Tf4k9OKqG4bJOFrPv8KSpxwd1/r1PZSaWtn2gc8x1KLIbQh3ZJKRx
pgTXXzeIcu73k5siaL4uySmTmn0qN9cQYpIEsI0x4iPSW8mP+erRooY800NOIKu8VgZiZXDS3xdR
WZb9FeaTuSr4JiHThzI4YL1Y7OIDmjiqw2LbCnJw/9MhoxrDqYzyx+qqlEY1sKHm+aT/8r/JyvS8
JS2Tiq/F2xfNLEhdMXJjvrB6QQ5Bq+ew9ge/OO6WGdGtZNSJcvUCVF/NEJKfQtj3kfCg/ZXNykfy
cnghyIgOspCNLJeaH6Wpt8ZsQeD9JQNS0faKT0JDlMEiRMkH5cGRkDNQdiiGviZRX/2tGoaB1wvT
zh/8ih1aJlbevZwuxSxefvwpUWqS069jODfA/1sGepii8okd61wp5hzpZB35dK3kS2Wm0jLLzt5n
9K5Ty73ZWS2U4m6d7+c20U1j8BP7crV6RZOSvw6SGKSMvJmJ2w38lBVZ6PRFZzwVpP443vmyQ/qW
kW/Id5MivdaoTNoDlNI793hkGJ34h03wjsSrR5Z726KZoF5wmW5kbXFeoc0qplp7DwLoEJTraMos
Df8gF7udmBgyQ0D7GoygR5rJFELl3dLkMPPPD1936Ad5Eqpx8Hly5Xc/q2FSnkI4IUSjNKodjhgY
TrF869W6njkbCcgRvxCcZSGMS5v93GgTQVGZT2sPXfhOFluXqg1NaIU4/Jr6aF77U800rjpCfDPe
Fep3WyDtwFRw5ZymOqdDmRxaxPgSvulP9Os3CcIWCHJhTGdIeygTLWlYWVpsM4oc0jek5h+S0bUU
EKtuKYbIavLCSPzGBuuWw7esbDAFLuuGa5neBAj4RlyUCB3hfO0+FY5ludYnKxVTadCmyNub0mL+
06ctBXERjjug9gAtTIAN5izs5UHXYgZ4PPkzQsejabj+LmwwoOfpjA5gAGUNMX+PSxinOTdfNgTW
G8MKRkQc/soW7ELA3DOLGidwDMsIikFgTY+1ttDttMUy3Qph/ZHMHe4VseHZSxcOAsWRPvPBlXbV
+/cOFXZDeFPUFUYuOl40hmt8fDjGIw2PjuU0wLD6P4UnyJt7FkT3+VmXWxa6jGmOKIT7c8ARE7vE
rAdDxcMS0pCNdEIxlEoul3hVpAFddzVwl+sYEz6sZweLhI8jIvCCjLbdnoBnZvTsZbyNGHKPEQwA
KNPn6tu1/96RssIPM7XXl9TM8qH44LT7ErxUROtmk9hyhcGKUha4oVCZa6Eql24X3pZuhVgIQyuj
aHGticmr3cW9H6SOvt1GYYbTqPis2WQhpVej4bWjRrINbKbrUMbECL419mRzSHQ7YKyl2MIEdt4M
MgoJvxVBUcQUuM7zwbahoFPLsT+JxA/3N/mwPBYaWKXFhT8VysPdyw0YmoagXVPex6tdU2KoCv9c
WWhT7Jqit2pVul3eLro3ESnQUUdxoso8nYwPz6v5WFnCcfWMZ3Bs6/3EWHFQr5u9/VhMtLGUuFQe
vFMWEgFlfuVYd2cpKNo5HhzF7Apq11wwh4bXCHoOahMGZa3MIshM6gb6HaVLLAXNRsaFEE+upbEm
d05+FUbE8+uZXNuQMrVBrNoIzyhtQOmQs26ht2lsc8PkA8sx/gTAxVeFvB6PkR6O2cgg6iA01/Sp
RRwZimncMjI5/uJUg+HM3Wr9+3eTRsJT8G1Qs+LCUfeEtw4fINriwUYnNsvropwtnk2SSsdbHKY9
iJvHHvrLqDYa0l0uY4Hg/cNtOO3oQGzCBUh5+6PfidA/1FFqk/8g+3Agv2SJB3lvgcAJvYtJDnX5
x934PrhaAKxKWuU2p976/eA/jpIlwLZqFGG2SNko/m0mStcRXpljkASgDI0KD2hWR4k5CJkeija0
3ZnKtQY3ZTCehZZWePjpQJN4MHKrO8iKZuuOT7ZMkY6Sw3BI/2Gi1R3L5hsCjtwdOHDTDKvmfuOW
v41ZDEIirtrAA9/Sm5e8o+6uoFjwMpUW2Ssl5tCbzx7iQcsUqQwOQpzP3FqmKfcxunY1sjkQXlx8
SRQlOQEnmcCT3wQ3NtfwZOS1W67ZFwuv71hIsyN+ubhYqT81f7bSxaSwRSeoZUEC3/m/ZFgdh8kG
SknnQ+l4xYxGWRzp4hWKXBhb4em0gsP7mrHGz3sSKKscvaihjLRVmmv14WuJxoHwUZGQJoTD55zN
9G0nzmwz2mq5W4HGwWSBOSd2ZMxpu/9WLcrjuIB+WcotAZgU7gFcH+FyveRuVP2pHiPJIcg1l5JY
cAxMycir3cIiBaueClNwEg336uvj2nMhTqBoEU68TERdhMOuVEYqteGKQPyBVkYgqBBBhFw37ttS
IWl+oA5ntjoNjD/UcDmBkz5FzCL0vSbDKdVv4+Sn+I8FRtf7X59TFXa9E1Z5QBQKHXJTBUbhoeTK
rgalQj7whj741WEstF6FlQX09TkhN46ObucGiFe1b9XKlcQqnewIvV9doepmX/9BO2LYrkHF73sG
gYxyJr/KmVVLwWq9ITXHjvjp/e/8ZBS/SmOML2UnYPzOdnajtgCYqKV6Pp0ZV3T+yT3ejExJ9BiR
MeEyCKXqIwPK6WGdiHz8JaNjxi42tYSAcm7tKk0mrEvbD3YOuyVDrBU1gdR/gGDzEM6l4+s8MdiN
dgOTmTD02HCvcbiFENsNcSmvJmPFflh+XCH57vXM97Ta3okKCCzXZWwlzRPgbMBi01pUiFGd1UDf
HmbiGWbhT5vzKI07BstMv1ip3U7q+ESArQlyN6DZTwCF3nPn7n+exukXUspx6S968TA0gxyFnJUc
dP7ySsPz+0crsDZIDnve0t3xCYFJS7lN0AReaQPWSFP5LX0fjHL9dRx7MklF6ZRVfhX17EaX1JD8
nF88cWdZM1N5wU28puavXXI6qdOCb+p/wX7Iy4OVawcuHtR9c1GniWee8mwMPLHc9O6yPMm0yg//
/pSszjs/BQ5Q4hdnqeBly+8TfWq51ski/DdjiRZ6qoCGPWuGfecie5YCOdWvzXDV/TWcJvmLf/tP
UP+bX7vAz3x5IQZBfFxhhq/xlKfOo0ig8Xz7xvRrcA7gN5Qcn00l1LqrFSBe1lL8Uuqp+AvLfD/b
+52/mSK3JJ33sQ/pEpilJy8c6d0OGUOmz0w347jrWLJ8eyL8qcFZCCpJZMSE93Ca7NPLHdwB5Prt
d5CqghcoU66oyBncNEiNJQ4AYZNHrHrT8dRF2xNVOkzoj1Rb35EllL83r42Cy9G5eAql92Ic02zP
GFIIsHSrFjIVfd6DVzoOvnw6AjS5L0uuDhOm5at+jNTd9C7BYxMOZB/fG4LtXFMHxpHGx/psyqd9
yvZSmMlQDXKtiqMiwwvqRu6UPp02OHETh6nED4vY7/vBpWr0kREva4MVXXbOtLkCkAbQZChLZaiG
kZHRWtQYsXN9/iErx5olRHSBjgNbNhwUH9HmhSFOCfWpiGgLmlRLQiIkuo2AHOeSeZzhxh2Gfe3c
agL+Tismj0hRMkWVcSz6iGPoujCmPHJjsJQcKbrPbTBHPSbWxiJ+H1JqMO8Vc/87ElT1DvM98aUG
e0tkUx6lI1dHk7wNtWKcmqapXkl+RiGZMYnGqWTCaSPgOqLen1FNbGaJZXRHiJyrzk+iH4VTsUoQ
Vc0ebCk9drLd7k0Lg8LKsIIx1Mh7+der19CE5Hhzbrq7m4/eaE0A4oE9KUUtwURk3lXPhJEVD9JD
AIUUHPHqU4nhYQdiAi7HnT2qJf3MGl3dxPzROKjKPZmP66adyLCpGdtPBfK4xNH9u3iMvveJSzpy
KtrswLhTaNtDuqPOv4mz0KclgheY3x7NkBLFopwFOPmB8xr24C41kpuCYeoXhp0ylysd94RcNz01
h2kwb1SKvr/Oum1xZUbKz6B2ju4/eE1dsixjvfKtj1O+KX4j662GMyDHIpV7bCGzXR5DkAHhS+kw
OYW6AhtCdmnJdL0oQ6MP4LFUdH+JJ9IBeWsm5PUPdXzc7qDZ7Yek4+HmUqQ83nS+pftdhlWOdwzG
ozkdyX2YknckQgyJZE3ysXebePB7seHxyhv96uAdGUSP9wx7dOYCWwQrib+xyqC8zxpZr7ms1GXQ
C/NKONFYvLen5li1dj/WyuWptzEY+DQl2jJptsUimWOx365vcVg9dnvf1Qs+vhE/sk3WY7rpGRt7
a6X26O+14vPDwUQGkUPQVfyvIefcYWQnguQtEW/ksoqpf2jkpNiBeLxR687uNZJUBZKEDDgy4GH1
RQaMEwN1tWekk+u/PlUEmbSEJfZ0BrzaiuaYvJU5A92cnw5vL+8Sxmwk0Zea0Iu+7pH3iKcrdh+/
WQmS7KjlkRfXqH/wuFH6IOA6Ln6+TZeM8HHnAgZ5LW0PGmAni/jY/e+Y2TqAq1Jk6awUZmSvjyO3
ORpVfzLrer7MWk6l71LQbJvTlVNcFoN9AIp071jwlZGGwllJMEK1xjVMmdOQvgc7+IZvkzCT34At
3R4+GxMcy0NWRY+dPynOKL2ofGxhab2yhzZG/qq/mqjcKiJK8C5k0gxK8aJT9tzpyCnBLkrZVost
hwKYn+vbM7R+J1in6MvOPrJqiUkbCqV19odl2DW3rXBTFGakxrshphPud63Uy0X9gq8ne7ccVo2e
M8375sZrhrYf1mRUQFi+UAoCFHTx9N2uzK2RbIzH4HV4EJ2Mp8I9b5KB6XNTtDUPEqRJu2DAjOoP
NtegLdBEEXOEi3klKWkD8xQW5s3yhtHLSSAEZsQBReDuJTxG4QHbvXEHRDO2z9hwZ3mFXqvLivyi
unT/cH9UeazAoUs9ELfOC+H+xc91597vyo8bWegvrLaGvdeGA4XKm/cCJ3BCg9nZJnuUyy8D0UgX
/Rl5wkKCBvNGWdYzaAL8n2kXo/BoPqqScLFUouxOM0QNUMaisbLQXAm3vT7zke0466k8sJF9/x7D
LB48yY/HOSpFVQ3vdXXuUIzufBaciSNh0l7FF5xiRjRgNkMIBXd9XJgJlq5FhOz9WA3rVwoGHve7
zCgMuo02PCfYTY+7zXY4L9Rgs2QKM2hhw3ZfNtneYdQ/JnGvwc4LHLeoPMr7GdjskbEY8afA/4xC
graB0gsxu2J/8wOU99vGAHMlMtfGz1pI3CA7UUGJ1mF+s/BcO4z8D7p8Ym7w3gUM9rUNtvnSjahL
yAbgrsJBqeLLQZfFHU4wkD+PkWCc+CpkeWgbYXsug27F81P3Dt7EIahjSLODV60firxKmQbfXWy5
RUSdACUVtl9DZxkxw1udshksdH5S4P35xSIRKf/mhJwaIcea/ayLk4hh0iaUjkK9sMitiC+E5BBY
rNF2x0oX9ltryixvqrcs7IqVFzhe6bjcd+Bu8RfObxqEXCUGYBZUjAFandK0uvqaQbHWV7rhQvba
kfKzYmypS9oUpTGAvCMBcC990qEHe4nLYYJlRyke59NTre1kG2hmqodBbDC7eOnTTZpsVPxgGctv
Tw88DoneGzwHirNVFyY2edeZAi+xnIA0MzfxlGHbXi8FwujSzslq9GZd725mUOIgChq/v6LfOtSe
BY3eUftTOCgipGmRxruVN86BU1zwXmxAHmo7Jo3CdoaR9BwAYNm8o01xInIcvHSMNJWVNXLaQrxa
bdFT1RrA4u1cEpFcm7Tjkmb/bbls4ge8M+Nks6SWxRdEMaVjMQdEmij+4FZkkzOsFeT3Qg0vT8Vh
7RfdWe6gzwVAnfHHlZKxWGiTO8C1kgMf6r6G9JtsTtU4cTxI+6r84xKDcNq5H6LGi3LbRAgwKuzl
5/tQCsdtCD0KzRlkduSKBU5yWr56QerpX08Dw/Zvwki+wD/ZNJa7rYr54KXFKt3P5tvzSpzfR5yT
diCQeoO0YkCAneKfcqgVHflMvaRxDzoi0wVsnk1SUeRml12B2pnqY/p9AVEsRxH0KXbyXD15oxRy
gC9NAAyFaahFFX2KMjX2rpr3qO5N44kTrSnJewAA1E9egQRac8KeN6csiYMXM2ZiBEl1LPmzH8XK
0FxHuijf9TVACcpxzKmL+pyXQtbnsUvz0W3OdXPT6992pGtamIBhszlkVSTnLwAHnUCPavevq8TZ
H/ASc2odO+89Yk69fvPBYkunq2I/LgL4rP+ITpD2MT6puBHvy3p+79J6itx9YcTAy1c1tMIBh4VM
fIvO9HgDUZPJQ0ilMyl4EhH/xqMKcz2Pqrp22Vy88qPqrPNfs3BPQHukWsAs/hi0IyBXKA/0uXkZ
V0av6aOQwcKVzCnvXe4IjY1noVzduMbeLawR/AlbvsdJfb/zZfnEp4Kzenwl+dNBnKyJfeNKeLIH
5cakPlYOABb6TMfGzUpziZy96ry0VzRt+Lb+A45TDL8Wj/7nl1Bn9khV9itPEXdX70g9cTbbzedS
rGxoBTqs5cAxWzMvmwSHqr+QgsCiLObMgytxygpxdf4zKJXu+gznaTI7pmbJ4hu3cpAgnvRMHNpT
fSBTtXDjKET06/JF1INHBCX/Ml28vCCXoyqpMwWp1606E+gaFtkB/IV1kFsILj0HEYrtBHZr8h87
EfwhN9uTiSdW/tbJLJaE04Dc7igbtCv2/9kDPvRYfGIOKxjzAnDLJrg1JPFnz+rnY7yo4VTnumku
kXdQVbmyWEB9vQv/7hq3TxfJ0BnYkmOvO3YWuZHZ68yVWJVXMeqI/06eFAEsVzxFCIIgyOh8qEfW
zI/ySjPUMYeSMtL+MdtAbpHvJHI95KfX2eVqREZYYE4r0QcKIk0jbq+MsFAodUotgZPX7eHwsFT7
do1A8zLfdKy6jvf+r1K0BwjJL5nLPNAAThEj+M5qUUvH/PYL+hHJB9BBHxCXCmqmuT4RZtntKwaY
hUIMQKY8Sj/WjrzqDm01D/muZWu6EfRv2BUEhcy9+s+1jxN5YfIZXk5lGp3OUKZ82R23LOUGOIwL
+0mDa95ckF+7QTXhgwVrjuwiaWV8TyEtv86rt3jciSa35oLR8kI3DFnLVAfDz33rh6UGQYVqFlFo
lOGEc410s1Zt/furtb6CF2COyd+roEXUhRK6cVEjW8zAhs1yjsJWYoofpwIdeMWCmkp2N1mSb802
K26JxaxK23oTSRR3RmtwQb7eiAOPwoF4sn2KFe8s9mqUHO0wXNkBd88z+wEY2G1pNIpp6v4EOUjG
oET183Xc4JjSK3xZtK32BXlDnOcYqV5nO2dY1TXPmnyUz/fzjd9oRMmve8DLCj0tcOskzb5y1D53
ZiTcu81bCd6E3vfNxpVtVh2nmxlyCDK6V90BtxXa4vm/g1F/S544ALTgaqJwfrZ80CpAW+Dosu2z
7foY/DgZPcfbUadUbXnyHzddKPPsmL2/rPWqYKIEV5WXCKK9m8vMKBZPzHqDwF9L7pmCMf2aJkN3
GqRt5jDgSnQmgVfmZbwrYeccs0MgkdHiI+X/qSV0RBPS1IUO8mjWLWFck3FRbFSuy07I/midhjwT
d+sljbmMaF+VY5T8iNgXTxAwoJxpfNxgqzZA6PVvCJNPtGLitY7GIosUnXoYeypGMcyqSoNHyQY+
EAoSnAHk9t7kFO9R+C0/KKeUhpUF5DSfYan4kLva32FlXtsw31+RmLZr9iL5Kbw51zhmn1b7LN6P
tEp/oDBLg8BnPfnUxIIfDUOmdAHZLGPGP2NHowWv2Uqur4AZaS7SL28bRc1rGCFCEXlMYLuNZAEF
RsoCvb6LP6ivZnjSqOVjuqLOn84gBWXJX8h1svUXowR3W1LCjSdch9BR18RcdqyT6s4TrROz5po5
jfDBIaSlpKMQIlo6ehAEsqDRe/q8vTvUC16eNCJgYzH8kFmKlj7d8P4Chnmu2O7IY5LIHvxRuL0b
3z+hxUCmNWVpfcdMIkzQOBPAvpG2mW0J/0DSZg6pOJ78KvlZ/Duf8X3Xkxsk8rvSGIdfa7wXHRCi
cimcDflzIjLTJrcCLowLEGYELRiZ9gvPCkf3w5ETif2MGVlDN21wmPUdWigDI07Wbbrm4ZnA7axs
Dtp8SSZZfXejdp/HvQL7QV4OaWhkttMoE/TdNy9Za0U7kmH/8lAyLOx43M/TXqQsPkaEvo9dYVv/
TJHKR8g3D72PfA+c4DOwGSqm6x9WAoNOCpCqDJAjXGaK5UnuS7Iks7hB1w1R/HrLDAuPu2wIAvuO
Rzj6jqOAvD0TDlNWyXsZbHyL70/PgqAXpP5f/MwBYyr64QZ9U0Nh0h6g5+rMDXnS6IETDtBwFa9b
I9rtMgbo5PYpADBn6lrBGHQiE4UqMhCH/oXfFHmyl3N3ooeBbFi3idDT9VbsnPmtN9I9VRbr78Oj
t3wLXkap8znS4GkPRCuDjtBty360M2vuVLWIj8iq7cxvWhRqYsY2LThJoL22wg0pLSmFOpxSMoCi
NR0V8rx1EHPVOJ3/CYEPcCzJfvoM3WKMeHPCobEMeMyO3gc5F+1SrOeeRhqzaxBcD+AVJnjQridO
dfhJ0yVntSi1Ly0J6Ad8ayzQscpcZLQnepFMtPKanlyGtT5DP0vhfPqwPqdzJ2DjZSN5MUh1T6r4
cF2aQFB0fERVbeqkTf8Pz+SrtR/VbiIc9spaZ4XN1v7I8pyvG6jvSrau+Ko2yD06+3kwyo580HM9
P5n5zcdlxUd0fv6eYPUajBqhtIY81i5FL+M1CEDus3tZ43X2tiBABdLPzZJOci+ri9iqxFW7xKj1
5IoczDMIgE9qSDrdb+0o0e/XwURIic/OHPuIEk9EGcCO7CsCkoGNfDLTl/ojw5Ftxuo7HvM03WfG
+A4HDVrVBxYnzXbg+84dw7vJuUm/QkBhLX+yg405pDPOndwHTiDMdct93oE5R8q9UpZS8CP+1Al4
zEfRNaWKZ924Fn55etru/wZlioGoClYD/bm3SbjTTEzxGqNqTuQ8TvpCjd/0ISfzIyWDWzJnt07i
zD+5wN45ekmDqwif7e1vXyIWIrxR8md+8B3bBH2of3QB5ApwgU3xAgkgCoqaGYw3VeR5958ztqZG
crGGDKrpdyBj2Yqy/XAHuMgI+NhMjOn6gSsZrr9EEAxWQhCRe3rRC4kuIisxA8J2BLJcSOIuoAGW
Z53WsFh232pvecxe1XyKwmCrnL0DQY97GXIAoTPIa6tMBE2AGsaOoMieSBCz3syKIAUo2Bm6mPSS
/UX8IMZ/BssTOLyDvAkMEyDE2tg59F5gchG9fTTXyK99Z7XqwAVoECylsjVXVGCugOEv/ckvvvQX
uFQdDell6VMCB7BW5Pomy6C6BzzSCgcMFWPzOAbKufG3zRjGuz59iQTjbZQaTROTrccS9VHa5/jY
gk5n+IEC77k6h7KxdTfDh7cXBiKKNUYRdM10PwL1M1ETtvBkGw96793ovwM2jK3yNYdpcvpcKMpS
Gfgm8hsPhASeG2gLucxj169f5hA0wfo/+nqVEztd9SDpIwo+TzSFPrItgjoMIDv8th9okDI/597D
zhvc8qbXaIZ1vpogowUeWPuNnmtyGETxP/Afbiu7c4mZGJiCDrOZEoOkfTdcHW3miO2Wp9XKNBs+
MmvMDHz9JgrdOdOLDgnvEY0DwOV9G1/Ma8TmcDCcpZXSeO/0tgQOvPfCaIAMiwoOTorotFLynxnq
aHP1yt84Fp7uNoAFLHZNf9e5h5DXFL+acAVRY3wV3nZudLySJp9MFxyaO+VnPyZuqJIRTGG+UMAy
SLlN10rQDWrrqyGlZzWmcVnCRv9/BwhX3V60cYgWfy4MeOeSYNLoJ+7HhIyIFAJuupSbxTNU29dG
yPslAZzs9Ykfkg90CXM+/87tmdsE+66UJ4/JKQTjdYJZWF8FWV+hPm0Esj+kPAsXL6bYv//bun5v
KbG76QtrBvVqO02HmAPzTIkC/UcMxYvnSjerosm51hxrzio1hQU8mOormyybRAjycj9NSSRgDC4g
Xyi6j5UsaywUcvLvxSem3rXC+ImCb+UVqQebfItPRnbJ+O6uEqH1yC+8hCCGXuBL3CdU1Wotkste
bJ3ZypCqhj5hZGpCnsHEeQusjivHMMs9XkZGxTA80QA+okvx0ki9II53z3H50/SaH53B6s4hsOtS
AbVJF5uYvUIFNA5+tB46QlYkcWwahfbq3hQJPz3/w/roUwjBfI+xhg48ko8yti7y18vbFf6fv+gf
o7NPJiLj+C/gWdZe6jPCmfkWdIE8Qckc6XgMSF4Co/mhkpG1h1FMYZfHCeI4Ac3Y5g+XP2CeyO4J
ypDOyjhuDvWHnNEnUGF0XJ9VAXTLrb/ZvQKQ6do2dKIANmAk+sG8SOtn+9ani3omsGKsLLwBHrPC
lQ+DuMxOhR3ecLi+9YSNdS+LrJX2VTFZvhqhk3KTGE0+R4xnYrGgBOM2kP7aC8ZAwBt0pMN4NLgM
AiKLJndSnDywNtpyhBT5O68kw8ps0YcPzXqzirumhkvs7bUvuiiG9aIYotfFxTplePkm0ooPxJYv
V9goU9PDFwSNxjQYh90Ml/FWxjS/j+EqnatA1nTnSPGx9OyevIGMOO+scFhTRzEqYl5FeO0hNFvG
JiJVCWGJMKY+lOZf4fMInxodaToNsI2oFprXnrBK0eiufvzQjfYAUPfsHkODBZYrdWmRMQOW2CAL
Xm+pICju2pSVm8z/A6vgKD3AOtYfN463MUjVaZuarXpK752i+QfyTIMDXUFVfOOc3Y9S181MqUXS
+og5PN1PCKGhst5STXLYnnbpPuYDLt8I5bEwKqpDK8M30pCohiP++8qPMy5XsCp4Dp+bfPPrPssl
rhVkbLAOQQ7pNmMQ+//L9ZLiIhjXCS0DxX/cx4VgtmF1Ge/cmTLiI3VbCXG9sb1EeYYRkbjgDi/N
AcQooHD6Jkj+xUglUcAiAkW+fbNpbPp1xyv9U6jijvhroKkuI9YmugSvr1I+UD4AVrerFh9zL+KF
t4WeDmjwWrpFtYrCZG1Eu9UOzqJW5opyeb3rV82yKrHLVvgdJ8/he8gsyyeR1Vv/yPKQNOTBLtrS
3Y0qdowfCLuTllz8Q45XUchSKU9SujPhKSRWEHrD/84q/3Nl/IbCnuT0NrqxCqbSL0YohS0X4EWy
4ohZUd1X3BfXjYesr/1h/hl7nmITMUqSu0eWi5bahlMdFbQfd5kT61ToGDOooT0Ie1y5TUhn6R8T
zg8j1ZaAcwqlUxw1ppHJxdyYdc+LyCA6tiXeptklj2E+KAQM1L4eRZNI3DZZ8/7b6BPYKgBktAiq
SGnIzOPBocUbifmVuAZr7lEwffN4d3on1hsyWMoQ8YwA+6YAUKzkVioXdPHTCb/s61uX44fgO2ez
pIJq5bruRlMgRtZcVuB8FFDCQxpN41jODXZKBAnK06TEdOZgEf1b7CCE1Jjq7VizaBlMJqLyw0gb
SmwmY3S/4eSqpCNka0UUb1VZEu25Q7V37dqcfcbUMEvp5mGyxODJR2o8Hyh7voEdqI+BnxDY/SA6
E0A8vuNUxobZxlX2zApdrphoguPHX+DLxKhGex3OblsDh3JnRsOS2L2MOfbnSHc5rSooTtYWg6bw
2JDPC/1Kng0lun50FAUTUXChMlSBqGgErhaXpgO6YGj38qNMm/1SnK3N+KfTpZ8Jqsr6AGq1r9kB
iY93AXAoiq/hwidz1AgU9NMWn2XQMHknsDOXGvvNumydaOvzi0psoW8aLZXNVlqN26vau82U0xwV
k9zUYetc9Jz78YD1KNHDeAzw9G0n8gCh9ON9c5sdA3fS4/NqJVY0hpBMt9Rz7xWXEA/Uia1xZJsT
fp3zukBD6KzRKMkxBRQZN82sn7I07nlOHKe6UT3rD0bDX/desBFdfigXzFL0R1FritpWHkf19Q9w
a1I+CIgZELyUyq1wfCsgRHi0d7BMMW19uZX/IvLKjRWQlNTan9RfzOZU8Qpl9PCix5W5mRHVQGrt
RVZc3n0RfXE2bipN1tmis10KTnjlkRSCTpr2TqPCMb+7CnIPZOZ6akzgAMIe47aZfboS6UZWIR+c
c8gU2dBxG5OwXH57YduKDro7iWV+/6VIrN2mtrEqOycfr2z7DrNH2Jpy5/EM7IY8MgWqAm0EkLgf
3r7abz7NXEgMSxyarY5qjNQ3WlKpoPkvgY1aC7oXRuV8KxH9X9cMvAr+okHm1fLLQVD+ckRAO/Ag
jFcuD89pasaiip+pWIHAQtnMon0jX/FKfS3sFGr5wFEgq0OpAIcEKRcUdtdjkEXg1Vp19Wfsvpqj
1db1Ao9u97DjnUUmuFdDBe2/7iSvI42kqTiS7qZhS13POiL5FW+GcMmF2SZp1tf+TNgo030EPpBa
vkx13Z+DOXv6uN6upGWJOq+ewPkShCeOZwOfpHC2p2kHJHEMIMdpuJ07lPrXsLOVgc35h/drWyoI
69Y4I3ZeyHPNxcnqez1Q/N6mS3B7aVPlBreEbgSdI1X3lR3zZmuYT/53NhNDLOA1s+AMk6GSkqEY
5BqT+GpPsVCPCswvn58g+eefsvviQGewf9okIlh3Pnpk6+DyJB8BefEKpPaLYnzQpQvAuCX5OaeP
60lclvh4R5hTiAt012JC8Y4Y40QgTk61siFFWQJyPda3FCO83+QMoD09yx027nKTl16Rh8SjPok4
rJDCTZwjZzbw8MpWPKqikbIiz8G/qlCn5T59GEeibMZHvpgVU783m+Tpy06OQaLXqMnXBLXslRm7
D1jBNDgz4Tl6mkF3sdsG3psQyDIXeVEM9I3GFDVjVZhs071c1IgNqzrs5i/7CjO547tkC458wjnt
t0fZV/URgdohPwSZqZsYgNR3ieJ7n0XHNLbdy4zW+hhzFG0sXR5pmh7wmcA9nZ23tALCsDhAMeaS
XHQ9h6IfihoUMIVblxqooG0VfLXh5/oNxj0R8Dk8dSWCgZE2vwmp+mq410RsDrRgwRNenKfZ82sh
iZxzkf8bVWJCVjB0pDLRpOnSWSzGsffjbvwRoSSykSCMuLuqfLzM3PC64Oe6BrqMRPABTbiK0ey+
vd8t8l6KWwJr28D425383/kuCGFMKX40i/31yGqwnn1floL3pllFbaCCVVyzzkUuFjWZ7JEqPeT+
+v6vBnSS7TQO97RUqw7IRPkozRz9DlD7j8xEnrd73ZXcLI3pOW8aTqfW6RmW3WdXHbjmkdU+0ifs
VbwqdNsh9A8eDpDI5S65ME4h+b7gqC2xZS/ti+rCo8jbJlIc8XO6zhTgI2Znud6v4/O0hB1xCFWD
zKJHMxfmnsVDwp//sTK8FPiAcdkEnAikxec1Edojt/9XVDMni1aBM9W4LZO9CqX2iIbtHS8eZHYY
72iN1N11aS/7TDwx0aKXadZU+TdLvT1I7mir82csDccgmm634AKyiDxqCecsnVxQf1CtR9NlBSzs
cxKFly+P0xtrfTmFoO3S0n8ZzPhh/G3+xieVmAOuQFaIbAwxbpCIEhUW4n7jP9Q0dkiie/0jQWLP
h0H/Cabk7SjTXmNxfWtgDYOZP4Jp3Rbqpzm92S7uSEyiTvEnxIs4gNqQOUtFda9RJVHxlPPWOdTS
iVaGOFWGtyvJMunIQ7AvY34Z24QrEYJWP+L6wz3jNOjDjmx1AQX0zv4DjdGPVh1VUp1pdBC86l1k
ZxCrLrkYGLU75gwnYfJgX36M7bBVbaNsZlT75dxlLEs+RK8RLScbLQK2Sv7YUCdT4PioUOb7RGQE
Lc9bsJBA9EkhTwdoRIh1JvKgAkDj9Fdq7ckvgGU0nU17wlIMy4OeOINri70/5tQfbrTeViXHtpu7
HTqn0zPbP0CUaZYVr4oyX95Tm2nY2m68ft/WR20BoS57y502iSQq/Y31fgFs889SZV54UcIRKRSp
igAmpnDjzMk94IuvR4b//2eKVMMt37cBHZCi6ZRKr2QzzW4NIRrEZUGYwokXLIynsbVweakZSTnp
hDYDQPaSOFVVGDcwX5cox6MV+Mi0s0RWXpnXR5kSSonFmbdTqZ4wNOCKwFcWbxmirVaSekDv9BXu
RRv/GqaXHVQRLrjIYvbRL8qurkIxwPl4igZJxfUlVxcHhtC9dRUL2rPwysswClFne3aowYEWrs6o
IBDREQJM1L782PP+yb9FD4kM2ChY6X39kDVguS5rxJqo5CYBNN6KyWEYBUcHnumDeVBPmKIF/MQh
hU+WPBalhYML5QDMaJDBEa6ol0AfqD9NOe1tWJJkL9r2h/bab2Qizq6fqAIzGJVjDP8jbNqVhkja
x+fJ6QuyESlyHKZGsW9UuNdcvIs6VGsQ2FBNpTmTyad257NbNpe/ed1NnCtitKsu5tzO0gSLv8l/
lMQ7KzmefpnOssBSm/1Z+/59EvdYhLWgaVMKkJ5P+10+0WaETEc2reSj14jI/EIoqSGU/yuRrxtK
1uhTcvZWPtao2w3W9Pk3vOv61kcwMgXOAGk/Vk1e8dL5baK9NeqHLo9s7byGyzY5VIjhPlRJPG4B
zr4kwLynoCliNNriRSUXVZQJ3fUA5+J2XqnZA5qvP9XoLnRqjypIdltwPJkqMoAYdeTC75xpSKCd
uOAlZd6G7LsLZxqeEWB1XsOqxYdsosz6sq0s5RkH9MkPQ9np2V1+ADnPUcV/HmSRK+oDYIa0UR2l
usRY756gGMbBFgGG/4+ME0B+K7++nw+UunrNwSh3VyAxvuMKHVV6wViu2tef6iYcj/E3BTvdXaOh
G4UpwiTXgMSPEur+RLOTDc3+mzJgGl5CZTghdHuweGjPflX7qI6Bj7A7Joe15LuF2I60fj4rpX3r
vSMRhF/pxK4FXeUIitBQboKsYrBd550JsSFmU/JolTshSbpLEz6PacoYIiBHRBMEJluA++CCKt/c
+m4C8WgThowEjeT4K5MLl5MJA7tnyIuVxema+OIY5Gd8bOl6A3NSTUcpgwMt2VHwFlErJObcXqsv
vql133u6GWOQcXlfYElOLZBohc9w2w4WpgcchH9mbE+DH7Vp7q9yqoInyqyULmvMB8ISOnMTu4lf
39rMdps0Rma8t8/2S4kD7jcGYj7uBLNAKiNbxWqf3K87a+LWyhDNzGx91iWEfCdRjKbntOhcS30R
mjaQFTYkI92M/vWcItvY3qvc+Efw2BK1CYlfGRbakXeRWa8uJ6GuySz5+SUFPbx+cRYZvXqugowt
D98w2DlhTjEUXkD/GpqtgyqZ1zEgS24tAC0ls/95YQQ8iW1LW50TRi7exTX1iD4wysvqdkTH9Gs0
VyhXM08senbNgf5VQZHwhTjDqS0PXd/YezKiKLncSAQCjZhrl30sBFvT1vy1NODX+pKwbvuc0Sqw
DZTcysdO5DhOUxC9injppXcYlQn0Iq45kC6HoETlVrcMNnqBGJ8je63kmhXc/iwF2qP9QCdS2qSt
q8fw3iwq34uRB1PUcsKW5sAFBJ1tQZVSfmqwNnUjVRWU5ss4dA0u0l+2c+K+xS8zwNMl79VBWYzU
HoKdX9cpeR3AcyAqKjmywoAWYBmKhY34H55wXE1E5ZQt6F4FW6xwmo3o1U5eH3jT7Rc5OESxP0NB
YCq0epRmF1W7IClA9PgBewiPWCRIKQN1+AM/9ee4WhiL9NUdiM754mWoii5smW0L5rMYzZWWcX5E
9mlB6uAkicFtFUuiu9azxM0qqJc9k+MPNEt9tpliGZioUiWFEnfOP2fj4dNrBjfYXm/iS3F+4zHT
ERSkMn9upU9039obzf1j2L93ADXjJVOVmNr1k9sMuuMs1MbVC3CmcSC551lrAlYnpvoW/KOxVHjk
bah6b21PEkZnEaN4G1hJAk4Ej2HC5h6WTvngnZWJMNJi2KKKvP76lCsY/Pqcy/z3Qed6Tf/V7//w
WhTc9IHqce19V8elK/sb8HpVRnuXKiXaM53B4fkTak76U0cevFwE9p05UBNjMremVON/3DYGF14m
b6eT+YWSoIs3BAwMqb9fB9A6iTqSiECqkZ5Qe8/f7O51O2ZdtcX73oXJWCOxMEMst0+4D5tihkhs
L4OZLCmmHTjD4Bbca9QK9yESM9nFGoOguc3zF+TkRrl7JuJqSC5OlALcGKTB+uoZwHlHoCa9T542
XCjSeYzmgb2nqqalePadc7BGpJhLKzDqihRg66QG+VtwKlcAGHMsh1OpxEvCtjHibo37mwc8tu2x
w3cpMBaTcexqdU4ysuyEf69JjlX+WcNZ/qBseMd2x58cjM15MQSmzzNiWT5ZSCLx925hzptzvQ42
EaIWQCJ7vaZm/w/Z65CjJvtyMLa0hgM12EfnGzRqWHP0GY3uE9xhrxd+o1Td3qWvF2bo0VjuTP0O
H2JNyzaYDDLnjLCXlcm/vKg436KYkVdpru/HSCS5xf+ldEjnfCut320oEt1X2qjmJ0fJKsc9uCo0
FsIKo7zrNRlUX2OjLN7T49R6GUugZ3cDwukxJ7EQFT9Pbbo1IWekamQkJUptGA29dud3S0GRgfZf
I7J1WqK9bT91cEinS/W8Xz5ITG3LVbwKHHl0/bOv4s62XbZUXWBiDSumzrT2EhXL6uCQ7YsiSTxt
jlWWSPcFKZymVDdIXwz7gNgTkGmcBPPBv/ZVAHnJp5fYG7tJ58y/djG18Q/mODX1yLPC+OOw9TLq
evmo5bEGuP6/49dpfhtDI+qbCpGopn1D1uFaZsYqxjITU6Zf1W9uGngZTeKxnk9w7zb+0fzI2dLy
7phRji0IRHoacML3m2DZbYp4q3hJxvY432zZrJ65Fh5zCFTb7mZM5S1ItumalianAsvnXvofilHo
Glo26FOhj6JwdfmyRAnXx3LvSgXFJB29jZLnMf/sFFZIDNeU7hynjgroicwEL1UQhsUtAru/g4Jb
xZ+SE0UhmeRxtu5DiLAcmdHAlJZgFcOrDjuiM/gzKFkNc1w0ZzIiJq0KW5GKZOk/roDrWkoqnoVu
vWbvFsPOdwESaZ0lf/qiUnufTgdfNRvqbiAJrvetOGZT3+bXbCSeN9BG0AgJ3gp1HjKtTdE5tM8M
OV0tFzIU8nCwYJBJwSQRBbBfhMe2L2cSAtKh0NnDwYd6qbP4vKr/dyyfe8eRK3Y8RMKza7iHvBmb
+7Ol/tmdRGZKFEHe/WXUM78IPjB1zrUjNPLSkXdufoWuzhHReiCmuXHK4K+3cLVhMKaFW4JHlKj9
L76JCKE1N/s4yyxa6gSzYmgPaQnZgGGmvQ6g14zZY86oQszg3Yyrf0byDv9qaMTpeONKcIKnF1Ie
F0TeJzuGYqRcW7aXqmdWA2pbJyo3QqLYdKFNSoS+uzZDq7PLzAjVRAGLcj88UKJiNUVRe1S2XgHM
7a1r/ATOI2C98VSMmwkONQmIL5TKwMXb8uWMEutieRiJBh5oTwK/U9hrtrovOrYSGld8JKXndxfX
ZRFD6mpoaB+qOXmTagpUGVAX9NaRUpSvoX8FY+9f0fAKDxwLUwIaetjxAyITn4tgWFmCKeIyFZVW
q30PHILQnXQU2rLiWgzwzIjDbxavp+WZCPYalgYm98iWuo7Gyi9wanm9ezTI2vJ6rV9JGxAPFgFG
ZljZ7YonDTVZ/vWVQP0dCCxmcQYlqMmu53Kr/Tw4SqPZeL8+1g8kGbXyplRrOPESL2oT6sdDoLH3
DGvAY0vmnAP7T4KagH7+ewc5DWuWoF4jMkD9zMELrCi+DZl0Se5y6v3UHgs78AwnyquO9n4A4Tgj
M8XAv1SbcIh8LIKjEySTADi/OiGGkX1Cl/JcMs5pymvyr7d0mBNHjsZR+AqoNlvOJdW7AL2C7eUW
rTMsE/WJHoH+MKcKn9CxvogBELA5ZCcuFdRhFp1iaAY2qJI7SSKfCj6b8RPMGRlAqEmRZQSRFKRE
BxUf2OPtky75ReIpqbMAyD+Wmb8cgppxUN9ItEDS/yeHMnnBM+XMwPnT2MwgZEMRuDqW+hCxcnqU
DRmwZq9aAMUbTHl++xBW6/CCCIj4EgRFo6BDyMxc3hdprx4S0/uRcnRKelVG9m6W2ZXx1kE/SEHS
P2M3tOfM9IHd0C0IdDgvoeuY2pHQEJZtylmXRqxFxMXeolHPqcLawlgU7Bawy+BhIR8iqB+Vbu7E
+J6jTR9ABOV1+eUEli3QHjn5psYvDu7vHtBeQ6hl6+M6j4UmvgnRFfXT2Z5P0qREI/jv4EKKjiLL
tDLtC2sIHavYIgtW/nwdudNY2C5XYzBwx65DfKpkwa8rxbKkqX7g4An/7xQxk95gROoMWtzBXgrd
me/hETBiO8cXzZ0htMSI+n8ZZHQbhsFsIaE/rCKvXxnyvqAUBiK2/jexSHrTwOl8w0CdD74as+bO
qhTD3g5ytyDLRYF1LGjn4mES2gPDTYhvHW2xDcvQ8MwW+jbvQgbg5p+ebk4NO8LsiS8H1cfYyL3N
QiIu/WS9ctJPWO8MFnWE8JOCh56CIBLSBg7vN4IjqFWulXWV3E0UEFh8WTU7DoaxboLPToky+GGB
1J5lhWNgu6Ciot3fsGQEA4kXXNmLbQ222ZvR0m+JoxcEQr4O9RdWaf4XdDBP0PMlF4l8cwYvnEjG
zezsK+nV8CeRnlZiOCvEak6zuoDVmMOpNUOyiWyrsVGG/q2K7M/P11NEW1isTfi7naq00yZrq3cy
pStfrKsgy0TIYljhX63n79wBfV+1w//bqOFGu6tAknbT+3SNsKD61hCgX8hsGk8HDsQzbeCtQYWF
/XqqEjVVmrrRjB/PBRdJ0tmxEh8jnPsKJ1H7Wg7B4GIiqvegrRVuadACI07sAV6E6riIPvgCXBEt
hxEPizfIMLLdWU9ZSn7J656op9yCCjgmrYqWHxr6ejluC+wMby5R5WiBEcgyTKSTxhg5l1vbqI9Q
HBIW80nm/pxQXE2oLGosUFrHXAvf+MbgCxWN4WP2KOEmv7PATZvLgl9ouiNDzqkSnIu+jX/mSVy7
pppJV8D/kqKMwIpQ71+CoLaaWztLv1jO7zXo/P+ayvVSwmT62jw2/FDo7XK6ydnlFRb8g+hmIht0
oszbTb5KTbscQkyoFGhWFlH9FfBtJxbLhzVsY6jcndPSz7fOS82vE/pgKf6pn1lzvoJa85G4ubbE
DAa6ubowyg3UDl85hDaWV6p4yOALARtxT9BTkDNnqVfTTssbcFcpWtD+rG9LEFbH3fea5JArOxsr
ziW2UTMXhz48s6wih9TNvC6Qtimg2J93X/Vyi6UYg6JJoBDN4bQEa9VjJ/QrbcQG6yNSbQMFJPK9
qxG4peGrk6TRNkZ4VEidSUVIEd1fOkUhZ9Ah4v5lTeWXa8lELFqI6xD+u5qgyRa2w6HzdWag6EB9
iwJVyZfe+zwaVINfiYikkrMYaymTgnhodihzXfimlRhvqYvs2i1Mx9Yl7vegSRlPa32OeGwQz72N
t92gFkVYAK1sc7GIkIVhJ76+WcHUCPLPwS3oWlGT0rLz0tBK/PV77m7VrAyOnMCYbDYfkEjyNr4j
Kzv8uQ7R46t87Ch6uwB8uxTyNWtVscrfvS5vXh56oOYjboG3T5zh9KqEanfFn52nUIfXnJL0Q0X4
Txls8l5CDho0hMbCKMBntGZZj3KJOV30O5HithbZ3Ska8msugjX/3sqWvAOPWSBVa+kCH8Pd4Y/9
GU4RgDt5l6dWrp96DekCqbpqft7G4jA9X/AyDCV130O/ZMDRUEONUIoTjLok9JNYI12v0Lqof/Tt
ItE22OX6wULYYJ+J07UJboGGZ5lGsP6BAa4r+l8a9K3ZlwOPZqbdDwt16SNQGphnf6wpYGOxpXa0
YLMFnzgvhYfeTOTcOAJX5vTM7pfiCSTVaQX03YDhprqsuqGrjoXjrNdDcKs6R9XAqR5y77aGeGoe
kdYivjt7TAadgrhh/8XF12k42zBJAOp2wtU49xuOlN04mi94acuD+OOyU6hCmfwS5QXfZAH7JVOe
K4jfNAkaC2wKadgR6N2yvYhPDhUAvTux7TlR/02UaENp9fH0jsw+RGoUXonWd4+V1Vasq5pTin2r
xzEpHbH+kSPVEcFBqqI0UYJbJ+OjtXOhkTFsk0ScaQUgrvcRjKWq6PdrtZZADdsvaq7ioit/iE42
WrDx78O8cZWJPrEDOQMiVtTmNWXY6m579Hq+H662n07rgNT6yL6c/gtDV6o2EEYdlvuuMFclsz2E
e11x0vVkJhHQrs/nCSM73vOtlv1uUWH+PleioxyOQVe9l/pNMFmCrDgl2DKb7aca2WXXKlMkC2DJ
gxWLIFUloEsIobDq38/8mCqnuuIg+aVYhBwdmppPZT/BNh9b+bOYLE3HWdu0J8Sr3aSICkk86p1m
ngOsFq8oix6tEL12jDxCbpERi9ckijIUBecFblFIT7BXGz1C/sfTH0K24VxCngIMR52RZaqWZCAv
4wfh9b1LsEAeEXobL0kX6ejPBLXRNYs5LALKY+OYU1fUoIEBAApugc8B+zD2RkS5HQnAj8dkyDT2
YDvxtmqKDeqtZN5f29yapNI6oGPLA60IZgR+HNg5tHY6wqaDtreK3ywmf4x1424BSDDtCeGt20F5
07OqdGmf3PwRw3ZeanoqzQENrCKv1Fez4hUjx0j2wVpE714RDhbqxfFzL6xn8rp4Zc4Hah7Qeszn
mlEWRwK/rW80MIRC678Ewh4Yz/3VVbXaaaDP2rCkHnR75xlyJPpLA34LA5dkQEX+R2y7fgHf8k8b
dlCHhbgbZIGUBRKib03K1mZeGtmyfPotSW5c+Pfqx19pp9Fx8dHtNpzdfJmlIQTzgZYUk+pKM449
6PDlcj38bcB1GVl+6Jk0eQ+gs9+bI/sXo2FmovO781ihjEGA/8B8vzVVY4IhzEGYJTcSlELwL7uu
XZdgGWE1hhDAjb8JO1YgrRKbxf2EboMXEmnUv5TgEdNrSH8f44hx/JoKPxaxJ17l6tFiGAqLo5PN
MxJboQTOUekIpxmiIJYot/m77aje/tjSB0L1Dq581+M+vDuAx2BQYI8JlWkUWWOsE52WM3LXRX94
VjjGn+j6FT7Df5WPdvDmiKWnjgoTSQR85mtE7gOcp90JPDoGBWO+VIcMahBw6DQd33C3wMxMqUzj
mAGFF6j3UZ1TcvNLjyFghHgEyw8bJRyLI0ml++1o54zJoKHR9/WCoV+a4jJe6GyfsmCDVySSkqCH
zPalOmGaT/x+06t/6pvllhUd64jo1FUwYrb+uKjH9vs2GszSbVeJKRpgR1z7XO2A9CCG2YNeD4AV
FLPoJiRzmLby8KZsX9pakpvasxZny25dz0ajruHBKYnLg9Ss4PVdho6NXyFN7PIN2xePdRSUeaG/
2PAvsBq+fGk5xWwxyUViWgEqcnI4Tz3hXEKKkghzqlBay2EdtXS5AcqOIJZ9zX4z2MEfKINvdsrX
VQKBINlZ2OnU3zGsuEADZ+0P0avIpuVS2Z4XJDcB8egL0FSqcJx3fxsDwEXRPeLzT8LSFvtSvT4X
5c+yrw8LhwqRCKR3xsivyfcPyDEIpEvU60cx68xe476P+ue84J896PaxtYtaBs8fx7YTMy2zM3Mn
yEkWf6fgXplv0hnT2zO0dlHeJJqg3JTPagdMQ1OHT0bzdtWSmQEsi46+n6PhwXBzbbQQ8BReQwX3
n28Axhw9QGzzRTGy/SznAI3RuWhi4sQVAvkwZWI+oV0o1JNgozpvHYxgv1o3KryHWtekxlbgkIRP
fdkjGzIXDFpxHRcu0aYfYP48vW8+or5Gw2lFQiU1+x7BZmYQEk5S4ZjRWFbRphZTuOM6csB3RT72
HJAzS1vaDi5W/r/nRnLwNJA97USbWjEQOUl9RQRUk5L8yc708MRAEqvJ3Hmp9nQSfixB0YmxPcTR
ztss42cafNbSc5bAoggLtFKhn0WIb0cYvOa9XyrElg7dTI6bzgcWwDcx0VWsWgeGpXEC9tjzZgoX
qE0spoetbfwD5afeIIzsH+DmLWtyAdS3jKVkKiS5KttRX6DolzvVm0QYecNdwM9wBrF29d4rtHge
i1sYnY2iZnWr6vjh1FDTmG4Wv5Mm0t6I+ej+GxDpW/F0rPVcGNLzYdg7zcMy5G2zD1In9u17/FqU
cNSD7YQzhEL3pPpBUwOPuBWBYIJ65Tz3SqW+VzO7AZiTAFhi/ppdN3Qk57y7heZ/UjTzYoAQWDqY
CQDqM8hXp9A2/kzBi/XUiWVBY9v3c8J6e5YmMmrSAN7Hf40w0dWgeKqvjefTQ94hKPJ6lTmvsO0z
ATXk+DUVjk9/joW8YqAf9+sj1OR5YHB45gqMOP3RflXbONRKiu6eO4S/cRXOpo2P7AmBDn5kspib
7vJl8GKs336ahYlXV2+tHULqQ8D+GV1dTpr2xhvziJa26cif15h9IhQC4GeXnzfMP0h7x3gCgID/
CBBd9PucOHtV9l3b3QabaESgeKB6t8ZyytuePNU+0H4Rv5AMVltIP04dlYnL2jk/1Zg3UCwtsTfK
iSEEbwhwFiHgn/QAvSmHf3kSNVUkH0F7FSiY6hu/3/2uv06nxIadR4mTF5gx0PiUh4Ni/I0N8Z9t
XlyhBs0Cke09dl0yFXytyj5e3z/z2xJR1RPcvHv8JNV5jV1phPPoQOqQyKGBdP2iw4pdbmccRfVB
wDJsqBZzT650QDopPBxUmG2zbSC/eMEK7F+nD9ZH2DYJIHbziR2/pxYmrypODg3mj/xPE5g8zfUL
21/Kju60fj3vrmX3s5R0oJIDyp7aA01z8XjJssl7wPLtmeK8tmO3hdk6kWIiYHTB8Sw/bVzEJbne
Xp/71mrBbBfDCD5M4SfIoAcjbaoBPhHgo+5hrH/f0ROZ/ua/X3kqFjoOFdYPhfPmIn4oGTMF2wzT
c3WieLVIpf2h65SSFCfHvGyCO5BPnDSasc1gdb4oz8M0GmmFjvB1hpZ/F6pe3Q9WBvqsp4mO5RYz
GH/QPGRTE3Botd66A8WlRm6+HJIw1c7qulWj+smc6fFPuOqT/DfLM4sCTS07K/E/L9O2osN6YHL+
qdgk/nM/+ZqbruWxGnV/+jivvbeJpcb8Fn/QGzmkuE69wsQAGjXSRRAmZjC/nR3F0cun/pXTiCX5
Nqg5MykQ7Wf6KvJpZ4kZjsStKRjF+s9tcIxClzSO81Ff0XVHVyTMKhZAKRVE6xgu+Lb3TyxpPLYz
OPqgjJ4/ujT7bUZI2OoEm0rMY3+3W/UXSkGm9wVFwAbB1HkkkRTND8QswiD2vgLcon4ned87FTyF
bCV33dqYG8WndcvqJjGq0foliBUMTw4jIPRPRonEZehibb3/Zfq7iTv21Adn5y07g7Gvue29sfG5
5DmqI3vEyRhSPxqhwUBnCOcZPodZ2QLaEknrsz0GQaPsqjrR68zPNBfCNt+Y0sL48YAJE7hLgYXX
ArnZV1K8Qz81rIO2SXa9Mr7oADduVCLsOUKCCKSpnqqKJAV6veg7nKKQaHcZBNLt9xSltFzF6wfm
fsFJnq2DEB/aqv65ekBcO3n+32Ofy3lAxK1eQO4kr7GB5vB3jxr9/DpRZxuIQ9O4o1jbDnyITj2f
Hmykiv3kX/EdMJDYGJ8reDcTAGE+/7/JD+wk3ss1zQcNAxeWLqIpeqO5LlaRMHUKRkVigujK9Uan
fF9lfO2uJ6YYGgFRsiFNx11Oz+hD0rUdp0B5Ztucdi7xxLIVH6qOQ+LMwR0lSJt1Dzhv/Mnx+SbZ
89+Xj/lIGmw4YyF+UOO63dxI727fT6hOToWsG3+xpKJqELOywNsw5kN24+NQ9HtaIbTl3xjJWXqq
Z/scwg/0ZMriApsmeENHuDWUIOfMsJGzXZH/gAYHqUNkc9OS/teJ8y5etDQtqaG+BQKw/RzP71CL
RiKpMs1+udmQrwBiNKSQ9J3OjFcoe52j8y3dtQtTKg6hd21Shr0QSA3WrYlqTLZleIBp0KK+e9y5
G5tGDasHArPE6+2/CODF+Kh2SyJNbWiV70vO5kgbb7BN8i4yJ35eNXZu2NUww+rqTf+r0pHuRalY
9VPESJYcsG7OmtjQzIuq5VWGhhBCmtuS5A6k5GMGB06AbInKVho9Q/dSKapBZVfAfwPicc/L0RnC
i2tylb1rbPj4IIWGmXRhgV19ojXZ3npg1hLqJ0WtQGG1L+QWeNprB17bssUT9rLFUkvLfB4arZ9K
FcIow6DLujfNDkvuRjA40FliPCazQMdZ8edwoYbIg7svQSXj+WNSyBSUufESUtHq6i6Lji/thQ9b
pLcJxzLjrto9G45D3/suUFdN3OQpWKce9nx8/vxNSRy6H3tNsZB5w1DPWpMEtRzcq3nKTYufmqU0
qYoJ4oJg7dpDNq7HzOFe2OWynMH9kz5htyzVVlqkV0BGfTs6RpF3/KzF74FV2tBseQmsmWYp+OpU
abSDjYOlHFfxG40KI68Hjm1azjp1eZCbw4jv8A3Ff+YdzhDEcGoMCpo1wFwP5UmlfzlT24NlKtVv
Db9saZOtkMf1C8ZYwyKnm78Q5oigldGoq6xr0mkeH6xuAKFGlUMnVObZYze5FQvhs0+9GQ7miSNs
P6dYIYBlyVHb9I/xy9lBBV7smSBeCK/erOh6fbggAhuMEsJusx73SZCQ5sbMNZHfFuuxb3/P7l+Z
Ce+0qBpMxMRLIBn0edNxyU7P9H13Be7rtVLx8PkIEYdWPeGq4yhnqpLncYjYwwcAzaiYW3qgraI6
rbK+N9/ZIIx4dYSEwv5TOt/21FefQr4N1o9cgiIOQBXzxJPgqz+KMAPERsb9Df6rHYuE3G/R8N8l
AX4A18URtUOXg3ZGEoI05HCsWWvUN5Jp6FQSDWqb7bgxfEZY/DGSgiQN/Q/HpwtfEWIAWKqtqxzW
gq3eWR2KgQnzFxrH05mrrrV+qcwTyxfGFAh3zoFvZxsFlMQNgP47hb4cx8mGkXeKz9t5VP3P3saF
IRYQ7u8Vo2HtUxxvxHdWxlbYSrmAWEY8gBQeg/S18YoXWh/xhxxsWOzKBg9j9OJTzEZGHfIEIhxr
JxjEe724mkQl046B1sJlUbfIAfdbLxv8RHVIIophRWvd0HxUL1v14J4yFKdP6KNWp5mUaKRQKkwu
DepzkjekHS8Sv9pyucZVMxc3UkGEhvLU4e7MqEGwrX4LTdfGUR+oGJcAR3GwEhY+7c6efG2n+VIe
lAHUKcsrNMZyPBbcfJHQSMeU7eaKmTbAmbmMJc3yWvQ0Wma3qt/RFwas2Gs6lnrEupRfERt3C8qD
3aX5Dzgb3SproyUi/uNXh8TO3wJJ+qMCFaikvo0P8mWY4NdJoQZ5KdZpsdn6mO09dQkVRUHl1xaJ
cha++7WOiu5xX05jFu5HGyg3xo5Hv96lJxNttBv5z8/rM43KAiqKpchGQs1rZL7iufIdCazM36bJ
319XaGmnzJa1MvbaUVUjCfKM8vcFr10HamWmmKdnnmUOv2QM4MF14HeMeRldbYV/F/qdBbkw8Ufx
CMtyuFHi0/piCWLb1DqJQE7G84dP1GU23G57b8laqr8QVZGPycg0lnpGV2PZzLxu7cG6DNnFEMOo
Nr+74ItuAuSv64oXgRRWyCTbu0cJ+IH7CDC99KvxYFojA8XJdAGm6OVFuIfjibvg7YV3711UZWdL
418iFlIl8C3jCcw93YikAYK4R5CG8B9Nu8aK0bZ/oH3vcLYmicLYeZsok0ljJAkYoGQgnD0UELmm
t9VINb7LVDU/3cqlYxIm5r6HuqfqvQI6O0fK4ChA0LFu+zUKuQIJQLwzMbi4ceXHOgsFoWz3Csg0
F/ynTC20qklZPK7eiyFBq6pFFO0LWURwtTs0KVxwtGkKlZjmhuMzgUg77eqKNB7seuqij8RJoGNf
Xe+MsrFQjwxAel5DbikwsLLR8aWR/EKiqXFFPzu/RIYPTQ2cnJCmqyzL5909HguLcBvX/RJCTiTx
UFVNYsHkAbHnWicJkR+z1uZmb1H31rStkj/QG7nFKf3/uK6QarhUZP135W3KgcP2tui4pUY+2XTZ
dFEAd+3YXk3i7FVb3eSDWEHuohWX4233nJ2z5zxY2FLiwavMbbrutYxEArRDv8DxIJqR+61k9+wp
AhjShNH2U3riwwyRocRKBunLUsw/eYK4ZOYeratwDmM+bvq1LMR2pHhcV4Cu5QR0rLgudzmhTJEC
hpJZxBxWxvKpiM+4smK7Evk3YmdZqF6mxsiMXR4WWqsE7Q5+uLDWYQDy48+0gpnJZcyg9fh+qfCx
Ox0q2iBHz7JhCgov0RM9vsY7z/Ou5D7PrPm1q2sctALYEJnqnMa4aAA2C1ZFjlLDVsNujfIecBMN
JnMXmP47GFRopb3dD4gCcJkuVqZ61GKKTB+fG4At5ul0Sv9Y+CyEpa5+JqV7O5wOr1B3etSJrTfC
5s5rrcFbQ2xQKC/701MPj1fAQ0zVzd3YCPPo4He5penMrhcn88qBIVSMorVYdJkyC1aYchuV45QQ
CoUi9F5AaFa5/MvxLnbyq/fs0QkWHtH17ePmYUiWLhbKHBdFKLBZfbUYQkNWNLSuqunVcLMR/snc
P8yAMcpBzaveD20gfeqwVuu6XpRnZHemm8RJyTNoa9hkh2fDUtv1m09joOTuH9470IxeqaWa9GtP
P0GupJORmudoSDojoh01j/LCGuSelmEgU6LuGO9TREKhrjaHFmujIuRT1vFi96h8ibF39Emnc5cc
OpzhonL3bgd1j7xBxYgZQTb1Y+Pa1txoNfe66a70uzyGOHzdSeYBIQsXu651lMbq0RTvFH2Bg4Kl
b5eQ6qogNe9aeBTnSPKlXnBHPw+xO5i4bGX7mn8iHm1IY1QAZfwMSv3zic3xFkcYh8HCGgOJhjHx
OPo1/IqAUPoO6EbRCZdB7l8oz1OTih/FpNqQ4vl2dYD8sd6pRA5R1615qomOIlXV66VCGm5gEHGH
Lwe9w1sgBqdPh8HFg9ZLwHRzXwFWrjiVwdB/FJDkXtEIvXkhggvzHWJ0zTehPaQv6NUB/Ix/WIgZ
lSPPoSXxpPX//pI2Ajuv3Guwf6+xWRvRBgE4tKLm0cp6/I+Yk2uuZVfIuPirC0It+wovUS0KotgO
+E0ZFoCgsjTxO7rTqFn69RZy5J19D+wfd/F0po5WhIL3i1Ith1Hr47I+tjCbv/ktaWk7h12BkXrm
jP0VSGy3njKOnXiYA38yRWwYkzZ1kBZC8iCiKKVoQCqD3hCnHP72YmAQI0pH6bGlvvVi09GdCZ6w
l99zfUICO8E1zzpSp/nAaUCWvlKmiU+gIKTLB89EsSKgBf/iA9EnaxRUSbZPWUSx+9veQBW8cE71
bqw5RDtzuzmkfEx3GqYvkNGiyOEYvhQZgoY9ujO2W0c3LyNJvanQAr1LSe/+z4Mf4tteDlVQ3FJl
B8g8NNlukEQKv+s1v6HJzX4srmbQKN9WrEse724itiF4Esx8vtWtSYf5MGX/tjn3hUWpQZKku9V7
qWE3+CL/yk09tkhIkFFlUaFyHrcKFtiBZaEIS5GT7GY4eQbrZ08mY9t/l3B0923AU4vgxiV+bqKL
2eB5caKml9TF/5UluknwBrNvS4UKNoo2Q7DcQ40EVQr+sXsSr3MOEcpuZn3CW1Eq2sT/zztalvmw
SY03SJuof21P52REV0y0CVPMpwWhMulH6D4VOqYV5mIf1j+PyMrMHuxhHhukxMK7VaaIRdwJDRoc
5yHlHZJQdxTAd1C9WqSSYMd/CvPGaZdwx5q9LrD4dq8huyKiK0J2yEa62tH4XRhNoLHiewXKT3Uf
RBATT+fAjWZE2sy26xnaW7bKOp0QdE8/8nbZo67JM+QSGwFbYUNHqFavqdWsto0XCEEWxou3NDHf
14y6kPz+bW8Iko3FZNQs/5PtP5SiFfz7Xlbq1mkJSfVQfr5mQu0LmhRPueiXJWPzt6h8hQq0X4Mw
dJipKbSleaJGkXyczZF8vd269DGQkcf8hzdKEnFv54ArbEnE61493Og2GWJZRbjK6zXU9fZKtCG6
77opF02zAlGyQyxe5dARTaPo9ROJxcs5g+dfZgHWqX4fkWwa/WNdrRslutvXxxB0xfxotsM0zr1V
J6GpXLiQLRNXBUTaes4/Fm0kHPNpY4r8t/38rQ7tJ3F76ccGUAhE8/HypNRmPzYI/1oBMJiGwHQX
NnWiOnzmtEo98hvWfVG4iXgpZssBuT5hPwcyXgpWAeFbMWtdzG9eMpA6z6tZs9GV4NYKLbnN2emw
quWL8vrzLbTH9Glo3MYUBI7j/vOezPG4M/rSatEEUY4tW+7w1tPsT8Pz3eAAXmXDG2rmW9yQ6EQX
Gi4AEhRY+RtdfuLKhUNUXSgGOXpGMZ8GYQsYmpfJWwzukbm/vrXLSNS24FT9m3ZndEJFuS8ynCfg
WTJ4PDajDKZYKbfVzGNA2bun/fZ25MhT3VFl5gwV2ANAHs6UejIvLtuQhur1lRYBihEgARdAJPER
1aT4iuNM3I6PNEwysFwmu/Odb2GRxeAD1XnbosDSSCxLLhMdcWAE5q6AtyAo00fqAzpSTTUqZfGt
cd/AQvWFpoUchf6CBQWkOXZJ+2BgnWZzu0xcrUjk7MHAMDu20QyVtK+VuceTWa9cdDWEraeiN7Ny
0vaPAMBiTHJ/xeBdWsIcmknkZqJfZWG3WDOgLc6+2fLWigolcnQurR16TquqbB46ZyNC892eh4zv
9t68VzkD0ANOG6yJdsxZk2zuv8hTdI4w9XAxWWiPRlQw6Y7SXjmsCbEn6tQHADM0N/wC2tQonpz5
PoxahDuO1dEmariDVdCFSeY10b2QAiqYgn+trFZ7Ai+DdXN/7AYFLEqpN5ob6o9oCz/v/PtGHMhv
beyJXTJIBo8xmY5u5lU9oiWCeIwtHSL98RNzQ3D1eUz6lljYkgOFtdsAby/wu/PfKIhVITIES1fm
7iJwD6dmRFKbeEGUzJzXRZvlWnEQtC6dAN+azx1uyutcQYnqamcIRrKEfp8m5P+Ey/tazxPmnGch
8jYGuMdJrMzty502qccwKAY7Hq32rJFv8dEQ5YtO0d2jSf+eJJMY3kUD26duyxF7vNG5+tIeXaid
+3GQlM8pAxVtJYBAP03lTC+8UVjdP/LfdKUFPp0qzXT3Xfcxf+zllalYNk8/lDnecXoU2oU28e8k
q7tZOm+on+3Y5PiDKBd/iXt0M9hCRirUqpsmulw8Z8WC1gqH61pRAnOh+IsP1N8f698JD3BzG9Ht
LHOzJsM5Y7pFczxnNfD1OKfOMbma3zoSEJ2Ho7IZxTKrnEdYo5VMOlnYzJ70CY9Lbr0/uM34gAqZ
S+nVw9TTN0QUVT8uHd1bpYqp5SQ1JW/xQXSDyYoFE1fOzde5PPRI3/MiuNio6IslQuh3ircM5oQs
ZjoWjDtmgy86t994gA6R7bR46miYzBVc5JSGzYQQNMrmOOTa+LTfeU7gnbwkI1ULnKXZEGRPtCZ/
6Yob94jgEsX4T+L+yZn09Jm7euq9t1Nqegf3aTrUaaiNGIkIxcldsj50EKPr3ARnxiDAdRq5UXMO
UvzUyz5wiFQRDSc9iMnoaSVYiMiT3ZabU5J87p9gQKGLQ1LGkxjzkhKNk3wKwELTVpBvftUT7byM
2CS2VPqvTOG7G3GMJji4xRwUBR8cum2ispRcbvkN1XrhJgPjGIvPdmYs0I9aoZh6/+eadw8Gs0p1
HC5AmtSf23XMWzo/D1xadJACVNqP35G+NEqVVFn+MgQDLHc62iBTPTBzWE4X0soYUmXP9/1lM0ul
OyS7twAEjY6qtTeVDsCS4Onk+7fgVep+jSkpqmfk8yDTGmDMz4jFRe3Uh33Xlfzh1+odkvXZMRRC
Ea2Lfa6lwyWVJjIgOVkRUgG9By3trNMpP/VW8K69UU3BfpPF8q9A2G+xFQTEFFAVAGMW8hV0bdge
RbaRSLo/Pa9wOeTDeQo12eFwQ37YH2q1SlrccN8yUSIM9c68UM8wCezkLTOiGeElle/5TFOkl37K
ZJeSwMAE72I02psSph0ZYBMXCmVOWoV3B5YU8QhkvmEwtPZy0cnjKUkfnw2TLXfO8JfvUftgxYrR
X0I3gk0W2sWcoF8F8/NmDLLJG2+3rDgK0Ex89DCuhGLlk3qn5BdQNhHgJG1v161VP9wcuZ6/C/Hn
+4UZdU2q5W/RMLQ7mK6UJPa2/CwWIMXgBiqhSq3qguM4mSf2V82hI4UUQiFsJ0ZUXc1fKylv2zZl
9QnTvR4IdvdNKeUhMPOa/NaayhdYirMy7jRrHfWZou2bLWlDDGM33jWmCFpfm+tBzzPZB/7cX8Py
ldoY5yhAdwaxUz6S20biO9ZnPSp1pGrmSv7aSHDNrapG5vbi3ecfcxeQ+uQcnFm/I8Qhomg0zrrE
5WUBQ2no2/VozNOKxdnfOENEZrdxHb6sjzzmFXHFzzFNldfmZvDcwG4GcV61HhgIke+WKnADJAFn
JVf++OOiNOFDzCqQNb3PySFIa8pp8g9YjHi8n2QXuCVbEEaeYhUgSog7T3XNXv1xIxE1TnM+7Oee
UXJqBysjbqqABooSxhzrR0jF/wTDPIElTUSK8KqUSjNkGkA/pmA/KDq9x9XT2XsSxizmTIqblj5i
ckH842d7GqFPRZd1RdMgrvvgaO/SInEexyxxXQiozYWVS8gETrsz3qqWemJ67KSn7XcGkDck6TTg
dcyDmYUH7OQwHVHBquX5981u/Sp+fIuDYUDmzml4jD0OUVzEoS3sWOgYAdheRrKEK2VS6EJFC4Xj
30YHSCTuYsQ+07PXeX1TCI032ZoHBvJ7xgnA10347ZZKAFMyLqxN19uTzVKFy6W0uFOsmXLwmYVz
4l3KkDqUMWUGc6Qtxh3kAj7mgwC4D03bXXz/+y80jEaw9lDzNBtia+nKfQtPlIneKJ+spHdx/Cy2
HY/QZwfUh0IaRbyLGVaRJCjUXcMpv+IPYZL/Gf2xZhR8i+3vcD0KEjLCTY3u2f/On9PcRvo/qA13
qhAq2Kqbmsy771cE02P+wxVYxaxoREz25ejD0MYBPYk6VxABXwp7rFuSnb9KJoLBUC3MgZocpSHV
tnhER7thWA5yLr9JvQAWCsOlbOmBWyY1ECRMZDqgGKkuG7I31wQjnWNLyCozSf0ILnNamms0FS9j
O0BphwZxDdhVJg1Fcevi80xsxK/b68R/Ah8vax7HNX1d9z2VStwWCSy+1spl28u7DrCFPcyebiCv
t4LCknE6VjQVQqwCCASlcFSBAdtx3l71oIYp30PHB27vaYw8FNPuqiTRLa+uAnZgc9U76b5V6old
dIuctvmgnc448WBcNjACFlazM9qIWKlrzgS2EUk4h9+TQfKkdtecZqB6F/ZZSpqtqr/VQITWC/5M
o67v4kJKviSnLwhTcqP6or8N4VKMzjeHc4CORChbha1mBE1XIllZzoRNb1rk2Ksm9kH4Jr1XkOAn
S0Wk+XqmVux0CwUhvMu0HtizOjcB9kQ4qCheWVAdK8ttHSvM+pd5nty7wZoVozcx2jJ8gZ7Sj+K8
ivR3qFMQblRjj45JdZ7t7tct0iTRyVtVWNPUkbMq0zMW6e/HpPO4h40p4+YYf4UhQAuzrzG0j9ey
WZcW51Cgfb/Pad1rOGmRDuNIMKeU5zglveipK+a3xYUWSwk8GMLlo/hjDyKkpeKJoqjoTzAwNdlm
pO3/t/JB32rBvJDQlB5dU/EXgLpixMTo7Yx1Afi4pm4akU0a6bbyEcak4s/2D8gslDaIuQrLaM6g
xzTJlaJFRbIMUFrz24GmLOKL6C8HRyhzjvSRhVNZC5rR8wBaY4j9GqMR7vsnDECCXUpnwafjs7EI
/bWHbzUkkItoCFU8OecqtpPQyblGCp937tm2C4m80OfPEEstjbApP1Q/5zLVQmeb/Bw9DyNqK9cG
xrBqa7B9V+u4tY4kzMxqA75Qu8mJlNSIqDOw0xQPtBq//HU1+71unwgRu6VlOxz2zFPlxAyTOfvk
WsYyalRdhENoyklRO6qSzo5JNEMuil4fx2L/Z4+xUiBPlnbb9dO5mpDpD63v/LLYWyVBqm2EsVan
HykCIUPFIMkU8xbKGQIVU947n0+5eAzks5JFr5b+4Kpl9v3LnxdxzD9sGH6MlJ3arSFspUNJ8un4
/4JPU4HomQZ1lWKdiTfID50AlVlrffF4ZENGID9DPU4mFb7BtPSGs+tkMlDSdbmLHjopwY3kvLev
wCLjy2OWwpdJYPEwX0M8h6iOe0GBbXvXikkHRh4uAzYzbH4K8XYOZ1kxYuSXt8sE7NmOUD+LEAFD
qu+4vByn6yzV6vvG6IPnltXqahlly8OD7XGiEy2AOXMfcaBEVMgjozWleBUC4fM650m9XAwV1+wK
64Qjx0uTRrNd4cY5PbAxJJ2jGl5o0vw9wd3qJNrg32oBq3urOVhyxZvxCxKHlLxbyUf5jIgg+MUI
LuDd8xiiHfOSdytFCeBl2/pbBipewm/H1xJGjnrlrkjTyl9JedBAiMZ4hSejN8dibbrGAggqqw5/
t6k/xnfBBJTqcxRGS547j8h88s1ERWaWOKsd9vyUSCIfGABM/xEfwWUJdxQj8/BqCWueLHRoI3qA
FwcnesIH+Appcsc6dD0h6Gyi6aRkXXiZo32BYnLXXfmPgccTSTL9PKj19oOmfPFxa2xO07C6g5Mo
hfbsBsBVfd/xoMhRBUEQh6N2whSuFNGGSzULJOG8TgZ5EzKXfkOEoCO3fG/M6tm01Omh5p1mLExK
ZwwMycmAGYfGrSL/8F6VHwh4j/xHh+lmnl3ceKibbGy/W8bwRb1kCJUyt1//iGI6yCqKlkobtmay
6dAYKp+dgdFUbddHvjo1KbbbQxCaV35tw9q3JgNj5JOMlAi6dRmPvWgcfxy3qVRGQn0U5HDkKprP
v64GYMqmUig2KK/AwyEFUHFOwO3/LPg1ZyuLBB/sqqDgo+7/xLZnE8qCjiHxX4DJzfQuiIDkvhcM
UzmMoZiLGjQuSiQb2guvjD+bWvehk7Mli2vQnX6zOi+GMZQ0AEkJVgfw3OBZb/Jbkpe6MXEPXHv4
A6/PPkRAmyqb2MvgAR1Eit2dbKWMEea/IwreSJR38I7q5FjXsN5kA1zB8e11l++36U+M1vAXaugL
NXpFV5JSF6L1lEVP/ABXEBLVOy2R7Py77yq10NI535Jn34U7BGMseo9XZDkrChj9HucLrYdQxopG
WbcYO7TMRromANvynYh2ccgmHRDpXqpBuJBK4figczuLdcy0r7uhHZrS43v3g/gYC4naGz1khLZn
pNkTF/l1e1039MjfqjiN9VuGtu9LI54KrMkrotCNe7gF6qtM1e1U73U7v9hVHd/ytiDsizR2S5Zq
sOrfKAjHxIeUyOyB9j7mzS3XYy2oGJSiyvxdEo4/fVpKtgxmYcSHuRL4VlRUpFkTJnAG43ScyfDH
qRL7QJgfbZQyPsqMLUQm+2QKjZJP0I3Zj0IM1JrvqJt4asksnIHJXob+0WaIP7eLYCBXYd1prU6c
b/r9MGuwmysLC+n3/ERGx2P78Na+RFkI0ZuU3FQ/yVMXq3XiJgBvueyRr6CRcQxBHgCCRsG9kEWO
6ZkX8bBLVu4xXlzOrGrHFnBxvxSsWkwD6aPHM4hR0/sY7bYXTdI1FpKw8RueVOlmx2iLQ1q3xbKI
ZFPpqPT6g2vd+gjOTH+WjCrfHclooohHr4os9YQzOEgzfHXhfJo9TSsCrTf76paXSg9t/l5HJFOl
YGrnauP+P+lvfgJV6gILiHJErrRiKDwMwzu3BJV5AQSyy2R6D2Zmt+qiPiRxooED4vYss8o6fWkS
J81PNzFyNF5DlMXh+CvohtvCvkFviAUcJLdpyh3IpIOWhXk4k44dxytnS+ETYHrysIK4zIyEIq7c
RiNzeYZpDtc+kZ5Lttuaz5pO6pa4emJ2nUma36yq3+EfmGyxs5EIK/flcPndltI+Oosoz8gcJVJr
P4pYPlG91RAdYnjtRkjY8/lt9/AAE21JppnnHpX2R8xGe1o9bsHmwYFJDRF44Ijq2njAeoqJQa0Y
8s2x2fdzHLMQBf0umkStx1ty+mQaTQYF3E6KpH9bD/bU6KuHv9CyVBY5gl8LqDewjzR4EDCzUjwG
X4U8NESMHIYeSNInLJmOCtbrxCjifpjpSw9IFtganAp6qUDOJc2DrABaXyuyjhVZCuN/N0TbE8Mv
+cYhKDOHzBB0Ru2wmNRuQ6XWUEANmiXvgwet6IDkXKnJIbaksWVkqjCjYwYJLJ+nLKFaaCGutS3c
SSNchObkfy6Yvs9wLNk9aFJ4MvcJEyc04KPooefkQQ+Dh49dMkmCVGhNh8jIwa2zgWSumGIaEqe5
h00y8Jb5lxbMWtoNDsSkU+n2kVesB6RZ7O+aku3h3QFIo4CBnbETjlvdcUuB7TAw0U0RrvKx825W
x2tIuPLKNR/Lvihod8XAn3cIUism79S0Rxupv8xBCzgIbX2uCM9DxFb24eg3/OvLz8QusJYEx0qT
vdfxIG+d7Dj91bBjR0wGdkqhw666C7pbUoOfBDAhMgM76IsyrV65/NUx1ICuL6YW3EreJfM4FqLY
LscAB6nZIBu43+ItRkdeRFV1f+2D3+NcapNvSxbzGeWxL1bwRckBIyEwAuSBEyEeZmckUBsT0aTZ
lKjdyFJl6vwVLKBs9HCZTRYv2GZzQ7+icV6PT+mD7jvXxt0cxzAaFJJv/g97gPycNNa9x/AHakxn
OKrY0JbiWozE/stoBtWwLTSHzT2neBrKzns8KYNJMw0b3wyH5I8XdhZhuJPd4aUeg0Cj4k01j6d1
BZFuuSRzUrCnV/plx2RQwFCSHGh8cthaWkCU3auBqAmvUOUqBWiMQ1U6TVAeG8xmb6NoabhYpQP4
G02rzr50sbfhlhmijfBm50FU7alO5pFTFh4oV+BL0gDCDNinKuesR1eu7DZjJBN+P8pe/7+AoFh1
WFLJw4a0gOt0vK6x1zYg8Gn20O5AbSP+jGV4QxeoS4R3mZCPw9j+PhEtTIPorObhQN1DoTLXYOM7
Fx4mWizF/HkPYrP3IdefNhdk0NeipaVXupzAvCOtFwPUSpG4si3dZppXNSN5SJtW1IJCVLRDe4zT
tJ3f/YgCSMW0PyTvLQp7rYKVwXw0hVbKwK/nam6044gpGOQZKzcy1ek0hKxcB105y5ZNXfz8C/nJ
XtEgY3AxE8ZWF0HcSo+x9Xhjfkywk2eN3wFHFiur19F58dve0B+PajEtvi1Xw4pFzwAkbUbQJHC1
2lHT6+YZAEJaWY9wp7taoAB8So3JGqRwRYOP6lqNA5D55xJfByaObr7VuXRERtn9sLqDAcTsky68
AdlJ2YcMtV3d7eF5k7sTNnyv/GL2pBtwPFF5kFLcgvsGNkRr1w+rRpdDygnW8KvXeTo0/0uHiDdc
V7o6kYjE6FY5Co98ummN/z0wMHbvR4ytVr/4/RkAGhDH677lzb47VZzNYR+NCf8CMh8Ljp2xlSRo
0i9pfz+K0eiCjSrEuyxMzX68UL/F0SO7iV0iejS0b0a0pIHiz3MvrG7lmQX9Bjm6nB5ZnuU0AgOn
WvPNizHB2dvzKgbSNHNdhB128bMp7TX3J5ymJD6zdAunBkLIGt6FIUGWDyIavqJZM49mCdGLKMV7
1bVaOOAY5/rIO2mO+yK3UFjrpn5JiCPfMSI0ypVnGzxShfN1aI5jeGiDURifb513tSWB2YXFZEDV
IDK93zIOf6u5h0wNVvxtl0Xf816+SWXmCC6BzUGZjIVUG9orFrMz23RUpcjCZnz+lGLTT65aGUPj
7j74zO/6sjvOuC9b+QNogI55Qk8ugKN8q7Yv7RXidBbGivq8OKa0bNEqqWMMUFS7WJAqlU95pjFq
hYn44bg6htW6+DjqX0Baz5rqVEmrpIdoq+SmKwOOXFJRIz33qS+7LHLugZ8N7iincsPb0GN8rnQW
6chLbcbQlXzusR0FGaWN7qr5vpPZvABgLug4L13f9yUXcd7V564XA251NeZJQnPxtGg6FfFlnqVm
Kkj2wsMuYAONf080Bpgla3WFMDWIEyl8SD8kAXQHEHX9WUEtiaoHCVzgRgMfbHr5EUH3gIUVMUWk
jaM6k4GnYcSzE4daHV2uxBBD1zI4iuwC+IoVooBhj+MJhM+Tl+ZsfdxKHvGl3jJU3qHfGRToVT/Z
boymolwZnGADYy53sqxvYDvB5H+V2AVOjRW1NiXj+MVQsw1FbAPT1mLhv9a1epeSvG13/79TYTFl
pG9mZ9bulRgECvPI9FEbca+ZjaW0CllGymnYFw0H4gXlYvSJF1KboUFLUa/vABAiJeVs9GmiKTSH
3uSE0OmaEXNVl0tfn9Lp7mbUcp8hXxrEIan0dPGOzhwl8XSunkK2CkozcoGgxatvEDb09AE1FulS
674rQDK0vLH29rc4nI3xFWZSNAfZQ9ywQNJfr63r4L7xg/Xci2dN1IBAVzeW7DlwaeDtmwuqBPsd
JZAnB+Zoi5wnY0qRxcqYKL0WfqbKVucy4Xs6wuDon56cuZDYVkvZakc45zaK5iFH8Y4q9IVj9KmL
0Ji7PcwblpQFyVD7Pe8t4FQhmiiklhEUMEGMsN7J+BWLmkMDVjAcfZGQYoDC8LKIzWalHt6dEAn9
IKSZ9AETdCJjxCg97979fmAp/NE0KYQQmOxKTGjObiUsdGUuE6KkNglwz3tKQq5C66DN091zYT7R
JRB2dQiieIPyR30rfzfCSSdGYMQ1Z79/ujX8NZBbGRuvPBV/rhdlroIpH7OVVn5Z63t1CIi0ALkb
nbL2B4kx4DyzAXbGjPN35HrN6d1pWaT8WsPUt/fnDniDWfkePOLAwXdYoeMGeEbvVvsrjdUfV9rh
ET0mqJZ5OYmWoQwvd3VIoHe0+WcCnjIQYPT9k+JjrQRitytfABCWkzhGx1uGMqxlP5J9WP3xXSGP
kGU9qOW0ONxqKfHX5o33/iZ2R2NYrG/SJ3TZm+onqSCQuBpYcobrNBBLc605OGePDvnlhEpRTp4S
S/q4IY2LqPsqcJTcpV2rCxmzELoMIFoW0iugaGPhCpneYkXh7PRC5sCaAk5F28edm7y/lOb/0fqr
EP86ISU9mZ+AHCEBo0ZVPRICSyVgqCIWjWFbMM0zlOO57uIC+9IBJzSCCHIGkQrfPoGS8fy1XgdS
RRKVwv+r3lL8rP/zpiyNIk5nQ+ZQShwnLeN/x9RGDdWp51Vk8uBZrqzPLIO6Ak3regyCxEWartlz
Q/f3ybZ6IFbIXhJ3XsFr7vrqxC2kzda9K4zTbT+TcU9O4UghnFRXqrRtiiU+6FbFdBo6XpClB3Yr
UuVjGIJpoHyy4EUKd4L9uNVYJK4RJ9HdpayyydsQg6JX47XFVVuiHmxaEqu6VcbL0236uZB8zWV6
f2f9IWIjUBiXMjXVXWBA6WVOOc0NQh6tpQuIl5PvRDhQy3FDCSDdOdQANapAWQOX4rk+KYOqRpag
8shRZUMjFSiGDQa+CeCF+yw5rfM+R2HYtobJ+m0n8YTlSZNcL2NXY7rONTMTJ/kwPNqgP4vzSe2F
S6eOyw2aQg6wZV27DWdmEb5fNlc4uGqh8xRImDGKr/yWmq9oD8R3yzwVWJVLKDuaqHC7eJ1WelBc
CmBM7UvqGUy59TVAnO9QFNiZ+TY7T6bUkFWdkhTDkRMErtRb5VHarW/AqjNucQPYvpkTV0MmaOlY
ObVyc2CcYW0SXqBQOB8gWgF76zmfANQhB1Z22A+VLqDc2E7lndduDqwd6WEptemVIaK+SbfhUAPA
0QpU3jrdYDZMz3PUKXGj9LtBrpkamz3kTuIyPTMfiAoLZup7U+sRLMdH9YrFuDzYkQcWaxzZV+82
ZenmtoTBqViQHjAtTFI0SMSG4BeXlRHRLP+oZz/m1SWr/xr9/nw7Xdhd7lvAgIfGxEbunE1SfLgB
jaZuwHtay8sduukvYTCA8ZzPLfpems5TSV/GZ33TEIzc26ze/TqPXSnboEhFdVwZn69MFDVg8Ri7
krol/+eOj50BdwAc92nAKffMoc4k3cONx8izXvnuuAED27KRcw7xM/aEdMTbep4S7zbvbakOhQXn
NNGXoelVN4nnBxXObtw2rsTBy553Rca+pt4KuqdeykCKil0S5BbCVB6Km/M1w22YiJ2/O04XHS+F
T5ddKRWGJLM0uYT1d9rgxsKC12PsvJpnVhY2nvOJt76+H9skuVCFa/fp5wzk4zzgBg3ZKJmiH9Od
Px+7zjL3jkY66eQTleuDURbef8K8iwfw9jqsj2qPxvt2p0DFqbN5MZG5ISXTZhSMbbYOcIJuwLR8
ZT4srbh+Mswah1Xc/5iFs7o/EzT++INglothIHNE7Gb3szerekCD3eOWTrsVGn50dYm9q14pNksi
Al3r3aOcxx5uCEc5oS3dNTOnvQq016rpA5pKv/2ACUmIp1KJ9Nye8ohpsm/RkQR74/e2msgIg9Mb
q/k7eQh6poiFrCnkfXao/2GnR7xj++HQIjUI/8HMdFUSW8yk5zrCf33g5YslwAL4yolhuol5IgpB
z4X0jadJzcQMnGWRx+KX/lxSMBVV0BXm5BCL3UGq4OJhYDYZhIjEbk2JSYyCOGi6TzM0DK6BX0H6
J7y3kKK6UI8mOONQaR8dgIlxQ58HS8JkDTJMBWB8my25V+HkQFO9h5K69yJfW6OEpslEHC2kWhiL
lVRf82Ze6PkEr3j/6mLQ6+5lqJ3rKxulkTnbB4mQPE0djvnUHAQ9CG4Omm97O0vtOG6hNV+LhhMl
Q+tZnMKbECi3BCHJeRKsMjBUo9U4h5zHkIy+3oJBQ0gIoWmuemlkFcVjz9/FzjSy8ESxG4qg2zFf
+EAJjbRu/8SdlbDquAo3BKQ0rWx3VxjwPdLCDT4xF3JfGQ0HxivHMApgeAl2EJsYS1mwYwayK+IV
veW/x57GCTVID4+TTMpmT/V+bDx3Ui+qw+GVki7dckpbKEcSYo1rTojsPes2I2bG/CZYNAdjmCWw
GywweaGIMkESQYaHATvnZP5oAXObj4BsRgTivR+SHsDjArp1DODqYuvtH7mRkG9Mb+u0sVfCkdQk
AjKbuoQm/MGozUSKL7PlqwuBLaZAYBiq9mXbaZeeWX1fEc32hxfhQrPlMfSmTNCSUIM1YkGJ7waP
p+nyPO9LZJB0tjYILOVcdcPCdaE7lPDHo6bth7gE9yFqpWdHL1FgHCT9bbW3bJdSk5CjwyVAxdeJ
NdBCol7/AUJBUaLScixhmuzDrusr0NmbXir6kJMMGtKxMUj1MQ15VQqPZXnN0D2ScutFFVRGnD7J
PPE5/JI5nT8E9S4bVwHvn2kPntMrxekfYVbgpyjzBywNatpXF7tsPa492pvN2yy1Lc6em4Mw5F32
527YLQxxkArrQyBkn3LRHm5HTSIO09r43+oMqBefNsGb/pMsXH3JuKKQdv85/P7Uh/qMJK/OC1yh
6t/65EOl1DpHZm0KVHruGyCUl2N7UIa//i8wahcUaC6Cpku4QJSG9KWQ58U/6qJW3QDxUISR04kX
Lr0JIsvmfr/QT8om7ZbEP+rEX3ju1r+IaWbsWPjpYIfqAh8qs4vDD7YBWn585WcMYZW6Ynw7OkdI
UvR0gPSMU5d/MnC1LjOg4lQ4IJ2IuGPu68FGFhTL7Z1/m1A4YPHKS6LyPy2zgAflHGjn8jY+TgXJ
DtxZ7FQP5aRU9ygL7b5Ht/RtyAq3s7eo+aUCS5pDBBsT0nEiOGYrolb3Qv4TsxelrM4Z00HYd3v6
XNAhkIB5LvC6y0XKQWtwifPuqhUN9uxhIoM4pW0AZOQ8B4ww8TYQMGBEgn1mPzIOA++O08TFC0dT
WBOdNCbwKo+3Ryzl4L6P1f94ZI++BBU7Kd/7Ax1GNlmXHhLIbD6MoZf2+xacDHuDpzh/w0LzMiQn
5v/wpDv+F5MrI6wewM7CAa3HdWBuKd/r4DOrdzMElcWZ1nsO2DfzBueSzJPFbPdngBof1M+ekCP+
6xIGeQ3sx8FSyFnizB9tbMZe0A7BLZFe5YK7jcAgo84YOwpCTTjjHkU8qV5E3WOK3+j2PNs7WN+y
Nnd8gV8o/KEbR74Z+zs1fbQ9i6PwCkhiipTlCT1X79asAlGnkU/OncBKhR97mOVsSwzZvUyF+NBT
bMhbO2UMi82Cy40wb4Ln1c8tS4x0PUjSfI1VHKPmcV+DTVkIukmvhBYWliYv5K0fEVfhppXy34f9
SAbnnyNcnfU28tbYSeINhM3s1C3kQout/Nev0WYojZX9JO/UbUvEZKa+WSEWl0qH9i3iP6KKM4Ik
DYK1c0Gf34TDFR6pXYkNz9fqiKk7sag4v7ncXEW+ULrhpzCX1m9BwToHw6W1WjagE/C8XnIfK+dp
jfn0jzCtCDoei2VPHi4sfSi+hr6X8Wf9/JmjwVDw9s1tqaAfkNn6cXrurslmtAHfXU5FLVdMYOr4
XGXBzUURzko14r3ny9kDzbcO7jfK4RAWaMwl53iId3ih5zY2zN38jalPlyHs89QNsm6YPPfY36v7
W+Q8Kkixz6uoRL9C1Wx12aJlaicBgRK84P5+K2B3Ir4HjBdDbCVjwgqm7GlZuB30i0DIEhT4ppc/
0aD8sh6gp5GqqE4obEmxxmWOcnlb++35JscTBMIabdIOuOfIMg5+5MfZUIEueR//5ohKBVLmCIUl
V71JoESFC9pvxLrhcNaydQnT7+we+g8twwuxnjXQ3OlDtJp6rM8GMImee6xQXtAl7sN682LkGAlh
YHgXEuQC6kCG78/iIwKQ2nXgrpty040fWjo/kxvAuGw05D8sK1iNCpNrUWUSXyp9hluRkpoyjuBJ
E3pLQOAGn8Xfyq+bQWgxPuojQybpwSlXCIDZpEFCnzLQohFhJtY4YaoxJvrHsbZO1WpxqjZEg7jv
GuRQkzxKWiOzc1KqLt64zNRyIoTaRRiLTZQmzsfB6PEFC4eRVT2cuHVlsGqzHAuF2fymO0eZLR2F
8gSAERTUuvPsdgFsFttBQPf0oMW05nMjcJJk/ieDX3TFiWNCld+DDe0Khtnne3cfsOMM8PSWNOul
mvtAfo3YMw2ufwYdkU+y4K/Xh1WhmTmLjqHnxq9VE4XLQUWbpbys511wxcNoxSiiSsvMk65sdb0w
R0lHFbmH+7XHGj4qilkAfaOKwOcY9ZyacQXbJpKqJQh+/agp7VaVy8ik1o+8aZn12kSc3/1XTc/1
4PHfqIs4pa+jYr95g8lPbYVGU5xKABe/DlxUPdvzkXaAVy7Ys/J0/COkVQbcfhkp4FYTY5oLiNG0
Ys95bB3q4QfAZJjg3K58lt1PBZ76UgrZzv8g9r0U18iI9JhMkFJRCW0PUfmS3dY22l6Z+YuVIvMq
al6KWymKN5pb69JQyW+gWvIQUCNkAwlyQ44NahfDWDvXFnZdJZcMtlBS1czNw5jvWE4pARpym9fd
D2llqogXKJxuFdbGJx76OgqDYwAHhYeKH+rUfjhcjIISJ/XOPWXeQ62HAbg2V40hzHkb852bg1k2
fWsB4evP1cKHW+Lj3ZDGJkl8L5hsXqbfpRtLlkWBOVLSb3kdi7sBnIofiCMe+QruaRoeU2JGg1Qc
tU56/gsK1fJ3S1/EPmrp9x717lpctAqIz9ToQvvMC3TuTdEE6DvPq5Y6FD//lGZmwvY5pThmcDiO
h4zfl6IdRMubiE7Q3m4NAJNXKRtfDkDml4ROoSxNGZVxfjTXpQsKq85hhTJaExqDEAkqO0I/5KDH
rfBz+g4zblBgpG9rlIoK+MuHV7sBGvuCN9hfk1tCEGAFm03hxth0vi+O76ZP/WfP3xCeKmeEBGjk
0dK3w9UTuGUH0/MfpqR4C6l5DIO+kKGJyshs6JaoaYZA8q71vZ+hgdkPzoMkDo4uPKd8SUVan5++
QpMqedDHsmx+S1vbozRMkbcXM4XuVPOnj+Xt13OgW5SjdLMEYPTOgyYSeLQm9twB1tOYIkMskDF8
4nbNhohz0fOnjvwrPGuMmpZMp6qlEbEG1q5Kc1gMv9/dYIgTx/3DPFbL+H+BIhXnZyZmLiDj+Qwd
CKI8SjH36u8FgQEm3NKoRX4gJWNrNvr0kT3XYFPmd9fUEbLOx3Ksu7E4yehiwu4uhQxEi3GpNOsi
bIF5Ns9ivGwnDSxIyBLcPY6fMLL5ZPFpSicjQBMPl7CCOlg/9q+pb33zamuxMsligCUsnq1FI2/w
yVkMntQElWeFxRrIXMPVerUZZNCCnosvmlpB6Rxg4cUEPaRnIko47m7VWf1CcHaR/KyLOKCfQnFi
UlahMNjbZo+12Xg+3HMG3GqtjlPNNlYdzCsSW+mTTa0uonLbEI2mCFSWn0NFfeKrVqrzx0qWLc9m
CRbL25v4AZbWXdR/PfdNw3Dj9NLKV6CzA2xSiYjYzaB09MRXOnUrF/PN9bP/5/IWh4qkqAFA8+no
VLglT0bZmFltd1W/cwvOHO7T2oxaWK35CXOPTn4RnIzV0vmsEkOLifksxKPFV2Dk+QCG73dKhgKF
mlCVEUoRHGX9aMSZFjOIl/rldwj2j6A+lJV6ldXf/hXsNya2kRFFHmyYILg/jrmIzpfADddWI/V2
s4XA+ABFvJUIE5IiWh0e/Mpk6obEzilAB7LiX7B5X0uZuzV8aRJw+3jIl8p5UiVxPtsqLFlgkUmx
6GRNEOZ97GU/wKnlyGXiwomyGpVkoiUHwa7ey3oHrZEXcXx8Ks875xnWNSNr
`protect end_protected
