`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nCvZTB6v6PTjPS0o+JcKDNAhBR8J5MXtZrwVnjz6aVUHiESzLvsz/MO3Vj1n5CWdMBmba5Vq2T8o
ecEWLFVYYg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fEepP/mLaLUAPmpxg08CO2fXfX3BpMKxupatPdTJFRP33reGY7q8putFqYyN0IGzjKbIaFz5Bk9T
6txdG8LggeRYG0RLCLWqVIrnST+yLGDDMCM20vwFcsLK+v5CipKSAb5Z1X6yr/upuusU60mUrEI+
GhOHzu/yCKzPGhWSK5M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TWogJ391sOUOiYPV8C0VmfH7Lt2OoFDB1ANIEqjQdK7RlTImx+9cfN0ASLrc1bgQO0Fa4GhJ8GaJ
kH5SNZ0UqTITV1dcoRqYnL2eco0e36ymxVIqXR9HugA4E4j6uLcwSCE6Cj1ehLRqf/ufvmn5X9VB
VSOceS41giDc1Mz7JeJ9o8uzSMDO3sl0O2bIwk8PUP32+Il2ZbMIvS9jX72s3mNc2texJHNnq0/U
bqSbDXjDFbqFiQSJDKYpLDZXVhCPDJY0HUvk88rfiZIqQoRkG6okTsYXNZNNjr5lHOAB6HzeIg/D
Wnsp2WsHWf71gIzfjdelQypdZ4NydJ0IEzLu8w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kcKntLIZHtCuGToIf0ZKpe2A5vIZ+qu+NfNs4HGHMxr2sSxeF7dOrX4CTntdzlZP8azlUvyxQTLS
Y9oKyb/Pj4M6IHUiOjIAdmmuUYFNhRjZ01bhok6rmcXtKaz2biqTfNOK6LSCBPUtWC2YbDC9rhu/
jvbe1v+EwAQpQpabsYo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LeMeViogrUwPr003VGu0u2/vn+NkJ8KNRR2p6ViPls/q5q1w9fjiAN//jia9+xH0QRZsrOxmE4sT
mlzIu2VTOCsqmeZE4bSH8wDv+4XUIN7PA7qBqC1jPZSpSYkaBRrvcqhhNBZrLe6EPInLYPGs4i+d
w+MKX2xWu/JSlJpPAv0YuJSExBDRHco8qjiE2kJNrBWRLc5i1BztcWTxQXcvt1S9sWNFIbU3A0br
4lBphESfaxDDWYrtvRe7MB5byApf968RkN0riH2z2os381wlDOaDZyzckOM3qQ+flbAhhKRCNRVO
dr9MaUYcdsLuLJS/f/jWAJI2hxcaGIkPqsE+5Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
tVAEmwHJpnjd605JiR6zjcv3ZfWzud8X2oLyUdK2qgwtT8zuKk18b7JorryLdsmJB8xtJ5YclsIW
b0SrJRTZOLMWx+oT3vpZfB1gw2a5koGeHVqwBc97WUfZEj8Mbs//ZiCohGsh50/KOWEtxLcJae2E
kuj80N/w2tMfWq/FmJ7S2B4IlUrwKorIcNgUs62j1x529o/Y0MtyiFUHUsFFzOPfMbf5On2jWp4Q
jT1kS3wYvvEUjZAzGONGG/yqfMbIsNIKGDz0By0UBi6ID5iSbgFP/BVnOxK65g9tJ0dvAphcI3QS
kHW0/kXS8S6hr15TelfZezfBenN8BcB0COpbKF7usOlWIp+JpfMN+r9gkndvcHkzcGKopDT7lH8o
udqgxJAFflHNJJSjz1I0lVkq4xJS0a5bvoZmuoLn5M/cgJhJjqTiLrC5tBhTwxRIixvL2qqAfcTX
njraBJh72F+Z1RvTJTYtG1OxBwNypO3EfHag4bOqJIMsnZGv25PH5vLwIu3lXZESL9unC0NvePpF
GtiDmBGZb0Tp3CccaF9zC3USZEv3/1+jyZ3vQcaZeQj4Tt8VZ60eCWyGuLAfTPir1QKl05XVXUNd
+Y23vCvyKPU/4aDuFShunt6kc9VixTifc8K+P8JN/4ef6JOFmVxELCNBXF63EA/spHgv9c10qixu
2qku+dGJBEygl4zDPvm0vDhdNXGbrjJ4/tzh+fT+HY7yEIZYUMAqE2W5C4P0GHoxhGxWC3qOG2tT
rilVIye/ZRZ8IcEvr2RZxAIba/VBFNYiQVoEdOj+BNVl9Vua7nFbWN+4nCtcAl7haimxP82m9rPl
nS1j2QaIn9JZcYZD8hMLp7sznuVKrLQR8VvlIn2eDo2a7yuLT9P94w4Hm/IKawjrqM7g1tIP9RHK
YoqDEEYx6rO5gav47ujLyaqEguqtyhvJH9k0ef88IvSx6AGBHFljd3uhan9AOQjmDGXRvLEFPbuf
+yzChMR3MuWbE+GiyTaHx1IetFMygz9uQ+nsUfZQ+i2KtJJGAGhVzYsvP6m6kPEsToHMisq+woef
c7lwiqDiqrafXLJwhLg7Lb+e3pF0HSUpHEnXZFNSR16hzbAiu8Bg/+XbMeh+yM5HQlbr1CgSmkIm
CjBO7zXiqxPxN6PhDz68rE/6ogu4fEkyThSeuq0pFRxFheXdDf7b9BChVDnBjBtJEklMOw6RP0Q4
hDO6E42gYIJbk+ooWRCWJ3+KGmVKsGNawRooHK468O0hX+mcbNsRh3vfb6w1szS2ERDvyHY/y/HB
2ssPbOqI+R72Ch6SU5+BOCOtNSs8TGomCe2ohFAdITi7rtDa8NZGcpdMNv8MYFvR9xXASyBeq+p+
EKFt0KbWDtgwjVMTaUHR8GfWPbPPvZ2liApFabJsdyOLwqmvCM4K5fCiYodSvKILxKIuKhIiVJOD
+U0HwtGRgTJISFm98egf2ZfNl93enI3MWWouCjr2bUIS0F7XfWQdQSuxsEZmP82I0nUXTOjy4+cE
nTyQGTbEz9uTBHUiMjWaz0FAYpEjjswZq2KWBKEM/Ls2RsSnOs3x/xfliAKjO2qOZYapSG7+OBbc
CS1rr7h6j2gBiCwAThNR73Lf5INjHK+gGbBJNgrSdmrug5djOdLsLXPZb5PC+Uix946//O6tmqBe
OKSqW73oXZHV5r+oDJJwluFr5CZJvPGveUc1Ib4oMvR6rkvTtS8mb0PNMZ9+IGndLbdX1zb4nXLX
1TQdUsXoIo+mr3aaJdFa0wm3WrYs2nVQwDEvTTt2CX7ZD0ANC8KrauwsKfnU08qPgRRmV35lcMcl
3VU+WUio3KzD8biBaskCkYPAjaR+8M13H6bFin61c624kxx39RupWZHnwh5O3oa+jFwOLKvB1nvV
rRhVHfL2C9jI9TI5hiyqYut6ONWXTFjTVpSpTYzoz8cJ+2zxfi/Vp5ihNe8AELTsXmRQ25x3k4mZ
W9TiA9kYiq4mJtnNerUAIa7/48t7hyi3b5w3ERo35a1/2HHUR1xlHqdrIQUzMXERJ2TI4IqgkwXc
5WCFsATnU9X4yUMBd0b6zDIxmXRJgxrsE3Jn7+yDa6zPV9ZkpY59TRYsrfRvffB0M7hWZmQeRy/6
cTdGoD9ij62jO7+Jr3KEYlv4eqAwptjHZ7mfG+9EuDf+ToMToK5t5ZxHyMFWtYaKfUVqtq90QWhq
5FE02kGq7UfAUcbnUJ4MiVQ0VNTL99VIsOrZQo1Cgrr0ClO8EENOqtVPZxs0qNYbNdYfwS4Gt+bX
q4tVR/TPbDfErF/AnhFfkje9sjo8+YYM1TyP7yLYKtnav+inV7l6YABpcN8Fyym3ihh1Z4fj3XMz
IAcnLEjkKeAbM8h7kxw1SylTvlskuimH6R7oUPgidNYF7tPntYb/qB/5qDmii6EOxftAspXx0uij
XPNz6VFMpkgzEH3lE1eBObRwl7ojbfb/nkd+16D7+J5lXbb0WkQ004fHGKFXEl9euh8N26wI5hyu
TFuUePmly1irvRiBzV2Aa21vEo2ggiEg+FAPqpkM+RYh+54H4nHfo3CoIgtWFzh5gzkwl6dWJGNU
mRZ7U64GKa2C94uP21Dpm9q0Ts92oNmnrfOFv5qbCT0hOxGxOZ0gr1ZJRCVK0ZRqUKu1kwIWBBUL
5IKOML/0qpmjfnFoivbnqMEJRS+41511NKLcB43QNjBdhFqOetM+p6+wczoeTc4NkItlBeaZZCNF
HqAYl4xUHBxJFONYD8h9p8/+4T674Ez1JG1KZHblNO7fwDqKpyoWAumL8V/J1xfytWw9jdEIQlWI
jDWuXjdBMlxUQ+id5Sx7QnhdTDkTNYzJ+HOh428ODC3qOC4a5Fe0ks8QAjaCUGRNt89UjKwNaCkh
2EPi6erLjKxFUsWMjPOJiV7iFBI3TvGm/RUYKpsRadk8eFkUeOfIxfFP3lGzuYVZl0r5GCRrEvid
MnZNqqqQ8eDHKqVV8x7CpKgeqyvIwkxb/U6bbIdIerj4a+T4JZx3FIPnXzKztXxuy53+emYbUKjf
tEpicAu7WkdNjqXxt5j4LP/tq6YhK2QnmL/Gqupe63P4sjsN8SyUvjdN0q+oy9s6ycAGPujQYS7S
YhkNtqPxBm5UUKK+r+M14YLIZLgnycTfuDEbEEXkMAmqApFjt+aRQTvqsZh3Hy0V/D4mDRE2LexM
9GMdTBhFdSvK+rTaW7pGpDdVa0yVtbLtwuuelFRYa3xGUgMLK4mL8tZZ9T/chEVCXyyXYinVeL2h
RQm6KTAjYgcbnLhP/jl5XhY3MycjrwKX1gtc0XgtMbnSegcGCf8lotaPEvFaTNwUXQ6ajxAuIXa5
/P4tElnJ9cc5Kkem5Z+aA2Z9UDbzsXVnhyCD70MQ//pHQNhi6OPauTtzweATKBWicSM0scAozNAA
xCgbJNF/9HphdcoRi02tej5Qkt+AY8IvaKDExZhYS12oMVJQpTID2O35BrkxfcJNOVzZmcAqzMMF
gTCpbjU+X2HSvmr0BQ7j7BmBby6fe19s1GYB7Sq06FkKvulhsLTbhlp+OnzyGkmHRVO4X42he3rE
V/rnWrQ2x2vHpu2PsqMaa19HaDf/rQ23r+iQjAU+Pl9VsPcU5ql2PCPb3WnmxFb6Bc7qajn+PwAr
x05093bJLFglIxrJBLRwIwhdHOixX90+ER0o1qn09sStXyD2DFUTwCcJgcOxtSfoX67irUzbwRVF
YaDieX9la37GMjtj0uPlOKEjTBBepCPuacFchSr4lP7s74+9G/4HBacm5jgnjF1JZpqWS2mqjcIM
52cz5wC6LrD4Xw0iYQhcqGP6Z79ap5rGCAtXK4Tw/x3AplDh1GQAiMZXQGxAEe3jVuoV3CjZ1R1c
HTZgbJcChBnYDDb9JmqdA4ZUFSKBOb8j6r9G5mr9bsbWd9n987T203Ij+d8DXZoekJ636KKuB4jv
SQWEAEDqUrig3HjOxBNKO1yspqE7yLs4WXwT/2YudIvsIvIc3tiuVN7Lj0F4qcAE8ngyUuCkkcat
UHuNsNQznBITyFW0vgo0IGp/Lp3Z5Bo8eoYKdCdhtUHMPmJgpO4LzrQMDMH/j8oDD5jDXjKeSu+N
zCtTQ8nH2ZDHwyVJMLdnb/dRhrXOqs3VnPXkvWbreY+tYlznkS4GHTC9/cg+3h3ma5aLult7jTxR
nmPv62y516+d1VcQcm74DFr3bpcUHrPvH5u1de8iU1VJ1hHmZo+9be74NAYXIoKMCZdaqZMSqeFM
LXLKwDItkrTRyhIb//eKWhCQIry9UPP0CekEWk/JT8J4Y1z2cAJ9vSKm2Tgdu+zAB/65/fuLSHK8
dZ+a5D7cqQLv8GUYqTUkhiWZMkbB050J0jpmCxi5FuPMl8MHmI1MkymkloEksZx/Mvlmr9AuuzmB
4HYTzvH8hE5T8ck3v3MY5P9RUmnzsox/1ZMa4bh25JfTev4ormnkrb1QapuWbYLsf3dnxpy6v3w9
33gB/2tCfLfTG6lyWoEtJuJX79NXL/0kxKFE/MWG2n9XdStKn89TNkMOS0nDmTd9lI7Q4JMQIpks
b5RPb9sLsMkq2nUEImIDRN+B+PquxGzzB/72QIvw5MeSI1FFJ9R3YmpdcoxQVuJVZiWHzTBpLli9
e+wUgQKexqPYt14d5qTRy90EVuBZ81+WIBzZ5ibXDZizN+xC+Rbx8Ev6JB2nadF+ex6E939ZNEub
utr+AA19eFces3kzebZcm081FOENbiP3i2PwBsS2MfGqB9JKjHFUL/P8W9QW2lA58PTF1LDM6sfj
0WBbcIdQGCp96Jtp8yWM9dm9f1zVjUCmNRzN3GmMvia3RlyBCgx2Agbkp+NobW4xzznxvMUGNHU3
ThYDJqhItVCfJB6BicLQthGBxQZ18prmN2AYsME6q15l1AXy9LJTYtgp8sSZEq5Id64MooRG0mf0
R+tlpfAjdXmYvFs2BTGAkLH1Yv1LFHR1tgK77MzwUCy+tjqW+VT45rvQsJPwXq2mpOg+Mx8/fDh9
Jhj9NruX/WcanX4xOFw6z1b3LcV497nCD+OvcMAg29YUU6y314HoqMQ+2GbMJdMZJslRFlKCRDqj
k/s6FB8TCWNUTU9mKJ6v8y4YlPIy0CORsvf7HVxSSaSkWRuXVV78M2mXh8JhzgkHulJ1SXa8KAEW
wr/oetVIzuwKoM+RlCJUR1qghN6vqvk5Ty3Y02Onhq02AJyzzTo5HpSD3fPa/UKnFzgcvpazzOtV
uNkRF77f5nNgsMS7paqYnWA0ZJ5wNRRpkY5By/4w3Fu468M7TvYTXJRZ4lr0LNf5UcfHBmWOB/f/
xXRAZPHNhTmV/H6TZxZKjDwxvSDTeVIVHql9O/pcXRGS75CK9XWBZoaUMDODZCYzDoWKCFjj3MBV
eq06JYx0IKwKhP9Z4SOo6xRhYySJEVq7m777ix2+EedWU9DBW9GFSOwo83iW1XGNKMaLHx15Emh+
MH0+IdEu6/Z0N/bXTmD0gc3oQzNoRkg8blMvmJCjyolZr2uHl6i2o366ERezWaHMvJccMNYuoXO7
7+f6dRT5HwjvsIU1oQuP1AaWh2gOeweLES86q02l7MX96wuHktjij052AE0j8x//yIVmsOkhRd9V
kgl8+il4f8FnfSYjdH+EQBF1sgvaUPAKEkpur9/3buU9mdVd9O2yaOnTQ2O3Nc5GlhMZl+EZc0xQ
AhmoVn9JvPUdgws4HUD01HyR2NVNvXe2bXsXfHrSOYZD3z4wRtsaL8/wQxWP0UPZcwJPuezlr/Yc
Rh4FVxfay2V8Dyka3zdetPOuhO4r1r0kLq9TY6Q4gt6WCcV4/a3VzO1Rl6CasTwDDkcntcfWe+g2
e5v6sI8rlZanudzpUNJmiKQ2nTM+ZPXRb8+Jncg2X4xtKcP9I/jhepNWBg47za6KiXJV5RHz+/gl
ZF/B4Igmy2IWX3/I9I2DdKgVcFNCbbYy30GOmVEh/3LkdrLVUz7waEq7tDBbeYzIIpwWP798jcbe
9GVkMOpeAO75mOd6wuuHecqZyoq6q+z0aKikMTwXQf9k/YS88NFJnV3aW13q7+wuCezLxI50qdAh
MEv2igpfpPr8q2hz9sQArfHvG39FkUQyioXlYJ94trmpfldPIxh2mPJZrku5k330kt/xKuOy8B0A
ZZwHCmQztmSMApBPzL++ZF/J76IslkWbGI2/mwKH1xd9kQRwaE4IngJHNegOx+SK3Ov+WBB4/0TD
TsfCz6CpYbLM0emJEAaSEBC4GQgctDF6A+IPbDnii/zBjxFZIgwF1x91Z6NPtgY/WRvMaF9GpvbF
HveB4LDuyR77bBt7KcTSIOLWs+f6YCm9VYG73G8r27zD+AbWVZyx4SsBXeDsY6Xy7vcOEbbXNzJ2
qZpnKeTp95A1ZDBo7pyW1WLR7Ne8dBwNJkPFq9DBv1F/CEQsJqStFxSbwWFepMlayTXzalygb1KU
zawJ4C4lHgydUgBDJeWmhgWXnQzeQBb16ytgGrF+E3v/BWaj7yiAdwWwmHw9y3TWURbmKuUBK9OE
kwRzuYhI0mg8Yli57FfGUC5IRQQ54fnydlSZdeO0QGBmITskYzL0R77SdvO6zCIG9umfXd9Dws8L
r4RTlGiDJsbqUBf2rvK3j+xW2Rg+GmXhwlXgGp0Ah31Svu6hduNQ+1y5dvTJ/Wk0f/iTpLx3qV4T
1NHRH9y4g0SJKOPoLbcWWRKrUcOM/UShu1eMPga0SoEd8IT7ZSZRdawa4rxnyNRYIcrOkvYbpgw8
t7gb0WE9TIoMpznT4CY64N3P33cMiONqk6PcCChhD7zbAhrbBqEAcEIrIZY1ac+Pd/Y9dj7NMPSq
KFtqEFPuNBSnEC2jQ2MSf3JfINm4kI01MWkUKIR1lgvo26OZ1WhFyHrv0Sn5zk0z0d/eAM0VrB/5
eJDsvpjv+tY/gDLkxS0Kxmn+rY1/3KOb1qXuuxpWz3NPq1a0AEKx7xPg86URPFisPhi2jyrd3+44
2r7uWvVRNjRdDkq2xsE05bTvhsemqDJtBYaWSekC+x3jPJMifXx7qpOecMcaBORQ2xoKva3ZczDB
ehmwE1pgepApK66uAqXjB6cqTcka1HSxi6+0W8RqABK0oNOVamalPFnhJvkjOEyVe/LVtZsIYf08
pMjABApLyRwZ95buO4rdl4UYa48l/ltD/EV4SSq+vJdDcpwXBmf4TZUKDtEEPxCKIw+dg1upYfG9
AlGSoAlqtEvTLmG0Ngsx3wqwI79usVMtO78c1I1RDCEMxyE0MtNu9AqcmnQAxZDbIdCVXgtpeqxl
qR+Qeh/7hyJQx1UdlMHPYOzAqimyLKHpJuaa0Y3+I2e2fAVt/gKKgOjt0PgFZt3a3e30/6adJBKz
HHpEku6KeKUaElvJ/INAoaQha+2VHvilKKs0MbqpJktcL8LDucPp1Jnn8NBkVpKk1zqJrx19DSX2
GuObYZknThapuHE2BRMfCMcTuGVxD9lX/r1ubFlvSkicyZ9Q9yuau7gJIluZlsOaf9w1NGfgYrBB
U+aaihk6BYWdLm5yd2A52WA+S+fhl+R3ZPZeMpkHcmL0o01LjrQ1EM7FbCrBJEvY4+oQdX3SuxMS
RxVVO00DSYrI/dFUoMyIKbzvWx1cFJiMwsWpUsLvfUvkhbikiqjgghuXtM6UacHUG3M8kaE00wC5
iJz3JKaKu3nv91FFQWZM/XiwZea4NCtlBux2I5nCmvixMXKlHxnptRutPmv2YMLEheylFpmuOr7K
mTv6RMObfK0vaTWjVCdDN2VGZOW2VRqU9bsWu2qg5W3qvl48iP1afPp3DgHHNjjjk6bnaoS+vhZH
mtU63v1YQUI7bJPSi4s1Rz71ac0Sz6dR5PIabEmBlu6jMBmGWIdepkYOr4lAdag842jR89oPVl2j
jFPySd5K8Uu/noxYQKBiWkbVTwOxMtVWcx2/+bHpNize/gB0gickn0ie97dtTKJ1yfvL1fZkEHvx
u0Ioqxcan0lcNKBFtc3tFIQm0bI5w1t+C+IaEdUFbhMrT0/hjaAoaCCW4gPX2AjkVrUSlyb88p58
Gnv3mVpuSt5XB+iG4Ycd77971Zm/vr38V378gDWPBtdrKE/BtW4t1wPdSiorjD/iwoZerOgJm+W3
ZeqokmYUsIVd3YWgFuMDpejgTQUNxLVDAZN7NObaKsP0+w+g6abwxAbY1mjJf0LvSlKGZztJsvZb
DmOOWPxfhZh1UJXe1Y/3Hi42P8IVyET6hlEI65fNtWOz6JqqW7AfYJVet3ZuSENlvmv6mirp3K5O
UdKNNxH4J6OkcDnvK6N9XngBdmMi/BcLTGcHha91AdgDJgyp1pxg23SyFg8SSrA6CeX9TkeQB8uA
/cjwVIOrDo2XxB2b4M4vk6/4SM7NXRhjR8O2RYGA/+rdMoY2IBHL1GK4pNajazJBjZCPcSNEWQcM
VteUZUW3Ff7I/toYQAVv9qcw6gl5rrO7LNYNCkGEfTk0dBIFgfCjzfxOKGTsHK1PlTrI3Rh48FFA
c3nz3NXV5R7yQV9vqJ3qJBbV7MRF4BhArXv6crIS6EH4t2H2XrgA0a9cLtOt7/sW5ZI0gHW4/44J
cdwa0gUNLvrRxQk50O9/B5h33IRjV8Wg6DcbML6BouGxnnHhPQWnpubKdtrggc0eNRXoyBdONeuO
8wOPBnNIcI/odqCBNPqMJglPKTkrtqHRcKpZdHIiREWBEpyFx+K1lhbG1B3RyJf2rdxDgSLsCnu/
5dXgV4c8KiyFwp1cKvrzcfrTurITB9AbChNRMw9gujqyYqIPGpC4Io1xcKf3UOo57Lfvsu5AsUgJ
31W6FvJTEr+O5eLUH9IJGFz4uVxtTTlnGp/vxrwHIbokx6EtI+aLRjmLfenYq6EVq+QbmoDw5gad
b1lEcTGTQIb/Qv38p/qSrA2aWm1DuDjLud3YgknbVcG5VjMwy/S0eeb9Fnov/rl4r601zK0NNEFV
d2wSYQf84aXq8QpgXUKBHIwt3j2uVpuBKj6Eiz3MCigpGRhPZZ/PtLYe478WRJaqTQ2dRzxT7bNH
e0Bv+3A5btb5A/IZX4DTeg7HERX3qFEFKDzMgs/UnvcqEotzpYc+AlGYoHPd/vGuY93HEQKYPUrz
oPZApZRI7nqPTHwOjR0qEH8T0d++GkIa8yvxFSPG/CBBnMpzzwdRsq2pCnfovc1l2pBqcTtQ484g
nCkhE8NhuywtpA/hofdfGzSKQ3ARJhOFrfRUod4XzeqWVYdDr6lest2Hig2NER3NWnklmgwFlK77
XIcqTNkCsbKMmgybMGhllGFVpE52K690aOTyUsayjwYWbdctc4j2YsQ4hyk6IPZ/SymWvJ2QswZP
ROLq235bl1LpJ7sO3SDvyO7RDhKdU9edgzxunNC5uk0vjCuKjhj6vwxuMTbZM7YjulsX8ZL7e8e8
tLEDqMMvdlop4JiPytMwePZCEe9S4Q85UQZZRPnxCF2WJfiOPQ2ZbH+yGrA28RVdp5DsRvwUWOew
nQM0aUnM/RHfjRoWEUIDlhugWapune+QIbv9QqnN8EN0jc4ahbJIGsF6yK37smaDJ5eizAtf8Eaa
jw8yiq34D6Fpn15woZZmClW7BwfCNEO91UyhilrcdZWNQXADdeioN7HPHPSnnPE6ILRb2Cu4h0db
zqB4T9CmBm2S5sBW1fF/tRkcTUbc0AJvcVQPh0HGRhy8m7iQMX2RuiL9aGiUiXzoFImykXOdDhHw
C9XURiWOc8c2y8ZUCv6A8mfRwhxurtiIzC8ClgLPKnhpni/c+Op7AY5e1t+RJ+MAU0dvTtX0tsQU
xt6tqbS+g2/pjx7+evNyfYc7SmKyLpo6WXzaSuxueOpTJ5FdgVHjcCz8rOJH+wQXBWpGptrKpa2B
+0yRJZKUYX4tqKbIWAhi8H47fOgwG7CtxhpGt+LVsOhwvTMkE/xQws5HqEfS3G7T0XPKYq0/78XE
93U0V4HB+ghobKAVoK66tXtVTtKZ9TV62mfxFPgLbwwjO8C7j9wKvBcZb9tEC0UWAnbnSNVhoF3n
78vE9p05aZ+0EBnLe43+VJL0JlEe8Soevht4pRVrXZBrWlgm+X4fMX/oD1NwofC/QccTEU1z/bGl
BJ8o4QMOWGMfGmhJwghDBxRJyg6qvzU0klHbh3iJekSetBqCz92g2uccjXA8Vs6ZOpw22TN5DP5U
Z2WKOj7O36wNrLXm1MG3x8f3tQYdGFznfR20E0AU/6qt1whKVY1ns+Ve8SQUrjDwGlHSOfUErX4V
HA9czAzNwsXS3pYaskx6amv5kXAMOW7TNKxMetxIEcYnesbU9DUp3G1xw5wwg3+1+ZcLFOK8nVKC
z6uyVqXv1ZE/ZdHAMNcWBbx5GnZzsKEKBM31WZGscOPZ6k68ZPM8/ZaL54/juUgC7UDRl+xiD3iT
2Z7Qb36Ml07HpH3pphA/GueGzSLqokpNT74ukmUVpvW0Q+DrKCTnmZJj4JiF4dzPcQWVMzsuM+Dm
dMRUXr3xlyrbHUpBOp0pE95gnIQWfmiac7fkWeNDnrKoit3UGqnOSFQouCxSRLDfN2d3NgUgnfC1
NG7avIarvsCwnQQHKVy3RSTlwIik9vRorEjm1rlpWTkrK4y5A3AkxjND+I+w4rRR1Iz7uKj2nxRk
qr4wpeBe+qV56kzL9QHD6bvb5lcYPHlZDMXuzbZ0cdVBFXh/Unx+0GNrZ/RM94RN0ByDpwKkYXSK
UA4tsSJ1nFLB9OMumUHWzuyes2WJSxn6mngB36q9/L/BKtFfFpGkR806KIM5Y2Fnh04EiDVGcXx6
+7i2ujDkl6jQjlcAla+OpEFYofaDtF3vEodaQKit1Aw7WUeRfEMgZlgLQjs7w/0snohOFRwMmCUY
DJbuaARxk0qG7hvydXgCAcw9CRTuSbP75c0xBIGyiWrn2dftMNSOFaDGoEUVRDEYeGpEjlyZnLhe
ysO+JwZ8vckYgq9Dcd45YeyoSsAiuLhIDw8aLZVIIW2i64Nyvg/DuOIBVQP1dQo7Ty84qUuBOIwW
TRfSfE2BjfDW/ehb8WwEe5UP4vDDIqx1fj+K0CPGBj5hYOZTCuJK8ACkHq1HOrIHtcSN5bG9qeeE
C3NvC9xQ9fMMJJH7oExlMisf/LFBKyPukfVvKEm8F8fZBOOoNDD89GFlkXXe5TtUWA3jGc4zk/aj
ZDsvls5dMdYMI+dsAGAAiTnucLd4jMlxXyqrHIiBN/EaKihimHSavYJCozS87M4RAO5FY6rJ3DEV
H7QGkG2jbmFfCUK57xRdLZCfrkcXEIC39eaI/gsIaKefs1n2pcEI6qxtRasHENRdyS1LwQNtFEr8
lxtkmsLYF2eavaW/sDJ1wKE/tYwfaMJFxmAMJ0hyiodyrCx463EagnzmCQamNNFWuxW79q5yTVts
sU7We80DvPfqvP8OrQl8eKCQD03tXllYqwZQ8g5whkTpjgjwCWTXaXqdMgasOSrbwzqZ98aEIQ6k
5R5m2xP7Q3GUAQZlsHqgLE49X5QrTuRAzam0r5wRVQ1a9KGMy6KYlyEGnhAhRz5YgVaKh/hSFjJF
L1X0ea3BJJly8uHhK6KhzjTJYOKI0V5e7t8pgfIdKwQEb5G+rLsQVAVpuWcRXQUXvNxujC9V7X9v
lqUzTZ4XW6aLQRkH7R32Z5IIPo3R07MoITzUavSrRker082YzJ+xUWip4ZQVyVj46qSSkdkUeTgv
7OyJg8daA5RApBSe/RLWdLlVt4TDDfIbIuvrkj8X2L/J75BksPzLFiZqEyQloZStdwvl5nHNxfga
CmwVENglOxquBhGT4rrM2y6904yXmfnb/OclFFIwfAw574hKmjZCCMt1aJDm1MwHvv6PkQf7JpbN
heWFdTnWbQqguAwo/YnZKqRWehVEuSlx5HdmzoNZH9QFuyqQY7Y7oBkKaJf7FcyWjyzGbbZ95R2H
zEUPNDfSqJn7SPvxl7606Jullth+a1cpZ1cOvXp0ANnGjw6TukiNQPJdClSB8RzhhbgFvwgE/KyR
RMbk3wiUBODwjxRNNGsboNDSnx+sgdOifE54YEi1BbBUDv1FGSdaWOeK+cDC+4I4xwz1TloRsiud
R7chdt0Rs+awxj5RlFuzPq0C2fazq6jOVhScWlqf/463aeE3ByyuPfGw0Y5vZrGMmEY9PuLAFued
LxKvnDNuTr8qWNhl9l/vKag7SsC7DoGtryjqvQTR5XyHtV9j5hrVXYZ1MUwlZWeF3ft7+o6ApFMl
ChsY/lEa8zRxYbLNh3WBsyQO9rEYCGJo8BFxOfpzz3kAcpNcMcpz/03bAdvYYPpVCnc0/GYQsPJF
JgE//njveFXkW61WUl/kavTl8QJ7oIojR6ZQ0qck0ptOtEWRxeer51T1GOfvuI0ZlDcoLAHYgllR
0h2bL2RnlAItlmDuWYX3j0KJOwDFQZXcuKgPJPh+Zn6K0oc0EjPcD0aVvNhHhwA0AXWcgaizdIN1
nFpFn+u+Rj4FHBFs3/iPU52p7VJivp74eIb3dXfnqLcgYYOnaI+DFv6Lgp4ohBbOCCPUE3ILGugN
vOwrUDloIEDSb6w9ziCJC0LNud1E7b2usCzCtFaKJLXk5c1Vs0OQMp97yKBpoWt9yRIZUX0b0iIL
O+9QsSym/gckiogQPYn4HY/0cVB/bBMKpC0OnYLitJQnILVmp2+/aI/RzaMeODuDwOlU6h/AeipQ
FZL/QNUdIpldCrAqADorZOGxXxq/83bwq7FnhcZ8Aun3tH8+YRljm9271oHEQTsd12aemz95sZHP
+Y0s6mwvcFds0vH7vV2Cdf48n1kYrUPHDDgU6KzkuMur3oVYMnfipoA1J5JxW5N9XSyxWdx9BBIu
fBPCz9HzJZvyNhtHnBhvvsvc0tjpbOKa7BKw6zlEk6h402BvMqHSUO/Kyzpw8jUBVOTCi5jAzDCJ
Ek8rabxbpQWw8oHDhPd9SwFag3BCfuLOV/XobEqWsT1mElsUNVoINit7Eddn34xbAsTZUi4E6myc
5fjHNzrk9holp0fmGy3h/rfKiHrknDBK780UJW+HtCrWm0zUwiWbJi6cZnR7JS13IcCoDWASRosA
DcWCiyMxbSiEho2AEoSV8nF8pHA1YjYJuqsLx4R/ljp7RQUKxZf9Ce98l0OEzfzVPxPVIFhaMp2g
vmk78BvXN7xKtUBBKkepaH0Fm6I9j77pcpfgybiyG8m0nShEF2w9DMPlG6spY8GwAND0skqtuDmz
kcr+jinDEOJO9INgfCKNx8S9Pz71lwM4sUvM/T76O2HnqHAD6czs1dEFXRkRoqMyFOjeTRtBayBs
gE8iLl8TsB5tdzJ11dgi5rpi4Bfi0SpyRgz5yLP9sggAiLQmlydO2aXkJqb5nJfrSxLCagGTBGJx
J9VLFIbuJSm6x/aP7T4L9OLB1VGml1a6akRpBia4USxUMW+cC5qwK1xwG6dVOwUzA5dMbIrGF46l
4Qj5gIO7dZvCo1Q58NH59vc/iLqheBmbBvfU2HoSM+xERsR6ltVr+iV540kpBWwiZF7CwKPdQe5C
x8bYql7ffSGuTWbXgdEQG5ca5hoUCRgolevBTZx8fHxh+AtM/amP8GHd+TUSFGOHd5SY8L2ykS7M
3/iHgkyYYgwk4pK5QidKEdfhH67ZtMUt2inDlZhAERRqZLDtudizQa3SlXs3l8cr7GD4zyBZGa0d
Xvl9dqBB8TbN+eo5f3oON56/MQRIlviltibD83El126MV8+X5Aj73B65vGYWwXrrfk52inDUzOzN
XT5RCBqWnW2hJHI7NTgWYaPebt4gu97+th6L/bjoqLHYMllXckEMmclS1XHYH4MwrM5R/jX+zLvg
Z/EO9VWAzvvKkjDaTM3XEU5DJ9vQi6nBLJBH9pxtLCQe35j7hHDKDCuPr0M5lL25fHsX0srGo00E
uEvVU/ZhPXPr/G41lcpA/CD7iPoCqGPst2rrszao195RUKwuKKA+TVJQByHK+Ig/l4poAt0MAdxR
geEvQ6eZ9bZgkE/1JeiUDPF09ZnbcSDuUcfxSU63VOBRTAvKIsu2ikvvZ2Hb8cLRYYIwfdn+FABI
XAp+ufJQC6XpcVuUOfvUL2JDdk+csfPaDOEPWw5WChSDov5nVrRadx/Lyuv945xt9i39eeVUvWTM
ESUOnLn47TTskEfA6m96U+lwIWqmRJXoPD/JbwIGNgc1Ajx/0DXlNPhUlG+F8wmmCvE52oQaBcGf
iqedROWunAjJjCskutJ/6eFArwb8abHEV/9ABr62JjRw1vog48yRAZfjqa3X14mHRK7s1iBJ2AnW
4h+3KnXynHnvjE+Bxwjru6oyqxF3DM12C5vPyzpJo9rYIfBso53Z48SOUAGmUrohYHZzwJHhhyBZ
d5Gnaq5dG9gD4WYV40NFctdcyAP/XnVOnMYblSAhnEfWL//8DjkxDcZQHODGtIR2cVxuKvxiB3L2
J8eZ7YIQfQYiYjYnQAhwY8tosccpc8dR9vyobgPd8OwI7YdsWsVRwib6j13TqGwUaqXT8HSWr4a8
Urx+kZIChIU3ht9RfiUirx1LOpITVGgE3aKnl5Vob5xvydLw2EwLJGYZh55z6Gp6alzKxTv/dG0l
2oX/oBt6UbsdBA0r6aGa8UJDbVjzrlfIoOiTVmjlM19rfanJdsRSOei/znc9yZxVrRbfQyRDFqOS
lEQlcH6NqHFrUlvkUZcqP+5ksAwFgdnv18ikQ4vunpo70QfzSSQoCx3q87hk5OwuwpCWPjokm4WU
16XaSpypVO5H2/9KxyIbR+ufRFhM0GSgPZMWZXh07H4xUM0p51pMbPgmgjs55HlWly1uUP5ht/VB
cSa6b14fEP0EpSbz8QHoJa3pwQpIXuA81+FoqqAeQbHL625wYqI4byvIan1nvzyeR6m5dUdh63qf
nuMGZGkQQeHUxwHa8LC+2R8pKapUX0Qn35d7Xa2pZjGeyAPE13MOrwH4pKz7cTEey6hCftdh6zKV
i4LpgCmyNAcfpASjkZiEueRta8HX3Zh5ejrbmeOVMA00/7FtO3m1Z6fsOzs+exiyidrriICQdnD5
pPDJbuvh3k1CD8Sy4B75jwef5WrI0bD8+49aTxNUBxFVgfKB8boEgmQNOy2OIR0AYfNJOixYJtaM
LQV4PNSOIji57gwZTVFrZC4kBtmsgX5Mk3HkCrlyv6L/+Fk1s02/af2UnrSUwa1rG0rFbCrEGJnE
Ecx2qShaOs3fn6od3CXWvRrVN+1slriAbGbCdKcBNAWW6R8hUD2KEzZBQ6mfmmZgHzcN2+AyW97b
ysQZT/m7ae1Vcn62X6VrE48WVax3f4QIwwvaOb1WMWSqN4i4ZZlL1N+e+YO2sNFst3eYckLrhf9K
Qc4/kYD+1yZHRpi6pJN6smlUME6j5xpgFQ4QUCd/QbSh1NYk/FjjhycIQDnFS6bOa1Bd0vHDZ/hx
3n9jejNXqbKihcEwYGhCDLjqoNJlLBSenUgHPsTbWbfZ9Y3uPKeQ7iDixj6OhIiJW4ZBKBQjoaWp
JKfJ8Y4f17/6ItTuhzoSKW/prReWcxl2vcu2CEdiQCrAg00gWm34WKvlgj5cRr8EVTddK1RGJ6IF
IqnYzJy4WIoYGPKDC82Lmc9exEsKBj63L8rCQ7vUrI1U9Lbzvizb8jqwNh/eqpyoGmSaKwR5DZ4Y
NvFtuXM81Mwfu10+AzKcCagabgKSksi27zrL8fyCGmYsCwip22wpVfeVl1HXwaSn1EG19il+Wim/
ulKUC2oWjr14zbR8qsG8nNFkxhlFCBWPpLic77PglGA6MoJr/CjTNr7ypcNJA9aWPP3nHirs8/Zf
d+vFdlfbZzgXJwT/Ne91qVNSh0C6kabiayItLPNnPJN3gYg1Gc3o0OTwczWcSgmnWHSlegoD36Lm
nayo2CZzIj9cgqNjbnxToPwutkKyPqTi8Nzl66ToYNsAmymOMx6IEwFXpoCa2HbAWZ7rLCQUvq8K
JVfRdgCJ0gEjkY+JOpYbGwl4r+3iwDiCGWNyHA0lR2MAvB390crAiESCtN0iwxyrH1hswcUzkP8g
N424iKKnKM15gewPALJ5XOsjM3b1PFK8J2IGlmM+Ix99fcNerjKiCGm1kIVfiwPd9IZlfUgN0mGQ
PJeYP0PUBpZ7ye5AnJmIj4XVXOXTKVT0p6pkoqeLHJ24+kSjs+mPXvCQ7wiOHxuCxNLu6y5X84Jw
rqcXazsnP0ouyKIhDHcOBBTph848YT8Y2xcTFxOyDRny1HVQobwOKnerP5LmORUsMeHZyh5lLhFo
15golKGdU+8zJe0ceeZ8NJ2Ct7dCH1d9yXNZzcF5t7n8RjaBnSwt6kFtYtrS2uKgGiXLoE3BBCEK
9WGgaGHUQzn8OrQ0uPeemqhPO69mabGOK4nIgnvUop8+nNSot1NXTmCfzwX5G8w2wEZ+CKSHYYlH
AUhFUr5KnuUGBzno2CgDy+V+E+OqvPACxSgLkPdLJg3bH6mvgzonzRkBE5WFjXAAi5i+M9Q0c5Iy
zxi8znkdb/mBjXUmc5Hq8749kpLj3WRhhj6wc903YQMJVUekgRNq7OJSgWfYYD91SdxmNkzh3QSi
sO0MSeN9pYnye59O5Y203xb7I8oPEGHEKzg5GynJlh0z/kJmzsOV9NtYzCs5SVqE6pdMfRaatPwF
ZU1wXO5qAr4c6i+mNqdpCfLEvUxQHkRnylQOEKvfbDD75nvfqXoft3MnsDlhYWT6V/Pq8/vGkRly
jKk/8GaqqBwePT5osAlmCU/dWDNaFdhnDvxMb9VhDr53vVQy34TgVh/LJozWm9W70/h2j4U9Ck0Q
IcgcvzI8jB2zD+w48zID4Plyt/LNu3B6fH7DOj+y5EUChEmtwxORK1PChOSIvsAIz0IXRJG4bDxM
PEb1Bpz9p3dCHs13NwbO4fzlvhZggtlrS1f9Fm8oHCj2PbyotWJ4n6r+eXX8tBztwbA8DhU6CZ/L
PUJPbPY7Ynj5KtvJjK63FQlqu/J5HbpwaECvjlVbS/onxxOvfrqAUWz8KElg9HVM2IoCVmhgdeAQ
cQ/IeO+PPyDJE+fiXdvS9Zoaw668TWIXzVOKDA3FVHbPpiyfW2PJu8aFm8SkMjTMLL7ESvJEDquA
VZnX7ndM/9v8PdLb7re2+CJZHRpIccPi1p+x6LJvStjMQsFe+G8jUmSt6in7UjSGBOJFIRRzOCpV
JNWYzOBZ3XDW5uXr2ECOxsP/+TMvJIxb0dBxcozlMgoVGAF5UlvM3U2c3tynPFGVzbUtlZHw4y7Z
NHHbezwGhahSjC+WRGU2ZMNY1FiQmxlgzUrgu6h2bPjL0JaAyaSAORTPNg9JmXwONfGxIBipVzNf
VhAAnajllBLcsxLg4yy1CuIH/IzpGH8LgsGtFoOSMh8LNnVhcLZPuHZBDxkTfiRYQTbAc04hf1wc
xHQ0V251/NYV0THJfAk9I+QVidJQZoxjNa/J1GnhknN+fQbiyo5gMXGlIthrvLyfGkuRpU+NV3kD
ap5apxMwb+Zxmylok3oxNjx4u1mkpt2W7aNYC56J3a8MNUL7Tl6nE2T1+lvJ/B1eaZGwGkGCeUE4
KXJ2GDzvr/y7o5TKD9pvzlDlcRza7rvl2zWiXWlfxTPr3cal9rmfu+PhpOjnp5Jrx2alErzzOjpU
ZCaWgLzxFyVkRHISWNJbds+E2NSAxFJbe5ayTvJmt3bLk7Px8I3lGuWGuPBx2+Vb0vKlWvZap2al
mYVi/vX/hhi2neSfBYGbYeUgdAo/w0+FZ6ekoE9QgVd37cEOiAZahfoLutJg+1NGDqPUkp4uzbeQ
rD5XT1ZO/FF7hEZTFA4r8ZIZE306cuOxK39vTs9cUI0QyRblm3tPDl++c4fScSKT28o4S5lwHYBZ
ynWcxkek9y0J1VDzegC7gG5vEB/sd1dFhQ4DkdpAvUhZLicvWt9MNnzmc7T0lfzxmG536uMOvCML
PgwEeF+wntHUxseiPvojnmM7Na8rBQhFAxG4sVxC8N03FQ/DYtGfn62F+W+WTaGmFzcPWhKFVl5+
cdZN339vmFncYcEkVa3dYvPmtcM/WyTEvubRzG6cvd2Gdk5ZLwVeNpEdHYuNFjW6Wn42CiaRtek6
w6fmuCt49n8zyHRDHiRofkJphlZzTHsZf7LU+yxIXUUtkAXxqOJqy955KhBUUkPyOVq1LBcxKr50
qENWw9D7p1jleb2aF4C8TqbkCie60rNC33nMJMGwgFry5m80NSWzLfxXAv2gLb1taC7cNmFpYex2
1QUKLSImeXgWKmp8iknS4KfxYdyG4MGZuk3tn0oQ1Jb2/+4uqSLgEq5tCs0jw6D5mI8fDghoekK8
E5C94IJZGXWlTPUQ0dF6AMmBHmoucDZqfTcTMKHoHWeJm9TKMF0GBlbxdwEnPW5+MvLfX7jNTsTc
hD8bfkrlfEhm9snQfMrV/H86ey77o6aVSiHXn/nE85nQALZUUKcNMKnrEvFTas2SaMWUFP7WH7IG
FTcdBMmYtA/KWf1JiTsvq0wNp/wZqea8nsRQczsPHCxkprPg4Y4EbqxbdSFPj6MAF0BNrXhcxYEI
gakO7nDgvmxsBtJrwjXuEP4nbkcXRbw/OphDGztbuKRiKazFGYY3sRrnuAXN8zMB4eJ4LtiEwKpe
f+er5mp84D8tguAsC95+KjosBV66D4DBh1BQXYHkziEITAYx4IaVpbBNsLqdYWx0+fv3ztchR4VS
x5/6FVwUjPZ+DxCXj0ysI9JqzKeKSvIbAMBbQeX90fo+G6f3fv4FZZ8ShT0ToWeFM9Re2e2mAP7x
p1Uur3W5/NP+77TgKxklI+zvWE9s5/rMnY7vzeru/DOhM5Eh8Rv6P1zEcC5n+AACBDvmfYr4XLuD
vbZHojAYefyTLoPc1BUGLA6+U85RK80AnH1/8SuKRUOnE1qrUw8NL/GOEZYMrw6m8y1fhSb35G7w
/FS1o4e0SpM3wbQFeHs5UjOT1OESTM85O3TlUKOrRWC9p9iLZDwRnJYfOaCULHJSJEd2BHUEXcS/
WiOKXnhr2NDTg9yL3fk78uGrjcQZ22Gm2KrasFh9koiD0qWYPZdOOEeVLq9vroYz/TUbzhqb13G2
kl653k/zn/UDL/7kNn5d+rS4L4V5UV3MCfsq1Hthq/uKqI5UvDOKRCN27nHBzhdp4kVR7wbikZRx
IMynI74k8WBKjF1tyt0nTzzxrHr+2I2gitPKcEkoo5OCGpfaDgQ7MCC//AL7bz9AWNHrb/sm1j0/
pDsp/66nKoUVXAoOsd+1wl7HkW2GNtc/A7tUo4adbmR+mkfUK5dyYXeJz3yL0oelViP5aGhmi9M3
0qfOhE7y+7tyVDAjq16avmO9h0a53iDUCTKL+HBQYppj+Zm5vb6dqJpWQvs1Ffxr4VAAU7QSKV5s
4qvsVgIWwixatepchxEMfZBQPw9RjXes7E1xNJvAelhhZFz/jnnFXR35D3GgaJ+9CU8sVynQTcx6
T1qwp0San6e0itVMA+iz9C0+Q74l/GMy4F3nCOx9MHKnanK5r24j7kYnfLw2SlfyY9KNB96B9kPc
IYVbZmsPRLLi1fhtTNLcQ8itGWlh6q8hQ37PrTbi0Rb4r56k21ayVib478G7Jl9O2+PfOB88Eboc
VYwP64QjEqxDwqRj+Q1a6i3AGCzjsKn89EFCENF7Jcvtm2HeFl3iNyBtZmqqhd9G2Eq3y1kSbFVb
pvagkHdmvQ8npSv4kxYB3AwZnB2Ti6+UcAhPEbfsSik0stJJh3sfcHf507uNx3NWMbVev9WD3z9u
OVS+iUC/nDKiUN0BMQBZW3eh9yYvY8OKlYzyJtz2hAsU52A/0kLXp2GzOtgdVeOYjJW9a6ciJEcD
IlveYjnAdu/TsoHE+yIYgc7h1Ctvr+FOi4a2QznUSgzBNa1vtMK+2+ZGK8eN5D/6lj+CE+GkquFl
zSyi4us7O/yrmj0HJF30Ge3R8SvpYvzCs2l/FRTTKEXHYwkqp8McNjMQm7krGOKqBK9LWCxbAAOb
bFeiN/8/sAv5XJvy4OiMysichCHMn3xnbfQBynDQbQhj9gNVF7VPutgrw05vBCs9bi0WeJgyo8CI
hYzRNdLd1E5iGDIjFzupZDPAYr8qUtV4fOrPuCWWyygg8eBVUFd4VG8KnTaAPgx4y/czmPsI6u2n
mLg9X2zsBgyWVYHKEzQSGmA2i2l7yjSE7meLd67QZDCrJLIyrzMtIjz3bl1bLOHAIxLA0+b5r4ax
ESY/KpK+vssFgXdQaj1/9P+TRVnpw7WxW68qxADennUnw0PiDpPkxShyUDqdxk9+NNSsgeofvNmM
bLgAIE0jy9JiM2YveafpUpwMg3YBsW/EkpIemjCDbNXviTHSnbsXLgkbEOipOxnxEu8h/6njimG1
NVHrq0D4TRDARin9d+FOkp4SnocDwVlqF2RqauYxonNUV4PqQm+6zn01VH8HPp3esKIMxEri7Z/e
TD8yU6vOmRpUURGEyxYmZx7KEQLrBDxIstcHSIJambGdCUvoCVHA8ZMDeQm0mRWTizpNYv1ITYcm
X2CvmfcH7V3431LbSALWp3usTrYwIeTzFIJomViafWkPX/MQ8nPxxIejr6uPeTVL+rcaPW+drNPx
RH7Xhaf2ZbBAvp+XTzYlhXm7E3bSZCq7FVsF8f0ew4G+f3q7a1L0tBnIy+ZuqOLipj6DCcxgOx38
mxbtmvOeelRd0jk/f0iFEFAx0+D4xOxqzexQc2nYDs+KL9W013uLSdQSlNs15/N532uHBlFc3d8/
BN7d7EWpASbsq6OC5I5J0vKrnVzNbTPzIRGazgpRb3jmOj9ItWWLERThRTCbKJiUnDflzOhPDuJ7
HrRugnSInFST4F6Az7sp0oP0E6pwccZM5pVPlZOjHmSaFtuhdcNpU4ruBVfGxpK+OGf2tpbp2DlP
6xtDlalKKWMTpL1AkoJvPMJKmYkNVcrS4wl9ngLcd7EVbwk8mbi3N3ZvtjenUU8ZTKQFdo1Bgnq7
7jDvzdqOJsYAkQ7J8UXceZKXVezIFeb7/lMecLqvfpT+B8t7wR/pAjG8z3OVeDej2FOwGdcvNq0D
0TIrcWPCCGjoiTk7pGTBRvEfW4j55VbCryVBc3jXPuxCVerPY9vkxtGFhmF6IcBJZo67sCbmm6Lz
qjhtELykff+6uDbVtAMoWWY2g/9FEPnzKmCi6fl4jUk/WzaeDFlBtZ//xOah9ll64imqxSTPEwys
1YCiO5Ux4UJP6zDX4bp6L1ePGOK1wBpxnKvWgE3oFY5vJ3lV5iF+4CzrYCIndFuJolUG/tBwpMSw
rnh0RNmgLpmRUDNUYIu1oywr1lNx9nh5BR3j1iQqjB222L6OECTV8gH3TDVXDY7dUDxBXnYQhqqI
SdNQMpfwxPtfXyd2AaNFIBWfCPO8Fn9sNnDU1HIShrEw9m4Ql+DcbQ4RuorStFwvsgIgsNK/Wknz
vi9Z83nfr3SGyf22NGvd20yKYxDP8DatQdrSXkuFFuyjeV0UkeuHgqPIyEeQcYKIoErc1AudxtU5
A5Lu/phwa3csEJ+FiHQjOcTU3jggBcNe0+xXJivzP/9fzYkadvIFmGjrYYzE3ApsA+bUciImIzmC
63SM0lp9P/X81mei5CcCqcU1b2p9h+bqXuyurUpDK9W3WEZkaCnwz3GkIa5uOcfRwRXRiODwYLoJ
iiJ5Ml6xrKGrvbiwEroWE4n3N7QV2+mTU3RJfMIo20Wfu5KixW6my+GpVizhJAywlMubcww3StRs
5jmvP6UFdCBfXQYcEIn8xVioCy7vBw2chADgF3OdtWV7wwc8Ct8HFkl76m1IpSBFAFfhQeL+Jfaz
mxtjhtf26qRCtHFmpiKYtBUHBnY7vHDLM3Y+sfP9wvEeXXy3brulavUqLI6rGw72KsFTQX61x0eY
cVC60MMVGKWU67sJSe3XcsK8JSsOYqz2i5jjuDf4CYttdYsg53yLPSUX4MW/O3cuDoYE9OKQWFmV
MKEhdZAZs96lirCRdg+zFjdjGw///uQWOe5Otq+lNFUxsXpWgBMNiiz+KOsL8zJu/fWfxN/57RRq
cAAsY89QSAI4g5X10abMh9ZL3hiJ999cfEC79s+Sf9HYzgCuBuJkxWfwBCdehc6vhMOl4gVRZO5P
YIL9W+Zh7544X/veDhzt2DVZtcWqNEpTlsSfsOKNpJLJb9KKvcuSGQOtCYdonZs1Wo9sMSOVGYrp
ZMs0Y4yKdRBQ+Hl4BbzIU/iMggzVDeohZHc9hLmMIGQ36VmSK7rJyS5IExf5e4RyoG34dfdj31Fv
BQspSazX3jRurvuItAT14THMxyZBKGpPt82B/kA5SQ+W0Jll+JPAiDkROHceWIyO6hZa9Qs4UwZF
CsO34mle9c0uSBFcLycaM4SxzP3ncOJRuddydwIN5hz2ZSbvpXpQ5+NPPqt44weU0Grtlb30l785
teBn4aiSwEnty7Z5NANxVlrJoxWR/WINvtAM1q7eZ2PtEXzBAqUFFG6T1vAjaMZ5sPQS1NAay+fR
3Kz+SljvwKf8r3Pf7927J2ieW4a7zr9UpduhyxAvr2dm9hVBBbhQmcRV0A7cUQVLpqQoWy9yEhzI
6Sk7JZ8WtAgOJDlVyE9FHTFB1dKEyyTwaEiE0mdi4Phpwiv3+ieTCONH42q44diQVJ9HcssD5YZG
pQTpjU7AV1GLc9QErHQpVf9UvDZPRDIniccvTTfIQoeDgqTq6Z0GI2RT+hXIAQoiq8jSkDa3+WnE
rrNmtTG2lJX/QMXe9nuDW3TeCMEosBFoXoC+kO1h6IEa6DyMq6F1NE3M/+D4SjlxfQjVJPqnUDpK
tF1g3xfygcG7Qkvo8yr0lXtdUE3EnYZ9sPJibtwQalghdcwRI9Erg7MzB7w2w3BrEKUy3YwEtY3z
s+nKJngsMi20AV4ZCm0g9d616Cl/4BEIlaPKMJKl7Zx2pZV5de3s7OVCS9f+SpfpD7x6zXiyfJ78
j836mDZrelFoK4bScT5F2NMBInJPDHeRpjJSx0XdrPPthblWZr2z1HZNakvRWM4ftnBiTVyKd1MP
PKWKBOsZ1nT6EIg8wvkZIPbxp4b/uzIffjfMxPhnzXgAt2zFE99z7SPomfjPuQRMD0VPHqAnVn/M
secDpcUM4fRKqmvko5ObWydcTk963RnUns4Nhfk/PvTZWtZ9RooqMWAKkQlUJdYAWOOR/atvpMbU
yKdNUHfzwNZ0z7lC3UnMoAiotCVbvFBICCNLP9/LNsgirCnntgtVSHDAAc+Phzb0QodZA8Dp3oOP
0IqfCnWCl5mvmHlU6LI6+4z1WJTm56qWY0K9owLtoMiGL2OlGfzgQO/GDyxPrKD6a8Ak+VmsSDuA
jY0p/sblo4VevqJqlQVjnh2rpGePcC4VjMPJG2YU6axcfstapyY2UT45ehOniHlBTRdnISxEeptT
sxb/7vz6pijkLebxx0EBakFUV1BaGdkurRgmajiWDDfk0CifpsKiTBDuRJ/9Iwt9xwNJlJCiIa8i
DJhYcka3Rhqn2Xv06v/zu4+Z5sk0GfrV8Mo5IlGKM5J3wJ4p0OjSvD2vL+bigjNEwDWMvOx8ot+N
4C+wqadiRkWCVjXF9Xk+K361ovuKLqFe8ezaHP873UpdXJdyF5V1toh7m31Sblh8prEuYUOcpi7/
sRzoprQIk4I0II4E1nNK95MtasAOR3KPoE2OBRTKq1TOKYwUo3xAkNmLsaZCYBgyVe+vYM2AJqXt
+KfINZKWyslR0pzA3BfaGqoXhA8mpdaAnXF0FJ+wkX+e8bZr/An7vpeIBUGjGtvNq6sC3C/dz63o
zaQvQNPgLRoEoHgwc68sdgWgrgkDWFngZ7TJqmdS+Lo5rpckODKWYE8vZu8HCATr5/oGyJyfblCh
T9fRfyWWkpbPyj8XzL51eYVteNkUc686SiSS8gD9ghdFDJOq/O4jfAIejgcTh1qPwspn+apjhkmY
5RFsQGspg30MVu7I5stCWFTN/8zTulvRmo8BQHpVAmSe02EvsDpEhkKNIbqQBcaWJrFHSSSggMHk
WC/OojjLGkZotXAqJ7G5FtZrXjpwJu2RtgBbZX0eBCJxlXQV7ZpGTUCPDQjN7tv6MPuxBa2hobzn
N7RbVpXghWVqYOH2+4OOlQn5BW+DT5/RruoEsZcYChZRPXvLSxsr911ykIT78G357MMFCJW09R6u
hzFlkWO64y5LNh4iNFtf5nPtuMJAwDx+g0IpOfnQnTJiMsEvHfv5qCWaai5czOgshv/H+t5+2ZzJ
Ws5aFzL8n0d0JMjGgoWoU8uKSaSRNUXC9e/fsjzTHuOamTvDrxn6vDPBnwTWzeNijFt2nTi61v+p
zgEZTUstg+28l4cbNeuPum8P76nBsj+1jDI0jgsxBPyUgNbvoBOewke2NVwcA5zONH8Hb2k5JyxQ
HKM1fvG51v95WQ7q3NgDRCRrx2ROZ3MmfGiOMZ6BDDFir61nqJ95Q0JWqyXJiXFvszuYrh4kkyon
jJXk21pXt0+fS1m3I7p3XYdi+vPmgyIqW0jX9QkDkSo749vNbi3PPohdH0yW7KizaZHcmV/U5Hc1
UA3taZKk4cChovIIo44MYdNe3+1uO5R5aIK6gknn5KJl1bos0iBItHQd+s7DcuKR2+Mdki5IwNo0
CzUm35ED/fUMHD4VJ4P6ph4txWrBA/Htq3v2CLfz1MIAHM0hLDVkooOHDeB5ixq7/2H1oBSHiSPt
9CgfnjqEhy4VwW6z1OMJhxeC5XAGktdTat3uIcAdBMLmw98ZzLFL3/vadP0xxTk/q38bwQ2NELUq
YS/nghc/+WQqmTBCWo4aDQmNfy3Mvz2rYe1zQ/6HmyrdX+h1/H0EAaT+XvMSoH8gU1t7NlzXPGUJ
sMxFR4bQlcnetFCg9Bq1has7uM1sTzABhkHkXVbfllvhb4VRsPsoUjkmcUE8uu+u0bdAogx0wiCG
dLKppfYvu+pDBBbYE9oJRM9YN9dnu1vtNP30FTk281JqHJvYYHpj04AEpu60aMaskIc3IAkgUkmz
xyLj5O7csFsTBAngXXiL3+hWX6xDpQegeF2P5nz0lfMzLswMCN/oeRU56857oGIPKwlwZ3P9diAc
tWmDb7CJTKJGhFVFFZVsoTum7mrshvTgLYuFZRkw7h+ibjW2Ef/P54iUTBL1HQdu9epPuRw7hnVz
8TIlCuhlWlUeyDquIhkETCsllLUzP/CNirU52Q8CPGrHduOfVaWGIDaiHLnucuthfOA/Q34BQ4ig
EJ4G8p8/7moB1mfnfcVzEwuAjjYXdlfow9N4yldygTdcgp+oyuJo368JN1Mc/3wXt+nxDXhAWqAL
Qp6V+9LPuv6kRdLkolBT+BwRGQFVOkL6qWGQtBRrCSlU6W92VqEjeR2KYQzwOaZD4tLzPgeu/+4/
4NIQq4eaV7/SyXxsElOdN6vSdTFK3U1VnAyTBgxAux2n+VglwQxRDFCOyWv6WhdS5Ko1dMF4YlEt
IJv68YUURC5IXDCX02qqGqz5k6IvXg6+3NbbGsCXR3SvxvS0mQgIvMgVF9/v5K8DCvT1qba/d7yX
f17Oli7u2aByarSANltCPVjsJdjvclfQUJ2zKdU3g4mu31k0jqORmU4yuMi9tKi6j7rJ/xvuym1K
91PGwyw4XgIDgsj/ttacIEYdWlId/VMpfgNNKsnMPDh8u5pQR+/evgcR5LvDQtn3ac1ZjshLAsT4
LwDtYilZU91zQIu7Tu5sWkw39U2BG/icvttbC1qmrTvPUH+AXV3BEEIvtMPO9mWy4hULR2XrAZTw
oRHnRBmaOfQpDDo5tEMxQqlF3Y+tqzjcEo/0ek48MgbGadwRYvewfVPuqZJTH9JGhG1/x9a/853n
nIHwr7vaxhq5WxxDHkagkRjmRujWG+tzl2YW6+L+CVpFY2i4dvKyzAg8NlHGmE7+7RED+m1a7Wyh
rteNJJlHxbPa08JVDJ8i3bkZlp/CetS73Dbo7NEWo+Xh1Eiok3DeAluXB4Sba6p4g8NYeO9PiyWF
mn2Wgc+kTxfBaZsr5TIp2zPJuB/8HQXLr+7PySbRLLDbkDZT8kQOrryeimeqKr7l8HAePgYAh4RO
8/CQ60w/XYe263U2FgJxhxCDsRV/d9WbqquZDNnUaX9zDcEV/Qro5Re+iXax4dyJODDS4xsTsxI8
Ruzorqk2/4YOvG49vXpOVaxzUiH1sggCKvifAk6RCoab73qONnVIIagrKjA0u9xIQeDBpwHjg/YW
QqKR7FgqgCyUWJwtvrV9oJjhRMnCvm2CtKjkKbII/Ix85zyhhITTuDF5rPYYI9haDgfAVZAz6exX
//TS3MVDI1sHgo9pLWZOhsAYRXiQfCbG3QmWcz93NCuuxudwSEmcnkp74zsBhk1fmjhZX1HD1o+d
4njAtJ/CyKHtYOLxa69s0uAlMY/RVhgecmgrBlR3IwlbF2F+QAn5d4fMXzX3otGFzRoA8dgI6tHp
U+viU+579HGbnqdv+0EO052LEOLfCHIExU/Ie7QkRSLtArkdHdTbCevvWNMCngDDiw9OimS1JU8K
6tHk28dbog2xL+6KqdeIUg73qA5cybMOKrcwV2vqhKp1qlg2WKtnWYO/Nz1j5eWaic9255EI9FpK
TjErzCk7kDboWBZmwIQ2rCi+8GweT60mtr2iJUcKI9PPxfRab0I1PGp4s/JmKnTzNvS/joS7+82Q
J3N3Ma7vvo60kVROwP1qEEUOttc9yQELE5cFkW0TzM5Pz2j0HPHgB2A/r7l7UsZqA/AGPlFHvCIL
ssqPL/4a3LyONfe++7DKBMLLh6qGF8oy6N72Z7EOz/ri9gswwdahuj+kfDmh6yQlZsjR42hlxoA6
ZwMxG/ll4X6lDGaFz7J/mDX+dg8AchSI6U+tP9tXavOZ7LFViPWShMC2moEdHNag49qH3DfxScfb
Q6uxJdvVOtNwgedMxeHh/e2bs3ouZ7UrvMoYaGdni3Bfjr7kyh2KV0IdNT3AYFhfW5hJu9lW/zIO
i/xnYzsiNY8nbVDi3jW+gwk8fd1g9FiTYHEYaOlS5p+Xc/IS9bvn8ZvdCw6gFR7NqQ5MBWTtArB5
hxLlBuw5lV978GFlC8TJ2aoib8xGS6cN2Qxd/LzAh89Mf8DfcZFdFNQ9hU7mWV7XVy9imwNuQWq/
C6+m2ojZc+R7UJcHHmhD91veYzbuxx13qygFB3PPUzz/CMYeV+Ru/XemQGWbIWuEowx7gzHKrSaB
zCbY+6WlqJBGi7y72PFQo83q/+RwGMzd6qmyt9ResfKCiS3C42ET06PxSkUi4DUT1ODBFsiSr4rK
SO9VpC8PvuXkROQ3HJ5OyVkGHssKzn7nS7tCvp+xKr3wb/APpmoetkuG7II4FcFoa5OfZ7u/6jE0
dhio+bYruqw0nU/o69qwPwNWaUcTJB28lrnA7m9SyJc3tatGXcFUBTixD5sHN2+EYqk90VBuDMNJ
fNFcVKEoGakSPRBc4YqKCljW68iTWFO54V20nnb+SLKXhxSRraNPRJVTuTkvGof+QFHTDgWR9Rwo
0HIkmq1nqVcy+x6RYb+VDcvvl3Ta7iZMMvWHymCpqE4O/+UNnAPt2kD8WNzVdocJHHULpDYo7hsV
47zcgXJJQk/Uuc/Mut3oKOLOYgC38S+WxfjmzApbSEMlDBeIiGX2o/hq/gkn+hYa+j0waBFN50So
w1ECa1iZFtSrx3u+UYcQ/Z9ldAhaBgRyQgxDNvgsQyqnwvbXL/tN7pnXmievoPdQ9nPvcsgzQuXz
aDOH0AJ8/eIKXUoCvRKNT0ooVLNbEgR3/QW7/jfGiFMedCberIvftVDXzByfSED0UOyjC1fLesvl
ghNpB+/Tv1Fsw3R2MrQgXUBb5n5F3YN0HwiaknRnq8i7cnGshAFkXv0xA1oksdnCw/9o6tCRiVl0
XKOrN3UcTAjm3nvG90G7hTJ0HmZFM113unTjRwt5C+C94tqIRTDbMC/cxZc7NlywadCuzIvmx1cF
UPW1E7KmTawgs7qsXMjuFSl51Jy4plZ9wCv/z5IE+9zLktmHO9p8QkVDdCDTiGi+sG85nxap8wfN
V5QfQatfDyIze1aztxKHFKp+abGaClN2Snzzlvs0BbHeJPAGuZ0a3SvTiedYaXmKZ+oSY+LlPQWL
lnFjbKWqBqQfvnmrcQxrpsT6y1XaspGlRphWAaP+OgI2S9BUWBTNj74CC523eOzR3Ru258GLS1wb
F8c1goUReNW/DX+zV6ZwgAB+y8uThLLII/tmYOKCMuSgps17vTuNuR28pQoS7okcvpyR5cHts9Ao
d7frlmpeZHUuirIIakuYTHI7uIqrrK5UHtO7Yc88obWCPvFPFawgkoTg6ebeQsCG3ysBfCSnk7h7
bjySvrkzEFtDqod4H99nFJn1M6gwOBKa+EgF3z+UE7FKnUMBUvJn5Yi4B4jOIuxyUIUnARTYPTof
Xo+FpIwBCl9Y/YiAHymX3LH538qTHwYfC61gyE9nknRmkBfd9BReLeMX3UijbOlrHxVVKPD/PhTt
FQv65NNCA44fQA8omWQILzpSacwdI7WgDH0VpnTVq6hKt0tswbgGn7b/zfOtlkHitV+JmdXOcc4s
w6qMcFc675wmsl8IwqTuPQrNJx5bbjXjbksE6CcViYwBzsHQc349y3KHFwgK09vn2SE1Rpve/jn7
VqEHv/mq+gzaANSt9hQsZsUtvx83vwCvSvMzXUq2Dovl3o6/etQtf9ItVCTG4tMzakqq3MK75YL6
rLenAq7+m3BvHqzvhFpWYzxti2HiCruhednsUCsq26NcrzYHBCyJzwPhyNlDlbd8AwQgl6pSXBmF
+Xb5em27fBF7xmjh3GR+s00cbMxhavN4wKAqKlK0rHw5gpulQE9nAVkOmzZ4HYKFOD/gVzFdCvCa
2dBu3WgJnVmcV0zVjepyyzIkmSIN2Q2MUPvyk0ctoqS/3Xz5yeaLlAPnjhfakSWoqVKZw3DPy6Rk
xXBB/Kis688bPDcFpoH7I/XXvVsM1YcFmFHk4MfYFclQxxqUoF35yeJ2gr9MAUT5267lsldFEJXh
7Y7V3H3gXyAA/bfdyXdkdHNoqQ0uDV8iqrppm1jGZJMCkuWUrsbfych1ZaPFJPL1XUgwn6+vSaWV
3WCDaCaoQQC5Q+G93B4wjrlyAbpyNMsMtuPl2kop3bLqacaVnViVZ+K4WF1UDnt6u9UA7uFqhsJf
0a3o2hWbCS6mVKdnlgijTV2GwPvkAW3tB9fiszSz5ch1x+xitiXaV8x7t8plo853GC779qzoKanN
RIQo+BnR7TAdaCgi+ZurcKKVmNN7bMbgNPolO6kl8Qn+QBky4hgp0pl+g9ul20xZzkpbl2grDPSX
OczW7sGgNrmUzZXdi9uRy62loQ1Qgfj1x7omwxiQA+Fo4qtnG4FsAUFZAAOtk+tGOchAOTCPjmKq
jMpCZSYyAqbSkldk8K3OMdiw0JG0dYewpdlqbmq6illdd/GFzArHoE7u0svIRjpnvGMdvJgAkO5H
tWssQEDS1cdd2kJnJtQNzK3SUG/ldFJHllqI2QFCePXSKUIzHq0tXSnH2ZEFhlzgDG4EExLCb5vg
bdaEBQKE+T0NSd6+5S4iYN+kIT9TJWzRZk0XDGG3exQa24lRbchJRT/bqwgHKAxfHxFDr6QgTuVq
2+tZf5/mZZ8WnuDQc+FjsZyKes3lPwnCgGgU/FUEaq2LYegGJYJ/qP1nmIdl+Auhpfz8/cv9ZrO1
ElO6Iqs0BOTEaKOcEBnwozTsxqniQZZhoHCPNjo3/A+MNc6/oR5mg6In9l49czrf0SJfe3XrWQEC
6FmbxLmYHL5av9IeYQov2YYrkSw9MrVy2tNceoKE2N3LyU2Rloug74Kgt3NTgHfpBFyaYsYf4o9U
nfNmT2awjdOkndn3looI5nCt65ZW90cg4zJNKFRbGupcfauJySN8CcvJwss8wFiDs9YGvF4BQKfG
enYD6MScaicdwqkQBQ0JdotMtndEAsML963XGVnbekyyE67N5KbM+W7jpXljqb841mYrM5TDjRHi
jKtGUjD6LPQow1u+CpOBn3COaMdHxJppb56wqinK114BMPPqO+mISJRCWMOhuC1LcDZJKojBlcjo
pc6UWJNrYRoGOL60iaT7AoFyF1UuljjnL3Gi5h2jOBSDEAvy9BgdH9jjHXEUygRPZe2yKn+i9rqL
M5F3W/ImgLec1XKXka56ckHGWErSLl2ofweoY250rsgqTwqdgVwMaijMfBZWShk1OHSpnx81Sovd
CXtPwS4qYWx7KP8nOhKzBTRt1TcrOroMeqfOUTKbgphpe1MaoQoa0VfeBMAsYDKxj3CHIa26Dmpi
9xSJn5OtiFV6mvN2TR529+UVBP0/Lk5gJEVNs9EvC91vxO7y1Vwb6aGzRol4XQU3jFzRHnLlGrkw
YQ/8QaI9S9mnyanKPWT0IbBott1yPCr5LYUnmd8IO52u9Fq7yQSrXJipTqJjPUNOiAHJsJKcO1bk
AO4hIjXPHo0SOh/HSConfRSa6QIu9Y/SFMAhiZe33WQxWkMV09LW2mWaevqd/ZA8Xk4mYJBAaudN
55Y4OOGt/o8pXaZEBk0zbJqgAC0GYKyFtX3Mo+pRQ8uCMxPOexXCKcW6u/GCQiyuNPMWCZxCKEqF
uOUoYrEHyDXozQ+6GG6JcLqEV3AooCzQMilBzr7C5WrICFzfI2+O+s7OVMEkqAVhfSr4t6OGqp5E
nc5q2BjMsq4+JjjIgeZtldPeRp922KvO4rI7mcsqlb4UuaIFWkc+3+TKAZGoy6hiuZKsamy6yle4
c3Xb0xdQ67fc4mDmCJbL8YCL2S+u0jRDzc//2lIYlZl+tMFSA03AOT4mNDdeJP02F28qxpMWCNFr
0iPXpd5foeOL07SrgLzLV+p1mRQy4MSxIHNUV4QADL5skLd8g/E+b8dNVTRGx+9ZTgDENbNs/L1C
so0gm58NvpeiBbXThqBKhPlwx7slq1RGIkpeWSjz05qb4EvKmyXASOIHneEVEqp30fPM9yMiQWn9
pBcq9+C5Af6jUxBbpclRaJqj8zhb/CorF+xoFfb2WB9C9a1Die8C2p6tf9y1cGDDmkCxpfboEsr+
kXjGIcrV7kc+nsd1+Gm2CUT09lHvYq0dz6JSOj1gHj/2HtdeDMbRJ//V7BwaTbhmCASpBu786Xl6
ixFceGi5E2nHDAk7TeVmVxS3Vb3LyJsawgrp6x/4gyBdOyaCJgX/hIfyBnGeOiWV0ORbIERsjOqp
nDMI6vhkBsBTSkM+uLCL5bmo1uCamRaATkDerXN63yvzM+hyd6O/UQTgnyNDBwdgb5n7iyAHj2Wn
iFpoSLz1NzNxiwaKPCpv6W6SDAslMHr81Kh3oVEuHb7At7VurIjpUlSQe3nTwFmTHte/SqoiyZ82
heGoBTmmayZbGWyKPf3tbXPludqmVA5x5Xm/TZHhvJYF821vRr/983A5zzI+40XUUmYuMmgh+pWN
Wpz5+HucfknWbnLF1iKrllumHPWgP314dG4SXjHnz83UTm1L+vraaaxtUEIf0VcupIuA8t5YcWnh
NIcKPAojdgCxWGgwc3fsmlk/80D7O+XSQE7niUiHkVgYtgwN8nz6QVUzMDH0JuWPr54XmxvG6Nd2
RQrMhlk1kcD3LAvrNb7VBwKQJMshtCPKGViG9o55epkDcmYZfYQehajx4MbNLYEISed4slDkFZPI
cWUH9TmJXyBvsugGLa478lmDSRWQMKQNMMDpH8dvEeVYrnhg1K/S6kaw6424OPs8H9+vwkWMrb2q
PZUGSvCDv9HHpcTSy8Fhd2h7H7u1xeWx/21XUJjwHmv3jUzqP6OWEmQDadfE2OytMWbrSjq+0m60
sC/GtDMKohAzct3dK23PRHd7yvcBLLdnUofU29igcql0ILJuwKJOSNjg0V8S0aHrZV/hjinKcogU
LdVFE5Rb1VsxchfNZaBaucmni8L4cJMYOK0ljW5kWU/oxJGjjZ72Cb2U2EDkLdsfSfmN8Hrk1eFe
hb0hjYUgtqivqfc6/irVuKQFBB2dpES4EdPk7DvRM57jhEjNWluRsynguHMLperzFdx8IEAr7ENf
vIP06MRFrQXx1ipl6vxaQgpVxm9C4D0py3ked9P42iRhrBOjBc5pIRvKki9j/n6y6j7n1ty1BAbe
sEPx+tRa2gUONol1zh62wzBR4X+O0yoETwW9E0M1S/Bx7CgGIrUfYb7QzBGKG0NnJrhf6mvKp+/n
Qd5l65OSukf42o4KP3QzhaQb2n5HaWyQq7DSY8uwgmtQ8P5Qc2ulPgxShv1EBfVBeQidTdbCrA6H
f0yCLguAMjc1THFJy2C6msxw60VNZ/kKFGheo14aHDx0QvoaXJKha7M/NPW3heYKp2VnX9wAkNDV
Ry7SMJCeFUwC1F2TyO+xI0g7X1z2ft+YGTA6QO+ILAIKrxix/KoiGYkX/LJNKrdKiNQ5A+A0QEBC
mEpkQqRtW9uuISONlmoF0pRyVhI1yHmZEAVGQfgtoSnuPFysayQ3ZcNKuUY1PoYHApLWTgLMDLpd
zeyOMMSxq6uW+QNulA23OIikbEO/huSr+069FvG9pIwtIfYqvyEoKSgyxnOILL50nUyuJWE01ONg
mkYO35fWYWOcfRcQFsPClsSRwEPOfKHjlqW+WqitOLO6UUec+6xmdHPkRkAfYC1laR7scxmwmiG2
Lu4czURYbV/PeuCNOGEEXZ9pIldB1hgxnehSDd42/BcFcH0C/hUJmx2OeRqJ4UYxxbhn9OGhdwHg
GqhkJPj5/LllLzxuDrWHCXI4KCip44bu5FQUIV9A4w3TGalgp/zTttpWy0CSOPRYGEx967U8QCqJ
Rz0+g8A13vKNqkdPnUFGxyU3Mm9AQ925p5mzvA0dBHE6XbJ5g6K6e9rD95RlsjjDVWEZeBEubVkZ
f4sowI+hDrRl6w+zvQtmpMDETncwFe6QN1A3hgUWAIp6GsgBFs5xLfwoNfVNcdtafCxcBlTSSj8g
mqFM8IOVEcXF/F97663TbnAIj7JJo412Y1PGw84tt3sr58R3ETRiFhe/cKiLIoapbFK+bbv19A6b
VAvZa12nsJv70+ng12Bp1BDj4mqzW1+87pGjWRTVmrVxY/HRGlJKZXESglQVi9IHXZkHgw0FMCz4
70mI57ZDEHwx7epJyfBohI/GiQKE+WC0FtmYHmr4SXuSbqs9GJnnhbkMti7T8m25VOeBRxZ/obV2
kIBOiRxpDbgRjOYWYSIKuMZhOQ+jXRF7pJQSEx8v+QJACHo1u/vvRepK1puwUvWk9GEAJ/CUS+OT
h7mxeFFphgB9EA80JBSL4ukutFTLwDkPhxSQYF+9zSwb+eAuquiuBJPwFMqzxVZPDUD1w0UkqKYg
JbkU+uuoDwBddx6iJCzGIbwZqSn3sicp4rII+j5dKe/pLVUI+uxRWKuKfjBP4B7SE4ADZkGvfs/I
FBSKErXpPOUBptjojxMHEPFZYbI2eMLTlxBfx3OlvIsc8mFMWa556DnoUCZgqrjS5c6lrfsPBIgp
xMCrlgMsPxojrNKDhexo4mVfjhEUViA4uCCTBljF9HyvIb6tKz+AbCUFobJegw8aI0z+WLlll+mQ
eXuzeAeaf9hzC04wXk/M1UgibPetIjE7V2P2SrFg0mpI9UXUgzyORcm/s52LSnQ1rdtJgsw5rMdc
xVcqSgiJ8PJVAIx4C85ARDXGiWP+PLPKrjvuMssaCc/YiLIxjtYGqNX/OV6chFEU/iEhPkkNxWf7
FEt1zLFqwnf0Ft8zUzhzsL5cczOxN77mGU4PZAYY4nEKQ7jgMpZZeKN271p8bCwIXd02ncs9+flV
z+FYg1i06UEh4FCBOe2TWpZWRL85zS73twAvw7CkxwkBQCMIQtqLq7uha9nfGkm6dV7jkERDVPi1
MHzC0zaSaIfnvkKJek/1p2eQ8xHdct2aYdSc5UMiGcMgLF2TQysYYqk9StRyJi5Xhr48Leq8j200
zfFszBYlbBRYfQReQOGyL7ZMDsWQc+xqniPhDW8drbdMoD/iCl6TnFFsbR5oTY78CdN9mnTldhSx
lVp9DwyPoe5qo/yUO3owO2VELBZ6qT6o2+NDg97mutU5MEVu8EgpSOymkbk3HYPtkkgLgYkTeeQW
tVWE3nkU/YFkK+zFbGhgXtfd8teF2fvt6zIO007QJYNqLq7L9y+omwLUVFtW1z39gQ7ArM6J0ZmF
7tg8d+cxtO5UdZNQfkuOMjipEo8qpc4nUAqmzkGz9rGn2U/ahhIRD/I9xtPv2BuhO22bEyQPK/ID
MOSZL8LNmcqnoazbuWKlNGkkG19aOXcA+6YEZWyCGayexFW1F9Zhgc9o9CyNatU1gW6tyFcurlhs
1rXeOFxDTvTY418Et5XzZtSfCb2BF2ot6bDW3U7nCotelU0EOSuu2Wy7tXGYZCH3MPrRRNDKr67F
p1VtPjbEjzOzEoen8JFYiYUGOhJdv9VeRWYBA124cAc8WhFXyeBFH67oFjb566ftZeZ/pgd6ZK6j
VBl+EgRyrcrEroKhg4wOBfcj4cdiptwRYn5K+agjHNpnAiQbCQoPx9nykgeHAPIAyB6n8PgkiDa4
mPVGLeRXFH9B5FRr2xHsn484zz52ur8uuR+BQdE3iWByR6iy2r6PZIsnEGmBueOXwmXaGPBCAtme
QCG1wfM+aEf/y3LkNtgarN6TcQL1bweasaDC6o9gqiV6RWk1isDyTWSRR0MuTv7pIceWU55UnFiw
urBhI85b6zh5I7DE4TaxVCnxk63vAtg0GUu+1AQPmtu1nQvGHhk5zXfdNpRmegxcKcxH1iI3mdNb
tMGBPl19+RDzIWkrmSOCUsf56Wp/YYAhIb+ahHRBCMaaXrA4jTtAz4W8vk0gw4aSP0xs5RAlW0+m
Spl6R4vvJtZI+0zTaz5aGXlRRvbdYIidRNpEFftQ8qYocZ/qtstZ14Efhp+UWeyHwyduzLMhMQvM
+EOoFZfLadrHLE8bNFgPWVoc+pms0LHJocd+iqAIALMEHbkwGrdDXNoWSeLT72ybD1fTwCfbSO2b
PHSaz22XGRE9J9LU7s7eFhgs2hrjMg5DxLPWP49iUmeKY4vSuYuUPV8AYAUeh1Zys8DkZdK7Htqn
RWtRVhR5YoQhQ8F0ozPQOSNlhRJQJh+PU9YK3SPkIH8dKSOdhymTIK42HqkfM0Uq+Ak/0MJALaBN
gqmO7ulrYSgcsADSnHQmvAuBtlEz59b/E7ul4oj+FYZ5kNIZ2mbjxZbTwrZccGWpGPtazDsXAd7K
9S4Zpxfx2MiFLfMLKxVL85tuB4MzZwNqtrMT9jtt/WwPSLnw/Dp7DGqqA/OpcWc5k/viZ92UCvFE
aiXfGpHEkakcNQNGB3L9ZFTZ3jLFEsNmR/7xeZxZGFcl9G/hUbCyGVFnEsvVqmN1vrLd/FQkvqqV
liD4Zc35FS3cOHCGVxX3icsoHd5nbxsCbpcRODAkOt+8906yXvu9skAh9J7AfGPT7gEvGfNYDpBR
28GxOwIukEBSmvU/zqaeFlsF05sPsOsd0iEtqOKjntWa1rzRNDRFx8QajMdZBHjdvNUerStVjLpR
9XgUwviIucIi7DaYklfPuabVXl2DkquUwf3ZDa1aoh8AI0ByUNiRq16Snm6WQtjF/9kupFFVmk6E
ugU3KxkJQFi8pPgbV8GFEIgKJP26tGx9Gl5vlNkNwbQlMHwUUw95Cs+C0lJwtu8UawNTS4n7T0Dc
ghsT3rw44rSlwlaFdumoG9pthZdpmvQw9e5sfa6HyyW4UVvVtPiKhxxlaC/rcBqqOUPBDzsUAVTd
5eTQ/yC4QzmLYre6To2SoAxd6MC+8BcKDHm5FAmJ7JQn3gDBJ+JC9Z/GPAz9agvi8d6WLk3APhRa
Ek1Z1d6qHDZ1P6IOMMYz39HuvYd1vn3N9m6O3C44Qa1u/Tqblf9t1U60ngHIIa3gwtQTGZ6+ZTK4
+irn3u3V5wJlRwOX7kdN7xVQPaZA/SnKHnjUwxoc8DEs9T0a9ipQWN+FYCAnIi5BXedZhzXK6NgZ
93qbTOjEXSzZebvAOe6+buVQV5I+W+w28AckcXXeWUM7Q5VzVZVRmVTESBMsxVeTjU5ddGgwrb8O
d40DL2ZhS9Q/cQEPzLSu5FKHLmD00luWMGaaYqJWECgGIu3oLU84fpD3vopQA5WziyES0HgiegqK
OG08EgjB7ijPY69umLjHjMFdJ82Ynb6Rw8l84se2xHs9QAiAi72sGVi/2jBAAT5gumQLc2upismy
gGLqPa9OqJ9CwEC+Lyc7i9zk3kB1gTgEqDW7PvCnIYSajuR1gKN0D2X8MaEYUcr53/sInw2/UZFL
04qzV+Kv6wvPg2g7oNOOhUSD8wmviah/vYtV9ah9N+BsXttq2KNCNFUdtvg0gvjFpR6GoSzksebY
GHl7bHlfhFY++G6f/3s7WrcExeuVm79VphZtKQtsJOVIlVB5dGOjkla7jsPhliM4Uegv1gQxXfe3
wcFOFq4dboZEBzAinGVymNItz0lDEs0OLE0GaDElhwtR3KzYwfDF35jF9AejmwgkrKTa8IxPRV8N
jKNigvtd+d+K6mSXRmRMBdXsqWGgeHQvVtn8bNKBTFHe0oyRzQt3CvxdcAylNOU5v3gNCeMIfSdf
evY6yxKpLskGL0YrIQQhZOpgu/bxcjHhUDBUqSa2YRKRdkSiWyqWUzO9j6GouULKZsagOkSOIMIU
zvnHNh25KETsi6yQQi8unkMRLjdyDLneAooYgzQPVE8SXLRs8jASHtlHS1nXZCQAX1qk5A6GphdU
/R3zBAveoKWqFB/JaueXTttC774fxB5rPXdHo7jzXCiD3tAqCqhbSAZgk/UPFBVt5qnzR0l4fL7E
h+EAdt/9qcfuX2x6gbq1ZA675JziFj5KCaeTwI/Na6IpNw8EMnjqtPu1rAiVgWo9VIsR/Lre5OII
spR+Ten1X5Z3BG3SHfFQ9cRnlg94Lu9ZvtKNnq/HktMsD/mZMVX1KaTZYw4jWcVbevTmE/bPVmtL
681f6lTr8n94CSJxQ2SGMASUpFNqR8VMMPhgrIXvtRxw2ELOtCP8Ck9lfT/aIapnKesKdiO4HAU0
9MtvayW0Lego3UHkPKr897t25D4+pw3QpS7oBVFaYT/8wf+9GLTrhE5PgnQa6RurPjjzWIiJC9I7
O7cR4Pbwf4dnV5V7i8NhLTj7YMWzwaU/tIJwaFzbdFcrgqn8Tb0kRQQsLPJtz366QLRkpFov5jhU
N42d489e3O3bigSl7G5TZIszS6Jxjzv0/E4OJjTKao9lnN48t/IjiEOr4HppyX368DrzeY5yfNfZ
4pDHDDxf1CnsOt5ZCSi+oGeGE/3fPHaGD4akPDwuZZWd8CCPA6STrXQKtoPYs6HY+gpLL7TdJnAC
TbxhKvIUiGwaezmCUsfi6JI4/DyRZdP0EA4PPUKMKE1tYo7FQ1lEoMCjGaZ271UBU1/iSXLrZBLv
OAvPrDoyxAdVT8ha9znATBlY5Nc8Gyejyy8I17FZBGYO386HCWroLS/f+HLqioAwIivQSjKt8tdp
bT4IDCgKQAc3YTTlF7HSEArhtNmIY7DfAxbynih94AqpZ+sN7V6vX6+KdVBHqCw6IQuo9XqE8l0J
zG9A1v6mGEHjLClYdDylICNnnYvw7m5ychLD7INE5HPgodIlJIWIZVr4PKhwtgEqGMfDq2k9iWe8
0B+bMIU+3MvY3X0qc5h8teHsMRn0076nT5DNbEI+jHAwHkEb3bjop6SkeAVDGKUc78AKbje9UGEU
TmYoHy97bu9omNvx5GiLNh32/CvxH7D/rmAWPdYR/WKUTbtO15VGnDZq2XUP14xFYUmU4e0F59jc
hLagfqoS/guARXFZYIyTqvfw5faAsL3uuGupXJwvDC1AbbHzTlaB/gZ5VuzoWSM1WD0SwDXIouLV
xlYTMSRBsM/elWtkakSs0ALdZezH4r+Ol95NFvhhJ02yN5Edr76INKzlxMQ1nl0fzOPpffq1S6pL
Np/Ys6SGNSytDjyeYmQ1cb5ssAzCN11EODopWRE1X2xfAgwQt4Q/abaCkkz29mJmpWHw5rxT27S/
AN9aFHpCCB9ZkKfpT8UGxLw4dqku6aIR+nGt+3A2sjXt9VSGUZQLWKJ0GEJejD+uEmmlov8n6yI0
rTnm1gISq5bCJr2xnCsYX3kf/G+togxK/EEvyDrC/6duZ+Zoi7qkbEOl+vQncJdRZrr8yyDFX9/o
ko/llswaGJxc9lgjvAl881DDoU7/hTi/d/E/bmzQ+3MATWyQx+P6HI8cwxMxsPFHij9y9bXapk+n
DkVinLG/4Zthp7yekVdSJ95N5j3R1IgtuyJfegf/zC+UgbG5BpzpnPWTgw0CRX3hW70StMo7PC/S
b8+h13bG+ie59GXUdS+FnoFGGO6MaH4C2zm5TMNtBOIK6FrjFmbjUWfVmQgpuliIlTVO8rBS0Wgy
jpY32Zyju38IjMQd98SIRsHhv/6CpeH5J9AbNE3bbf2Rhx1d7l/m9FmJ/B1El517xOkDt7C41ach
I/Ds1ncphAajHuTCI1Wi1cIW5vgvM5VHkGASHPZ7zc/QH/56EoYxrJ8sMaZF5wxb2QqafCu6drM7
PkHp40+uADCkpKdH+OthKN6UX54S1LpUw7m4SBjBndcz2v3OCMEhzXoABaLN4To2yqEi/2vjFr2B
ptPqUxNtrd0aimHBIZXEmNhy4XMELhumtDsEs/Pup8p8R3xzJyoDImKI2kAQU4ymfnogay6H7hJZ
oAW+amCIRdr2flyrlIkDCqMO8alGwjclHAo8RhNl0QY5rbWGB8u9kduhPgG+8ur2RqtxXBDT0Fkp
fmS8GGtFcP6fcS6W7TbBzP28OveAv1c3QO410F3jkholB4Iaf9xMM8yi+1ASvW/1vcM8F5YffqoM
sKDTnkkEP1fptvdkrShuk22DRFPwo7fYo1GG89Y+GyTmG1c5DtJtKiQ8Dhcx3slWdxAqy+lsjMzG
dPj3W8FB0xBGEUY4qlye2gpE1qaBd7u50/aNPUCEGV4qOep/wFdPJRdsqcX+KgGeQmMgTbJsem5/
HJwrEN2bNNCcA0V8mdMqXayO3916lQmiAbyWSV7fbJuIFgg9YBokgZOypdgVmHlMcZGecrfM/IAE
4xbZlpxhyBjzwr24WNuu0hMunPe5Bw731vvR+A9Uty1GDmvjm4EkCwveATG8vj+z0Kfa+2nfPfWe
00SQIAIHYa/Dn+clnuBLbyiK4SwgsUmU8fgksdC/A4tbCc8pels0b5Ir/i6AbgoZphXsk8/M2+Yh
VKCynjtbYWwivEGGPX3eVLO5p5TuzbQQ/G/MX1bbvFSOIZa0EftXySYorRAYxoN+orZxR5ZxE4yI
j+at3m5EYingKF+ufnyQLx1nvfZ8lLX8G4GW13eTUngY5mXWj5nBxKFJXxdkVKZW2GjNayWMAjmV
u51byxHdZRGmm8BxJ79U+0XLrHzd2v17Bn1/Pln5Or2tkJVwR3Bcpuetz77U7hY+ww8dkAZoOlfp
KyANzDorbBmso8sSHG3k+kJtUc+nyZVU7C0SuR3o95sXki9fGtoMOK52d3mBfbVxFJeewG8qawJ/
QZ36mvhKGxKsfpqmzKyj0LldEr10XKzJ/zlAg5X+yNY87efNmFby1hMKjrTqeZxfFHGG6kjUxDDn
iuSnhlJ0b7gZAe9O8wLe5d1KPnlR3ra1FEILji0Tt5ZWgjXupTdJ5FuXtMYzXCHWnh5iHhI8a5Gv
/muEirldajL5Ynh4GZTif/HrRTB6PARoMDscQNO1aJmitJI7vjBGOtyLMhn2aajXkxrDklLnnXlB
h++Sy+SZ8W078JohytJAHzeq+E9ZCVOqP0ooQaySS+BPLjTuBAJBMMoJkjfZxPIlFDvukj1/E8VY
d43505wvOvnzmVjnuR79MqLS2SvxCrQbeE6HGvyeudVAXEWrJ41uNtrZ9741HYgzPBXTJZ7ztfCZ
G8jSvZOll3r66jcoMqIaQ6IhDMLUP7hV+A1Q02cV4kWnLmrt6YkJ5qF/WKsBYhbyqKiGwfAorlDP
myg6wRdM9wmVxmpwA/z8UgDoKFeQKv6/HgpOwCJc2qJMS9vyOXzVgOAJQvhQJvvZ3uL2V1P8f51x
thjmgf/4WXSAYpFYs+IghccBbopnuJj/J4KiXCEq8SFz48VHbVgRIA3fyOaOeFplTO++I98KUat2
yhopDB+NZ+biWz6Az10DIThSjhBDX9bSEipLFmmX+KJaN69VR6+b4tzkC45j5p/JoqpB/NmglTS6
OtPhxcgxUI0RuOSii64X02Bc3rorSVKIuFolon53IVoXZMpAo4IEeWTT96z9m69MVYwQ9O9ie9z/
hAATkuAKvS6nLOSvHRhTQh09/Qura1iHZizdMhkeBIR2nT8rqUr1Rn9rBmPoJfG+H5CrERTAqp9I
z2H9gzyjt/6UR5gUBRrn2dvNzWIr8vDqsOJb2eYqpTGHRyy+Cl+axGiBU69KWsBZ7mpcDqTbsr+o
fEO9AnMYIg52fFD7AET+FVOnJa7YPAx4T8wNdb6+RwTY94KCwhvIHFfUwfvVoDgSOiht84xgDFl9
nn717TSC9C5Y8s86zB4TwxKUBDAhoPswoZVWXq3roM9wDyfUdUWLZmaj84crNn046TTTVmq0I3LW
EPOU3elv5wosdtDs1KaXzWVcMJKtpdQuP/j4mhgiJZd5AzzTgsZnxfKhFo5LsGWEioLX0aQWDpiR
cJgnPppK3zt/1HLqkqIblJdw6ih7oj2P6bxrBwgCxT2IPbJGIwYxzlwalFIcDDmZBT4rXDxie3sy
f31Gtl3u4Tg6kJ7bm556WOdQh0XemXS67Lmwrw0L0D5r3VMafdd3H/t7O1icwC9nnaRUMqyG/TdV
UfuzH5A7p28zRirhLARBzxoV/aJAUlGLW5b7fzEyMOAKB4/lKrSsIa1ZmjEb+fVKEWDtndwYXAbF
ZBFeg8xfIMgUpwinnJt4TDBFBO9ZzrrpU2xGvhQEMXEmlpOn8pF6RoaqF9SwoL8WmenbhqUjmtQm
aCHgzOJ1VjRkE7YIkp1Oq3pHCPPEGvQuLt2dFjIVu+RBKNRiK/14POmSpcDHYTXquJgb8t+gNzb+
cwOYb94rAfwlK1lqAe78U1XB3prWoePa/OUm5eUqgqtBkvJouBwmumpTP3Ef6C72mrAjr4NlUMp0
7ADut1N/P2o2Pxd7IPVWCiYMQFPF2E1/YswKdGM4mrmBwm9Fa1/ls9QINhFgBoormTw3ZSnfmC8Z
ATXcz4VfCnR3z+2uAvhINdOdC6P2qKPWe1Eisy22lWZYwG/MPKRF+c0ErcRTs1gd8AMAhr8FQzso
WaYAEuXfI7NBRombQaoYyRcms101X78lx+JhbQfrFWfOzf5CXvPzzvczogfcIk6cj3gjrS4En263
51sv3g5zOS/LIUk/FxCAdLja0Y1+jhqv+dkH817XhF9ibIdfDloH6QVlR32yJselwEr0gRkN5vyu
nW5thdBkvkj46GaP+skh8/MzpDGr8swQXAtfXgfv4YMWPCkJMMVRLcBFCbKTmb7YMwEs0seOiT9d
nHX7zcNWVAd/4HtAPZOqYxhFZPD5PJ5RBTLTqRXLB99HyxXHD6otkHEoSTNK3LmDXMUG2vr3ewr7
s7k+PvKNaXJs09mpPkfapBOfE7rCVfFONNPyeGUvms/6c3IRRjBhHrc/3+XvB93+w2Q7dcp16wsW
a11B5Ub4PtYT1634Xqn8ojowSkiTQRP168s+k8LtmmK+t/DR0Knbqn1rO3as/aKod8MAc3X/t574
EEezBu+CUzchilTMQN6nMCAoV8qv7240lpL9OgUC3tke2yTbWgMq+cqeUA4vtRnI2Q269jWi5hYW
CNZ6s+OdtFS/r5T619UAG3xGyuFtrTudnXTLev6iAuEKW/qFiLuFf0tT1PSCVVBoofhLC5lysrWh
LOWp6ytUU0iNjpBjPQ8XrppURRz5WiQlZYITuvWrz5VRWpKWEwmKZQDLTcnEH+IOt49LPfmLgGUM
HJkPBgMktiTO8H24Q/s3JBnDVOxp+/YDYCtcDDfvzF2rwHbL4czcgLN3f/n6LVzZ5Tja6QUPf5U0
OdsTlADAluHgQvT3eJj3gA415YvezcHUR0OICgB5+Sv0/0OJMT/F4sypYcBfVh+AZojwFcKgd1TB
ARStpwjaEt4QJCqWIVuZXSENKu8P7rNFoXQ6BzF08F26Ugc0J7K4vATQyDUqAWW91iTt5Ab8pE98
4+uMVcn+bf9Io/vUHY/R5fObFp8TRPj+vEtu5wHNXyZF1H5J2QSfF94harcmSIDalBS9WeCpOLY/
U4suTqifloYMVkog60qjf6f/5Ir8HXMiXwNKemKDXYHMLE+sTtoMQHLZMw5Vpoi3XgJ/37AV/Vwg
AlNnN8e8yMyo/qRDbUoS3nVT/eEFLAsB4hmSn7WKFPMyDtx5s3HVf8shSBVml1lk18sWc0yiVMVg
BswA2SVvITG6emPUnAAJlLr0QyM4eIxqQ9BPUdrj0zdjzN/zcp3TE/8+q6iAihLZIADJSGJwDHQP
wZM7rm8QWb8w7t4l0izBT6TOuf7M37anSxkZ9sqqyVoj0qfJXWgOE7EP/fCXZ1/gxVmfj6vA/+7h
TqNaYYsvLHnTYm0MWCpRDqIugCfzSV060SrCTdOiNVwThZ8kYlDCgR0l8KljzF6h6TJRiy5E57Ak
8L00BEtq75kaRHL0pHM4YHU+2nZ8NVzEqsyVN6AZy67YXFfpcA0eU+PXuZ3ZXm9ePL9ADoQi7LYG
WUBqYFDkIxQyPWAZxD2xMIa3BCKBI2yvGczBWpMrF9sUpdJYiuatjFCG7RpjU/Y44ntdAaXsP8Bj
9jq5xpe7iF2idl41fMg1L0foNdvRQwyQQfjE/cBvss7XtqR50R3uc0hdlnBeWWq/ZiiAv0xOqD1j
DPQoPrm0sDNZnfxSYWYGa3/BhM2RUiY6U8umisVFq1hrDYH13QQ1YGQ5X7yb5mV2N52dSo7yeQX4
Q8ok8YJEFmu2OIJlPmUcc5Qiz32mMYNjy/AlMOdkF7Vzzprerjm6TiMT3O265jfLhfgReyaMjzLe
xq9zH4Nia4lFHQZAVnfq9luJPY1yQ+CpN8B2eG+ATldOGSHxFlm5sydpNwze9/khc7jIGJ5JtiRc
fl77SOe6IwungC9UTn/9sQoxiZv7RJoPG5YDrJlz497mQVhhIzeqiZeJAH9RaZ/D900T9PT2oiJr
aazGUs7CflUy+0DMy8ePuSQMb1O2c4HUeo62j2YWyim1J741WbRaxHIhjWJcozujPrXOivaXEm19
6LPnDr2RqIV75UJxpiEItzer0b9uxRWnP/AYt+gQxrvl1pKjKKYveztp/wcLLDzup9IvmtA9PN5Y
qHkYpdWd7e7laUPQZFyza+I3j5MObnVxiPdKOgAXmr75SbxNs1zHVoNFFrCF4IYQ6vrcFIKeiGzT
7giiDHSip/Q52gZP6UKNCAj3cYnaoYdgi+Hgot/FB9yfJJb+cVfYbSEhq37g7oXVYA7mvbGtZrtw
Mx8AkHCw491fyskL0p9AAgz0ZCPjweiFn/y8P2CPan+wUim+ciXRTMbAY9ydAb2QWLv17PEhvJK4
gOyvN/04SthbDt+cK5YC2ydMRGiXhhBe0PAAF59pDf2XiHRyfcYzhu35/f7iBjJHZPMW+aVkMUUZ
hUJaEsOVWG4y4UYIPckdCDqsQmXNka2xPlqcJIabo08K3uE0bR9RFBkXS2n+QsCqeNn4mNyf+FRw
IV0o0kSktiDkjmY5i1guaMU3S2AMz2w0xlVu9R0Oeo4HZ2eZBXECsBLGwBpGwoE2xzamDiaC7lzU
3MiH18g+rvkZBqZdaVKeRG6j0iVy2NJk4Y7l2RrjyM5YUDEjaG4qFyWmBDAk0az2dF67rD9Omv+R
YQ3xQxgbSQLjzh+ctV3CRst37Ea1wd5kz2xOWLixM9sfrXTlOXAcStqNqL7w44CDPTi26hdPFpLU
BgiXyKPPKWq2yDAd5+9s/sEooSWGXuZwFso3kKrqnPKtEa7SRyCKlB+KrP+1oRo9rh8kB4LQoc0l
E0JMpNg7IyiCrcSJVaTGPNBdKiBhvc/d0dw/6f+qgASxmOk0YtUsWMIzWsY4kDNxjuB6b6MgF5Ft
W17u5QXqKoYe06jRF5V/eHZZw3uRd8WIaiotL3J1FWfliT8BitJwxZ5NmLHdMNqMEpy3Id9PMd/j
t/yVZcWsfad/iVNN3hBgEoXee3EKCe4x/ld/vckfZqdpOQK6ayhsXujE7CkrNfTaFNcADUlviY+2
/I4Km+G+HkEgBjmskOC5TRqUOTggcKWvfCjIQLJ9eUOjYGoPLVuHCt0ifMmVKEe8pMz1inWviauo
3zmJUf3EMuLYgeQVOzIxP0qObD0o6iLIkwLbKaSPntW1AGcvIf8pXSMY+IUk+vgq+AUvTtFM5yht
nROVgVKijZo77WvcWzxixd7GlL5iVlKm0Xb2q/qzcrKK7J3WuZDWOAU7RmcgkaO4Z8RwIIhd2IO+
EmCAsq7YuPtjnHQ2yj3nutfkrLEeqThflKspIjchAjgSv8ONTb2I/U6qzE22yzaUNzqZugSPZvDS
FJtxyVY5VcrBlm1E/UivL5P5eK78dFxRz3sQf1vnlm01QA/eQClrMOMn5gxfxBUl2IG6H/iRl29a
nGxE4YEjdg3vXTLpNBjOyVezsiPCPbocXNJ9iewAxqEfaTGUUbDDPl+OWh2Uw8HE5cACBtf6Wdqf
cvfU1vpvufxAIgpGQV7c5HrdwMdthiG1bC/YiGEzKqbp38Asw2xWggoYVHiM+dTh3Py27aU2RRIE
i7SITHg5rLVYLcoOEkc412mKco21hrkXOnfa6QQUnWIC9zrOXz0s7CsTRUxO9n0n/cE560LMlsXz
HaSVEIaRjdXHhcnv41xDCY8zp93+zeFnOX1FRB0ymhUlJEPVfMZ7NJClW+REQsrvpRpbgpaXMSpC
J6tuFEKEwYQ+VpItpHxYKFXojl3jiI5BRtiC53SKk49xRfupRu8bA4geiZxFu2YdVAfyYaHKlQTp
3dzOeAi8oHuoQcuQHDugFrOfPkXD0Ai+EM+GOioQCtlbOJzwPy1G2ff89s2tiG08loFvJus+K/cS
CmJ8sX/6LKu0UZa09LUPeKMR7TDohjSDFCcZc/6X1exOmaIBTuLBbR6wrzzXdTavyNVk3fWxvNKD
Vn73S7/RIdalrTDIqvb9v07XEvcnOKPqHHs9s+gPFsIwWwTk8Smvx1Txk4oXDQo/7iasM3M6x5q/
16GI/VufEo4Y2zPMgMYnBf39aSqaa3Ji2pFx2ER7vxSZRASqNBhYV/UNxLtwyTujDU/p2TRXGIwW
KaEuohXIK6BT1aaZaFM9NS23LLzOVGHB1z8QDyMDMQJgk4H3LoDxJInKn076KQPU6VilvPpciKuI
7dNkXEOUGVefobyRD2yXUNUkq7i43jI6ZTGcOFssy9ja8Z36clvB7evmTzs9ZVd9jy+NO6M1mK+5
7/ouoPShJ6YmSt33iwikXNJe0xX7hTQSy5WZ8EdGkQ9zSPyx0DFu/IcfCp+ijP5eppVOy3rsipHj
vg0mRwpAmw7Hrc9/rwZqRme5oFLzMYxEwWOChfid5YTPQdIyzPYH4kx8hlOlGrx+mo7vgCpfTldy
FG1CBCes6ifsG2FO0goEADTzrr07Az7hMp+yFZBZgedfiwpXznhKhIK06iT9RPKcPTN+X7fNqmMT
rHCu8+A31D4+9JRJZhO/S25LeAgKxeAGdV0OpuNlVz2PLjFOy/Aj7elGP9QuNXXVvZbEz0TszVin
3cVS3IJAELzW4/7u1/SiMQp6Y7n1bTzVWjl+US+g7w0CsTIU7itmiUQ997c/eWLclsefqeetkTsg
PQT4gnGLwb38yw2M2D75cP9jG32vPAQRDwlKLAVBdAufQCzGvfg1rnfGEcMO/MiiYTwZMUVj9Nn7
7QkM3/fN6y0AYnrSyhdMN2y6TVChE8z9+0ehCXUpxbb9Kcb1S0YIuAsEgyBZ6MmRcWMEUXdKQ2dk
IGApF+VORe7sTNvmGfdXjZojIDmxkgqahsxDs6ugmGamp7tWTS3cD5Ns8LQau2LZ9R8+dw5uH+5l
nGf58rLWyutJ3NHMs7s8n81IPHHPMqy/NKjFwWtDODyjrhtUDZp9jUvWHksTPHYRaiwYuiZwiQ7l
XKtG8qLPjtPMqfwcT1nYjyupH4VGOC13jiFBxkZ3f/6KLAzLX+2lxXPB2qePKABgx2eV9AA4Asy5
PFatDMeCgWZ/A0Sk7eyXA7jZ7ILeHU4i62Ii5bPVqatoPweW7ymRYIuq77cp1J7Zx1S/n1N6tZzh
p7DmuiyhpYW2p1DDVHw/HtVYQs+lquIlJzdV9tqTUJ2VybNa8vAwR5wxFvLtld87JvzkJzTYCkzF
26QOwfhWhLe0rB0KINKKWFw5ocwyA6H0Cs0uBtJGaGJD1FUMFMrVQGZtJvUfHqdGSfkwaxQISdFj
QGSEPIrrNM8Or+2K8wEZYgBJqKhBzqG7gmsf8HDL7L+eRBGWI5sek8C+dt9shmdMghnkn4xv77zx
QfppkYizHkXj+Sw7db5WAvRwDAYrQKQ/HFnEU9z01W57hPwX7OvuaT/GWaUuYftOx2oAbAOWOrhz
P5Not1izZ1eYErE8iSjmFWku34ZlYZMo2Cl7Q3JBvDmmr2QwxPjex385VROenczwM+y6S1fROCEE
1nxJcASE7huHgD05bC4gZG6i+gF45bC5pXx00WpgFeEXGq56fc2Sa1uRyb2o8HlOdbmdk2nayUyI
O6BCi2tmG8cepuKSkBW9jKfChq+D8bN1RAD1ysO8pMOClVvZcJs6Qyjz+uEoy++HXTGtoS1zq8JL
EtJTjDlpw0rpsfPYvJU8Omk194XNQ9WPHeWN9/YSK+fZ4oWeiZ540OBn1gxdk7XfzbYOW5BYJ5m2
cc7KXQqHq3NBicP3BhRJiu6t2Tx1W1vYNSM61d9MOYDzWZn8g5VPy/hbUWbCK9mnE2JFlZgxw1c5
v2iXnWvVIL/CPQxd8B0KnZ6MhJc9+KypQ62W1U0SXtcAbGaJW5S02P5babIhNADu9o1BElV53n9Z
yLUrCIO5rf5szhPWmqz8atiX47ZlRF/E/CCTVODuLdm32ZsMYjdkofhQ66xAVXtDv6sfZsDAqQZ+
oDmfQOht8xOGhsy8gunwIVBYtzbjf95YtrWeZ/9D3UG+jiN/wJmbtFfHIz2Pc8B74vMYjhj2EHoo
BklIB2N/wrDSfKfdQZfE+56WD/AY9tmK0UqRKgAoY9CCXBdKKnkaJyq/Rl/iaZNTHXQnVKk7MbGQ
0AfzOOu7nXvqbB5LdFXZYkcsXor1LhR+8LYte3IAkhoeB/wcdBjsXhld9OqOlqPdNjGJqo5sWWaW
BmpV37Id+xCwTokEKjq0uRjSwf57Wp1RoBM1jZnZPER1rcJldU690KZLA+eHv2VcJo/F5zRWR8sz
IhCM1qgfjBqEXxnEIKAAH5kqUHgD8CeIb2ypsYs6a4vPVFFkNeC4FWK2LhnN8tlRD4NyITToPn3Q
kKP2P7ulnkHcR17+EHGPSPTYIZ7y5mZw1Vy6TcPBmgAf19P9VtU9unVTzd0DfrKx1nPxlLcepMfh
yVxKE7P75Wz3xvyN2PR950LBFSpDfMjUDkXCMqj5DfekIOThzVSXkLrmRwZVZdyeVXqN60EVVNaE
S3HDBsuZs80XVEj3JobIVNWGboYbLZq2gZ8Ax7C6w1JIdaRl7aI/NOzvRarGC0xK5lwY0Y2SxOMK
/hWWLCJigh1MViTZQ9r5SYdlilisDfDOP83YduNiWU7YvLPXysA/vlyYR0jySgNLz0ZfFZALVm5V
NaCq8wO47om7aFfRhn2InltzLECSncD/yXqlHV8kBC/YVqbrr/+sxH8CLqVQX9dd4Jax3RK05VW7
LjgqmpF4MHamJVzyUPizh8yayOc/BlDNLfprhWgdRIVU00JYTI9LSMi6OeMPQLfS/WLklJ5i4EMf
92s5epRd1vI++Y1Mfw7gyIaZUaJPFMBJ5tKZ9XkBVehflK4Qt81zzLGzJz6yhrYr1d5/e01ZbaUf
J7ZowEKrz4mTAxSgl6PPQYkx950A3rsMMFYFlhWt989jY6N4FHg1usdCxxcwu/tKgF78ZEFHyXAs
u/vx99rbsfCwMrDK2Iiba8w/oqgz1GB4l4YvtN1KzRJQSkdRH36sfnKcWFGeotjRmnHSFaIlh/Mn
4c28Z4xEPM+rIsSvOWKp+blqOm1PLz4yT83xIcbE7SXYqEFEc5lvEDGjF3ClwluP1RJXMeQh0T+D
1AaUmUmqS2GqhU+ZbOqUjPtL99Zpx8B0U7RmLx4Cx/DqPMlzVCTIaGB67SbbddFV0feXhaSb/kPo
ujfVfw4xTnjzjxyRE32Pqx6JDfOtYUJy2WLMGew39TVAQHt1pw7FBLoOF/7rNHXLhMdyyXTQe7Nk
bLKQCuFP3/DAytrU9Xl7WW7PnJVg0JBb1V3PN5jQoHIxJVVMoruxucmYNl8mkmPRWicQNav6rvhH
6QMiyskQZbWIciOKqHH67P06GMQZXfZ6x+xsBaOdVeJ18+QocpYHQDGFwHc16GsoZ4mn02kIhJME
u1PCMSb8E1B2yQv3hZtTXzh9rNhfudAno6oFaDkXWBGNN/VI3HWY7eAP5JhvOR69aP7oswbv9Ysi
RQ2M503E/i5wJbF8/q/RjqeIwWsapoGOiUPD0Ko53khQF6tNjye2zAX2w7rgdDMAZ97BiRfxZmw/
0HLKmcgQ2pX/Vg42o/lE3Yak8BVYfQHgo+WRvU6ZJ0BNcu9M5jUmWGZlRwgbJYCDS9S5fTAC4Z2s
plFzfJF1sLI3B197TFuH/jYvpV3VhkSigtQO/R4XFvVx+IVA1CHO95dcnByr6RRIsBVWrVfRm9r7
9DI4WAs0qfVA/1Nnm+yladjUfFfUqg4cTqsPmBXoiw3q1/2VcxvY/z+u6mgbQZg5hV4lVBd1Tstr
NOL8NVmOK/KDy4DGLQp9hlmPD4P58Eey55vN1tOp/q2vxEj6IssR2v7aJyAK7pEtAKOx18oE5bYH
ZIeedaSBV8r1MaZq+LBe4i5iYGSG0EsFn0Wq1kDVxDKsUqGGX1FjZmeDeQ2oGdNFteF3u8McM8zP
TdhsJ2YolT8lFFVxw1eiUbMJxru4XX5LdxGcJfD9ZJaO7egQNOirxFQDVxjSSYavwKOv/wbthXnJ
sYgI3Z3wzHWGAnEZCEz2Drr9J3juj9xk6CcqnimMMokeZrJ0r8vS2BdhH5yB5nBOK2SU0lHB1cWY
hGkC6nFkeUosXbFTUF/THzzeDBrBsy3THebpNK4qnBP92nPzEd9069HIEDxCi49HQDwOyQaOhdlm
wsxVuT1hy+dVdhBc1thW92A/rftYbuzA49s770QFruhlVw6xCdQShFuvwN6v7WWdMj7Xxhg53Naz
YUOIGIeneIzVHI+7xXY8vWVbyN81qfSK8lYMtkonX+pzSKapPr9nNUnIOt7Gg7lYnCBAMSiFxbP8
+CphFsNzjJOuBXfCwJVg1iYwoMIuwluFEh6BZj0iBCx4p7Sadf4R7N8hky14Q5nf2IUzTtx1EoHx
x5hMyEGVFnpD169IFKVwg4wRUNXzKsLcEn4DUMSUtJ4Bs/YYN/KPpOu6QDOlMGtJM3cd3AFlvnfL
il3S9HFAl8HXuHHN8Z8UzSh+rXpzedTo/EqtwT/v86LW+KPHhfY/lvS03kpaPgOsefFCU71x7lXf
xji9jngOJDQc0ekxI1/L6DjSg4Sx3MCgD+BTRqkqLg1oX9zyGn6Y8V+t6iyY6MvVUTGHv9SkNmmc
EM+ehZIZZdg164H29Pg8tpIHn7PX4lSuQ/lt+Bo2xRPGCHzaU5FONhb2dk8aIpKdA90fxOyDg+yr
Lo+wU8vEivWs+ehhlpfskemuPJiBbQcE1H6tAIyqIIxiqs0XlR/bMxh/9Fs9ZersOmsP3cHzNS5V
ndA7K4iJ3iOct5UhUcCoR2UCGgxpZuCEpPJKlZggXktNmFZ3YbTKViErgtMc+rheLLExq0tX3Tsl
qsb8Vluisu3y2pSJlhdD3kgS8qi1heR7pqv4DUiakEP/BMTb+e5FURdukz7oTP/Y/5krVi9n1wSp
xlYJP7jX59RHhCJF37RDKHOmE/RsHfyvdwgQnq83pLA+WF0OVQFDkhlz5CVZf2E0Lx7Ervyk4frG
5KBuVX2zfODncQcK7ATHDDjsYI3HUd9ErpNwR2CeqUG0o/EHSta76bv7TCDWMapeUCrk+j8HKbGF
8p1/n0HdE2Cm0VlQJ447uIMGmJ4BgZL+k8b2yJYAuYsH53t30bWZjRnA+haxKu9f2bLEoCz1UNMS
or1hwdYxoZDRIhOwywzXCsnXVtlp8MCKAwmLOGamqnxI/H/TrAbY5QAJV0OiGKuG1ZR0et9ZS0A6
NTSz1eXrffSF0kf+eZnrMXZMv5aWeFgnUCthtftUkzwPyIugN69xWo2aT2wDFJRBWSmnQ4Ymq7ZB
WyOgtvYhtOUKLJPsoYwSpdiBQUY8/56dIrsMl+s2Z9/t50VDvrytn1ozxT15fHECdCFw2bnny8vG
jUQg76BWceY/1DBkBSMJL6Z2l0QPI9ph1AdP9gli8YJfhCmf/P3yRmns3tREmtn+iP5VygA7OWKd
Gc8GXiPCsXyXH9ctL4ofsV6uEZO3VFloRt2kcEEfGZtAsK+YYok4AClPjj0lrIsn2AwNGrLTzjMz
mE0afh6DjjeaVg2iFUxzdQtlF35sMjWTPXzl8PPLEI/uDx2bi3m1FdF98dgVJu8htY9m+dLX9xB4
Q6upuQg8xdKfpLOeSsnX6LeUcv3toByetmvihKY9jBGsHDTMS+RB+8B/v2HQCCU2dyNaJaeSQuvr
Ovvhht6EsMyBSL2z/0BCHITEhS4lkGsKCOww+sKOruPImoI2cYfzav9naiwwAVL7inXCyvnBkolM
q/ARqBCzULQ2OXZSFPtqZHCDrwwEcSBHS6/GzCp44Kjku/2H8L5R8WrWG8bfsS+iklJ4w8cUkg91
scU6E+BBgoFXE1Kz0EJRQfvJm1i7hfGPE2iUBUyz+ICQmvZ7o3UQNgKx4ktLJJ8LEQq+IFUjtnq3
Z6K6n826m1qdKrJf0pag+GAKB3xCPBtuLN1OGBkNYeGgmvqX7vtxpErkbIHgOi2NPTYnNUNojnvs
fyTmYeTiLjo0W950bffyL1Bas2YKpDBpp827owMHux05lJduUNOJoBrReN71oNqAED3b/ANleGkY
8BcWr42hMghQLh0LMngLW4qktWLT5tzAzKUK9yvEeeOtC6DtPjoak2JJN7yAgBPYg0GBxVmgY2Ni
OHljknxSukh13ISNdBSs+wkq6kVsgkJbOAZoHJig4HeVXOr1u+kJl7OcOZTa5s9jJEVUaZIXJqxg
HZPMV9kvob1YOheR/DF72Ne56NNy/W/HZLeh9sLQUcPW7XxFvN7wK0n5iWkmJYcq3FDeF1c8v1oT
n0s7BmxwpO0dzB2YK7hU/UwmiR+EXbJSblFyd6LfEboSUhXJoxfoHwTrp1aPzAhqIyksMoRCKGSj
gP4HIpAObB6U2f4yfvlLg9D7AB5jISHvLg3cVsHH2929ChEIXa0HLZYR50iYNzzB19QwVpjJ/URv
ldL7djGSfNrTNfe8qBXGqtq/YhTmOmXEyT1FT10GZIkgxQY5w/CIcHur5RWxtayDuMaXWWQ+/L8i
eIFl7zP5J1WBEWMqi+y/FskGRHlL/cPykwaT4CBpBJf4eoEQgYeMGOa+SoLSZRVK1nKRhlRBuUEh
QyBvVoc0dszniDvRflVU2Q1+N+nRoxDPvDCNoq0HklHqjL7W46M439qHzxLcWmbaXpTJb5Jam0e0
yzmCAU1aOLkC67DGMdeQAVvRGYr/SnGlJ9eHPl8MT4GGnGcNYsnhutRp0i5O+QpMVXBdOOibqXH2
Dj60MZiiAuUXgTF1okB/5TIh5A6aXxyqJgl8rp2RmRk6MYU3veSNJIq+PueBeCp8B9Wio7UZOIqZ
HMVp/0NHtX+JQEhbEndO3PR8ii2VHytugszEvRno55lujM86Bp/C0HwmP/pQsUvvH8PatQ2mo1DL
U0PnXAt5r450sRiKx2fBCt/kvNrLqLn0YX6WvvYJhpQtIn6Y00FNlcsqiDKXaX/rFFCHD/V35jHc
BnLwX7322P7Qj1jxiKe+W1Yc4zgbWEcUBSEYXjvUhXZ30x2Aiwn+H3nupCYb8V7vbRWezpgykZuu
fEbtuX9iuhBasCl8SwShco7i4pkXk/ikN+Tgf1cOf3CgtWGZMm59e1GIov61vDJrYRmBJHjP24FC
H4NDc824ObnO69nrbEi/mC7vYcuYpW+Ivr6Q3quCEwvJhmjpa0tbJd9Oa5fyOleKHOLWa84brA4G
Qg0i0XkS/v5n7Be42YsD+B47IboRxeT7DSDNMAOvvADMjUPbkIS2iWzcaoyUT3oOosJJ+DMI1zPK
ul8ez1w07JiDqylwFRGfYzxr78Fvcc+FTlegBLDdyoh6l+H5LwUJuz4tp2NY3Eq+tlJfKAuOqpq8
iXpZur1O2+mBK0JURdwGz1al5a6JbPMVTRE+FuVeOOFM873WFTIqrgvy1qcZiGSNhk1RMywfWQO/
+2Lwk0I8rUN7gP9Fo8sJqcad2A1HSTZu1v+bwn66QPgRa3MMY9zMO5ictK8BKPxLtDJuIHS5YF/T
YXYMstFIn7HsqD5X4la4atD10eBDO2BjwSZf6PtSRNMxqKDP/iRgTfi4N3Fw7NRdE171ko+rSyvP
ye5MAqp3zjdI8oth7/eKZVtkroNLxsLWRGB+AoBMx8FPjrPC0+zENoww1mHD5oG2BY/rybIXLPRc
B/WzMJZ4dLmLBt4Xwde9Fdy9ZDWBYs4+GfZYBykSTG6CDBFUEmXSnMdZPaIqc0iFTmy4BhS6oj8b
noZMJQB1BTe6gKIGpCDpwHJRbzN86mBIDgRPM8bXcGBVrnKbUXvHPLpqXjJtM9f6Xsx3JPqBdxp7
dx7nvINBtUEko2PTRiqM6sWEQ62YA7fa+cxCMeFYEAtqFpovV7/Yk9XD98r9nJviUQY7NtXGt1XS
JACF4Jhn4KEJws01CJ36SwoCxt7f0+3w2zFi7IiBFQ6KZsca7L+bGpnuGJ+klGqsRtSMoGjgkeRn
mq8DBuSmEroKW3OGBkJjEDxGQ2Mn1Zj2Pq34LKTi3+coDSiD0wODGgRUVROpAf67TQzaENU0GJgx
TANnVbHDZs3OMaDRtlnzm9+k/SeE7PMRAJM2XBW9KNN5yh6TYFEPoc15qUzLF8PEPDEoLouNHa05
rkpuu085GNih1yfcjekI0RxE5hBLgS3Ypunsm0d9eZUnOuHt87Ie1Aaqci95jrR68o/IN69j9NEC
SvYewJpt1g4o8JDA5NoIFHhU4giEdXYKVoYSgZtleE64abLad54hWItYAwXbtG0XQ2QMleyYcBEp
B1yPOSJKxjLjFDX9CVR5Fwli37y/OWgW0SqGoKDTUahmszrutoo/TJqLThlrkrAJv65XEsEmT4K1
lNNktTVmxgYUeqweyvYcko/cLFuNn6SQIxpmDj7sfTaWDqM0HIIw/IwJW2bsEq9jNzYIu1eMYLAz
1MH3hW5P+hznfworcwU7r0Az7fw+oIWwrk0xnGFijLYibBewuaF358gU0Uk40VQEB6nudgoi1dGO
N2cMMLZGDas3uZTt8Xk5qKH3+hg7EX77rCXL4dX5M8KRomoyX1igEQjrKQlOkbawC92nTrjb5wDi
6LXirT0rITm0BUcQsdlx6H00lp6MnYFcoVNTlg+GRJvE6dpDYFKZev+bo5SwD56J5gQAfEbnKEMC
phQuLfyOnbVCW8DCwo/pKvfphMd0lEe8o+97md4n6Rd14hsOvzldGrJZxBZvs+XnHxI2lKRdietB
DyzcvfRrHwKW3igEkXu7CysN3qMkiC513jk/JIsYPJegC806r/sKorhvx/B27DBxjy0b+8eMU9Z5
SD0qeWtx1+dZI+2PzMMahgYpRE3TmX1o1dfHZnv7TmAblzxXsnJ5LryzJYo8Sjf6WB9KcsBO4OXA
7BncIlyLfEw0B9HvYzCR2taDkK3h6D88HVPopHSmVbPIwDqQF4fbnaG6aH7VWCTCELiqyibwl03H
iGn+aPz7AGIM155OZ1aML3TD4jhyXY6l/V2qCPK3XZtIJaynuN1UDeUfUgGc/9+zPrWQg1yyU/W8
AmVb5JxU8z6tlD6jNn8zmEP3icigbg/5TpYv7wxIlHJRkz1AyHf94ABJaO1iogTQXe3Cc4mhvQNU
GIHE3exIKfSp9oiCY2mUTP4ZBZuW/+N5kaPqxYK6XcTKlmXGHCXV+yCi2X8qpwpJ6aCC0cwQRyqv
JVc2E+LaSan7TOSx0/Ethiv/H0D2kxvekds9bHG07bewLgbBcZoTrZouTi8Di98YIpgDbGepBXbP
U76I81bmhw9yw3MFXdZwkbGfD+jq2Txs5BCl4KBBEf+tvgDPcIJ+buPCz4GEStu9RTHZwNXRizJs
aSJ574q+UK7bHr1B8a3eHXvBhcWH4exdfBTJx55HZAbHE+qo3i63uIq8HSt1nnF6kV3wDehfL86i
Nm/i3Cz7n+p8Dd++Gw2YME/YX2zCuZygrjhov3mOK+5gExOhAx5j8imXhjtOXYLGDs1bktA+EIrc
YvTf58MMbC5jYuM20zes+g==
`protect end_protected
