`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ahrhEGUHHc+Fv+y8HP2i3fkx+FngEvN0bgNvZmnfQxIzEsAtHUZBLc1Td+0Ub2L4YMFezul5Mftc
00jj0oWM8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FS1H7vKU3gUQ4X76cmM+FLJ+EYreMRbqqYgm8Im9/YT48Jomn1zLPmS6aTBuIsXLNw7aJFuf/AHH
QPDXJkYJIKIYp4Acqr+mT1vn2eQ/+Ce/OAZDAZbVMIOSdQkeTXIrjWchoQV34jDNOU/xckatDTz5
RZ25vsVdAewWvs9lKdY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q6u20dAFfl2hVymFft+wzUJVneYgakGEIM9nM49sBxYE1bBf3FwnwacN3Vt70j9UJspgl+XKT5Dv
UFY76qu9M5M7KCsppHJMeiH2aMzfIDCmtbCPrd6krlxrGOuCxfAIdH1pft30WiA7940JMecizJ/W
HhaK+ozAsU13N+qjssN5m9pQHiaRKf7zd5RGSfGmI4E0I37wAiX7beUHQnEf2aestCzp6FvqfNQP
rNRaIjkRBXHnrvdXhc4QBpUGTWa5gRsMwVvhPS1LEScIEdgxgKNgKyIktkxi7+y4ScPdmpxoTbPt
WsDqQpduJquBDD4Xwm6KFhjVi3N8fPEe3TcEJw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HFzKvrFgBdSqhQmcvHkL3buLoxr2sQ8snAcWg17b0eSelgutgSYxrGDzNGGS7M5VVdMnaN1UYG9b
EDjYIf5rBKsHKf8rePYTQC7W5EH9f39VO7AwWmKqA0lWlyJZk73qClW/3lwfn8Dfc/Mi4NZ8baqP
qRohp7GXPJcKdHXku9g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FzWluHb7i7b4N1KjeJiFC8vRTJfOWkJDrORn68zM3oo59wb9R0kfGOELPIou+0ucpcLHFrH3SrIK
goE0BIEAgpR9kRXzKuXq+OITYR+NCJ7sxBe7jGNQnoWIlVbCaqyxBhCswa6PS4QnCAqm3zOFBnWZ
qeBR0pkWLoEIgbFxdWvnWfS2u49tu0GAmpTSkOj/VbFc8njdmWNekfA+dwJ7So9G64Hrtouvj3jO
cEDpufnIiLAMK+70OCIQiAikR2BcKXIC90KwK34D6UHJc3DgDBwvjlh+j4z0TNJnGzq3/twWeqE0
7V250DL8Kt9VFDXEeXrfzod263Nts5r9ajb/Vg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5728)
`protect data_block
MKRLFvyieNYCkUuHudo4Ejf8ZFXRA9a1QQmSiTIKeWlPCgqZOpnOVbWV1MtNI9cXwTAL7phPf59V
ZXqf9cM0Wd2ikCdU7HYC9iFL5vBLUO2Z54Cpj/qyMiBD1Nhwt6FMPLGXMjtQKSVuqIpuqRMLwpxE
mQXSjE3HwJSWFMSyH3MXs5LfHx+MhzGbeyVKEAUGZIp/bPQN633cVBEe3U+BGDFYbUnaZVM3LBk/
tTAv4YoEW5p9Hc/60cmT5GoH3EbmWH7Zb98DTjgWhSkistBJuQp8TdojNKqNV/aLBi19h027VEPs
tSsyoK5y778pCeAplPHvLjghNjRFWNR1s7Y6EuF0aFRPeRAVypBhu/3QVi4iM3Kzp5gGj0vgQU4s
CJQZTF9Hg02QQ/Dkv7nA1PkfHVs1DCNvGH1W6z4LmfUC8EA6jpntE2qbhk+vsNwz9+VRhNV35Uv8
sSYjyEuSmqwWBW3QAY32YSKRYlNWoYs3Bzzq8NQNtcAJqQLrbShpBKROyd52eqmz6k1PKZqYy1yK
zSMKPpvYOSRFfgYHzPBS1vWtQ3jCHPcVKKXHuyqGuxVklvb+pWRCyiNWRUAX/wS8wpaDdBiZFlKd
wBjGXJDMrr0fxku7T339Ow2befJlFY4wyT5ofBjDPsInYieTP04nz4nB67T7ayl4q0OtF3touu6/
YjkQBnvmJx/rB8qpRyy5z010fKN01Emi5TGSBR6ZmAqHikMCBrMqAhLqjbBznCPOQRXI+kFDcvkM
Pe1zERd4QhoVOFF40txe9mNelMxlPPBZEi2g1+dVbB9SzqWazktgtvYFIZyXMryci89fbo8omvze
dHMzVIuET1bysP62bYT3LQmGInq1SZxHYbIHVWPtmwCUfSGmuPt9jB2h7PrasoMVyXXeDAqneJKU
9IYobeTLZRQjYbVp/PCeu6Uwa5v8t2gMV1NaQcO734UZ4jU2psRU3nX5O37zTfy9JNCOEhRl8ejW
oC6E68fsKm+4K5I+CAkdY99Db+SbJ2RsOSYl3QTziIwcjszMe2WIiLkS64NfnvWb0eV7+RvXaPZr
HGqjHwt4iGKc6trBhg4JwYCH4LxmfMKQi70q4iWtff4odxhKvTdrEe+t5pl1ufAypwQEUZM/F1cQ
J3U4xVAfiuNiGgax0Wa5KLVLu0zJ5apDYl7zqVrfp7U7aFLNsNzwaKUKX/DMZN/Lf7n1w004nnD+
CyhcMe4HwOxjCPM8y6KOARHw6vEK5E5PUV1DtHrQaSbpvro6cMvSVuUGpbKQXeWrrtQrPj7pw2AH
JsJFYVext3Q/GmyB7f/XrW8tT30yUtDzqcMZZZLs2Gjam4Q18jR8Xnrhe5rYYakZqOjSW/Pru4ol
0sWh0yynabqdF6pIwj1VuGtFZ6gO1R43Bdz4WM1ZDDkBBj3X970r9R8kvusRNPn7qm7Pr9om+Wz0
upOlxoj4wYlhd8safQer8//vCjJWy2R3x8OfJ582bMjQhIv6xOSvYTgPC8qafXvm1ntIj2H5eKXm
dd+sReENT9uAZ/G7xEmdLjrXCnehpGvsv+LkdR7mBulCWDycNSTvnMD8JxsTe0WJNjoUxGN5TCfh
ulXwgq2wMCm1bfzaO6ZZbo+7tf0f0kSKHshxE9Wp88SgX1iRvIrlIJdUaTGG4h4TFZG7zxBRE7ss
zfk9OjuAPGZ+c1PcsHGJNtL+qvvyGLLHzSytPzOgVZtzVtTD6eJL/PrqdJ7J8ThiBvb6B/3YInz3
esu9LLSjWUwCc0LtATGOxoNC7JC/MZo7kQF/F43oztd2QyzqvHFaU4jsLLcHZ5n6HjoZA+SY8nPj
e7W+SdBn3FXfFl/334ONYRXCPB5lciN7iiwwCFbGKENK1TBzA390dvjFsmyGlvKIlj2q1UBU6yZa
KPSRQYjDsjA04uuhAx9s4+Dcnkx9vbz3n21VKg0SggahpLZaRZ6558AML/f8e9g2Opm3yNIh0TSU
+Pn8RR01GSi0XtdA/oPewAfPW7yH9+AnRuGylUQB48SYzdcuAD2epslK/aRl5dRfmM2EwnF6EwmB
9xYzadoIuyhYJYulyzzYntx9H7zR0XpHF/G7OlWR4K1ApGwLSgKTNpTiVJFyKclsJe1co154puzk
/xxY4SJ85fcjrBrKG2SvH/74H6VoVU8S/ZjqJ2ly/ieZlVHNQS0yTge7onskn+wwSOKpvVQTS9u/
gi2ckx2WcVbVkgaQ6qUccdwzPLFsyRGcSPVyuKPtC7PzEsBS5ZD/ubLihb9UGsDaZwBd34b4Jh0Y
zrpTAwqldc/xhCkv4inEp4s5m7Iq/btJ5aC1r9BalOZRFAyjHa5VCcx271pdteXZp++es58XLijq
29Vy3jtGYk4Q0OfleKUBmzqlctJvuElGJ3hx76v0/kTKPGcEfzFeOESvcE58SbnavHmQZ315pHqP
mUwkXflMvVkyYl7unlUfPVuQEV/e81YJXYGc82AMX9mOh3yXE6fcaUC6VzK+S/M761nJP1GwFVw8
J6fL9s10HuzdUJjYs2pOPKT5hFUY4wygYAk6Zd10Do+xZ8BkjHmhdy/UcUYE++FhpmJfydPkeYLE
Sgov+IfmRxRbHACy4qrizLTblPMxm9me501r3E2VamPQ9hcBPILIprM4ZmBdH8N4UfDLhl6jwvTh
Dvb0ytd5Qfh6BebbR+XHdyahbhAZ+a3R94fnFWVG6rOiktdUXctR+qyOjJFXTpSTx0TxFt7RBlEB
McE1LbZ6dYsl8v7xMEr8brGLzHEvDIJO1DRyPr6UMQVHqYAF4pnxGcyERvK4zpdKBUEk+4ERT/8y
h8/MLhNwJNHKhkC78xH5J0XDV9JtnfhcmS3mfDQtZaPEuTciAGqOYIclqhLrj2wMTbcA7qeLNnH5
LG/udbS5dcBXX9N08P23R2Z6x47ipgbXiXS0iSIo2BmSM9Jp9L8IEX5xwQ5LMOQCtF/wXJGFmaUg
f6TQ+/iKCkwr7+leg13a///DdmuEE4QwzgsxWsuk3hFBTwtR48qpuZBmNEov3seGDguQyzv4d1VO
bE2Be56qe3PyO6UMrD1SA4zWgzOsEfeMMlWRU9cZ4hHlwURNjLyFFAIx0pd0orVLres929v+R1I3
UHueVQVpw1MRakRQ5QmQ2fgoS5GdOuxhOXiReeTJ02i/xU5QsOe5AP5kDaRyjAmsojkwpF+Rtv1n
ZmaGvgZwrnL1cPxXpyV8gutDg6WHJMzQeIxV0zNHPteGgAbFkSaPmmtvS83l7V37HD7fHlioRJO2
9kITQui4nRkPIolQnRq/PCvRmUTAuy+Zv67b2eHV2ye4stIm/iw1hL7P3/0WAX6Kx0hdZBsnzSEk
bYt5lVMGkS7WjiiliKX+CnrtNLLazcUgjl7QZWgrt0gmlYHLiYdUfW+ADtE8u6ztBheQUSr9ziK0
eV4RYAnOoRLN/T+LvgCbIAreSvBU4G4hYWJT5D2GmSEQfwSCoPiRUtRlI1hq4twoSujTAbY8+NW5
3lCdWGKi2cOBU1/lfUBaubHjwLWdp9syUnjv87GPqBZIYAmRAyXm2+Zs3U5iTrjDa3jGov3o95Cp
dXZT7xpzNtl6pt1oNgeXiZN4eiJfThzL6q4m6tF69nJbgggBOBXkFcybS7aHLeQ7d5kEjQDDOitk
6668QFJ/FoiDFqBptX6cVNrI/FrfHloMYYlsQ2BsZsYnLwyUwKy1+w1+pw1HzQRQO2khgV6/KeU2
MreRjJ2LvUXTg3mGQSTIcg3+P8aFS+jcYEy3ior41zHOKBguI8NDmXXTRVx6h5j42R9OWXLZjOaX
/MR2WhonfZT3VvdlXitApq02FDADmQryLA6HtkodCJaGzN4IR/wSwr05ndga7M6++EKd3l6CgUh9
ep8V/dw0qFDhjQ0GWAI03svnM9CCgLNfQhPlIpZDWHtJIQ+WUXc1bQ32EFoKtoUuPxk3sr4nDY2x
dX7WtTCiVqrMvkc6ZtLii9CitODpmHzIj1IgsBe9/1uxH2vqJ9i4FDUJv+k287u90MlJMFpnPtCF
1ZTIpAkerkMafQr3NJ8s5H1oVbqK/HUfiBBAbg7p+CR2FZbl4YfqATtvrErfPY3z0VnyMmNRyGP3
Kh4Ev6OYXvo/O0kY+advs0atDrnYj2K9zrEBsshZhws1Fa6EeHkQJs2JstVnvECEKdwVTz/LnWO9
Dqrl6bz5R+e89GADGu1xd4FLzVPiUfm77djmi+OlLALDe82B/UidaD5YFw6kqccVqUT3OfdLmrMq
mwbqTALoqqyuwX42L7vn6+ldzVqAYubqJjiu13baN8LDWp8PTr84WlJCKZCTnGHznYeHut+iDSt0
HeflZHaxBXPiLkjOJ7xOFAKaCYKT2gpUCLQv7Gp12OgTY4SWwt+xjFll9W8eeNdICvzk/N1xUW5q
xJBqJn+Mzi9nlSrs7Alee4EoNWZJmL31Wj4/aTnUVOENF867nwZENCM7/i7tKAoCOfbEhOjBdYuu
Y9HMh0M8sL6I3tW3hUlgy8UqDPbEN37IozJIOJZrUVWEMgAnTAuh09DVEtGu7w3I4jvKM5XD6NCh
nI28x5uBJ2qYrdiNIXYHoEWBn1MrzuGpnbneVN58TNu9Xn1t71GAwW2T6+ayU26xolufXzcww7Fs
djLbTne08GYiU9yj67H3h7FCm0WDzqn+nheyp10dyswVf93dEeXW2kEeYbEy5CSN2VPBZQmEW7gF
JJOf7eiX7qZoK4uVVgFTrZKTwLImKiNvM45KIn7u43yOd/EY02FSLUa02GQz2SQaQUzTxXMylqez
wuiM82xIuOySi/RcEP9mrOs4QBzmG4uWuI0PoFa5lEAhVcLFfNuEsm/EOqpdlOP4RzVG7ITGMoxJ
0Z848D67BEfDrju5IFZ8tNwWFak2Hc34+uulEiDZkyOvta48jgw02InSPevTKvrIPJePkNwuoC1O
PqVNhiilrDcRBVnIhwsySuuB341sdnQluQ2XqihytPMTk/nFUNUypiKtwuQkhPbzPwEyRep0AZfx
ndvvtdGFZkM1l23SeK34dYaKIy8RFKtUViq5HjdBCiMLVMH1bbgyfn0QxjIpKJSO2OAS+K2uRI9I
fphrJdDo/gZ97/sbK1tHPDu9xDgxULNoflAxApxFWtK8kSG2dQkMrHmsqgIVus82JgCuPtc3hYpw
pyBPP9V6K/rW0MC+VvVoHu3O1MPrgGyVi2P/dPDscEH7zyBfBkfNMGnoIiq5vDHPY5YKu74W4Btl
T/JNy/lAWYE1mRkL3v3+Avyb8apLsvqZx69GlbFexs16U8Om09SZoQKG2OauO8wZiNz++QSnEZKm
CrEvOf86J+/eyMPCmTN6zkX1FPjG7YbYbV0aqyIA+N4LlMdS9YyvsQNIAcntZeiacQ/VoZR0/e2z
CWeV7mno3fLNFugybGdSLQ/+Ra4mK/0/Rb3iKflDLgjNBf3X76uaLNlLFW2JJuMQ5tIWhXEkpxSr
M3kx8ooQ56/f7YO5WbOmBvNgxKHXrcU2h3tIU2ba3W0Wt3TBqEATPF6PjCh0q39/6Ay2QspPSUoI
N4rCPkYdZmPxEu/gkGgFe4AXRzt/sLJIp8kzj0+IAyTRygCfgX6M+fQSrB5bvQuAuOsDd8h8cl34
bH+Cagzm/+hblMwc3PAnTuvGZIIZRDPot++pNp86uvsFNEDowRQ9SPMuFKPODx2GP1QhVKtbjk2K
c9zsg/6dOx92G8PCjG5We0QLdqhidckTqrd1LsdooufjNpEePRSxe0NluiMULItolWE420uwyFP8
0HLYb+Ly4nQImnlRx3OPS5PnOnMzjvgJN710nGa9vxObH52lWvwb71ZVB1hvspZcPtYplH1D+DtU
COcjnlGojL6D9xkUkoAhA55Fetn8Yxrd1kPt3DU0XE/6tYCLAxEdvsz7VyWfSd+/jqq0kqOe1SAv
0eLxEDvDGYdqt9q4+leijfA9g+5anbsmRt+tSAwO6u8lxGgv4K6qq/E22AgQawtY7q1IjRGkxfYc
uux+wWZ/uWoixTG2tqDzKbQ/pz29/ylgXjJbjBvhMbI5ao5Qt3pyncRmr++tkSn3uB3GS4Z0eFKc
AXsv3lTjI2LVwkbBdLBThu5h/04UfWhX+IiOncXviVKqn71uld3JTXH6gOKGIe2KGuMx+7eiflUo
fDE5OVaq/t2gRyKyo2fDXg4zN2hhtRoKeOFypcAvC+BS8brGPuveUfYnRenU9B60JHnlHin7saJT
ZF3+RUNQH4qeNuKgF7TGarHgUbaojwcDO0SgmijfzfnXMWCgnMtmhrF0xGFWv2deZyCRVH/reGMg
wBpMPTY3K98hqcS+bp/ijyQjddb44TfGLJ2rd2a5MT3EKmAiuLPl2iIez3chr/+ji3Cj2cgcr7Hs
vk8zYoGGzs3JJSiv+q+1yEJf7EPXWIIXS9Zh3C/Vaq+AfQGMqG0cYRHShkcBEACH/XHWreUCKPsq
0SplabHHdTQ6eTDtyG3kE4A/wgW1bBZ6Hk6e3KsFAWPFZeu1jXo98rrTtA+MK52z+gNhMVHEwpdN
/iW+HiBzcaqtlFKsFQA2mf8i5W8r453pLmwIVo+8LdwXNmqwK8nOFRHSKczK6/WOE+Fuv+M7Op9i
c4JAJVdlFM/Rcba81MdaOzGvTmQBMWYXgHp4IIsOLZIlZNiCDDMXDnGeJqkJUdgHjI2myclKRAXh
PaNRr6FFzJjGT/HXKpj4qZ5pOP8EqzPj0BAvgEpgqcsPMFE3kpoZexyI2NUIJxq8EvdJce49P4Vz
2SnqcDkildOGy5wRUoJJweNDmiOraengnN6OQqQh8CSpQY5dxjgD5UMhx4kQIuvfpvEy5afSB0P5
kbQ84pOACVgFancsVSoietLC9rtPbFkB6rd4YJOknD97YZaPf1WDcg+wBjxLoOnl5584G/yqTQVv
HlgkCR2ppgyY5zVCdVO9fjdgA+Mrf/cCyDVuSGC9/LbNbDs/sg1Nas6d07wwNqgFpa3me8+QhTxG
Re67OEyQiyiCq01UEJIaI2bmmpTVkp8C+HefYuuph1o04BKeUuV+Zkx0Rq9O+c1JJhDhhYU9+sUF
+iRCQo/f15ZU14/IiaxWN1sJkvNN+NxT5sOM62aDksfmCLc82drCZkr/INcp15zLN3nRnxnDdGmA
n7jWpeAvl7btCogHqrVHupBwbpG2LuvMwwxVXMjDRyRo1lz+a5gAFPcNT/xesCzVnL5POB0NU312
fzHiDsH7qmup74Pzo5hx+Zbx1F7sYjHJNbYDPKzjgBrMH75WA7hNUl5iZNdZDAmb9QDxtXuU/F23
ZdJAkWPbLFdff9UrWXFRo2YkcbNmMV6vknMy5l72GFJ63Mm9PREZebzQUl2lsF34vkOYTqnkkeD2
5Xt1fUIjKLdWlHwsT+Mj8B/qYo4WrxiF66820uFQleqDcpDsxaeBKzETCpGIo0x+zEnGSczSdyLb
hPiZ0SOoqLEuhAZ14jnBBf8r/BANDU3XoURfwTtvIXWg8/l+QxPL+LFnCh/qpafg4znWNYdVbjU+
tOtzoa6su4j0vWE1gyLxLfUgfrT8qhmPN0IyCXqUmYFg2eFxts63zIHsLGZWhgzV316BYQ3SpgeJ
yrRmb4dGKas0EzhsbdWcYazkVcQmrcL3o2B98g==
`protect end_protected
