`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UqQ92sq8O2PLALfIchCzTd6pHPDxVs7seWV6ITsyVFBQkI6zQzhhuRIlQSC4EHKO3hrtX4/o7tcs
8DDz+334Ag==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RoH55dYloOZl6VE3Y2nDIHNy4u5JHTyiYK70GCJNZstc+DC9a8BEmzpBUoB5+tTyr/05laUf89mE
nE4lRyeQcZ5EhNrwrXwJTsIRGNJz7vEACNqSS7avZ0QecPLBvJCIkz57aArIA9KcmaFZXJfR7vis
CWVWJM6VVnDt1OHXCkM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
piEMpctTyEx02UiAycYfJGhYavnnsd4pZ3ocHKiZcuUhRc4LHifDtzUXassxXTpApuE0ZGfEGdY7
QSYgGCMeqge7b4ox2pjeYLcwRElo7qo6VldegQ41b6VnKDRry0HvBp7wCwmrRtkNUdBwlG9o7z2I
N5YreBs98H/45gGlYk6tHdxezA/BjvxLuXqNF5R1WY84GlX/qU6PIg2KYwNWbTeGmMIg/tZOK/QM
AUmO/xECw7LlIvNT3v3h9MYxFFcdJPsGO2Wq0/FuvfisPSHCCQnj+gL3dq36UTFXt2YoShhou13M
RLM0MCd7ND65ZXTNBc3mkDW1+meuy9pMG9aa7Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aSlX2m6QyIrEOjvZWkr6dta4tIZxWbcqaeLQLv7goHlC9LPk4Wxc2zvmCBJszk8nhmoTaVCC0/B0
UEEcGAZ+gVOlseZG+QHhypFSEs/0zIuY4Aw2mhpT5eGI3bbiVeiFNaGgNk7PSkDoS46B2irLCbU7
QCTDpq0mnfWihVTfnM8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iuO9eQSHI8OkvExftT6Tj9X+QURRea7ZPQpfNhgQ6myjm8HE2RSdLbcjiVfeSEcK+nAne1OHs59h
tT1ycWmryfQDTS6TNJNK4axCqHfPFZ6ZPgGeFA46QjQ2P3GkGPQQJEUqybAD5hW+vTACr3kIqop1
gtkBXtDqnqv2esU9CVq64jJplO5TMBMWlUv/HskBH5CRPlr0iNXue2y5iqTY0LWexi3o0kvdTMs3
W4V2f+TZc5qz89AqskRUbfSgq2HAucVLtYLe7ak0fuMG3pn+e7hx6pqCVsaw3ovu7tFgzo73rKii
rXgA8qNfVgyiZ2g1mK4/SSRSRqQqyTxBJ6ToKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 176256)
`protect data_block
Tw/88eOt6LT32UiCSD1BQxxhKDonQ1JF9NXP7Z/qrfuEDqmIms5dEj5ccAoii5oXUbXgKAb7BbT3
oPh5s8K/x/Rp3tiNWu2lqvPYZGapfgcN68dkZinn6vfyu8jQ/jZ2xBwMczztESxzfnIv7dWhjkvo
TzO39FyahlXX6IeVq6nRCrO2zhQZ/nPfPmhFZdNsWYtZft4C331BEGD3P01QstoM2eWJA5vE+to+
Oj/2CB0u0zV/pE3QgRFAXgZEKDPMiOmD7cxCqXv8Qb9fr4oWDjOQ5doTgKmBQk1D7vnAuHFU6Slz
glta3adABxu/1MkzgkbbHKZMzx4PsFO+kiJR1878/wk/FKym6kMKez/C7/c+YT7x2o91mi8qQqrc
0Acf7JD7pcuU3HZf+U6ECXf3+gH5ZAThNkws5jdHYk0/nN1W2xk8PuQX51Y6//teJoC+uD4nK67s
YBwwJ9KSCc+EoSwCk3v9CaBR4zBwJvbLYUsczWGW2yCwPK3Pu1VXXcrpdY14C3JX8Y0VqGXtGwzJ
SmhjDX/bmgD5lyRoClHKpmrGFTCKXh3Ed2O6Ju7yHHZ+bpqiaySzBN3ywz8XVcBVr4k0DW4xA/6N
a4cXMvffsMMyN1cUHuhrDntXU1yjK50G9VGP8cSZ/+QYVbNLe1m6HbU5TORPFzpXSyjguC9HG3ND
J/+/17TQIU1VEgDGpweRAnWb7bzg1X87caeaRo+5Wqw/YOLuvwXwxmnZSK8MxIsG1hqgQQJAviSY
Vg/2g/OyiPcx2i7L52OJzh3dv8NmmTlid2nU2r/k1irIDE0Yx3EgPRMr/bjCbcRpSUYQYDOebXeH
5Vk+dWvKdVbSPxTYOpM1b/1N8aaLYnijEfVINWopOkLFajJcvg6hwLHxJNToVNGFltOYpAytu1pa
Cu+IbLIzHuSXcz0jju+u94N5Ex2jl6X4a/69os7OWtzbTE6tSXggWBTENAGD56Mq4ZePXAkxwv/J
wVb+NcRFJc9nDBt51FfLEEeZDX0YVHqeew6Zak7hg6Jk+5gGTh9TbGZkOrYbqH1pdWtXIs1yDbsW
ZhyQ+iXcWct52BkA6FVxhTcbSfjrBtOZPXVM6FWqV2Xy4GjKy/bTCa7x7HIB9q2eu1oyfFe9g1n2
zZH+8/r+5lwuhYQ3qzStkhy+iakGvO7OUlyfLb+Kl6wd0xd5eCU9Bx6jLzntA5j0pyZNnpefHXrN
nUAzN8U6ifdzmbiqbAXMGmSn3f/zKwHP4WqAAMDHAj/sugzGXHOFXrvHmwt2v+yPAWp9mPAUETCT
kUxKvIrv3MJ9XYxxHUtS2ZBqtNiJtOuJgkDxKVsYXuoL/qWNOCX75c6ghzUqoFJM/FhyjS22jB1N
2cj+ZOFXall04tFX8Tja5VTzAhANV8IoXjdA8vLuTWospvYe6VYOM4qhPecBulWa9SHt3Msklwjv
CPv8HtTkPWF1huchXW/ODVlkIYTkXSZfgSrnSi0IsfIn9OmDteCBSPZ8e5rC9JQbjJLNUIwOB702
pHI+3Oj2K+PIU3Mb2d5lg0/dvWa2929GEz9hvzBCroMDe5EibIunVsJ/FeUQ4yDkZuFWEQrUCZ9X
miKbH4W37CmnnZq77pCcknmQ2dYODLgCnt/jJZlOfrvM6imJmoGvG+cmMGS5HibuTEB2uwNmXWoy
i4FYbmZzkEFwc4nW/Ua4R0JiPsndUHI8TL6FxgK4BFrV2AoQxJ10CXSlzmhnTLrqXteYelPZLrQo
wzqD4Ez+2PRozaG291/HNT/fkE0WKswMkO00S5Ty9Cj0UUpkPRtcDFAvk3aZvOfLLXO/s2yoycRT
oABU0UYjPJpzlfTtw1ruDCNjR6s31dUEalrEoO/1suN1/JL6sHgFF2TV6301qmlfzx46/d7vVtcK
Ru9iDpnpnfgRyMuAADa8cpGxP5yqIuCefbYVIN0kK2/Zr4GqyLOUUKFNY0Rkn9ZHIOwnCXsV20js
jbdGyYKm81E+Sx6i1L3rJSfLJzoJO0YyciLPtsTZLt2KSa/TbDSGboYdKiwg33D7wN7QAEBKWgZa
zoh0MCuPqA9m/fZbjWx7tvCxI1DwvX1gfoTMAB6QQrWGoWjcBpscDcXqYqT76HmKQIzKle8OLJLy
aYED2pLuNY1NGK4K4NP6XrwiN8HuRZ0h0bubAIih60Rd0XBSWdi67v1gFo8DSS+J/b/LOjzPg+KH
RA3M9YC7B4GAgKu8tjZQn94zyR34sESDzKrnAP/i6qigFlm313KcfjZWj+ULbQL+eI4+TznFfb8f
I2SaQFwtTkjBkUjWMJlCrr5qhhxz0BSYP+B9CFUeU9iyq06UprxRS5CKPo0srWIzdo4oPF1wDvmO
5CuiyhbLrZZPtnuGTtEAHtEp9pNU6dFSYht7IFXdEeznUZmoS3s0OEHuXBYRQnioMKPpIggizs+m
tPqM3koqnBqtPe0ApN6kMs56Qw+5IGL20V/vv5BgwNR/c3Lnr1Kb4Ct65XAhzhVN25j4S/2MVcI7
fXJTzg1UR8mfW8p5Tj+Q1mZnsh5E6O8ZX3lTbjp+vGjc0O/vaYbUYtnk3g7AggPamIEQXKxhyu0I
tHHwS3VAh9kty87hK+qZMCzlBZ4t7N1Iyd/+0G8zimZrr0XEUXRj3SwqZYnx6mEySd6plzO9t/n4
MwNvES6R55GAy8KjjjzT2j55DokDmve05vNyyJ8KQaHeIaZ2XgyXzU6nyl2/o3BQwvO7PonbkTK2
HKq9j6Tv4AAFbu0PCRaqExnm2ofuMnHDsS2tfWAN5aitBupS/NsRScPQ+cHfKyNRCv//3hBBDrJJ
OzsCc+Kx4uvqbfM7f6LCMAsAjsBcTfjur5dp6jLFsYwbivZI9NUw+QTzhlA6kjMaOpH+Gij/Hnuz
SFDiwXK/yL1XOpgeMoAZJIYe7ycCSrhHByBotWHZP/ldwKQ5yhFKrhqTnMc8Ca2KKjUNaBFJepVQ
b2d7FexC4SKIppt86Hl177O6I6JEXJ5qi6m+iYdEQe62nmqVKYoe4NJHS7aSCHbxi5GEravOrm9q
D1sZOvEmq/ByPizKiUEx8Cyk4BXmPHPsfSQfCPcGCNb5Dh4tnpsuo+B0QthMVfZACKki+RMeaPOc
CCKmL7sMGB4NB22WgY2eX3uIpw0JOrRW0WmYZjhVfs1CSzy1m/bhGSRn/qlyxTGN5Dl8PZwoNkrn
U7Bk3Mg5/69l8yM5O64Jj1TiLhA6Rgbe5asSAmnvOP/IiLW11GCD3np46qDMJDhYNFB7sQ8BrmFZ
g/g52sFjjFou9hYqQe+tQMK/vzej7azUnafLEPGgZx3cig5KkSYrHhy12IKx6lgM622x90yhnhwu
p50jU9a0CncP9uXMB8ZjZky6R51mPUqTYsROwKVrR6H+YhkQstZUJB9FguOtMb+fFZpA0FNeBGJz
wX9+++jixwig92F9AW6c25XugNSVk2ajq03cx86UGyokJNEo9DbQ8CESMiruPC3xc3RzgPkJLIEN
Kw9Dwkhave3mJl18J5lkHaiGlYj/F8HC1dJJ+TJLjXOemBlDc50Pu3L7kgarebPpYG56meoe12MC
7XdsrbMEbLudZdnEmGaAaPlCdKPNwSN10rEPAPwMYCvusNHqNqMIPEIqowEuM4NjLzXJUzE/uZ4g
utn73cLAWvzIUFYFWJubnWrqH1pgpM1oVCr0Rhio8H5uJ00wYKHDK56BVHRkdsvpv1P1QHHCUm2j
w/h6t5L5l+zBn/i0rMI1WPEjUu9rtyBjDUsoW/d14gHQressw4sGi4G2SYKy1u/X88WAx8lfAU5Z
X2aHNMvrc/G513eq45Pqaeu4Afvm8lqZ+KqQAbf04G9SAHYI9KFhgkgrGCn4PGYqqNClTf2XckBT
gnnauXRdbFGmqUOhxnTQC+vGr1b7UIvv3eocxR4Kz9C+8YZ2EcEHfkVBUnIat7O6FsOc//BG+SBT
tanZOZRh3WZb8vB5L/H40xnyGxD8D8L2RKIpL4i9Xrm/h0T+aTXC8oAom/W+Sjq7SY9PcLZ5h4KT
uv2TlRrmOQU9XBCUlMFHlnTQNMQCguLt5k5x21piEwkcN/GfnxttHJ6V+QF4Bj0yOo24FBzFSn09
HehDNlif8mldYwLEUhNqJe1nZkR8Bdz7cFSBdlZhqNxiPC7FzcaYsDBkGK4iNXlp48M1H7qlwlTy
MBk+/AfxSStrtBMSoBHWVcc4hzkosiqhFFQbw+TinokY/KnUYRRBzsZp/zxc2ag/nCTRgGXy89yM
H6Z0Ly+Tku60G2eb9w6iXgXaQwdJHuQ0iZ+h2cwR6h5MKqzaauxv4pFWypJChQmrO7Y52lLWttVz
ZXTLLJVSKZ7vZKTF9ZeA0mmzwtZ+S6g8xInXEfdYLLE8TDHaj2EAXIbKjDtcYYcgbmbhAOyl00sw
ZTMavEA+Ij4AKrAc0jtvjuy2zN+2uEyBrFS+Fvx7iTQNF1wIpnwUdMRGrJZFpm2uKUzS26Ti6mnH
OkM8fapNqktTZfpZCLM6TNfjyo3po+RdbrFTSf7tfpTPacaabvIDIM6sBm+tFroFJ9BznjNxLt6c
LGpuOAtik6OAH1jWwSOzBVCinocKdVQ2Z+RKnwmBJD2MIXwUfVNVkgVrwqWC7oOJHzesvpeQeZ01
kgkrOW5081hHntAW1HYK62mSMvDpwAAu/VYAabFyBDo85wCwVXnBqLYNni1fGfc3Ij+nDOHbcq0r
DJFFw2r0WWYIg4MQwmSVN1ealWrfetRxX4TtOA2jauk+uaoJYP8kxl5Py2f82Sc0khvEHnbxPfK5
hS6H3ULNoEds/r9vt9XMdQ/18wK3l1bxWtOMFyzoVegZ3HSxMW/sWUX01O0U5AJLV4IxQSUiPY+J
tPRLaG2PTaazQSm6iU5O+D0GvxrgBMW+CuxcaExWdV55PBtPKP3t/Iv3yzbqegENoahxhHVA/YVr
SKWeRBvuGhE4aH4h77zXUmvN/bDT8nH/c49STdGcQPbjBgLW5mPNkqSvHQTO75oWs/Ed2vjpZvbx
HKDSW8tUVvJEz79EeTB1sw2k+KJJKz/+P41hOfnuQcwvfgyQ1zC55eAWSEpmldKDERucIpJhmj4D
uFHWTL6ES/Ib6+JDCLcUeaPH0etmKJ9jV65OKqPraNuSZLX52v8sYSQ1LOHgb7hgCjf8OdAbQq9B
n5Z/3xHhFNNUrwq7qq3ORDFEBdA8Qk1Iex5w8TTSRdZR+yCmp4366IMH/VJ985+LK+dS9qXN7BR/
1oBePe3E0qWG2FKUiMzb9PWerThS67EfXvu0fd9eqY+WWWEZxrHZ0ZXrCoqxINEHeHLwf5fF2jnR
YmZjON5hexqPwkz0ROvSBTrQUL3l/KTuEeDKLzb1Xg98s8jMv13cF6vtEkpizGdJWCd1tZ8EHJ05
3g/rtipUIEeXMJo52T9yADOEm3R6sHgoyzEL9GZiH54zO4wQ9ay1ehfDjP+mxrakP8KW24ecrhXi
itNXjXyN//697DDqkzU+QMcZQ6L/GFyO/pEBnzITZb36WMznZmdzLPd6HoMuXy3npoSiWteNmsn9
8BM7BjYOetsEhqJeh/y8NpMTn63GPjRX639SHQB1uTyBgzQ0DWITaAKhbhY7RjixmPy3+qAmEkVb
vq6nUNCp+MjivlIrTKl8wP5+6m4K9ZrS5w9tywLyLxE+H+u4/UBWD360rr05940JCT7+EhTPv2ha
yBkXcudGTszsf9CrXEgm3g3ThTXFHs8xW06fNtDxnuJoOkngSgWy3EQEFWk4p9q02qvgpXIrZYk4
3EjLSLgk7j68Ymh9R3H2WHIMS1yXBaKY5Km0mHcmFRGNok24U5+NgRlRryDqFqkYNJdxeuSvHBOu
wcilG2bf8seQtFp+FA90cupt+uVagaoMA4oo15rbYZgx5v29Ve1qcpdDbnB0fSvIVjccHtnCmUpI
G640AVuOSiE5lf3h3DYEl2rsNBbDhrDnkOrfuLOTCB/G/nC//Xk70YGhwRaggaHhS9EUFysBQ4Un
PAWtv0Rel7/n8L3vkpDQCaieOfTuCexuTYm5gkiG+AqhdUew9d6ufNGRsAJzg2EJMiHnqjqak29Z
0ho/DPCVV+DzulqOtfqEAKHcyz5EeyXwSRktlx07/jFAv6/KadXj5Jim3tUwt5z9MuvMNEchV6dx
qmOsgEXYaW+33fdpq+6Ovbm9Id7/8nrsXQBIGOsSYHMJk3cJwxfx0G6DVcwnhJEgJa37IKJct8t/
D2/0ViYOIe2brFtyROnHnkwA2piM860vg/wcnwu9sxUCX30G6NY2GV/cv642s0UP5hkFAQjD0Arx
Ec7Xqr3hUOcnn0XjtnpBhQjzZ/VwrVBWPVldhSN0mRl/ONZlLeXJCK7fvUiBhIa9QUaZxjyUT88b
EJildwM0PMsYAyrPawBfPxc2b4Iwg9J0BgJRowu7DlHFq9oBm1gihIgqe0ltR/rWSjGpC24Qx85X
YPJ0A3Xj8JQz2N81jheDzRXmW5VLAUa4ifTGRML4zSIHBLahEFGtsj5r4R2TNiK+yvJdIOmu9R4t
CjIaDNAN2VKvMaMjPvZNeEvW/bbd10qwIxEY5ZPqA9HFeL1A75nxVKd6Sz9aOxYtsHlQ+zY1FQJq
yUPPWx/vmzkzjH+8BQYilT5Y0kIHzhYNjHjYqY6GPJ1SKpB8FhkFL2qDxi6475YaRZrZqJupqGBO
d/0W82seCkxz1FfDzVJ19HC7k2i9p0K7xRhF53jhuisJho+CYejnWRtD7Sq0WzaWteqVdKDNeJB2
ELqqDPO3A0QZD2yeRuCVNFxPi7jSZxbsAetgI8cxN3wGl23/CFlPBc/ra++N9LABHK7NAkG2KsFE
I+OaUBMwoF0A4e6KYYm1qSCQhQzGhFI7zTyF/aKC5b22PbDLmB4vUq7ZIDvDCiZGhmDNsP7py+Lc
2eUqKDVwBZ5cR/QyJqL6qymPghGtyloCx7YFDOfI3L+6ewtZNKJ5FuuYYVhaOzlYRMpyNjZfcMRQ
Q5P1elHA7ICobSbJ610wDu3mEUXXJyV9xkAV3IK3N4U9R2viGpb8JEvc1f+ZyRuZjRH4bv5yloPv
ruJDlwrNBGEIibBz9b78rNAC/kNqwn3QxSM7qCFDxCz96NxDQJ7j2+1FF92cID23CYSY7e6Bl1K3
QgM6I2KIZTKJpS/oZLZXlhyTEV92hwPL/12R9qDQZaFIqy1cxaec1cUAu5f1MWIFydJC5ZWHnplk
x1PhbBNN/kVoZcoV2ZrHNYjO1FB/rkr+RgKKwqTKedFEQv9TIZJls+MtKhVyj5dtKqyc07o77tu3
QqxrYm+LbWUciXU/n9wC7u1oycPyQ5NEKfuExP316qER2kQW7vPieN0v1SDz874UFOoxysg5+ryb
RyZSpLb5b6ONdK3zHePOYa83x/7g1R2v2MIRNaCTabsylaGHMk7uG6/LAYwoV7rHSaOMK0HolLFb
F55QAavAraTOHWjShj8CoVtvCwdoXhaVlG7jDZNdJ2Ssy2YO3Ne/dEZmuXvrhDMYrcfARqJ2XxWN
ri0JmeLb8QMVmoJ2SDKssws7vU1bKbUKuUiOhGPpHJ2dj9A+uaQwWMo9l9w/4Od2rabWotE6NeXF
TUZKQ2uhKBr7IsGP8TK/SEZ16PhHgecQw/pWwFsS7ZKQt0kv+0PpxTBEkfQB6mr+LAonjhQWSr0+
jnV5/F4w30ymSYPhHhMY86oxP4veKCWKGmyebzIjjzXb5pyR4DuHKEkyLRKdxT/a1R/qc4d/344C
M00F9BymfjZquya5IoDO/4JVT1lu3JPAmLHlNd5vV5g3zmDcNMndK4h5P+qP2Pja6gYi5kpRBdu0
IGYQ3WMvaq//xa/ren3jVmXhw7E2xzf0KxxPNggtVNElZgLts8/eT/2ooV+3uV6n0xabIw2Ko+4q
jVDormm/xAgE0NSE4tFkYWbF7se7/N9aA42Zp/vsjL91ToH8qYnR2Z1L2B0gpKBzG72DTx92Jl81
TEG62QTTBgGm8Yl4xUU+HXqmrqdU813eGcgZfwpI02Xf6mufZhKC2++mpXH/ihikuGRRgsKfiwxD
2HwnawAXXHxJO5DYx9V4MXgbbuQe11iqwyr+hdtzzesE9BPcvUCnM/9VolA1OTrw1JGgdElXeeFF
r3XMDyJWE0NfVTBNTZewh7HmNE70tATzK6JsJVbDOllRitMqpp/jtLVFJA750bjNEJgUiLTvWBbV
zkXnsZ3qx0tOoQBr3noGyzUAGrc7ZcCsKl/STzOiX7Q5Yr9hPql+/9iiEpEZDxLnyBfl3bhDCwuv
FkqXPk+M6uyM3+GXQwb0d3OXNIAaRuPb9ssoxiGEb0+6npskUAvWjpf7/jeHkhmY3MhQuYmpikP5
l3ip1/sR7RBVGgzVG+Z6XUs/fu/BFD8DXjahBncINQ/0lxPz2SZiVxePqZ67ZhK9JMnL2mRUIJtV
vQr5vGiYZJMgwxOCcZFEO5ivaIVfK8ItsEeFjnO0w1RevY2a2cbj/y6gFR+ahHWlOKct20DwMr1t
32x16mK/93ipR073rC7mnVI605u/ic8FpkjJPg4pQbqOcno4aIp01/4zaUPMz/mGz6aJa3ENlXTz
9qkbPj3cAqBD66k7gOixrEttKycUojUcmHGDWuBpr54hvUcjcu2rypNLRxZDm5/3vhDWCaK6vk5p
BV051/kRsLCbyvFGtgwhxwOuRTYgkDs/8f6CJLAZnK1PeFPnAUOhsYDn4L7CuaqcvOhsXU6m+RVv
CQLhj0aqFq3lqee5CWPhtuZ3NU70wzQK137nCDCAErTuaJuTLzuttVPgrWiuRN46rm1M2pAUBUVB
m7cH2fYQmCz2FcUJGqaZvk0Ki8koXD7UuNkFL4jTt5xMQhIoiIZ5p1wYGp5rZv66Ugs8ejsDN5QQ
Em0VGJKds3l94nUdmxIP8Xdaw3mCtvmTSmSsjCIN07S0FtRlxuTALlJt+u0yLJTAdgW1aniakaqJ
w5mbNWJoH8/WK15Jby1pLag/UwOWLCD4OG9j8G18Wbuy/WPdgyCEbIdix4cCW4CGd1h3+wxS254c
g/IpMr/hzmeLwpW68jfozzuSHSKlaR8CX8J/p4338KYQUlFc7MIjRAEwmLlm5E04XEHM0nhpawie
KYWgYCzb1GeYdWNxaeJM8I8nH93r2YnC6Tm/EM+frkIDpLpfo1coTRfpPfj95DH6VCeqcPCn8WVm
U/zpzDZVJyQr7qUyONyY/Bn4x6mhqyAPAz3vSEj/bC2m2ZXiXwBZU8uOXeWJS7E2ahKHpI3zrAyS
K0s7Sxu+USz7yKHk3qVy+P+UiZMysSHglBef+BEouQ2+h6ztz0rJfApU5CIraDlLBr+F4JKznYbh
mFHzf5w91OP0yDOpThM6fjgjWX6YSye61lv9mjeV8QMcneRUq1L8aYtwMnGRIkfwnm5MAJkT7ZHC
9TExDoh5R2H3jW9JiPsKoBSeltQWp9CALODTw4mtsynF7QtngjX3IhHWy8+SlwBtplh+jnZaJ65Q
iHynPn8qGwADpJ4dwoGIk3ItqVjfNn2Kgh0+ZEvSI8K5f0AJj5o/usZ1+l9zL/PFj+QxPc2fewXk
EV0svH2G6DI4gbLl1moYBvhcyHT4JHhi1URVygJNgLcefFMQrcdvzJn0U0f/6L9jUQFLwiHe3KyE
RFA/oKnCprVMv88KX5aCThZXqX7aE5mlEURDlx8SK7/mS0yFzfrEcIlREwlhoPnGCx+FDms8qNfX
7NYGpmnHpcJq9TKA75kd58yGoQ8Vo89O1fW6oGpANjslNhhPaw0b0K34JjfmLovIKyR9CtHAWvgY
MQrQwK5mGESwCScwzSlRZg43vjsUCXgCy+o8pcuARtcPs+Z4wV4WKcKTb7Be7NRZabiq4poYPhMf
vwFFlb0tgwYCoYspexyke8sEA9gUmZ6bntp5sOCS5paSyQ+bnQlNGQ9MPObxjVNC2vwPAxHt2yT+
Kul9qJc5ERc8UuroqAE4rOxMn/AcDLcnRPvxuOTibF8lY1iZBGWHKyEsNbBNWTU0L07fBNQ/ZY63
C7a4lX6Yb5mNPKQ+vh3+O15lFl+kfiEKA4smt/rQXN1+Rasfmi35+DqH3xBDv9TaDYxINnpfd26r
NwSvhQB155545Vw0vqdMsEhoCI100BxUyQHW63KlSwG0xtwRCJ55y9Hghz5F0uB0OtvKy4msQ3zc
P0y5j7btNXLWF7sxktWaQMQGqmpmc7ePztFz/n7PKDOOJgBNQtLO/fa9T9sqrqaqluUBWp7NMYoJ
QyvJwEGXA+dOpIsoUqeL90YJnFg15lHACO04GmoBovelmmvaBR6j4v5nllL1njQbOt1+9FB//mxu
kVJoKE7fO4YC82SHDr+1WD0SN8YDwPK5TUNVdglfPJnHZWpTt9oRpEX0t8SlWQ4DTQSWnrfWPb9P
FkyykiQgIUciOAbVnSR34IfJWuNOqbF6ufVprgML+RM5eCefLmkFuo5vFw3pqHdz9jOxM4rELbip
ckOfHrwMhBQdqOY7CpAUKO5VZTlKkTZzVgVcFdNPvEjD3GU6gsel567Nax5/7TRpobez6lGVWX/h
/6ukawsaouyUvW7uePBqTUwSF3MK/rjtNDueTp38y/xPrFTszSv8B++96iaOi9dMh1EQRsNMANgB
FiTuFrzlMkw+li2v/WZ9GvKhq2rGbansi3STmRAagmIN2iihGfRHF/cgxvw8eWY6gBcB+WpqvgXL
5RUSExPdrnZwrzQulpF23MigeBv4au4fboySxxhD2s79aHgoF/wTIdcLuSkIufNnNVVo/7zNx4j+
yEAVOp9sPSljR98PbPSBi07CvT5re24Br8Scg+b9C5xPrE51yU7NPEWJeqlaDbtRDgLR8VjRZa9w
r9j6P3a0tK4H7S9KsOkSTZK8dSjLAkFwbceL1hzbMyYOdqeacYKLvGQ+jGU9sCg9By0BiMEQdVZD
dqaCbxZA2fUptOmdBxu1w8E4OFhrUE8S0uxGw0Z+FnAFSyZijBaXfvLJlBhBP0nF7xddE3ZLhrCu
hAJ4FujjrXLu2+XL1TjvFuDr2JKUuTVr44Ve/pf4RuvQjfVax8VdQ6RPUOq7nIFTCqkAdzI8YYmy
+jL9WZ6I8BtnB7Kksv305PDpjXv5ymgS8QKw3tHtk31TPYovwbLryQbdvDasTPcUL5vvGwU08HGO
ZR7h6+23r7Rh0dbM89Rdj5ntWZTnnQH1UI0QoiLy2OC7waCA4+Ufmk7C3dIkixVnICz9krBLC8v5
mSbO2SUTAEZUaWIxeMBjISS+Cucw0ZqPYioTrPWNHQOW2JQEVIqKPkVpNLPAczVClMF3rIWHW53E
c0R3fwBzb2RuHnFlC1EPFHYMlNkHFw+g5RnqzcKNiAFMCoZt2Ej2pqXnPk5cVaM6j6H4W7evsd+1
PCRGijou9tIo4KwtGhEMVsU0yTFXgh8rgGPlVnM9VjqdfPSrOZ2cWvy21mekAHeTLeSAiIJw7jDc
XoScPUa8UcwFJ5ukyiaiv1TPF9mCytOWQG/EJyzbIhogpHtXZmr1rwfHDgBOkycQbhVZwpDep/9K
TvXyRVaxILvZKakzDqr5vAImBbrUZQnKODxh/iVO5Aq3+8WJVEIovBnupjPZsy/vNnebwYQBYRgF
ywHUDVrLIzDwfZl1IGJyq7gUUbf5xsHF6uVHVi0eAdUbBAoxkUxRvBV7Q0Ih6DuBmK69HtH985M6
TeL4JvRgxRHg741uTTyhUQ7Ja5bjw0mJWryl1bHpxJTjSOGuJSA9fXJnWq3GIDX1CJmnKDKU+eCm
ewYvqeRxgwgzQvox6BK4dVaYBg5AJ66OGS0RjAuKRwGd4tS+JxH6nWnlwy/97iLkWh7NVciC9Sg/
/gnJ/NQjsgxMpaO4RzFmQ3NaSNHLWJLpXbLFV7vWRdKYOJOhCtL1KrUlIpNVKPf2A2OKrEs+VeEK
gNclC6m90PWqmCy9puuNYRf6jPD/3VZQU5pgwFUjCniFbloyNUSDR51L4+1yS+AWu7PH34Ea2Yfo
56sHW497zIlIkR0yQA6Z9Ry+k2sdR2IebiQZ3c/BQgD7ywyHndjZPdA+unw7xXwnUfnhMXc0PEof
9FGWVg30b+F8iOr9tenb29tvnNmmCyU9yT1RzQ1vzLrN26VbVG7gOA0GvmtCFU71Y1pC7WilBTcC
vz/AIiV/GIY/b59Vb8CllCaw6FbfeB/q2tKSiSMTaJGcgXCrEhgqlwpPmYsJOEsMJ14VGBjEvHsX
dcGGMtzQsFuI8mMRlSz7+rWLq6hfYfPPyhNHt/2lqgqWVMJczSzwv22CzRrgvsc+s6oofUlHpLBs
HjDD36v1rM+d7IgkWjVVhdLU+zxJUxj5tj0dKm6cCs+Rwe0crYH4wUJO31TKixfl1TrUqQE4M/dP
5XLyp49ne0Uisj6Z9V99xVfu2yEloRgLVPEgku0QHqqQGgVe9rEEeUSsZXyeB0eIYKi4vUuR+KlQ
k3hmI1anDsWYPGZeUYN9AWri0DgWL8/RQ4DpbOYeSs34bi3VwVbC4dNtYeeBqgs4BOBeqUou8ifu
Is5LEmsGvnoKh7U8i4lESahkG2FicW6gyVSthkA15ATsXArdL7nNipCe5WWq+fi8eugvkmyRe3yu
cCqrujeAQj/eUm5/YYSmt+TNAgkIDyYvaij+NgHDsyiV3ougNfhS0koUtNvROF8b5Yub3K9VzYqj
yUuTkG96YIdTf8AYxZ3sn+wUYoEmi7WDjVETyW3UfwhvlhgpBJ4Fza3OXZ0cxR/YlURnzPXsDtEy
kLTmneXIFUO7mp8Vv5R14KJDMOSuGiiXWi4vzSLvk02nbEZlh257+6jp+CFNBGGzICOhl6qq1yda
O+da7FX1z+XIvs8nglunws5u+hJAh33H/Q16R8YWqSCKTs+KQDaE/E+d632JVvD+0TXMUI0ZQzDF
K0uIdCwaTJlgEZ4WvqiSi55S8EvO6HYOnN1ETGuKL0yM7uXbVYIF4YyKQSJPIuNL1VGBYABYX1Z/
8hknignTNiDOtZK8VtUwUwhONxsmkYEy8yWPsZI1b96ztMn0PSQAHWDrzvwA0UDXyi36D/F1IebM
LRtG3F0iJhlVG5ITeKO6ggNmNqS8djatFGp4+P3rvP7sWo1KymCXfLnWCMH3Z3DLXXFMhQc8DDu6
ozi2aAoE8KhXmMMjeI/tQXE/eAB9T6CU23zYOe2Glk+g2X2YWI0akaWGojjpv8Ec0N1BTP+Nmzjv
crdsIgYyzTAkIJUIUoy2Xjc/MHkERyqLaNsRd9bxN7rKHkwhAS57/hgw0mSzi4PvlIt9pB018UoV
4ycjOgvA37ejDXHTaoPLz1+RQmILID/KoKwPjArKwO/0+IREDCOhd1LVtjfDFEu2rHpQ8pGkIlFq
TZI50TuQR/mw+LY6S5Kb+UbOOv7E34iCTsI5XL1g+NMnL2X/dJyD3s1ViWALfuLAyVKFRdlKg6sp
g2yhQCPALUTSmvQsueArqRIB5mZEYYxg88KU824dVHGX0GLB+vf1HbVRrzF9/4NCIoVYvOkjmoCk
YBEU+VCQ14vZyjDhPY4OVPeZfBJRWP16xaJAUXzsmvXcFkH6BkqKSkcw4qMUkDGjJf3H51p0HjB9
vRhvlIqYM6Fcst4DwfTr+pTjz2x+/ooG+0TKIXtRHqIEeR9XH2b+8jTqdx7Tyzwo7NKhjtGcxHIg
K7q97/oZmZ22fH39Iw39DTtS2Hx0xBpn4attz/CjrGXv7Kh1J8jGYQs0VbTBlrQC8+y4k8JA2SgX
uDF4uAyY4hb9n57InN4CdxRCr5v+pU7LHWK78PUmGtW4OsmDyBAp+ovywBpkFX9/pYTrHFJAYsfm
QELWb5feSJ7DT713owPQWdyvlicA7klqrkUvMnt9Nw/jcAhRilxuM7aK102KuRo6NxJHDGEBSxyE
uSuTG9Y48HA3mUIvpyRSX8K6aX3trFEtr3cSfmjWNfrS7X1b/9EIMzPaDVBmao9jAXiQeczUlguB
cwmBGtMv209eH/bapgndX3rySYt9KPnMfYi8DI6JgIE2zOfRdcIBviRu21/tAIsXZ9vHc3TP+YQ6
1SzFvZ8Re5jx2tH/miwZfJb2RjoDYydY5HnzryC8eIEPle5UXCGqGBJAxrY+aQ7tlHqFE2QYhjfu
ndUrrtdlKgqaOJSiRsAH1mKRF736OKv/e76O3rYzQS4pbeuqRXfTF2BL9sDw98hx3g3ibTm98lRz
3WmBAm7A4Wug5clSfaOKDSws2Fw/1aAO/nnvLcKlNSPGKeELzFLKEKzm1ztK6VayZtdMnl7rtF8p
8sKhQ8NFG/AE7BCLv7MBFb9OmBGXJQuScFpmzRMYBB7IHUCbS7HbSJ9PDxQ1qP82gfSqHfL1vWnE
6k3hBpTXpBzuz09ECbyfz3xdxPauydD1ceLe99H0Ee5ZKkDxQTpaREjTXWFmmi5xEjAWzaH1woo7
OdT38BWm9NBQSl2qOXvbi336sfAhYT5eaK572IdLqPl45EyVckxB5kFuUFBjaJP4+em02anDYPtP
/+BEjw8T8/o/yTnoceGO6DrG4I01QV8EzzCA1wmwulxhew00fhJ9lpjII56jFJy6dP3kTCCWJHDL
TjcY0AYcPgIIm4TEUcprjAPXPxbMIMerzuESnXrSDdAPKDwWa289K19Zz5PN60+KoJqdSrw7zVGb
RZLET+oRS8Zi3opx3f4Zb+blFH0teKZbkg0Z4V3jSKAAbtieHgrx4DVn6yKHdX6gez+cALUEyPYc
txtpksZkcH0rVGFrAJ1MxPpIy5QF3XbMbqmAiLJkcZp9NKpGyKKKTtnj1D+7pVihgdlHFrBMS9Zp
edX771f+C81uewPth3KJgGQEE6TJlAGGoYl/cZ/5gz4TDRM2hFK4L3+wweE/HDrDrfQ2r66hpyeh
/Up336S7w0eoKdQnlZQSpnryaUubIuJe+UyRebjRHx6MuT0qAbokrPGSQ9a5oIPFLB4QxnCRcfpN
vu5WubDnbOWaZLQOax88Arj783Bcy/ukVPCmsPXZQsGLZuHTLVAO0as7r+z/SVFKQuw+eeHBvTEg
h4beulX6LJq0vv5Rr9mCShpwrhIM+f7gyLd3yqNGhDAc2gXHU5zWlUFtmpoLAJqAqz9mSI6QDTTd
YKO8pdm0/9IdtlSS9fjSq7eNgaGc/oWG+whzYIEogEtw5RVXl8uqfL8eV+vihp4lH6ZTzoaAZwck
6o6+zszb0qfxeXDSGHjLaxbjfZT0bYDZmfGO6C2T4uoXTm/knMheChYk9Ds4RSvDnTuL8hyGwhIK
OMfmk9Fougr1QncRFsAriTA1fMJIFR7K3nP1FH+mQkI55OyILFvLq7Jc1E4+lBCZrinKu349i/0U
eOtZHNUuI4qfd+DJDcen7ltv95Fcr7X8h8PwRCj/ahR9BL0jhrLZiJ2lmZ+DMKiyibCgSYotaWnf
/lunVt0uP5BZ9iB9+5IeP9TH3SJPu5xWAMcgSy7i92kHyh3f3KhFw8lC8rl7K3LQxeUPSo0lY265
iM5CFbsTkWnLJXwsAa+VXrV5ygNqMpy6k45BL2e650JDThZtjK05O94+RazEYdNFCXtKznlDM552
D7ESZavfvDSB0AkzvGNIQJzh3rGhqysDX+ytywSJpmF3F0P+inMqd9K0iHLlVR2dGqzqtGypdFcd
l/3XwJ6veCRL8jgzNvrmXJz+iiwefJCem2d215fmyfLvRNy3Qs/P/UFIbLMxxqVUOVKk9Nak8+Er
tfBE2La9JTRoPihht9mElXDzuXvw+t3t9h4iZsQowSeBao5+Mz3u9iZM8dnZCRe+RZPB1CHMfl7W
QOdv4MCJmEjpBkCqdbeXx0TKh0ulw64POXBkyaTkxqlfPi9sP6xXHzg020vtRzSSRc9qKBEe5nGZ
rwG58pn1PEsuyk3ymAJ8zSdJlGpxp32sAt6ua7yTS2mVVnrkEC7pEaf8oqvVWqsJaug8b7a0ECkq
oqnVyRfGH8paxA8biCaUUgXqUes4FgsEdYCgR20nV1eQWIEK4d0W81tqmTc0jeiuUlbV6zpKgVjN
aYPS/2s9OLZ/shYDeGML+CwMvK515P3k1OqamlfVzXqSNLP1PSqiIS8h06CPubaRWvr7+dq5r4Io
xPk9xUd9gfUJ5UyTOIvmUmZ9hpNuJqI8x1aE3Jfx6gsR0onsN6Mjz5B1uiNdGyH6S/zFbmD7HjYH
kadjEJ9fdK7klg6+qHVijUN83PaLehFQUyxayvOYLnBVAThigmyxSctXy2WEZus+PhgW/Vvq+x1T
aQYka4LWrHZrLXNJEV3buJiQng+9jVqe00bzUHUi27msW7GZ2wqaHxPW89SBg5nWDlSYpgSQOrGc
M1zTUXXRqd77I5ebSgbD4KJpQvVnSvxAMLoKC9B/B0fFnq0Gv/hGm6uShCH1mPrqh9IBR9dIPFuo
TVsnsrsJxrflRDLIqUUxzAdYyIm1G47Mv2p1g1vRNtBOb+W1grcvGKzDwNdpgrT/QmWY2kY447pX
KxgZ+ZeK5+92NJt5zlr7vL/7CUJT2FuNllH0isGhFeQ3yL3/mL8b8cIjy03ZYmvU/62W/W+89Mk6
B6z40Iqm725wK73ujY/vdbtyOcs2Eaxd7sJCpR7XxFOrfs2WwxC4vLTIEXlkPbW2y0N7iSMq7gtX
JV55Cc1fGugeTgsxgkFmdhYl8Vwlx8jHHm76+ypV63S1CeaGRgT15s1xQ/mzbYQt+jie55Lqo+Kr
qe6fnkq9w9d9HToDGqc3bvbmMl12PZlTBAAbhvzNgh9THF16uBR/4eFnZ56m6uyn8dfkqqUCE272
OeiRY0j0XnK+6G9+lKJCKo5WEDyKHZ2zzumObokBrb8NGfCty41HhJtg8M7P63aVndizfZz84dc+
m/V11X5fW2ytGWE/v6K0Q6VONj1gylYvau+V2xwKAJMpxADD29CSt35M+hkPBIOo65Y1+eAgpeBT
vAzEnSDAobgHa0Gl0i6XxvquCOtX3xgyrl3BkXirMePNbjdEmjVlrJydg5J+9k6dTeC/t0IWELD6
SuhzOsDNKLVh9hSmKIZF0fDKcYr8jhk3t4lOngegt+48SAZtGP2o3qGaFLS6PpRXpv+uegZE4YME
T3jY3czUs4bUj+xr8WRZPcxvPRJ4oHKHeM3n+t6usrywWMYwjztj/FTGQt/sYx3D6LsM/8TERFxA
A63umYaWI0BGiFp+f02u4Mtdp7o/IXpcVTGiQ5LBs0nQc8tJNb/6lkj2QGN4hP937rM/QPY3nfYH
u7lqSXZHZr6MRTTaCwMxa+eY15QGP/iRJq7FyWizaz4SDCODAAI1P8+jJpXs1TkcVyqjEoAi2Y4L
V5+FaF7UvedHrqQLouSfaHjq8jjAlXhXNgflWUxBMx7Q+6xbQFxwatsnN/FFRu6gp06Hl/UMdJ0y
xLy6gB7xlAEDz6igbh5BuvlUoRAT9qDNy9m5ZnaF7Bkv0kozfSz5x//5sRGR/mgjDRxrz9GAbIUe
GzZAkg9U+aQuMgVSLhIQi0Law6Y7bX5L7D0VI3RsdLI4lYTMXcezrkXOGXys9NFyVQQGayjQYQ+j
ihwXFf7S5iwAvHRNt9btUCVeypxY6Y8W7sP6jxaMYnu7bIe40AKKiIA0LVPyxrVTKeYppcLesfwk
/HlbYIrjUwwrIql7ICWU+bil9gj6yNEr3Vkt6Wo2BtVHcWwK94AJc+GgdpAISX50MyW9tyFS36qb
yeIrdOL3XDmeYPN28sXhZaR3ik0yfK7qx9Xann45XQqOFA/h0S6Hb+2BEt5AciTO8F5xM+orYA2+
Ey5uxGtlQkxgMCoIEeeuwYgRe10wpqqMOFyXv/A8zj0wo1bbtuq1etazry9Em6OlMGailtbTwEiH
7AO2oYfXYuV7eTODkwCLTGa3vJAZrxvPxaXb5I3q8cK4fzz+0mBssOenNUc3iydqxWZX7q1h4n6s
+lNHlITBkiccB99lV+ZuGh5yYxTt1wt3kdljxI9nqUSyQxTdBDFm6KTaYkOqrJ0ZFLw0bLGu+hey
oqza7N/8HICaHHDeYNflznHOzGYpHJIy1E2r6B0cPhydnJ9Mzw/KyQz5hrNgnlfOtJicLxV1P8BI
BSORzj0VB5QlG7LZJZRjyWqZUrL5BpIp31TFmvAROIPLBGCwglvuXFQk4lfH5iBk2FeX0/vnNtAb
YpWgQNKd6E9+Ev41IdYtNrqnYAMy+UXEzxImB24oxjjMhCWdD6YTR8TN/LOvlEBz5xQ8DiViZq2v
itwKjR3PeamoLFx8DEKPMWGZZMGAFOsVWoW6Ti+cOXkdRM9Daw5j4oIRgRYOVLjG1ifktwRq/Z+y
N8mO8ZwhZdaPNOfmzxHRwvYi61aZBv0O5erpYn35My7rY5Wau5gjRuSDT7WYFkM9gQ4avjL9H0Nl
Ap0KAsmKMyzC7+oFHrwAHhJfJwikeay9vEB5K5nYV5xjCitXrSWZnOUkpLzpuDVX6/O0xd+4ZKlY
5PGSMMHVH/pAfkCFq0rMnDHH+Y8jaczQYY/RpXHYzYxnTuHVXUzM4O0kviIQXAbTYyy1Kj2YFVAT
TU7sRt1aMWRdf4WbfDwVAplBcLCj1VJBk9P2+tIBP+tL7OHeZ6MM+vkcqt7CO0eDwAuqcpnlc97B
Pk0HxdpiMNtibreRo75LHTdsSNF0mLDZS9i8Cwdl7t3avh5CrbXJnFboEIx6j8Uh7nbFaI4qWFuy
9e8gry4DtH+RsKLwj15n/QgUCVkr1JVia/bis6MTPxRL/KMwaohG3AhCqnObxDoFwGuFD4ZB3Kof
LxjChhGrzJMdxTpfJYCpNTRG20HUL5/t3JeXd1D07YVSpP4X3vBr1bPJxCQb8QXf4l3tqdHG3491
j7UxoUmi7PZ5RLAJrH5J/2TCv86m52YPdv2LHC5B4PU6mrcjwOw6lYsWlBw9RuoVVPLFLLgqUnj8
LeK/CHMnp42kjtZhdaSxlI1CzGgRABKmL6zJ9QT5/agQoizhoqi8N46XywhCkxN/TBKTTOzZxMHk
Ouji5jTP5WA59Mv2g0orttBpkH75d3osqaUjQTK65slakGjcknuO35xxk3oRSGRFCMtWyweVen+g
2PuogDhvxhtL48RQeV26idcY6v9iK08GfIgFjC7FHnfBdV8OUIxxIa5+YfQoN9cjf29/93Ovjebs
2H0sd1fIJ8FDOSIi5OtAV4G/m33Y6/6/q/O5xHJ47qNx5d6OwPBIuDX4jhopwkQXm/bU7rqS7AbB
apiszlVYTgzilMk3dt9PFWvwd/G1fbGY9iOeTCYqgcJ9yvwUZrSygL+sDdzCAxpW/4B97cFgHWe2
oodipcjuWoIpvdODEE4J58qBxj0wfbAv1hPXRL7FckyF4SuggGqTtXzmOetClp6pyVSrDMDhzEuE
XTnktxoNpRGQCkrYsJ8TOEOE5DSX+bWPXeV3T+znxOF7KKQ9byeIgvMMrVRFs9QrWubjtzVMNWmy
mgSKeItshdr+9Mssd/tYB/qKwj836wdv+UnZEtzWp7Yk2d0Z2Cr4GoytmlGqElDGfNY4nsaknVqw
Y702CK4ZqA11TUDeoc05zNZVTpWScbkTT4lYNRrBUdL37HS5me2dRkkvAEn/7lciRaw+pVbH57Ib
dfuebYKwprCVzzAba7y5e4GM0Ox+eMsW1LrtE0/LZbsjGHPSNIu+6mkSFi4vXjib3Sm694QigJAM
UoigyCAzcOpf0YWb9r51bzcQNeVskO83hc+D1+VAiC87NW35/6OwE1Fb3N+MhRTi+BwxJsHYhi+i
U49FMDu1ERm4m91r8yYA/oLn0nC7Om6vKlIAvZMk9BknxnIx/cY+qDDgbxcF6xbkPVwfPAi48mOx
vIJkx6QkBVceCY40kVtDtLtFpVrhwjL3qtgR61LGl3AvEQvi4w18Q8HoX2jai4/2eIyfkbZYUPO9
I6pSmF4VChgfPXRDijbU3mpdKhUHSDo6C8yKokvqLrRimBdTJKBePL+d0tYHZObqYZCitgE1vbdN
IOkKv0865rqQWMsWpdCRzvRCYBK3wOvpP4Glh2eCGERWbDQzp6PbTCuUAb1pngxgCIU0FrWliBir
AlAYPzUXYSIGJ8eqDpMIbzyh2X0SOlNSrSohSvXjQny92T3gvZT3x9wt+gvZKPCEXvGC2P01UrO4
mRSYWuwP129Tz+cy5jlo74UIGuWXSRBQZSUopGkxrJ5NPwmK3oYUbU8vjK/Wqq5ctHAjZ0MQ7d0Q
b12wDP1Er2g5lys1D2vUKIWPJBs0hLv/XVlOuL31qCPl5ZyrQuW0tAGAyz0E+8+pu1Si2rTX7poh
WPf10UPaEkZeVbR0l8oJfWq0fmT5Z+vVSp4W3HJacDWCpilIBvC1JqvFNsL/LzBSohgbx7KfZ1a9
5VF4Dm0O3m+KruKhzTpZmu9TC93ScxFMdXh+wPv73MjDD9+YIGFNQnKudeUi97FG4y7oTnQFikOs
6OzbgWUkr3G7MaLs4GVJNu16zeeoCxeTopUUZrOEzFj6ZatcgOZu6a+wSYQX1QZCEircr9piwku+
Lw0LKCaUePsmWtmIyILpsRegXLPUWI1s867z5QD3kGzHURx2jjZZYDgNMEDMGs3AekuAPrb8Y7Hs
Az2wlt/bbpPxRKCz5D9EB8T6PVcrZG0jaZcc46UvEQqT3bKkqzfV0I8vB1HhS11nexhTVND6nKVP
/PlRPPiGEA6RRFDD4fpk1lacG4bXdikJtjQ7bJXycEgW8+vaivt7jS6/7xSjQzx7srIvmQLl1m4Q
5d9u6Pzhp3v90hYjAI9tcptdJl/sgp4D6gBqVczC6h3jc5a23rbOhaHwP+uIMJnoKCvIha9FOadI
p0IO1597LVN20NOXxfZOHJiWUDmt3o8X42VgfchNHrkEihoQDs861ByTnbdpv9ZCTSYhpyhVZ+sD
TSgC0cbE1EJA+FZYZMIEocmCKGNNdV4By/LuocuaL2UGsw8/nv4QDTj4+vRIDFxDZ3f70DedJZpk
xSM9qWpBJlAoQ+DHVKE9VeIxcnQiN7jhEiRvznTqTO/NLVVyPguNPg34XrDMNw0oYP9mBbcmqE52
Z10jrmiFksqoqblRb76YWKjiUL/PFsRaLyOQlIzRB7n2VgEuaMFYDHMXkp0q/PpjqQ7HVBdvuoni
/4j4NyMKqT7VR2urtDOxg5r6kuA4fL+CwfqwasLX3vedZApKAuKO1I54MuaYtqHjcJHNYNi7RzDZ
oEeYPjXlWZC+DjZCvicBYiT256mAlrPmJ5f3zpUGBzn+jk4egTIG7HzNjFuOne7Lvnf+62XJUEav
WrmBSOwv3pPKPGs3HO5F1m2bszy09ngWyjr1dFUzesUQzEOqKRbnt3rcE/pO+PuJMm8OJXNjwOCd
3SLLbxdi8GC5wqE12vAYG139k7PudluL4BuGoY1JByFK456OfjSoBMmDQ5UjyjTNN9Af615gCNNu
o604xDtuSt3MsxARRABqJy/qlBnwy8wm2ZVECYhbemnykH5YPrRDgQlFTOrT+DLE4BSKjKxbsNmm
X1xMIrwfMBBk95dN41kwk6yGSXV9+6s+jUHdSxqHHSzWzdFmOjhThJ8ael8Kt/aWF0CC4OWJGS8U
WNWe0xuDpse6seX4T9D6QQN/Y1zGC3KJNP3/xpa0KCkmMjF+/5gp+TBXJCzXYZXv444eBs6RjDrO
2Bs/33HqkZl5fbKiu12A2fAulrcl6Hz3HMPixa0sS9Vdq0f21jOxwQ/YvvHOcwp1+BXvaOE8phRG
3plX/zeRW1a3HciRB2Mk3a571T5A29nQeKlsIEbUwuzlK7VCXwFzR81yj49tLH775Dzpufp41xpD
0WQlo2Z6Eg0k1Fa3u7+iEo/CCEVTVPzyHz+nu7ujJmYPna9iaH/L624X8ofo2ZtH7HCg2JBBic8S
BO8NXroHMhDvdK9nNLuGzO9uxR78Y82+WHDPbeq0HXq8HQrYFm3AldhP3y2tAOvXSDkUzs2OUUIR
9wbUdfzcm3GWMOCjAdYMQselYrw4sHyB2gB0oWtBC3DH0SIP/BUjMODyNxjMD6w1yucF7TzUqPN1
jH4DucSoq2H3nLe+qk66lvd45vyqCRtqLr+OHH1WiffIdd/FNU64T5J9bVaIZ2btNneFOzjWot3G
MP+7VdOelgu8zRkE20ctSOMY75avnSOKbV0fbYNx7IbAseQW4Z/+KaujJChad3BA9oh83vS+qifG
GQw2etwAJ5g3GLD3CIEE7BgkLHwI8y6vNlnRQ3+Qqyh8yzvvatxzqXnSD/uPTyChWt/FFSySkkHA
23kvrwKq6Z7+DSydf63EGhMMGkXv1CJTp+p2gq6/hl6ymgom5EOZ0/PBitVtKHoITIXzoj7i/LSp
iXc/RNphLInFMQyQD/x4h6ODHE5G7qdLeHJAoq1KopTOpFdfx1ZhIYYtIjhPtTcXDdodlBvoPLmq
lZC5ts19QT428n9w3T6GNhDyVdae6cWyxjFgA4w2Zwt9422tk8AKbGeBqiHZv4ma7uIDFvR8v2jn
tKm6mEg5rBhy2j0QJMZiVbG2ZpbL5tm9l95+kB1cPBOMCZP7YL8uwpsnOIYXFrQH61gQ4xBPbjd9
xTmpiT+XqWiytVLtnvjci9KY8nAdQBcONtHNJCRfQ8owpmGVHITOIaFi32YZYCEuwJjkNO+25cO3
MCJI4qDj6++y1tghKCmq752ir1Ze09WtmY9BNNFOuQYyO/4nLCW6+K23zbpkWdow3QG3RzV4O3ib
SMW6ah9ByGm9lmr04xmpnYMIg69Z57Gk30gZmnnfoekLjZ3IO6FfraSQ39e4Umzv+mg6FUY/9cGu
+O7X7tg45Vsv8sfJiM9PkP/LLFEI6Lw2k4omhxni8vi30TeV+AEuXT43sx+073okwMAiIgvcRwHa
sP812wi3JFEkL+n3dTxunDqnqbuIXZCxmB4Mu36CSIx2p1MVcNMz9TwWh4Kan/F9pv2LEjYgcZUh
5Fahia7QOr/TWLhaWTddp9JaBDI5ZuTM0URmtSgsoDn6n/MARQDHBjKMYLmR8SJz2tH3qJse1ldp
lr2GY6cwQ3LwP2g+vHVWLY8uoBaDtO95TENYg432Cme+AhsG+exJbInFcBXkfsv3WiKbMuTTuok0
GjTdckIg5xk5subfX+NP5LMpIuji2pn26+Oe4ngFbjHpW++N+oT/WJrpqqS3a0Uvw8oZVUgmRkiO
O46aNOWas2YC7VMJWmvhkuQ6dEfPfB+mLDEwOu3a5iU//mKImEdm5daH5faPir+IjH5RShNeI61s
VfGyDKgvmEX8g0CpGLfb/yhwyq0Gy2GTJiaUXe8tfgamd1uRuRe1J9/el28nyF6QDn8G6sPSM2AV
RURkMk9xb6mB0hXRfRguzcN9fi4orZt6RDrCrI/CxizyxJIWZie9qFxLpNucgNYdj7IBjre+I2v+
skidoT91/EkXie6Bx4X/SiuRXQfNuH91DCocoPUymgMwhG2Q3hkKLph0ZEzYYqD71PV1f1j9TW5t
7m/iaMiracvwRxW9IMqG6Z5TW9tJNkAce+iWLTZ0pKDVKgQkRBDfgaDgcNBi9JWH3HPITqYi8adO
CE75iansX8RcRiZmPxHeK/7WOtAK9XZtzEUT8tHMg+FYji6HMx3HlHzS3qNjGDW5jo7G9mmdBzBh
FkzGOJ7fSV4fCZW3lS49bvrfXaVZvMkp3ge2S5+xGCeEmScwfauFHzWL+LYpOmgueMWlShmbmj0S
V4cLrq+cBcmdSwS+XGSflc8WZNdUSSJHuUVqFt7K2CS0g54slo7F2I+TuXyLpNIUSNgYsHY85CRI
7U8swgBL33FJXfVfoLSZoQH7OO6QskgNtYGfFapW9vLTHQO/RccW3QxhU9VfRmO+mjDPH1NXbHKp
AKeb2GhbK041+CceyXtTAiEpxkurfnHf4zgtKocf/D/D0XJlic96SS9MpEucHMt5SR3ytUbJrlpS
Ye+LiXqPzQO7iIlFdJQGP9EfBc3jttU14Ov7gPPMOmTFepbxslJuvDUc6xunrfd/1G/5qYZfiPUI
/qlRtR92ToFK/fdV+FnjUsnSu0gsNUua32aYaNpUf3er8pwR/740OCUDKSeGcyRElGfWudYZmNKQ
BPP9Jz/o669c5xZVSxjRC4lob/qCDQuX9wWob/i3oe672K13GTWjj52bXvWu8HXb/niWzG0b1vVs
R2DO9OcCC9xWl6CDxkMiXPuC8tKmpsZf1RxCZ0obSAHHJ0b70H0CYPg9FKh2t+zI6VHaqP+BYjmz
UPb6j3zEZRfY9v6qkEZ5EZdEuJ6gIsSpLBNjlehYmB+4JJEkZ3KdARlQ5qApToYUDPweXM0v9Eat
1Lz8BrJcO9V0rZtlUZJl5qL69l9cXG5z/ViqEYSO+KF/XTbxUj7P7l+/7EPuO8DDDgv7o9Gy1R57
ERDAYI5WZTBGdLgU9yqutNi1sHdDE3E1TtS5oFjcmcCZSw80QJ6sItBIVHuJBHevy5QKuQ2kWms4
cTeNUs3ygyH58XvbA9SQIGxetT2BlVu0xWiE1thZHC2RgFZOJbcKHqe+WWXi9QE6A3zleRqdGGrU
QvDR6E4Zm0h8hDxo+/ME5I18Aqwm/8JIUtbUa9d0vzFh+wKDTmR+GKyHj/T3NicVY51X6BxfaLtP
fGWSsaSFRbj4p8MLVrU1A1IqAKRtVPFhJ9ChBugGOTV9nj9ZLbIEpIVCfaK0MydGQAanYAHwDfKV
aPghqPdS4ys6Hdn8IQO70pJTosMoUvHWjv7nt8Omegycy2N0Y3jLi+G+EJozCFkJ+TxgSMSvF0pi
UvxILvPluqpboFjENIOpNuUR4ZaRBUHXzSeQ5ongQ2GdoCYUqRr5KansFn582K6Lk6eKxGOy5SN6
yfnM642es5GNOGJDhkYxkmrwWfcXotWc308YtH+QRYNT+OQrb7fXXYOCoHlXJzjrvWJrwTJocFnN
o279Lvhu/ywppnslVid6NOjph/cQJHE/p97wGJuQIgRe0bTqWUZVwxc0ekh4YXEKnlVorFp+f5Hg
usAMeNdV+vpg78nNQktf7K0aazGY72DRq1+28SnlVeMqQkO1HdoUQgVLXcvykqG9uQnm4vladqmY
3BlHHpg5Tq5CWynnXoGe7omwJ116/MYWdY5OxKNRjn+62tXf8AgFuFHfPs1/KnSibz/nf5BhF+HL
DaBHG5fUaL3NdjrbCg9Eafm/NJ0/+g98l/ejAABcXJmP+DjNO6GtVzVvyoFOBQ4uocx/ZjzfDezE
1nmJSf5UQXlkcbOUspXKi6yR70Z6eyo2OcGUvf+m/jGrMBBh5seoGMR1ZJQGA9n1I6N7qfQDU/xV
u0Y7AwYeotX2xltHRsdzx3Y4S6I9ccaFhCpiAO7KcKY1z7fL2H5EBD3DLC4s07aV1Sdel7yGdEZT
wheZqUbDL11mxag6lZaEmv0bwDKvHyqFo4BpgFFNK0/NO8nxYPK1IG8aPJDvDVMk0XlIOFjywYym
NPUy0WZJskWr45R0EI1oBwIfPHgmSfh6ILoA55smQ0h4Vi105wJi+hIZNfGwublNfU+qN+wxC2GU
GyAGvap7wQeCFqx4dAmD3APl/J8PCwLCZDhDcxu9djzKbkZu6A3MPTg2elJil237CUWJu63b4QfZ
W7l4qWxBSDEKCtIcAHohw0D6Adhsxguowq66rF/sKUKBOz4pUHp9IWDaXb5Kqtikl/FYRk2GqQeQ
PlNnRqSne9u6ExeKWbRLXbysZc87CSIsuCZBT0mfvDGf1uwHTPSfqmC1ZxN78M3KupAAPiCtSdFU
Kx8u1rypjox4xqYIhd5F2kJQE+OjY//3Z9RJ8RFJAEtolWWBj5P0YuquqSBxuclsEAfdZJJWxE0e
u1kHuf22hJoXaDb8NihKEsa3+Yuyn6+zktstC8ruan37Wfm3IKFbkjHD6TxQnUvJ5NLiIx6BA+G1
6CAqk/Ngs0/aGSljVXqQJjO+iwwMVfd+W3RcPIQoVMYa7olLLLAy1dt6BG6MZ+To7NnBdafytovD
6ue5MgxGlStekONmajVbNlErzjpEAlW6tfwZ++/07S0j7u6UZP4Wg0mnx36gqHX3p2peIIO/50Hk
ecuzOewtoInjK3iwI6PlInz9+Nx1L2B5kWTRpTemT9ZlZsaxrGaiVmTDVGEeqx0aR5MqpjTbzqNf
L55Xff3qSPZujSjuMbHx7+R4XLcSeauBXPuNJST13bVv3LTwkdW49QgILzsR5m6SwpkNghKFo3no
CiWrLHn/wZe1Z3AOTR/yeggIpIW+NeMImqG1u/KFXF8TmzXYxCuT+HG/i/8k3LKXWbXG31TTrGnA
Kjmms4q6aCZGa13GMTlWedI7MhcT87znj0ClrqVlV3lQiwFAgVuQvW42R3C0eoVN1cGyyNGbo3KL
x3Pv7XY5cXzNt6WJp2rEWwfCexAw4MdWLSQZJ45BBjUoSw1reufAaRneSOHe27fGsq0tM/zPki9O
sJB5Oep0Su6nYfaifkXRCELVNGPX3y+Q4Q2yxkwGxYRinF4Kx/x/HLAwlp9OY0zeDerH3EFacD9t
65/goihCcecccY4qKdWYKTWF8Ng3Nz2ZSaRPbtGjff3AQKq7a2VMfd5RqDbzLGD99l2FlKWeFLCR
iBsx28otkZNTYaBhNpuOKX7J4f1TPWnnJHch1uJtllRCfZNB3Nh+hcEYSeytuVHmqSQJNdVrLa6C
hnKNcRt7oVw9IkheUAgSWoQWUQN77Kv1Sj6z3qZaeVZWrlWEMTuv7Qshj83GT4yLOXJpk0FXtW0Y
j35PJDCu4uC1VYcdTQ/hTNl0YatC0tPSZVbGivgrVgJb8GqVGcOXf308gMlVGqW+kz2X21DEH5oC
LNyOZ9lfb+FeRsufYUb3F9d2uo2OaN7dnGGs0N6EWbXusevi4/FaEqGuH7Jus3GInwn7MoMDw5Dm
H0ilCYv+5zI8WDzjFS6SiFoRIvzsBY3bqJleH7BtwJVQ+ySL7J8+CnOC6sSQe58tj/AzmOvl2u0E
IEyLnYT+7CzTnttihB+Tu2BQ9DDxnulAJRJHj7kptpZytUk0vqzsZRQy/iFJRvS1OWlU7IhutyW0
ixEg84eLzXYWtpDXKF5lotNKBQtc93v4yZQgfI+c2c6x5mthMsm2MgeKeKeWCW9KW8nHlrvPmdcn
0Ocg2XbqXWfoxCpYjtt8cBkx3EUeXUdlYN3OoeswKy7zEuqSKXiXenCLs7VA8VxlYp9fCgMjbHMU
c4BZi9wCGkoUwHN42x25NG2/lyg637sarpvG4o/NxaqbqlmmluXBhyGqH0lV/JpEgMwJjhU6XU0G
ZBz40Fso93pYdQKCEUF1nc9Owopll2LGH/gOKc4hXhR6d2zXl3tRP/BOW+nqJ1slqoznmMsSsLgC
DOkuntsRQH5ULRPDzL/TkCSPUiWL1dcj/W1Az6AfSqP9niRFS9RSWeynrxdgH98oJqyDPQAGEjDt
N4l3hO2uGvfKtrfLdSbDmiGmMrHIyqvTx+YMRDUV00D4WlN+A8PBjMFDE+gVXYqEexuLVoLNIqOg
OT9Dpm9WwsLwWUK+vOTm4oEmel2bpAcHrUONCNOqVNPQhOm3Dq8LaRCX6CY09phQ0eNMDc7rZqMG
f3Lf78a68BcKo2IeU4/azoxSWskOiykVCo/GVhuW6tsIogUiI5tCBqIVY9RWD21nhVAZgIJY07SF
KF1hhnGSQeQUlXxxtDcrhsGwULqQ+PVTlH0I25pb++SDC6oqG5L6H0M0YiFmbApZp5ymLufTfmon
YL3k27oZdLXVGMoIOQ4KOdM79EWUGs3tkiLdIvX1YFHeVOGXWb9SwWjfU83rpR6G+lkXtYDy8LN0
4GHKIw7p8qo9YRYCJXn2rm42bBZdQ+jZ+csqyJbQkYV8N9daBfxQYoVUkFnmrDKP1GDssewbJWFt
/0J3dgZUBSFAPLltk2E0E/GYZ37DpFRfON5wohyr9qlDsZXBVTFva8W8jMv0FmztUptfcMZptEgW
vtYlRUPS8M6O1tMCDmR2ffQw2FIKNjUGEJJUSM3jr9ldHsj4m80C5TNykMaXYcgo6eHLgyq8WVUF
ta4kv9hmYNCVH7/k1eH4hZhOZKoJ+j+tL53VelZNP3jNawRgOlmxAzriun4ya9L0+pTvMeD2L6Ax
sf7gSdJabDk8BvEKGKXehnke61QjtbtrsdTOgcOT6kRStXCfMjmFQceLEJNszaaDJytde6aNzMnL
+nAhhpSkHi+sy1/A3f6+1k8fN/fXOp1nmV85FbvscdG8Ns1WtjqYO2kCw1eNKu+r988ckgM07Y4V
PWLVGsJTV1BwZ7bgNJtS3PsrZR3kULuoR3fLFvZC3RBnxDjAm549bEpZnjWX9K/09Q0tPgFNHB4m
jhBHgDf8GBexOsReLwaJQeVMLd+qG3MdpLKt0esuz+hKQel4fXoVxsaeRj763kn/jyUJlX9VkDH/
ek2SMZgN4KlIiml3ttutQXVAXdBLqInlq9aXu9k4Ctk88b/suO+INMxUATUee7z7qbvlk0Jk/u73
hHcZP6adYAhQ95NTJ2KqbVVIY7Fj4JYBxDANrxKxSpUDRF+IalOZpx+rebAZ/5SPmkvviqzHvSIl
hj+7c4bkQlcnBWGPWRKYU5EmKVu2nI5MqS2Nq8GRgJplNgN9a7U/Q6FXWQrWF7KNZkPoKU4tyoL8
/4W4uYaIW+hyy724x2/fokawlSUfZazW8txOLSkcSr/6sSmHYpK/FEZQRiC5oqhcCwwAEJ5Ki0hE
KjobYCnnRgTWExC+N7pn/oIcwaR4ZH0kIETYhMSWcQ34tgKDussjXHT4z/DihyOsaXXQKTJkQDbI
1XQiRlvA3Tyz604XePfkxxM9xThVK74iTvv1mEsj6kgGR+Iu0a8tIsulL+wEzNnj5EuV0UyOHyrj
uKFxaffLIdR+64yKiKPfdrdMzMgwF6O2imT8UDeTKcZNlTy7PKzRw8EDUgTsR8zg/Ojy8CjGlij5
OtBQSGdsZjOkwglX+WpoLTpHitqre8+eo6xcPrDUaj7o3QcCr9uGzg5XeKzNTBc8aFQIrHp3yWlT
ywWW5WXJEneQDSF/hZVNGBA8vBdJ+oOo4Hkp6vgaCOmutF3bCD50GJrYm9tIf0TXwHgBiADgMo0x
1s00vax2laNWzKpoEAfeTXVUSks81HCNfxNrG3+ElXZVFgA+qAf3f1QJ5BZ3itZgcSSMVQyaAHLu
+zbskr0nct6Dk4EUTceb5XQ66UC58wXWE2XU7uNwBGm1IwMKs3xb4czoIvtA1eIYtP7yZnAw+FAU
qCQ3SeZLZuQS6QoR8uH1CroPqUGdxd3EVR5LXrllneN0onDRclvmlIq7H99Cn3CaatKC9oByc5hD
iCaa9TNMK/R1vd0oQhAhvhd2tvf7r3aAHwavVfYTS3IN10R760Le60/ZOri4y7pglF9sYD2/kH8T
FIQ0Y19VHwVCT3Yv2rW9g/XUYDCgbJoDzo3ARuFfWkeHFW8CGqNlp8MPxWXjmoGw2Sujw4fukTcW
Wckmzh6Hmq6bLvX48RsBC7RiJV/LjivGYJBV9kVYoMrZEkXLjR6dLKX8CEbXYVKFWr2L1eulk2OG
+xE4rSbqeIw+GMNNwXqIqNKZPh9omBbuqVj5cqnlaRFfjoOGoqEfa1CDbeac6ZkzqlCAG8aIiQ4Z
KLCRL467DXwMMO48GquBmG5KE93SDmnGELFf+nzvBFLUvtuL1gigK40rXs3CIbotlnQcIXjm7b+/
M0ZEcutNaYktMqo1BxpiZhD0pSCa4/0AqZ3uoRx071hIveTnRHxfH92HJcJ2OAhElgGotPpPD1mm
PEISyES7OcZ8Oa/0207kYQ6CswFK8Rao4CGaXtEtWjNETY3GC5MCpJ0PKUBlo6QWVjInygYCuzkR
1zy/t0E4LBFO+av/hC1FGQ0zNRoXT4qv6EQutCz/O2Ols27feyQvTqTX429lqMlSKuLAk3ZdmWJ9
+aeIwVe4o1h9p+v+6NWxG4Ct6lRBTPL5d04N7E+VhydoBdqj6VuRYon9FDxz22kr80E6ZfDBbsdl
GM9PqO9V6jMvaN/uyTViqBdL7HntwnHa46ZXLDu3Afb03WbkPmNB2PvT1tQMU/4Hj/Lg11nSnzVd
OlY+UQyvm1wDV81XfKUfcQ5Dt1RmqYhGtj9zcAs2DlhPUqly8tIebThFSurbol3/OUa3ftU0hVyO
Amcs81TcrtmY5pg8iJkqsOBMPu14svMkSWwPBX8Tk6rpgJDm1mQL+X8JyXELzVV08J+m6usj87pY
D5kkvHMHpwDOztsmm9C0D1gnJvGf2rHyhO8+dWr9fAjXUFQ3Ff0/feYPRyXEVEVbjdL96m4PKJLa
u8dNSk0pHqciw8kP+kGpWiJBZ1eEYnfSCizOYnRpYMm/NiyeLP+kU8QpPlS2LsuNWxA8pS7cia0X
P2Ef3tlUNaRLGerp5nKTOf9IMSLnX+v8LnPsylt4gEQQRGLdLYOTEPuho8XAEwUYo04ObJ63e10C
f3vdGfPPN6hR3W9aoWy7dtO2qfqM6ULjA1gjufvlleOodZ43uHvDZLRe1F9LbJ3uGb0ud+cL/tz5
2H2dq/IegZzmu3XsJ3fqMY5LdhvEUskvOTWZbi1asYD/7pzqL/bhh54cVrsBRx/LhZDp7IUxVske
8ECEnSuWR5juODJbs8zihvp1r0dd/+YnveLnxHOGDZiqOFLare8/E+FDMLJb2txO6nNj3aynJesV
x2F+CXh8x3+fMgLNthfH/CbJdcRGjVKj8xtCBKQwPs+IlmbW/vMb9+lLTUBLmL0ig4POK6qK3TIB
Xzh9fkmK/7jmu69qoMfXoFa1lBpqygbpCE1ZTNl1EnZEgIyiWCTCHZNUBh8qxDU7uGRrRReqvh0/
TbWULLgI8Cm3leA40qANRXiJJ2ChN6+akgwZ4MudMcbSfMUM6p4JQzucujzYcu7aTYOtrfSqcef4
NVmxYYyuMROjDL6hWLb3qFJQg3RtaGA/8c8J2IwhiWD+CtNevEUDEpUvmFJnN0Mh0AQWmu8y6Na0
3O6SSZN2LQTVBRJl1RhxkADbaX+AZnq/vNuMtqRZFtUmDE53HSWjqCUNDD4/HoNYi8XQYPbQF3zG
x1xdOoMAaNi5dENG9UC56RXpKi533ftDjptzprHPsE6BWG1n+EvkXjA9fFyDp5g9g8qk9vPv3Dol
CPMJU4LAtrt7yMCTrPxJnbVT8MH8/YwuwIK/arZTfd+wnkFfvV8Q5+k+XYJ+Z1F7PYLHrZ+Lhnd8
fnrZnFccupb+BjrKZGyDpC0QjkwfTCiO82/47P95eLsvg4GG19kJ/dhzgJ1BpUAL5hiLWqDPelmw
EfAFdUcO7HWWXuN9+2+T/RNbUAu2rrKszEUIII4X96AG11acK1JuqCHIls3Ew3DZEydU6+YbWCtE
oa/yhlrvslCqeF4SIpz0Km/Oav2VrUPfT2i9YcQZqJIbVJhr3NiWID+BOM5usDpCImJ4rsr9iMV8
5hoD3nI2yxLwazhA0GcEonhew7ZcN/bU1bZpmXQZPLdJrFRLf6MJrWzvlZI/4LIYjovdScRlIS4B
Dy+xkdjBNF2htPFCzYSTeg3KNsSQ2aefN4nbmZ0/P89VMw3xnDAAtnWPrnVTaEfxZD9H8gfy3zfZ
Tb1xQAshdIId9w/knnI7MTrkeXjj5ck0IEwQzfvbZsUFX1U9sycLQtkxHSGCq5O1n8hn05ux+w4i
CxoY35bPe+wxRJX2AXrpONQFwoJ+W0UNe+2tEvI++qWvimYP45mXqOfoF/5WZF8s8u/wgN/x4P9Z
A9uN5K2xG4bvjlgUD5kKu+8ipdmMLk5MSsDTh/f0D4EWBMU//uWxw0U7VlhHfLJufte1KGCC+cYf
5mbyHdUq6TZlaRdwdzuUv4GnHNr04Najd6HDHqp4Kyfbc6aQtG/lyqKKah+asxd7qjjDdKfVkQVZ
G7gAQBb1csXMCQ9wAmVBBYw5eHq3o1DvfD51aqQSLTWI4vxbzjvutjvSNxl3zxbmuUqduljqBkcb
Y1oTxVZT+z+r164vmdwMFgxQC+/q/uLGTtsv8ccRfNwFHQr0phc7QwcJrxEgEHyF//KuBnr185sK
p4tI3ns8n6WtshiiJWOa0pWFjK+jAfhXv0Tp90YEg7useF2XYUDyQs5GBhGpHTZmuOYSRtwZBGeV
EEHRnrf9e1Jc8YyyGXLgHZsDnFP1xYh5rCYR7UBEhUgV8Xk1JSWJPG6IkT6NftV6fFXe4qanVWDL
JqngHvOstSRiNzxMkA0SIwxi6bNJhR6KCFCDOYN9COnJRUc1R+RszAMFL+UDzgkO64uMu+0glM7g
Egmqi5qGfJX+DWCLR1mobBS6xsL45hEyoajJDjMiWlS0/040gwR3eVmGrY+AlP/OWW6m3BNrKcyY
sZSgbR3HM3kglc3TVoeVKf65aDXmzZHog1giJKPxS7HMcMm7nKEbMYGwMVTke5f5A2Li2h/QaeZL
PbqQoyZbRMcKkqyal062n1eEqkFBL2Z2CddztwCwk/YcT8KD9Al/ibr2U8FmjrcP5BpxteNKot0V
pX64BEomJldRzN+zcBAtPr3hzAx511zoGtcmo0AIKliHKPGaOg2TsCe/BjWZpMrNeneH0TnqFAAg
jzwgA6gRySZ8zNnDeDRzPAFSpcok9JWDmMRE5jlfuaT8v7hGCX92jVEmKVMGZoQ7SvfIpZRglr8s
pMTEUnYib0q/LJSuthGKSUgyhcVVDYgwof7Z+QtPdIpJNpwSHvs1I/LtwVBVryglWqkXcyfzuHRu
xnEBotjoPDBsiIwWS5N4nNjKBVFln6Yfuc+EwR9ewQPJHPCepejPifrFNrvDSiBqU5k3ozGSIsfM
FD8UAdoeU8iJES4dHxFdK5/QF2rrzwt5MXwoMqVMndoHgi+sUcIRuBsUYEHw1lWc0Rq6T8ZIIetU
UIGOo2NbtsIokH3f2xo4lt1F5JrrOlo2xWppnQaOjNu8yzpUIl8JbuuTH+YN+MpB/Z954hfDl051
b+FzpG0w8zOKtPxegE8pcKHt59k/CstO/jWX9x5kxnSFi75qEXSRXGayOaVFLgZISOZrtJcS9hXV
QefsIqAq/F7ce+yUWikgHPZuW4ISNaw7bbXS6eZU3qtYwMCkIME/trRLgv47706Rw6bFWEY+xyB8
FdwpRMYjYtCmL2Ny3bWiTobx+MleE+XgD2DuDasba7AJ79DYH7ItASqWIlj+Vt7j2W2apipsiBZY
9zMqq6fyBN9X0OS6chnmFdW3qBzFjsbwDlDD129UzAWdSX1Lzo/Bj+7Zjr8bexvLcw9ju92ODTqp
u6Kc/iVqLsN5ghLXQ/JqP0cjzkYRkR2YjTz1uSeqQ7P/ySxS/BMjuoko4NgMDlD1f91mDeR3I2Kn
XM0tU4Cv2zeqXcaf6qaVDRvePV5dAJY3tPHJ/1Wt2gXF8xGmz+2H/EPnZLXFLtc9U5KU+lsNeOvD
f+pSE7zLGCoQXpISrAz0U/52HzYSeSDcUKozOHEJFS1YzhiviXZ5NZNS54mTj2QadrYTnOUZL+3s
eAmBa772A0rfWJGcXbC6kb0oKb+2sMs+3Fij0gctKu/bJ3vVvVt0iLbV35o1DA8f0qhbKbQ1oYDY
MGVNY1YXQxWnV6pzABzcS/9f0pHPWILQJwNf40npsoX4CcAI+jjwSa+q4thkFbUKl1ThwSQkkVnX
m+EwW91em7iMfznVc9z/ibgmz2XehiWNsu7PsWeJ8/rqytI6SikPkdBcsSKcN+38U1mrXRalTjsW
QEGsQZ5XfDQbyEOTIWZAKNK7baFeDwyjxdQm++I7MGsOvuqpxeD1iuQvKD854405MRCDhtt7cnFd
Yv5jWrAK2tMywj51cYuKrpOkvo9szZ3/UIZ+n+juHM5Fp5cLKi/sSw9Cm2d3IdDjSUybEqG6xZ+p
gcFcVyIpjAmJ7e3luSVwHp8v3l03RZu+nra/RUpZUPXCCdOalHVy8QmqwDEm6qdyBqeUAqdV5jcr
VbL4scQ7DTptz4SONky6egMO6NNzzpkCtiJoN4ChBuJ3G2yIaB5zHBQ7uzuYSjUlYy7aOCcM5Ggt
1tD/quNsUlp6z0tIF0CGFTPp+ADTzhlnSPrDhdmPVp7p2rY7Tyvujn8TnAL/bG9iZUHIDan9ys+Y
452AlpkE1GQSBcsODuB0sBLWsw5bGz3o8fsVH3Zy8PXbVvWZOGaBZOmy9QSIE+UVbgJDFreRSG/y
g3K7nyuLbQnKjwn8aNSMPtHmT5gWYYocAq0D5TUZUZgqbVUpsbxJ/XqcHv4iitkoY/7vZaqdFgqf
Wq84IHFlSUADADTGB7tymfsfwpCvrRn7jh6H7m7RuuKzaYDME1ADnA5EN/nVDb4e+lPwAggy7Nv8
tpu0/uBeMpUA6huh1ETEn4zZEIcfh6qQOoxCL3EdLWMtfdsFUR+GofWDvECuc7KB0zSvxUBtV4O/
0vqdWJ7UYEGPnANyJVd5qYBsD76Wepx/lBDfBlCPVDiDKngj2zvYnW8/Cz5mfQxY6nDojb95nkvT
1bgF7bXF12eKFPQCgD77Ujb92cAMq5gQIilsT9TYaJqZwwY1D1q3BeCMHlgCle914RFc2SZEr1YD
z1c9fXvNorWPC/Ca6dOb50yJ3E/U3kN073Ikxj9LM+7r6g92HHxQGlFfIvbwaZPOVWM3HuWM4Fd2
nMMjKPKQyIBFYhXLcheJ08LJ4izIe29OeSwz7G4xKD2J06Z59NfFC7WXm6IY5FrgPl0YvIBGryYw
hdxyq5oeBniKNoBwE9MVcqNR0CClygNZP3yqb2iv1oHM8sMokarnJezM/hWeEHhFtYfbCEmsztID
pb6M1mDt++tCPbV7K7wtlWcjS6GpeSDzYJzRqEBzTijnreyRv72sz93keHxwIG5qSvmvdXfdohfR
B+Z4RvG3glDl+FTOj+8droNaLCgwgDA22mljR/qiWis8TzVYVubEM6Z0qaqppOfssJicDspXj+Lj
o3mK9c5hu9k5E0NK/eDSM5CBfXCvnGf0imB/8GGXIFHt21C9DJO4pDscivcF0CTut8AQnFlUwjsA
v2ZG4CQPCAarrWbhsc7/i90xykxiuXmUGTRMKWEj+jdpWDP77N8PQyJplMYnulhAnt9N2q5X/B4o
MhYpWU908Cujn561vVEM35kFISy7xtc5BOAa19NqUbeycH1U79GedsAeiVOyHvpvwmiJFgdfDnWg
ykXDHV0wD9RVw8GbDmEI7ZRPV3PNBTWLhYBD3dOL/N+4YlmYztijg2gUMivA5DpzH/OUa5PiDHyo
pEsG+QsbcLqexOPhx9Y+AJtI9TVVQqumHB8hq7ykOg/+Z90r4kgUtKWtfKf4Kih3qpoQLASbOiOc
V1wb203OpAVP4wZW5YIL3qNx7qsqgptuvoEnchqHG6XRupTBxnkm01X3Ehl3fN4L8xeP633X18sB
O5xsNOTg0noq8ZkOb/P5TPr06s4lULWFlrN1OM1ADGAAXiVLACuPHe9cBCfZUf5kb7L3JnwvZPM5
2lspNK9cS6BZfdQKfwHa6KkQGCTr2odm79LGRXl2rdxOy1n8FILZ6Xg1cxF29oVBJRNkf17lpGUe
xJgLJyrkgDhOYmNJRJs6LJQmgfXlgWLTEIeoZSZhRy1V7HP8DqsZfJ29G5gpCGqcrkkYgT3IoCcK
RJZXlzHFPttamefbHTkzISzNnLf8jZNb1pWN6f9MMWr1I6QKyBzUvSZsohatgdoub6wz8ORDf9kp
s3IsSvkHR9o7qcN9I14v5iEIOr3QQxiPcFJgOTJRBgFJMCKBswqySvF9heTaGWQKiHHM8fZie5dL
HSmxq5jUDXcuMsNcnR6qDbiAi7n/21fr5PWakml+onfrjj6q+xOLoCk/e9TV2D/fVuW0lX33vknp
MMHhB+sYXkH9IB+OcY62tgkru7W2hSROBe2aOAdp1LtzgQ4eAvCXsouLrrBd4K3dYRY5jyozblHO
AlvSAYA67HpS17OyfSVZgF0A9JymFBIkjL0GbOUdjuKUzh+LgCjZ2ds74afDlUbDAztangV8DHcJ
/PSPCfe8Pc+YhkYkolHn8hMCBQZ8Q7XTzDi7TuIRjmtcJXQoeSk8pgE3tOaFuFol38FJirNmtkt2
ipgvmbPftGHAPKFaTyuL4W4uu+he7RHGceG5AGQ06ysN5NBBg3FZJHyAtIpzh3gjvg9gOiOgpUIL
aL9RU2MkWyLx35k45ktbT5/ufDbgOI2lYqRV8FK6fGBZ32sTNWJNSKKnod6h3cRKQNg1Y7CZRuoB
GFPF1v15rmPfB+CYLLFnO7c7dq3vcVrhmGXlVUyM6vDFkMbpaSlO5bomTDjvvODBXjIstk/vALLX
Lrdw49XW/m7EYSOZ8pRwprRmjL9eEyrvOdNVe5NpE2VLmJIetCrcdVAEl+IRMmMalOT52d0I2sYH
l2n0OST/dngZxeNHrgSaWdGk1jcohWcwnYAYET1Lc8Zi7Ux8RCcZckPnRLSPxzK6m5VCqJrh8Es3
BlDwez+wpSaYwyoKjW35tcM7CrM8rHb+g/+NozaOpvKrqdVpoK4Wc3abkX2a9rO3WS5+d8GenzaS
r1f++gTS1/xWPnKfU9a1Gxy0QYgvtbUZNFBy/iuaHsywPPNaCsvEriYtBnq5r2Gi9iLOpgYaf6FQ
2zUEKRmzOmKLaFODX6PS9UpPufqtJYToA6MH1H16LEhVq/aK+2SPcObaBlWWOIYHAdiWo855NreS
D8IndEyZx1WYme1Qkgt3CUT92aVYTiVzOYt8lEn0QBu+gj2o5qRUVImzCzvGNbJlv+8lEr6DLx5E
ddO6AH0/UB/4oEy4inxTamCb4HsWYvXHlVux/2Omk4gZSF9z6q/ZbCh9WWI/6WvGDXm+kC938/1D
8I/+CUYQb/xj5m7c6dOzbXABKUSc0qO9KrRG894OWsusri/FD17NKEG3eVBafqIb9lBPkVokNx1J
rgF2J6zery6pFsbYK/+cYgdtnftla++IX7e4IwWc2dZbaQTwyl+NTK1qtTdPwWe3mvZWpUVR5eTs
GRg6axYXY6dga1cY7r26HYgmcmAlfV5pQM9brT5XCw3pVM6v/kMVSeVbJStzpgLrxJLhIISKOdgF
o0lPjD1q4DifcrmYs3OMCi6aTaD46C26PeyBka0WPFVRHNogtfcf8xyBRJwQCuAL8kN1LK+WNP7p
G687mfMvWGqJVj85gYAZCJm3yRBGb0Pmj2v6su/BsIv3+F9DBoUWv3LU3bKOndBjTH91SXBocILt
lxsVOEPsYGto5zjLEFSe6BsMNY6R1rrVW8+USTNpsLTx93oieNo6nK1WWwY5gmd63fq8kuBTU8oX
foXpkRHMgXnijFcsRCmL8+B32dSlbp3Dx8dy9d5nEcz4YUe1P5j87ZyOuBAI1obGhlDGEJbsNWTh
LeeQe11aVoEGPtqxyKuD36eF6gbKP9TVzHre99LmjjG11udaLpZqgbvPZtasLUlMhI7dA8FBRq6/
uynjMj9PMuX5S5mtXwSAjt0HES4G6QRzlpHFRMN2ijK6BZAOPJ3MOAEdSk0sYK3GGrAtnX05qIVB
yUBJnM5aj/67sQaVArLx2oVX04u1d/NpjtrAWwfrUfIFR/eUSNbPod98WwqawvonxgmPf05d79jc
+RW4pUsKCxQv2ja/4ShUJScCZhf12KpYGJckpfQyJk+mhGThOFQI3y94NDTN7QwWuq/RYRz8Fk2n
dAvn65HhRXhERM9tuhHYjxGJN+7I1JzR2nQ/ab+ZOnVkgnEuVMYVXPRYlFAIGpsDnViAXHt8w4Q0
wztblFeR6NqmT2xQH9ay6fdEaVROB9YAuXE9gMVkLgsc4UUQDl2kmoAXE1jHuSCJ5KBInowVuvMF
KT1X/uTyjjgBk62N7vrJtDBJYLLR9N84bPUOKWilXwK3INi1G87VWTsPCfMx2AJrvHnUYF4rxHnz
KyR8gthz7SJGZV9O2NV+FHTvnUW0Cyo5QGWN40JSHxKCS+3yiOS8QFLQaS3GwqtIF376WBvmUXOe
Sj3B0J+4+chloxCLHlecxdvufo0YAZKYLjVXwLVJVwkKjWlibpkO6Fwk/ubdnvQKJwzA07ppM8wg
zP7LXFm3Y++Y+iwn7UzMSz7JdtK28t8aGTcIiKwZ0+HniR6D2kHCxBa551pAceHMMomYsXCpb/OS
oSoQS7P9CUlMFUeHS+y9zyd5ic0gHVV9Y0qI7RSU9KWw/ELTgl/T45Jb4Th9Sh+1a9mJdLvAJ+yK
271R8rU009ofK26tO9N7fdPDZFQ7jpnmhEp+3vJ/R80FVTOuB34u9A1bZ6tKTBshcQjto4ydP1ZT
Hkitehyq4aO1AS+Ttkf2wjXMMkZuZjSLLsfNuUA2v3+YPi+1rVAWGLAdDN8QtTwoyxzDd8h6Pv2S
NRcWPI3372kLsnSejyMg9J/9nI2FkHCc1+u4H9E9CrdLHIkxLVa4El9lGA6XnnpEqErQcoO0+EMf
giDH6O+tBGfSEq5+vW9E2ooqYwHBII/OxGB0pM34TemRLLI3UUx3/tXAsmATm3e6BUgX7THKHmB0
JtPmSe/Rtyna0yTKwnGECeT3Ro7AQZyg5HO5Eo0G+JtBf2akEUpSzEwxCPyiVdOfnT5vHv5OpWDE
6UI554GdZvz4aO4jwANBBdm3RPH5eaIHyYRTl1/61YR5qVFN91VprrkWpKHad4Q9nfTaTs93C+Jc
IlHvsSJPhh9kcofLFs0d42sgm4aVjaVfpqIjQDklvMilYrNojfrfWlqxtmODacxNefJEK/NO1wz2
sACy+IAds6ZVyNU8rQCK36L34L0rCh4zTeliaiVfFJPCcxYPNmdOxB93R1xHjiqX+VN2Ludp6Uw7
14GFuBUptBrNFZUTVEQ+8nltl54TxYZIYP5IqnCpiIhwCmVuqTrNaAbggCgewCNQ5zUxcax1Toha
3I5zyZGndhdEZNGFz71+JIzhSpSK3Kg3QYwhp9uZ6s7LrkbvzDQkaWgKryNe2dFHP1Xi8uAK/7Mv
N+U2uMnZJBHpmvVFcaVmL/ZFiFnVYxX4Gjd83wwRW238ZymLle/8YA8cHiAmyk/jXxcSjjIJV/Rd
lycmQe+1fNN0U7WSBEJ/Sujp4Pp6LOF4FrFOV7GzODaB1oPc53dVmS+mJa1oroKA0aRQjFquLTL9
UYEvBL3HpFoYEScXB08nOs4zTJxyBeELyGchiBRY4DPl7Zv3+Z57cc5Jfz+l5EZxcxG8tmi71NZn
BxyCSUvDkZBeiWFN4T0VxUc6c2YCvDnO2+AeG9cxS495mvzJ94k6v0f2lX9uTgc4X9cRQPPfaDCq
Kn9GmaHIEGaivHa1xfwA+QdjWKdk2hcCw2zOoSKAwvecljFxyuUXMmmHlH6edMCQRSL8x4zPRkSh
6b/p0Ja9Cciwco3FXKNRbGNf08rQ3gPzAL8DC2nEktJmIRqEqq2Tl1DwbH03YEc42BYqdu6qOebx
mJ5d2uGQAGWiMYOC163D/R819JLFVSAu4HALFiRfHrUMQm9BU9cSA2ChVffX7oBrhH+0iIG4hrmT
3D2fx0ovYL1XRLmVswOTGJV2Eov1yp4KOdgqGpy5dJ0UhxmBbjhxxzsysb4mzSD5++XYlfz5u9kW
9iU3bW5VXu6RigePmjAbG5KjjHesAsq+gSrO68s8YXHZ2CNMICduZjNko0Bm4PxfJdXhZx7V/KHe
BS6YezDUaqAbF+64x11V83Y3OAyofTEaf7YhV4P+gJMmL1blsjnyN0fP1ZVNZJlpQeQmMBZ13/r5
sO8dWNuhwaxNunRnzUgR/2ZbPVoo48zMBviD7oVOF3xkZh1rr7ohWIV3IKsMERHHZKYWOeVvZDJ6
f+aYlij4KOg0qQv5o9Ws2rutRwQZwQ/fU6uU/UpUz1Oui4ck8hG3wTuS9bGWqwMYI/nFZQqRFL5Y
FHsEVh/MOfnHglbv1PFrb/lFcvZIxdN7F4kCD5ktkkaqFXQH+hJvczuIeBlu98mTHJlpR3qIIQfn
GndJwtvNlAc4V7oIKJ7Sg3ukSw67v+ipFeM4jIciB3Q3hcf2DqGe87hZCq7F+GwFoGnWmz+3+0sR
ox4QXqAjrvwyuUmVPkbRONizmFACQ5z9J1MmW/FxyvKSuGpgsubftoLH5ig99Sd8rVbDUWEi3YZw
3Pm6sfqDT+1grTMEBW4iyXwJeEESjEkk7uGSg2+KcTYuE9LK8TZy8c3wXSVUN42dL2JKHGG9r5t/
X4KqtHzT/Qu04dredeAkOZVe2rAf5ngF0ycKwDyaXKTyDuWmqwS9mvV/EvWR62PsrYtvbkdKHan/
XAoExVwlNUBsmI8CuFi5gVb0Jp69Npd5WpZjT1qNxd1TSVu2Ku3tEcueijsaCSKGFoIuRlpUAJSB
yRcAMobtmVTwh01TxGniiXZUNqFNRK8sXfa3DCrCqSP9f8U39PDJuUO56fbjGxoGW3uhOPYshZtQ
wQnxbiZo3PahyqyMM5Mc8Z/v7an/IeRURpy1ODGmdMXm++dymE6o4GTeMCyRZYrBmeFkv8ksNv50
bbILLWUsgUfWEZPQ2Sz/B1O3fRxFamRsvW8p3romN1sGPWI13fI7PN3G/Lop34PNWTxOPsqW4fyj
zw5px6mPXe9nkCT45kQN6vt01unz8rBe2re1dnUgSy6lxG5M5CHZtqGKpFkdoy2eqV4CFaA6MF4u
NUbHImPJw2owDh+6eAdxM/E2bXPygUZu/PUjLwOBi3ET/fQDXrHQ718GzsGr4JmuIdO4xqSmLAiu
CC3Vy8f+aszK6L+3oboELjsODX5tyV/zG2coWiT8Cruq1tinq77MjzdRZIqUi210m0YF/prfCVO8
/oCkJzpHn5xa0JK4HwwdP7oV/ltdudr7+pe7JjXfPhTjw8/oM64A+H5+ZVjbtT70SgtpldTdqgGa
Vyo6IDpruOkLGX93i8DdTY6qRSPFgF9fMAD4srwc2Vg8TU6DojJ5IQG9XKDJiC6xdc9R0ppdo2zq
J9MUqNiIqhVZzY6ybRLWTlp48l267CkQEyTkeDNGXwTEOj2M+zje50huEbLfrFnyoaRdrm0Q4P6/
/82KJwO33VwkSWuSd3YRih/+uEYupZN+jD31CPm4A8JmXSp7Wv34kkz1ddoaZY/uJqcylfANOE48
FpDFVhBSbeNTLXzUosl7DGK5mwZSMCUYGi6WCvN6gPlbHJTRF+vy8B20UcDmzWWTzBxQQd3wOGUJ
I4ufXSAmqTMWbu+7KJATsBvx0/i2f0gxQl7H0pUMoEVRALbVtdtZbfL5+eCJ16J1qpB+0ZrtvU9i
vVUxjaXF4oN2Cw3XXWpfFw+WbUcPxAL+9838NkdLWIpNTDUERh9PVDdUHicgWRoNtLFBkfAiuElr
/qAJBUuI3Y4hYwjJg3KTQyqyB5qRnyG4TF1/fjcrFQmG4zzJW8TrryHMMSDRiZXDRQ+5IafC6sHt
TNktlSvF6n4ucuMq7vgW4fU4t/8G8mLI4gab0IxX94W6bw5h1/hIKjRsmYe/+C6c+2sKRL7rR8cM
lmUValOSYf26gfpE1ItVxAxVIImVVNnYoMZbPLph5hH1BlmgtbmTaX/yKjNE+ZAVIAw/8FSv4+Sd
JLoREvynlfnl+zvjjQv0lVnyc9AgnUbaz2Mkj2f/VfLeeg786wfzkYJpgiK8tkpG4cdPVDJwdODo
2oiO7BItanBWhSoOFrbd0ncd3zTb4fs9CAEGWykxsc718rLyhMwj+QcGDjXq3o3r+CtDgbGwIxCy
VdDFNuf5poUAXWW+hRhdofHzFPUKjzOnl3QIPvVP+IL0tg5beRCVFK8VvGUtfJvJEryp7/vxX6cK
fRyQW66w5xx/ZG1XiR1zVybUEgh+FHZDDVtMtd+w0YYhxPdN5wWY8QWN01eU/CTYb4oFah0S8U92
lktN4fBfLsnMzlP68ICdRl1P/+Ri56jriKf28a2MuAJddkAdfZpt6kmmHwbb42VEMU7Lnb6oDKK0
VTmdwuSmNS/rRdJ0iOTR4IKvTKJU7ftP9oaoYR2+Eintv1T5r4cdc8Q24P0qNdkjvYxrIMCeFjqC
k/1W40JYJR3GSLTYzCK7vaF9JbzYCCK8RKuIwcicAneaoh/EMhuudv29BDPdMAde40Emalk4QIL+
zU7hGIXaDdWrfSW5sBUkU+DMhBjViN12GiWtLMW5zgX4l7UhJmtn3dKiPDb0pOBQ+iPNIZtp49v9
3KZCyzVRL6yKGh+XWgFycJEAWYudvKmqQ7AGztw/g0i6fIyVrw//nDSlEbBblynHWlkeDrqegLwE
OABROB7l2F+IEhVGAw+fCmwNcUes0JcfeexVh5sBRqAsk0/pdW+iVF+EmJZifly48wY7nf5XgcHs
KaM5yufBz2wxezsf5sPfvqj10zDL8Z11KH1pc/nR5u79SdQrgVXYX09rYPVsnidaZyMVsH1ippXs
Z0pMH77xc/JwNkDIQmPlPsnBHYGtyg0YgZvBtF3eoM/S2sfph87Syz/ynkYFb96nOr5oyaL1l8Yp
551nKeMOA0TSKJzNyC4bie6bl+Fq/EYs6iog9V8fbro24wUunjjZyKOnD4A5AJ82pDaOptcfUgoG
hHw5H4RQqsZ4uNhz7OOGwsgUzVKT6ZGLwIMODD7ewcvBIlLpeAnCFbbM94OPA29XbEXibf0J/OaZ
1h0u+SZZHjdqfW+Zyif8L++zZt6KffIVyGx3p1ZNB5qE2LKKnCBmHoE81pkwXo1vVp0/9ZjmG+cZ
tkyKPAqDuGYpj4mmEqr22voy1+6PuU7N0UyD620tzwSDKONVUAgkCg3AzDFe3KVNGugCmN0Msg9e
7AvoKy01cFyq0snUQiOYOuIUfoRZNd2lP6VlGBHUiRgmah+Q1Pe1nFE9xzMiY2k8rfiozDoj0Hox
UMtZld2Ou246Dib3xUUMpMmfVpGC3B1YHkWRoDsmHrWQl6KLlEZ+2yx/jdjpRUy/QllXOEA2AVjE
8nsvk40nja5VA+9SSDeC2gde1p/5Pn9XXLm5hitwfAIX3xBLiM2fCnhkwgve4QOeTyvRw2q2FixJ
1danmLKWKmdOGbYFgfugjBQRTv4yZdNam0PAz9kEJ1vkjooT5qUZzPW70bOsQ4K5Yd4AB0+JX4dQ
PpZ5/ZozoOWOhfrTIbsv0BR48jQLu4VAx8vNVwNiIlbvwCMNv+bDWb2Qow81+8xMesBpUSexvzdM
hJR55kPIH5hMC9MsUU/bFmJTGUrmowu/tpMklFAh63au1XNw87uKWpHtMPJkUdGdruUa0QCqAp1Z
R/Sj3wIyMysOLP9lw9n3/paSzxgCXiTUGw35Ws604G6vFiZLhIteU1vkDp2akMiezPVp1zaijMba
eIKtpot7GbE1ITh6N2izprEnaj0X0J5M606Ml18by+HR+WQPvhu6cNdT53muNrfW6Xjaydde6Lhm
G5HzhH8ubKzYRrj0fsN7DtPU4Hfx2V303rwCuiz20+3SlotGwZ2TOIMIg2xnCdSOXwMigaQfJmtK
FT6TD0RNXHEPtu6v+Udpn4+b7scC16tkpHOlgPnwpH2MphtOUbL0f6c1ug5O4+NW6ijOKvWf7nLf
8vtz21rJfY8WsegHsquxLMHW3izUYb87OMynPwqcsy3qxWkEidKCT2PURdvluv8aXChFC3X6JXN1
g5TKVy3SDIBr99Jsp/50TmSG+9DoPHHDa9FSUHPHsrMvxVBJNSDrxC93x5U5jBRkWwFBD6GoJ2kf
QdmqXzyU0YGtt1Sof0NnSgDQj5FB6/wXXO02vcuQbADfktDXcJeaMSj1R61frztSyUTknbd2DXxG
rjQ6CyXML5oYYjzaPQeG0od73cllgjOiGLCpLoTtv5cpLo/rPp/MFCvmIIENWLIc7j/n83epEgG/
8x8ykl1ZMOXxPzC2XLGyZgKnsqqbrF0zVgMCuFhF2Ydv2z/pSwcfybvVXY4xbpqt1UQY9ua6+VHS
5YGzxcRB67ErN5JRZ5wzAmswUoy6Tt6cHA5z+jc8yqaFJqm2tCEOUiWE0h6yeUL5EsmfHN+mUQlM
sKZv3PVdLZ2ypPmUEwO97GPjC0XTJJT6zUd1MPqQLh+RpQB1c7OGAyPTCWjRLIGrqxIi8g50A+Bw
6i13zDnRk75Tf7FzVc6AkToRuRxAR5GTUvlhfQXyLQfLc4ao/gH4ZOAzyLwp3bKuvTNVguOq6HdV
Wcd8gcTQ+5WogUzRGTIFzp88wgMO2OX3G7jQPXzW74rGhvpjuYG3sNpUP0JTU56Xb2WTjOI3kWWX
ivHjDiHu8n7F2L0OPGGp2eWu70XpT139Dt9ioxOSNwbyF4dhml7BXTEMSjGAnbyYfzjo5CYOy6Sn
jHGs1Hz/k+aASRNEuFRh3lGvuONPtq1AzLUvk/xQHSHunFpH830QJR2W/uJ5gr02Dfq251nQEfJZ
WdG7jXIZrdJh0LxHL4wGvy8c58jFsbBUyJSIvfIPqGMG1JoWRIBWcxqdt2cNufNrWuj0Zk0IR/Wo
B/fuh2/iGhbNyH8OCsKQuoqFbu2s2d+N5k1DHc0apLTr9Zwm/AGE3S/cbl+Nz7itUglBEUZQNXW2
CGeJQxXLUAJ7M5YeZWw2sU+jO0iDYZ6+DluF3zN7eucFJyMqxEkpwDQ9CftRvRoyguK2YAth6G0v
VCaVmceFbSwNv49DH+TJ2pkVR8JIWR4rPxf9S9GcpTz1qM03No1brcMI2iVx3mF5FqgRhZpsAvPH
joVkDNh5baDtr9IAxHLj51md+xky53bsfUxkUxU4QJdCOjYG5OBFTMgtrQpGSGM6P7jEsFWsHwoO
qerd8zff4ZjXqDRklNuC1CtoUTC9UdCIt60CMS8Rgx3b6HxKgCa2DfTK974BbeNoiKpuMlmuzEUm
Xdm+fQLeuvIukJGw9eS+dEViyaBZ28DuGa97aFHJCah0iCC3AL9BVyO3SFyCWzwOpasyf6q1QJKF
FlnW3sMy9KjLirk54iR3o9qUiEY2c62MoK7GNzfkktzVayf8M8OCHQ/LA8XYXns64wg8KfAcMsl1
bDnNpnoSwD7TjD/bqK1MTrt8oEL03SmzC5MXyKJ/btMD7eKfLogwGUnWA8mJBFp5j2wGV6TQ1fZe
bSYw14vsjsj5jQZYAMUceS/OhjMBxSLRTSbSChCz04vqc6VliikpfhKDBAbhNWFZf4kSEL9MgnBY
SZzBL6+16S0K/lWJ08MzEg5YR8RdvWFeColx9wPYx/sfzVtJ5rAcnV3kdOco5gsTwZIZa9BqOfDK
0MLs12HNJW//D1qOioOHSMyyQXq+Rpc+/0gxNs/7MGW1k6vP2OTeYvohTILtSgZSuvD0QsKk78vm
SKxtESVHVbDWWMocK8AqTOWyEBidQHAxdUMFG//2f1FqmXzNhTdnLPBth3RBIgNGY5HMzSKy89dn
SlHA/DItSyVTD9DPBo7Sx0SH1+I1tRooaT/NAL6dUXD9UfE7HCxRrrn2LRSg3541YZklkFECabiV
aWpPbgPeReE0Tw8pdLnDlWa+3cRbLuyF7XK6gb+bMevlRNHMl90p0YXR+VInptPzol0RR6s4uxms
snjppUCIlaiOb6UgCvE9kZSTbgMIkMxFvdTQtBvbQBqmMJrImFPkz/ilftQZRnj68yXt7c/KjJWm
PLkBUQn5pYcApvn3G2iu7pV9vum63/ircYK8Dhtwf5pRUEkgJkk5zO7v4iHDr4hQU7fOUbKTXcH1
KlHfhO4rPOR7k2O6gUms7RZ3vRvDbpm5ApDVazsPAyjlfHdBVUmbALITRFDtFa2RPR+oqT7YeNm5
rQ56NQva56JcvelQL1XMC/YinjFKteNQzSD8H/YaZzenj9/Ps56jwprVZPjqXTJjcvslt/DKoy72
PE5maPm5TEvkByae2+InLJ1JwspgY2S20siRvHvVdXl34d7RVwTYXOxFxVJlWZtqA55fCTgrUT2G
FSvrQwH8vO8chRjkxPC45U5oLxjymXblvK+DBRUSs7Yin0AfzHghtGTn4P/kYopwglRTVUbGL8a5
RyTXxEXQnUHlucpVqHV9C2i9MVdFXQlwE2usjtJIUxSuvURVQoN2IMQN+Go2/r5vAGX3G9z0dxaY
0y4CKsGCSxlUB8srm7eGIn31wgXek3WtYm+4Xybn4sgOdgg/p5pLH9Rqu6ik5l2BcQm2qZVlltlo
BtTk5TaqrzmCrb1lIxfE6z0trdzTobYp81y8/RR301EVEREyfB4rzwqFtHDHxFSo5Utx5Hr+J7EE
6zzcNqDbJBbHYg4/TTzKOJUAHOKsbAxEVUTtdjnN2Yv6wIy58hYctrr8k5BFymZTyaOpMmCZhmcd
FWs6N+BBWG7bPfC3L4xawsr5IZFgmvXglI7W2fE1dgqiE5tTpeHjf46jrjtA+8FJYFv9SpdC0t27
0xbaO1qmq14naHAhT+nAC9UwF6ipFtss9rXSVtxe58Lzb33mA7JVv8CMMrkydBIDVmP6/0nYD2mY
njVM9O/p/f/F0Kzyb+fTRjwVU92WBq+Ipg1Y5JuMWxDIKDIzoq+dXOuWPW5MFw8xlnCePTUw2qq7
amWw8yYEwG++5AcrF1xkarUHewyjT0DaJa3U7W73o2N2+Df4Gz06R0Z9dix/Vuu7tvnahEkWEJax
vs5AWDhbMjGUgjBT/umo1PXXI3BHWxyglBaQe5AFx5cASWBias9QN+BkJrCwQEoY6JqpQqVieOpA
8Ib0enDxCJHYXYjacbnL8+g7iAHhloDqHF0cvG9tyDa8Qvv9AE/rFm73l9Y0hMmEosvMcAT0Eiwk
Ew4zrIIIBkWYsA+tOHwhK07NMsQ3nKfldz+Okjr5uwiQzb8Urzuy16k5cbBxDZYh0j9xMekvqeda
Ovz9+Lzr5KCddcthjt5SK6stXGcZxHhtUteTKSKlDzacfCMQG4mJPHyuVqqK6iDqyRtmooPl/kLp
OzrJLgyGWGxg5wxCqyl3dBgcJ98cMRHl4nI84IoLfsv0R70k/ttpvTOiytBfeC2cZXaZIcloGzsE
zWTGp8lNLJ5s9+KJs8qvpgcUPZQCUpLrfG4KGn0yWWo8t02KDdJIqxzBVXaipGIhXULX4WzWlpuu
KOFuGjjQziQS9Vg4lcwQ33pj9CbuMK89vHM+RB6kr+avboKthWyLL81Idnppbfp2BsD1eQbplHMW
P7H18pgzeL2/4ojhWL+Fpm8g66A61zqRYRMdcbxAKwuXGrcld316E41kiKU0S+TuQhkha3QF+ORw
ssuVp/s59IlX2qlpnu+aERcksLWCjY5d/g+DEoQH7IaAx7jp/UP8FVJB76zO9BOrbM1fbXjYodFZ
Fjk/yRII8F4Y5FvuZ9vHvSShsFgQYLFjIP/zquSH+QxXRtfhWVu5aI4Yb5LJ06+cvmC0EHYLxDv7
sZ3D7wJSqX7loksFfQCGMH4uEX8Um+fNaccAtTcck/k3IgM5ep7Xw+3I27+p/eQ9cKANWS8/LaJd
a9NKGmtwGjNr3b9ji1M9scdohPcIAhH4fiCSeFp+pilPFvRlly3lONmXFueI7llk1LX+6pyccRvK
SAC6E3vTqdnc67Ly6SO+toe0mE9JHbt5mdXzOdvS9CqvZ79a1LhaDjSVnQpHfXBmsOWZabatA65v
jueP1kegT6yagrH/FwhzkRHsHcVOL7xBGDSVpzsdqZ4mjvoNqvk7DaLIdJaVa1dM2GWgKnF9nWGc
/PcE95NggU0c0P5a/HtJjQCo+MnqH2bpdSz1EjXluSPJ4/Xx+jiEY7j4KYmcAU/9XAxhCmqs24UZ
CApXcxIwa5RDjuoU5ttIiC76tQ4gXKGpEZxZuFQD8DyJE0ucA4OopzjjBrgFKQwi8+wKvRWa9nwI
RZ3VMSAqAcNCDVxAwvciOlWVMcF2xaikiXy0Os+m813mzZUghxVtYxWbJWGC/bXdvvcpKMxwQwwF
oe3Fc2+ostIS13E1tDMuHAqltgNWWrW4IOoCdNiac/EdpgOEO8gkORIRVjp2VcdeMGsZY7kBVclq
6pgRefpJMtbo1Nvjwkx+Cso8ckqrcgwHdqt3BS7DgSCo537VcrVjya51YAZoMgKri9dCO12jjppT
m9O+ezjP7SYTVNoP/fXy6QKevMfsJBhPC07EmJhZwOqO3VhzkS6cQsCvZ3wLd12diN1NJyn81RMI
kYNnKP1EehMzP2mkoTVfP/DCH34I8iOBQZcP/SahBfkzn2lQI2/F6VW1wD97GNY8EXrWdqeiQcAe
DDUFcEBk8SP2OE1sBGYmhmFAjVBsq51rJWNruW9lbADMRKMZLuYmimIZckBB4BpURq+keEZ3i7kU
kbazIz13bMUWfBWDxQk9U6j4rKD/QiNtYEEOzRVGPuwRJGPVAJp9phBTnlk4eFHukDMnBbn7epkT
PHaboP+rVLzO/SsJAww9KPg+l/NX/QM3RHC6jsIejoctfTyIjavKOYcFbRcqwZC6K++y41GJgeOy
qpGsVZzWDPJTJGGktiWpYCqszOh6OpS4/H7QtXESXpo9+fpyI48zdBOk/cXf8Yh64neWcvEoFWRe
bLOCOwYYnF0sWEc6pyUoS9vbcTa8KYjnsRDTa/gMHFg97XbRaI1+e7RblcD5lqTr/2Dj82nb9raN
P7tmAwTiRFntU28cGfFFYgn9thp1hEvM8a/cEXnZ8FRWw1+cXQcRgbDWqbiUBQOJnAGk6dmsVqVI
WvSyJPqSjWUth029kDXZo+6YrNUaMDMCskICMpjYVcVvIyF4rGKj2+SgGZkOUS6qqapkA4O8UpCx
ryVb19fBjY1GXb00/Uaipn47xsbs5p1GNjqnuIMImvaT7Kyp70uOEwJu9uqkDEyt+HgzWL8Gwpr1
huXbTG7Ew5zZJU3cBPDBft9/SuWkBB3m7WgOD2pnC5M2fpwPk1txuA1HzAIxPUgtf9MjX4lxaS8Q
1xZ1BdZ3DquhUEyFb5MlKe/a4cNG5vXTCUzHnG9d3pOnM2iNyxCjgPLWkth2+wc8YqcBndexgUeY
7behakqg/+Omq1amIrb/qc2F8pTm2fjC//A70SZuQCjKuNcQk2IxTBQy/1/MUkXjpxWDO2WjjXJS
P2u56dGeiuJy30LSBfNxs7m8UrA7BAN1YpF2KrMjL9JKbXsg7M7Kojblf5H027Y1zDjXILxPT9fq
qatcATq/mZGgic/3oovGuUiveIlXjTvBMkocJqj+1FYnUdX0aygyYVWKcjCCZdLADAuvHmmjmazm
9Rj+SgiZwzN2n2PuluispMuc9bU75e+MJv1pr+KkLkWRA3cKurdUouqSa1rrJoe2Vi8ifC7LQVtd
LxEk1C30XQ5W2YK9bWEhqs2Ab9nC/mAFw6Mo4+tfbyydNhJaTXPrc1fydOe4pC3tgXU8ybJDwooQ
mvq08iaENjpmytreq1At9l5o04gZ71HMnY47yq5RrovPc8S/aOc5V/dVSc8sN9O71IHgZYvj0iLl
TFI53T73teqmg6Xs7tY3iOMawsLhZ8LPX6kwFMdt2V46CPfFjEvwqL6FE3BHI8RHGVuWMw55UdX1
09VWZmBZlbPCePR2w/vfaWn2oN7E/GkSMpxEGg9bb8bgdZulnqiGgWcCTMcocgoTy/gQVJJrHp01
PL/1lNeaedJxODdO8qX2nwnzq11FblsBmyyNsvq2euyo3sMgh7pl5XCtOnOB8ChufTFvtYeHIPse
APOqMMEIMAC2OHLwudktLNekW4eh05wdJloUh/iDbLksJCyAFVH6pboxeeiyTdfRYc+U6lGM2xuk
e7jvgburcLb7l0xmrxU/8C+OXf3Ohl8HKe/nSWHdqdy4QwtKRvzFm++J8YcTwmzuUtUwX83Rek68
SUSQxd9TfKvlbaLjEngWMZEfqWs3skwU1ebuTpVpmTm+KeNBDyblyfUo1G+Rc/4uX1gilpKSTPg0
Gk/RA+5vQ1PgnHyQ2MRrGfROqX6wDNxaYDbdkVEaRSf6VOcYr8QT8X1ysMN5UYLGDZlLsFxe5Syy
1EEWGF6wsZSX66/b+EPMdnx3Rd/WqeLhiXb69ipUp4KiViNBqFwuTMo39hish2+kxOUBqVPnBWUY
mB93pMNpYG7QPCQj5syAt4jGnnKxvV29lUJmmPZqTJ4OwfmHkp+D7xQzZFGqaAfJSq2FZdTGtNiA
TwuSfVTQXNB5TzRZgFjm0usq3KOBVUoppy26TzzRntjJawAW2eu06VjS3VEw6sJkpy6PjUNc/tpk
5EmNBVXa/lRMymtaUhUFmlSZTC/s73lUQREh579Dmb4qPXKsyYNPhLGAXKyMcXqiK6ch93fQljz6
yIsu3udGw3Fee22yZcH8+kfn4j/+VoExKSto2eqVVeLVXyW5yssecDl7Rf5wIIRNtL+ugsntCAXR
zG3YcXFU/F5E7sIjUVN1gzRlS/nju2qoLc9WqLTd3Sop7hPHD8sxgVVGw/8A7fR7Dzq//SiqogXD
Jw8HniCS3ErGH4TtbfmVQWdWaDjAntRn7tPY05YTaMj7A/bOiw9DM81HzrPo/1Fw5yVuOqZjHTTf
iWYAnQkKEONQtLCyYYb9S6VagoTmg0OcH4XqMKCiNvXbjOtEMKNNszfjby8gG7meUh1cVx3J9CB1
9/x2l1pg3/uUeyr0iOBv0Wycp0vx/6NdkWciZbtJqvi0t21mBPG6LOKOxLTvhNtj3ekNDQZ59CQD
4KDJ0OT7p63kTsXOccjYGjfDciOl267tJHARe3ZwRclrfPgHkKEPZoq9im/LIx7OcBAO4RX6Idad
3SG2bwg7N3YpOedPbDZg9KU2H/UIx0XKYbPZWyN02S8PkGoaJNJJI1Cj7e7YFzopuRvkZvkDPp3d
Wx29rXoz5ebpBBBenbdFHFYrrZ5bQZpixCSB1yJQYxor5g0uvWQ0eVTpJpzQ4l62cCuWPP8+4esH
FKUrIT5R21aiJ+sijnoMaJiZzXJ7G0DyQ4mqIWEbCVWehbod2qcKRm1Dv3Ju9hyG4GvE7JwHzr3f
DyR+pPlrGauk33dmqIhjDxzM2GcgynIdyYR7gLwBEtAIx0249uLsY/Rtk4RXrZvv8k9O1mqJCDzK
qEnc+K9emfZc9QC9eoT5VmzJf3iVGCyVne330k+IwPnjWyF8wLPE920isOA159EHx4JXV1ohWnKQ
01jhe/W2OUcnK6pGlcLJgigiZAGb5LegOd970KNbAI83UpmLDcMEu4tzlZUPG87q2bVqQrZVLmE0
DH3KvRA9KO4HJzwxB8sMAnHeQfXEZGFpEuF5TC228eI8+iBCHBqhP6U+qqbsyBM88sA5vH/4HCMR
L63fD222N2ARZrZkjd2m6/19xdTzrYQYhx5dHVpf7flHcpAYVEcnSb0SXDsZZvvf5qJWoyK5CIYU
iWvtHak/B0A+7LxWqLrQa3H/k1OQRfNi7qm0BHr9wLVaTKc88BhMeP+0HDy0KEq1GvpKfNsbCpeV
0zBgK0UlGyI7/A3dULp0OZ8qrVL1WAfx6ELRwNn5ZBgSWASde/WeRuwPYvm+SBixIXIkNO+WXLul
r9AorWETUO0+TXtMmId542fR2jiwPLHuAn4VU/XuK21A1apa4xznAd7PstkeyBhP7on8od3ORRju
xYhmxb/r4IlL5HRWo/wZ+uu5LVHGRrVJVByhroHM+lCG/6+N4NOo7T593gc9KL95dshrlxIWdykA
Zg4ZNN7SufDvEbZ6rWAQbXGAuINSm4FK5ixz2oxRnW1UNfrPJJWqA5dGRnzKTQe3lDjXb8ZKx5dj
M7X2M539NyKiZ7vzJVXIS8+SjbKx2GWBm51viupEMGHLCAR+DZAMDP4zWktOaamAxA+laOx/gpWp
j3rdGLQ1bGuwC6Y8AGvBuEdNy+lzZi1uUel1au1Fve9GzVH+ekmJ2/1Irt0p4GeNP8cdgZBhByUo
vnRyJRE5EjFXBcgzGeY7V7/hFhb0CQwXPgLOpE3bKfNR2DJPpIHjB403BLJip+DuxgaTSwZDxWUX
37H7QsMLKQFqUS0DNxFxhF/Cb8bM2HtsT7emU85+VotwzMJkjePwVmrKX95LplYLQ2wEY8zwbD0J
+4MXGadQwMaiQUsPZsxa/4265XRiTKgd2xDj93GJ8LhFGmB5gsVubI9VrypTaeFTMS7IXt7SxMU3
WPAuHWJulmeaKSv43Y2g5kzbMjo4nAHXKd9n3sxgbUeIhbuxag2uYfL30af+8iRPv/4DLsrnmFo1
Jts3ePy2RYRd37GPHdp1kIKCOsnSCcPHhcWmepNYhoBtHl6mp1FBz71RB6xDiOpOaIT4rkVHzeAJ
bSZcHXi/br35p8XW+cLJAlwe7gBalgulMMKnvgofMxYzjCJlBVdWZmI5B03MU7EPRWQWYyfkrTCH
EACOPF0MkFFLNUrsN7lPwEYziKjl5M/5G49eUdfsZOzu73RPRciTjbYH5foCrKPzTCpURa1lNt6Q
A84DMGyO/ht8DF0sHr0UuyX4SuwnYcSA2kaEDBlPf3a/Ip3zW2H3yap/J1VZ5Na/hxNtdSA2gwIX
MDF4eTR+Ra+vX2t81p8eWReD4xPmak33yfR3upx/6jElRRTTLXfxWQeQx+cGU5HFZOHwztHuR+nX
9wp05/6zBp8W399aykMybbccGOUNEe1zEv/uhwYs73l6MU3JUYq4Qn41rTSCDexhBOar4QPZbIby
znMA1RBzhtTXJY+3l20v6l7yfBEFAkDilonnb524mumisb0itTavv/k96wkjzdx89Qtr1rm+nSv+
DnHphV24h50aTb3Yw2VDGZ7qotM0b8KJxrgOgUR9BwffhcPkEQFvUCOSrn8ylqGr4aHYc+Q03iJo
eKqSgurOUphoB7J9UXwOWPYrIYwBs/3QV7UynpxjEi9SYobNLF3qLzEBAEwQc3vHuCN0tVu10C31
rMlDjVHm7LDFDWp9I28o5HG/4ZiUXfwk1GOGmTejFLCFycTz6C+gDjrAQYRS6bbQT+3OXrOcIwgh
bLaQW7bwfmwcsf0/WAxtvaENBr6J8RFmRThlRW+rv5CxVtQSTbqV47qk54GZ5BaiAxhG2gF2af1r
wGL1kXxC9tzWIxOsjvocU4BbpCAyuWWHMA1kzpEK8O8sHGMxjgyADqiihARx5VO3H5nAAbhEhwwx
epqA46EQaN0MieYtJ6yHwcXSmYkKHohYk9zFfQwM1AJmZuUfiCen61H/eDR2E/XeUxnThD4QsCCf
IaAoVYXAYA/k4smQpLM+HRlCVpjZiDdx9JGjUCkFiTNj/Fbx89nmUPeLHSPF8WFjm5aONn8TRguk
tel8DcmsegMUDklT6rWFcduwwwh9YWWG1OUiUsOD8vRd+P1fOZxALB86k4xwO5QxCRMJ1+SnjHXG
rvbYtvd6F6GdXoixcRIkLuoyofgow5nMd9JkiJv664fD1C3eo8TaobI/bWWTB9nrBO365SBbEdpL
Hvvcjw8l5EW8YEhvBrh5PFEpOCKkLm4bcn2LJRIb9mfY/XalD4Dyh7FmG7lsdtEdx7CkktFyAfJs
0UPMKh5g6vjdKZy+vrfV+QPXvWZw44UfzKo0eqE0js+yW1w4jCQ9XkjYZdzIpTXUwhEWNA6mR2+M
GEXUvXdmdECHexeI4wq/UUOooPHnZhLFGH2hIEpZQpzBiZu2Rgm8YoFi5QYMLwbA+iGU3/MMto3f
t7H6LbX7mHLvv3t4ZmxycXT+bETzkKNDz57GNWJKaj9Pph1pB6kRf1Vbk/X9A8fzAncmaTqUre9U
1RIg+sqa1eYt6AbSDzP12cb5FCtsI0HSHXQR90qqvxw+CAiXK6VRtX3Ff3OnY5RrvLQvhsEszQsz
AUF20JnYhrc6QDBLFEQAV1TjfM+RDo+CyB6vBRQ0Nd5/d0Y5C7a6Igt1Dq6MgPWhfgW7W8z/ANS2
KAZh+aQPf48uetnQ3Rab7lNbfS4Z92N1jK3pOXEruxIlHSgLSHzKr1PVu/+k70HV9Gly1nX8kXad
FPzTe3NC6C4vID8jX5Cw9UbUMjm41aEWDqxlgYzxO8ko44U2g5kmwOTe7xMKS9zoY8fEfgSaXewU
5mw2lqFhXYvRZwaycHf6YIrD6PWq89/nNTnRRpEOeGoR8Eokte42ceyhJUfqvr9NilEOcH5QX04B
/xsFycZK3yoYZx2xYdUsSXAKpMEjSgrnXaBOMHbYeQrCA8e753T16W56CGr9IN2dROAkvzVo9P8N
HdXU5Gn/7tqzOmr7wVusrDobUMoan3K1pnUIXg0ahIJrdBHoe14iXX2NQ+5qQl68rDOcV/cQO8GN
IMw+L6abewrOxuHSWyBW9hk0KI7cbRtYyCT/JZVppfn9MJIrtPUKgW2vc+B7BvUonIQfDS21RrQJ
6n5icTgLDWa3kQUXShNmW2DvmikRRIvLWn2rc++4cbg8nGPJebvuDj5hCmLTVGX5xpZNmpVzbiaG
ppdVhxiGjOu/UdLK9VcAAAQjAOOwy30LqKcjWX/H2NsHcCtruWIk2wV8LIRewTEyEV2VdvOx3Z8X
7vb6AcPe0sVA8cAm7ftLB3HRq+YZNk/sYR08V6MYFKjKEXMcZsB3L5InM6St4xO0uJzeUQxM0kao
lfpWLGW1UCrD4Jwt1rsXCEWB+h3v2YLWel//Sr4HO/9bx9mZSGcAuI3+qgt/mApvl/S4cc+U/DlL
71r6wWwE6Mvot23eji7sVUczBhjTDAccY4vcY83WLXRzRAPSPrHGqxs0jLqlLI38MGD4+kfa9jof
C51vi/q4187/ots86wN2j4XwExeA7/lkk3pIw0D7aL1rSsTxbYF8mTdsVFBMSS0OopQgVnIC4XFD
6at7gKUAQgRed5FHbrjsWL29FQKCK9tIhXo6lA1CGacXXVCiZ1jFzC9308IBs/Ned7no3oKP+bp3
uYgTnpmVhOYTEsPjRTZYqUA7glDMabTPsPVOFday7uxjN3xtdXIBfH5P1Pr10M13ewDgUNhSHzS0
YZVpc+feg6DCMNBNZipMPcna5Y9rhxqL+/rwhXLMd59qEVZpJD3oFPf9Aw8BKzCnki3NpKl1FZlE
Li2m05CEuc8OCSWhnwk21aolew+7cPl+yvwzRotOOEHk5qpbY4fMFQljSwLE1HGdTAmW4mE19EEH
SyE4TwQh02m+DudMpCV5Xm+QkIxFxl1MwdlnyoZAlG+8yVcOBiCJPnIENVlNoJoYwZntraYQbM9F
6OHbaxz9JjTp7LvOYYTM6tXe/c4vWOLSs+69hQvUNll6FXkx47WnIDEv9nZTwXMycXdKMWwYxahm
hBPLJZ0DzdDaoV0KrdNuarPm3gh2QjhyXfBHj+xNAiAqBkvjQLPCRLNP644oCsrDvBoBNuKyt/c6
vygIy5kVyP3tACsOCGuobaUT387TYW/5DeCnLPTEwnE82qaVnrM5uR0rK93uf18Zqv9i0KzdLLc9
n5/SHrCEmYj6Ze7VlprSSkUIBC+4q6pZxSRLKldMWcFA6E9NUnWE47ha+PgzXGWUlFIST08TEHSf
PRs6JC+Ua98kXVvUtSVaR8W4AVvJfzZwET7lNK8DPRdYJTlX9a9PCtcGOBq8bUKudpUBKIkBiSZB
J7KNGQ6v6kbtKBaR2AMuHBb0o33EQ35q8E7RS6j9lCqC6P2koA0OalEn0M/jW429D8xu+Ihhlg89
XeaXbrAJcCjLM1d4gpVgJrgCOT/+oGkkhfy0hchZAJSSpVOtDndasFwW+HvwvqcUFtES9IQuKUud
nZvAp//J6znlhcRMeKnk/86D/DwL7RuChacM1Z4b6EuNYPzqWbxo4myvkkxbvK7RKxfswi+67J1S
Sn4mx1jyDzGgYDgXAYKCH2QgDPE/ammCs4Myp6pMZsfHGOxnpyl2IG1ieyu1HxuA4Um9QQdC0K7/
x5mZMz3O3RnqH1Bx4Tjt9v52ByP8mNpk1iQl3oYgxlkE8fbjiGI8q5OzXX00LP4YbHMzt7cA+lMk
6eh1vjyIodKudULeSfTr2HJ3RxzqQ4eCRnRu7tY4eaJ3BmrnfaviXhh+aFntBwrqNB5w4Hh0M5sF
xuJ2gkBqr98WiHXMlW/fVpsL5mQ1bve4T/PMArH/FRwJh7Z2/KC4pSAcgqSOmarQ7pBR3x6PfYAv
oQhUf863hYrLLDMrWML5E6EsqbjOuPX/3Ixz8AAb/61/omOtHJg55KVfl9sZW0chWayn2pk+gRy2
BnSiT1FXmuj8SiuJatJznbN7Ypqtsa963JNqJgq4ZjEcbkG4ds3ehpo6/A0T9CFzUBtD1ZZtKj9x
r/cUm3TNtbKdaZWfszO+P7iv0LN2R5GwLz0SY0clWi7VbHyqhEGU0OxrGcAogkOMTGvNY6njCaA0
HdAiLKFz5/LOSQxL5aRa4JLGJmjlt/6iZvCG4hROwuCEZJedVUxmWEZZXiB2kMaZ+7/wQRPVonlp
Ii6wTmlzJXVIEq3/EZqD9HF9pk8JNCZ5ko79T746Q5LsgsyHqH2syEwid2ettGHV5uL7rF/tA9M/
44zZLkTZnKKrahK9ZIJZoTPbDmLqKKWD6rvTt+K9xsUIITjXPSz2TIIaWiGb1A+vGxFKKFrzj5y3
+tKsMKztHsFDIV9qHI0K8yTXo26LJONZwlCPgsYCZVafHCYYcehmgIHjaKVFQgdpZghfBZ07qyJs
ktlv3iP7PFVK2yGJ2CC81+EQnueFn2XWCuhG/HAPX55jGxrL00G+scjlV8sud0GfIH0CRrQzEFwv
tPzBsmioqoccNxqZkEvJyECCQqnyB3SJDTwPG+ZwUD6Uj3zAHNUlOtp91qiCgiNqR+TTkUokQ/ya
UVmsCav4xpkjMBRz7MWxxt8q0n0F+E1/QSayusibBcN6lGsXplQgPB/nikY3x8XguTCVanbbxKs2
nkNMU9jRNOWhwX/DmAJQp8G09Xf377+jESwYz38ldrqXpeth6eOzeaAXGrL1JD9gkLx8dOIUyeCH
96VJ/Pcwbun50BngYFlYPNG2p+isrTt5beq5vv6EZvVxy1Z7Chj+CNvk4ExT3asG41nE8rQYU8nH
lWH2dYL6ns8cXvXNkiB8zTNQlhnQF7DNCsDQF2VWiM53S6jsL/M/hh0iA+0+EAq9ZoMxAWGt7u3Z
xq6uo3gRdpyTlu7n9Zey+S06gEQfTPBTOHY8DAmGLu97HRrCMZq9RpIvfc+mR7H+7yyZKM195pt8
JWeW/1lkuzRvWHmRL2fPnC2zrFJdY1Ro3LQjp2Bsx3Zk8j7ehmCTP1EaaKIwN1PsoKIlwonIhklM
snzefnaZLARaR6SvZefZmYMP0eqZhgxQepuehCr+OC/I55QrcWBdslDDLFO9Upqxfw9riiUhjI+B
K6dpC5PABA+mMm8dQ7tsbkqlPWWSgbONugau2UsnDjUP0uiJo81OdJjjNbijfCjzxHpYimGjv42X
vk9QB9STOSD8GGjfE4fwC87biF1CSiEEyC9/lKgGYg4Hwy4KT96c0hK3twOTC5U6EEv3yFOjmihn
EM/P8O9xdEEYOo/Wr1YT1LTu8xK21he57Dw1Q0EyhFslmOlIIKsozRLvW2qV5ew61JCtI7migETl
wx1vP7ynwtfc3leopTjn36P94F2gbwNAZDqM8w7dC8jK/pU9cp8piVTTui/CnbN8gixnjGTInyah
z0xyYd+NvwLNsMoroOS7m2er+VQLwgDVgoinL2okxzEgXR978xcwsp7rjcMR9hnTcV+9Lnrk9V2N
jeaH64lHgaBI4aoTbK/x8+9O/KfmZgIHEonux3MdGcZMyXtAtz1XolzCYuGpIjUCAaBskEK8K6ca
ILUzb0zJlZ+8XxJ0Yv/adVtAil/o+zj2WqE9qhUzTnrsWidzVOv9tz1Fz1cjDS6iitrJrp0oH+1p
/4tMO1UlQ8vpSIhmeVi43Bjk4Ryt14PdOk0rdsqukVvBdBY81TQlc3mHDSUiLdPBlgtoDvgnHdT9
o2Kej7C0DXZiY4Ui6aAviYcj3DhVNvkmOe/MRpTnezByCqxnvEjZDnEvwqThLTumWw4n0mRL4bFQ
eqZY9ByxOFTkS1LrYmABrhoW2aGYBKgZKdPej6PBF+B+fO0BeVMmMYIX5BZozAEBUUbjY0sluaza
j705m5j031hkHmgZ/5vbNgAiKeu7dv/3yIopsVvNoDSIwvD9X4SGNq6x417nrbF+IhazZRt9+Ef7
H5KapVra779qVREO9SLW852EfA4xQXz9MoHGZ/gmoCN6JJ+cza1mTamYk1k6WBW+zuV/24UnPJ+s
2mgcD8JqjY3AXUIOj9MNeBS5CTJwSRgfFwKBe5EYe4bU+RgaXF+8y2VSoS3xM98602yTVd2b8j5u
wF+H1T3BPA0xD5XS+u5PzMKjOZMiJA1EFPv1r4QAyyDRureqQQNOhesIyk2ZPVVMX17cjs9PFc7d
5/3+2lps0SyxrRi5VNKEWMzOUBy0JEEToPGrNbhHXHi5yM8nprT5f/N3ugwfGVxI8rFWhdfaJrd1
EcU7IYDm/WFsKkayt0Cfp1SN03z5Rxg7xvQVwrjxOEPos1/LvcW8lYyFICiEIaZo108QFbJp/TYj
vZgHE7a+ynQ5NNpuo54h55nCxwVtkQ7vqkCQ4oUGTdO0TfnwJ87awlrveD9B+9exxWbm5AYUWrrx
7QoSUoWdRLq/g2AvK49GDPL+W4X+FoP2K9yZQGb2zNntsH8mPAv6WjYJHZ/ddZ8/YF2ChmSYi7vo
j7SCdEwnPpiT0cdD1t44zz2ONAy16ayWORxhcmK5UZtwjqQHmAzlL1QoSEY0qZQC2GyEHxhH+0mY
LLLpDNdY6R+yBhgbvTNmpirqTCHyV04ni+LDcErOushO6PQKmBhYZtNUUKovsdJOuXOHRwOxyoqf
kqkrPFd9W7qRxJwUXBOQ0gCCk3wTI5ZlnDHOvTqO6kC1cvpjGt5msu2xPEs+HvXqno3DOL4xRxUh
iDJiwm9v8RC90IDkE8xVmAvv182CcYe9ExCNfTAUr+PvaLYEZe8Q6CEH7MOZloSqwsKFauCPsQGO
krKOQ0fRyouuONd/ntqPRtl9277yRnLukAfBbzb4VwJcQWaEt1o+07VykejLAtDFdEwQPiijamZY
pwvXg3p70gXTSXoKTBekpqEamMjfcufksTEYoElkVFspZIkBqeG0TvY6M6f58ghYufMjoFq6OLoJ
cp+Wd7376leyDXsEvf9o6iwkqCYk719Gy2a85Iw71cy834M/JRSHLogZz+TCA24X8DV7YGyzp5GT
1GrqkaAGLUPUvHJYn5sRbxnwX6Hk919NVDpfvDkAh4obsP3eaVrfgG63asxxO0IscaBGcOFSR6DX
ZccDZW7mVh5CCOt/LiqjFzlW1KaU2LPsIUVk1skFvMxtiSpQdtghnbmzSpwbJ24UTaFqrM8kZ9c8
5sym0zY+wMFztl6LlTL2gGyfbmW04Nmm3C6czVzx5FqNmnEjsw5sXUIVcyWIQBaj6s3jlJb9XQ7R
6TRonUiQhPuTpctRrvfxC5A08vqMQQU5q3j4jhwqnVpsKil71im+EjAyaPoCxfq3oIz9gNPTVfo6
bytWxbWovmTkQzeqoHxi6aqSsYp4RtlqtPSPRliCrHAVKGIunXy5fqQjWONq7W7gq35I7f/nSZXj
isoxtxAsEeUrv9zNxxIlQ1oNFAiJPMeGfB11mlpxGMhhs2FFcdnJDE7Wpan40nt/BWyB5+7yWrzv
utDvjn0eKJBpRySSpr37AhjQ1q3ptW6KppD7/wPP0cV+EI9OYWOQDqy3lMGNPlRAPQ/2egcBS3mX
0ArRD0AYy1oB0yt+igwtc5+FHrcZoO4O2uF+QWAtWMH90M08N+XakVdr2ymTYQ7fR8T0DlU0TykV
ErDn+CkrDPdzBtH0z6f2SLuzjjUNhYi9cwIDFhDKHHpSoploHVGOMxWRfUmdVVb95tSnWRog8d8W
Snr556toRQEElVAnzk0JDsMyPjM+DT4kprMxlae7WSOgvogFpEFD+R3j0nc7EPNwrdeWcqAfeogt
OTpTHmHmJnGFrZBupvgPNy6bl4GTAI71S59tsz2//EEVchhs/b1ha4C74yXGpiKGUK8riARo85bF
Hk1X7DNnAi/wdPQK34mxH7g1lcZPhH86vXtlLu8YIik19tdX6xqmurQc7CKXqHYfTMcll1kVrLJ6
/VxC2cIWNZrP62XiMRZRw0ND86ejVJD08snzch5KodNqoC5i5qB8OQ8JN0SzOVLqYwhaOcSRoUcG
y8O7+WGeGuhXUyAFsSlyvVqBDTaMKJsut5jl8p+o6dp7KCyGFhBwRaKSEXIlL71wPMLYZABOA/oZ
ijjOsiEq98Ix6iNjmbgcsREdyhAItGY3olL6fQ9ry4x/n73rECjL9ylIeW3IJBEZ39521EWv4F6e
6+PnT7QRdDa1Ey91fzjO8Jytnewd+ESDIcDM0vyKSbDpXTOVjK0GMkqZ8KzS9mEhMENcKEpz6t/6
XmPDezU1NgpJMDppYVe16EeKkQ9KJS8Lbk7aKf7sZlWK3dky15eVay8RjrXiaByhNuPERnBIexhj
Yp18G8q/n1H/FsZ8bQycu9u2ORnbyNkN4q42E2GlIab/ghEFOJo9JPnan/2mIUGm0vUoZsL6Ngzv
iL7s+KYQCA6XCDhb7CaFNFu5IzPmpKl6umGl4KnF0VD+PnMGX/+HvJZFruaMbUh1DvEM+R+0I+fU
OBuujGJGc515uossj9nwJkGDqt/Hyz7rdLYB0I0F5WVyBCr9uOOYWiDTP5OU+8oyKx/3F2DDBQl1
mXYNnem2nZj0JGDmfvlexoKe/P1zX/tYDPt/hsxns6n7z65y3nuJzSBRAG+joMn4b94urthLg9FH
Ia64zdPeuCkDJW23bsbaBBJzHyYSUBf5syC5WVijALSpJgNEFTLvvCWIb0LkFU5yBTxvp/sxbfLR
8ByPoTwnvGJIuhAMcbrs6FMgw2nGOBfQyS+fF3jvPQ8pSzP35JJrHs6Bs3QV7CPH5zGanFQNgCh/
VbKaq7zyzib4lSwOnUI6SzIEPqhqWlnBdzrsDBJsyrm8HcgAQ3PDN+Tnsa+T1MIwv6fhkVqNJPlo
CdQPkq1SkavATU+uUl8PY9+XPxNc9oM3z6BJ8v3kuLS3vG/Ly4QrqZlOq+Ij96N2/By0h3SS38Q1
872tRvbpZ91Z2Rv5tgX6BC2lVvpPQcWDP/Pw1lKqrdCm/xOSU/PHYbZC1CiJ3uA9Mcds4OWG0eNO
zdcoZF2OhrGzzGa21xC7FbaRbbwEvdLUfJ6YLAJOo/amyuOznUYObjSVDfcohedAp3AdMfgHGnH2
zCC3K2P0ss8Al+x2owdbKLcxJnt3nlG/1nt4zf21onftgJtdlMIwtCdqn+UwXVNSXMceS0INQ8kq
k7oYWeJOy9abFVf4h6VpYZ/zLivGdD8DIrJ5lRCFQGLqsU5hyyES0JdEDmAY+EraYrLN0YPXoje3
KpLBQclmc4ado2Ia69ykmJB07FPWPr+189bmKI8mspDNgW9058kgAAIkTDv/bjCIreYIfyeQ10f7
GunKdo/6yOx2iSzqAHsLGR93TaKDk1AL3otT7nlnhbqGydhnamAVBEgpGOxrEW7Wi6ZVp+mZowbr
6F7wply/SujgkPffYSm/6qqthmsp9zlhaDCwtATpkE/NHNLp6VhOYaAxCfVaSwzmC1WGBYnmDyM8
BKscegh25wOD+u2AC19lyY8c5OTlwmRWZxaKh8p9vSkCKs175tjZwR+1WSxOK5xCv/IdKvURAV3Y
Qqn+I+aKkjNYFVjwNDBAw1yQOdsPJakEV46HQUnHrvrOtuX5NK+v53m2kC0ow0+/Sg0XExdnRej4
+X6cp8iI69YXdg4tAVORuafeJrjlaUzy08D5C8fZnhfLoBFnep7TPoMLDOyoYPHnErLTkvHV2KzP
9KxrlDTGfvAFsXyvXxRH1QtoGNf149chekAO/CxwuLPtilds066giru/hdSCupNzFnjrvRftb/xG
Ys9WdeUiDQiBRvH6d7Vt4MMTtPED7O2S8tbba/K4BT0//cnpK+Z0G0k3BQYAfAx5K8d8gaKCzBlm
UJScwG3ZsK1zDo2WDvQMrJvc3t7KLv7yvRiIjhaK+Bj+F4uRaaC226IspcuOM2Eo1N2HGf51mlyQ
pKqOwab/j7xxOgIZjv/9ZexKzSQcgiy4fyUhdarti+TcsOwt8mGSBYrrh4+xSiY9s/E0NO+eWced
fWRULVS3CjzclcxQUR/AIaTUz2axYIWt49WM0EZBnGSc2vP1+3azLo01k8waRZSjuQfy4xf2ZKg5
eOvKj3ZIYMgnOw+hR3fxQXCWkNkLVCXszB1sVX2M0UPw7H2SO+xFkGoVE/jjDiVBGFj+Yf69PVZp
rk5DG6+5KZDAb3kTT5o8FX+/Fn81ep0Tny0J6U1eQTkLpf+jVbKm489oeJBqyEdPyXVKAgH5bRfP
w4a3eEHMeyVqxEFvkwtrcVxd7Qoh577Qb0DkzeaOJkyBqc40yWqjM1v4nOYYGPLFQjpexmRBb8RE
4gNN+EOAfZvNVlPSlWBVVVBQmduSV3IWT0HxIhzOrbC/PYncoYHs92dbo3+NzNGphWERmlze+DKo
UOt1jXPFEQd01WRw96QiuDimVzY4l/o2y4IukCIkHcihKtDoysynO/oIVXINMGkf17B5pkZ4HQVb
HtOnN+XKPvx0dvruue6Xub45f10Lccpr74YIwMNjPpixGwzHMYnaCpqGcvKUNQhvQXNK4baJGltN
ZUT45ED/L6iAjkQU0al/bK8Vqap0nCTUVR04jvOupHnmnuaG3/kCwqQmAfbjgIgHyM5P7PywIU7G
C09p0/7U9f+/GWne8bJA5R5/qkPAVBX7LpulCbjRRoy/Vl4bDNjFsSQIcBV7O85RphJHg4L8r3se
jMeF9vaHvFLYMEMoj/etdE8CE2z8DmiQz+I7u7+FsmJVeFDU4N//NBZcm6AHyux1GDln/hQ7JG1e
gt5EtI7WTDPEdQl3rcTNxdZgW5nVepeg4IUTkWWw/2PNR9KgNp+zoIYk6vmhp1WBJsoTcvmQnRtq
DF8RGsLDg95C/76Ccu8v2E52Z2X1fkc8XhHEtmQpoAvn/pytjhIQmGDiay5aZwuiQJwl4Dj1iEtH
LcghRpo9Ufc/gG3qbBmWPHbeVyD4Jk/2gGa4szPkIq8gepzi3iRRNFims0PVoyehL6G8Zg5VwZF3
9n7O6Mt/UgWRaP+6HsUDObRAuxwaE1FwkCyEkc+xwOnZgYqNAMW47vdBN4UsTZr8oE2SeNoTG7Os
49PZn2hBGxKP6C4/VGPnszI1/rBhfR/HxGnNeobzPNyzwbvBAruWpx3mBSN/oE9EHPPAZMT/4xcj
WOvQIBRgkgDs850NODVc9Q+sOhou31nnISUUh8q8QiSFGluWeKtvB4DfRhOyGXgzkpUh5wGMdmCq
umMxuwAPfP9dfAnmHM1PzQX4adlVWUffH2ReC3Wx2eWizpw3tcs951Q+yxqXHK78D1cmAb07bqe/
uF74AkGoU8XgXrLhMuApMBnUb0ocnph2/lOuIfIwjIw55cTPT27NRS6Z5AzSw1+QFzNFbaiCZ4Mr
+hXc74OMt500ELlUDWMQM3ro7WdNdgvKRE9X4Ox3zPttzLZ5rtR/Ti22kXSPZ8bWOvdWg0KLO2jP
XGSjS++0oBZ+fJ1fw4gyf96gKbw1WzRRxzwusdvNdkfDp9Lahiqd5h8IlfBZNsjW3w1Mv32zvbj9
5rfc8J6UnEt7OCTFE02SzUj4r5fIfW7UEh0lFGxFETdoEvathC8a1xMnoqyTxL5RSMlkkHVbv6n7
9ult7xEuEjr4QiLYBi0fNeWbrf8MR7B/iAGxWlVRwtxRTNryw1Zfm75dNPXehi2aQYZdbs8TkAO9
20uSsEcPt6AMasLhwi2Av525A05qVr8cweaNy2wYgR+Y+Jq81wd4p4zWIEMr+yhMgKMyxGaeXlBK
64HHuDlVSYoGgOpg0coN4dD2Vl2E1P+WVYRwntYTJXw0XR3P0szyDkFLjW++WdoWlvgPDIWTW7J0
t7EbGIYOFOUXPnc98vTDR+4gDYiOrta6unO9b/6HMABAiY3chV1sYtKH3c/8zDED+fjrvp9DTjRY
5bTTMzpGHAeJVakARjqd4qDGnlsK9lxlb7yFBRu+ts2o81L3KIRxwsDjCzp5RyEZxDkTAqY1kzM5
FTKlOLFgdHMp+WpaivZCCuvjfuBMvcui9qkiEtLcID37Oto9EEpQBE8dWIsBMQ5cv6OZJToRCf3u
fWck/1sEcskqw8nG1eyPw5xRmMmr2H4lfo7y3EJ5eb9cZ3Wcq0Lu/o5J6Ng3zDUw0S/+KNl4+eDr
5NBoColjx+P3B+gh4W7q+t57CJEm6Uo/sNAKNBC+fUDxHDLxEAyZjGA1uCb2ym4ixzgf4sk8e/UI
gt051xgI5HAbcbCpLvFBY8nfNSdDozYmkxIpYzLCH07JcnR33zEutsXFcSl1t5MACCWvRp2OxAfF
XmC/eUwJ0Wcge7AEdZ6hrELrGjCCmeRvshrs4tr0cHI1kXI/VgbmqlGpOeYaEA5jLYzSc5fJoBe4
NnSLQCF3VkcBHUOi3MnJvA7wXviuDwRBBBl5wOTmdKUTJj4G9fyXqgTroNByF+fzx96XPjWeTGwn
xqvxQk2DZgODAd9CPxbEeEnAciuiC/gxwWFCs3dREy8nxRWpn4JiBU7NAzeyIEYk91oWXjcdQY/8
GRrkRL7LAwya+Amcg0w0Cgnc3+YCljdBD61JmcVMqH6OBb/V4LiOq8PP+weNqGLHWmH1hGuQbX7J
ZSr0izpSxw8l+trgRyRsdxq2EnUnTLnGNb9SfsG8G2b/mMiTxAXkp850QJ7bCN8IeEVjrEfJ4JYg
tDdSDXXy0VUsfNquCsI2YTWGG7fX8mslwjj0dfXkAnoYJel3z1arXkDtq9hlTF50hkq47flUKNcJ
05pFaP/FG9KZWNIXZeoKu34B9N97nKPL99s+Rk6qREprw2PfXQFz4tUenuDrInawMd3suOGWqpuA
87ZVeLspTFOXqZMxUdBd2RkiaqbtUSwauwDqGd/IPtwFAh2J6uFBZBedfu6hnuqI+rb2tyhIRqJV
ibMXtVt9SNrX/aXKlYXPAZZ1G8i1TlIJSAOKB6LDMo157rEmukT5Q5Nijw5F7tBrlKL3HUo4SKiM
fz3A35XsRUesrOb7p9mshH5QEu+PpeE5/trfqpWD1vUaALTjD7V/20fNaB+pHNtW4lNdTfpCi6h5
O+NczYtT8sYVI6Q6o5tCpHseVp98Pj0Y0PgI6p1/yb8Ejr8FhlYCPw0E6DXH3s21muP5OfhwF7n0
gm7+L3LSNI6IKh+AS+xM7hEbOrhAY6B1UbqOgFE+FhjdpyuOszyg6gKNHUm5nrJllIPVvUWIPcnG
5Xu29+BanfKdkOL+4TFvu1zu7evcp5TI6EXH8oIzwVMtSjyTPEdOGKjIoMwHJiQzuecF4bJrrVW6
KfLFUvyqGH9PTalCkEp0UsXQqsGPDZQ1SN54fdtnfdW4QeMQPgAeI/cFC5tbQ/T4vq/jDED3OmV/
XV2AW1mhF3u60lat7syn8GWAju5GTjBGUL13CfSeD+iMGZgP/PtMzlsNDDKRcMHBU67wxfQ1bbZA
iGeAPro1jhPEq+4S73uG7tAxlRcI0dYSP/S6tmfODbZkqOmbrj3keI0hpPtxfbt71Dw1PgrXylwR
VpSDyTzFVybpzJ53yIgvnzahRe3HxHIbpXK3ku5B/nX+ucbSy/qNA+4QMtYq7XXJOFlpz02nIkDN
SZpUNrtOtRa+CCwTpqlEXj1Y16gHkMoB/2TgWL+T4yodLXL0vZfL3ukLMuDVy/vQ8Q3fJJ0scmDo
ut3s9ggdOOHKrHXc5Y+uVEEOjx1Ozd3OHX3HalMrbznQnmbDqOjrxuazgdoQCSf+4ebapB9xcA67
PKQ0mqVw0/yiqs27WJShIi/9EbSTP2QW9DlhjGQQWx4WR9Qm+zyy0MchfjeufPF1lDkrvX4JpRvi
HsZjRSRaYnZJFA797Gdovlklus6toobkki6BtLFZ+FHGT6fR2ylXPKiDtdIB9CZ/KdkVHT9nT5gu
U9jA8tryM9g1SvrrytXzsn0EYEKZltAfs4gbPBi7ilR1CogClfUrRYho3UJvReBUR72pH5GNgQLt
OTRV8d0mCNrPiHXYB+taeZzjSZWQ1MuBYbBVbXfjAUCqpyNth/O41deXED2de2OUR6nPj2QqDHS4
SOiJ9TOGHpUR3Cw0LJmMeOT6sGF9YLlOXczxkIqvlFxTCTIuEifoHEB9h7G8lPCZDLLn2I/vDeGC
jjiAmsTvrRBk2aTC9nnRfmtX6uTJTSnsJSoeyALkSmmq/FqEyCZB10Ou389oUnwCDmjEXfTKV88d
+rrNhNZYnTVlYrnQZtqBiic7gO9Wd3p07f+adOElUHt62Dwyn439U9o24v0wouJab3bWWCWc1qUY
K2nSmq0PQTsKSLYrDrvfMkGPyb4x2qD3SNTJNVtauKE+fZJpDifY27uQrU5sL6CTqs2L8wl76gmD
nyp6lnypYLQbVAomUDTPdgkl9OGr4QJ83WlbG6yNB2C2hcIFJ1MHMRqdpqUEdTn2nQb2+TIu1HES
nvo4DlcWy0WR41rrK4mOPSZFm3SoDkDwT3JLS1aGlyKy+YiZLNjJx6LirgUjj0Pg4fRcQb5JaFxE
Pze+oao5SOb2xivWpmiU+Q4UD4d9K2/S3dBcIgmBB8cY57u2nLb5CX1Ps/ngeS9rbLjN/KaL5Y5C
h5sErQccWpny3Nn/LvSUT+/3d+u1kxHEXrqNyG82lsolZBYeFIz6Ng10TRqcLC/Sgi4zVPAeYvRM
ZZKDXeP88WOG2G1+SV1vU1NkBh0MwmXPz0dRq6lP4IQmiK8d1umghryc/mI2/MCcnbJYBdeJZM9K
JJP23tjONV7Xk+fC+5+XaGs9o/Oo+mCVvbdcaDv9GdEDDgoBxTauUaM328fvB8+NKUUtXhCxwACd
kGmcPJi8sgl9lL/9dhM+NNReaQGwuXUY++vb8HSIPBqnxvhwFebhjJ3db5q7DVjFiq+CeBe5/zyM
XGcqvfkBC5NLUK3mZ3bm1vvbnzPBmRGxEwxvJLjrSIA68QfFVVF9CFJp2vC+btZMjz0ey8ALk+Pd
oms9Xcw15RIJFbS0tJwxQmS4tuQ/MrHyJDRj84k+x1JF0r8mcL1I9t8Fe3Yxz5tNT3c0aButvEWs
+0KDCdoDXKOF9VdUnhU59mp2BZ02NaosYzOWOHlY5t1/yXOMgK1bhxduVFWqNSxucP51MKgjRiNa
1ZNol7DieeGiw8DdpGb4AR1AdObUacAh1LenzzB6vyYU/9lJKy7YPLnOUS19vIzKq2F77hl0zmNg
zpvfqK85RkJm8Z58kiEkQahN1VWWI0qT1/JZt+YdgoqV3VXjwr8JmR/i2tjOV3VHOZRjegis0TzO
E4p13Y3kZeXTHCuMm9vIHpKKfbgv2G509O77W/G1O1qUEDMMvGVHVeaXGQsNV1eAkO11CrOBEBp6
lB5+q1bmTie4QukTYHvHbOeX5hZe9xfYUXpXH7Peb2X8TwUbvSa74vUKKRhs3Q92GRrnsZXMJa+h
BPGTkBWd79WUfOy7zi52z9oPHgy1CuSZ+Ue2mow5Q8HQbsqUtrYpXpjrsBJvfT5gZSFhaHr74ozv
2izq9RTez68ddUYn4CnXNFM/dfsn7mhsTsoyK4VsQ5TYXi+4ueAc3h6mg0zScQl1hqhSWYv7ifcY
CpyG5OXWBQX+bkNSpuQ43Ur3S37je71hbkNo2SJQwcpA9byY/OmRIEZFxYoiKfwUwTGs+XWIw8KU
9jrg/xBgm7P4ECx+qWbs6HPGj3f6uqLD+E6vM7bE/zRG4f7VEPn/Fnfpq3o1VeOmsn3wRzraS9S8
CXIg+iv0a9d0kRujH/BLGxr3E0s/yoECe5C6k9BwViW+H1NCduHJwGHRyc3RY0nrE8uoIo1QhDvb
buU8kkKNCy3XDmYrcnj4TM59r9/tl6P5kbY0GW34qrD4ZrlhJyaT9n4rvvFa/zqXCP4+m+PfSU0m
OXpK3RmVWKejhbZaXshukFN1bZqU2oG73KAvZOUCPc23v/7BvR/VlJo7VAnP7NsERJow6+injY4x
4Ie8ZDHibZZyAItyu74O7AE5/Mgvlzu1tZRx9Npvbs5PW0h6zNUKVVRN2zqBy8FD6otTWG5+q9Bb
BMEAB/I3QgfB6VOKXUn/Rl6WNx76gL4WDgh9oivIfm71O5MfPcp7RMsxxp7rpN3dLAXeGFn0sq6L
9Oy4qsSIeiACgkH5raUvwz5HJMTVFyYKwgkbj6eNvLnW235pXwKWmoIAbyKjGD4X7yeBeh8/Z8Gv
C7ow38fYft38mbf2D2YxfKZIG9IvKB/Dy7B+47wLgas87VYw+rcX0GGCmtYycLPFw9IuS/oHsm6C
eB+EEq/44XoQmHKK8rgDk1MXVF1CStkCZCgl6u3CbWLH1HcwrjvXdO4eWQFPIWnEU1Xk3xBaDYAy
44maLPEuB14thS0lNLmKLLk6kfpj7U64FNWrjYdhsgNcKslRobB+mIOSjycnV5zSmC2MSJOGo0qY
ixgsw+KkdagkHQGVahLj4OkS6OPNUSwDfnzVz66C5FMBmpoqooUXM8FABFoAcquyaUluUPhDM7pQ
xT8ap7vFRy3Jd71adxI3rjEM3ARUGH35Pdi5rGa74P1eWQnW6Y7WhOiUMuIkZTvE0WhesdLnRQLh
9tN55gJhN/aaQkLDGssZVJnvn//FKN32PxZ+8nX0sBErT7eQcFDB0jS2UeoHXnKepE+Q4nR2GUix
jzfYXYm9PBTU7pFeoPBqfgnLg9+8nzHuIVUcQMDgJ0TueJgHe9RNWmvUZTHWWJhh6jUBBpePyDkn
0rYDucEmHchyZppU8zqtjknqaoscUIKLsi9g4Xp9FU/SK2pm7gsDcScbmUCWTwj4XobFHX6OTKLl
f5+KUpaRxBzPFQgqIvgaHD6HloyNIBl30Ewf7Oftw0eeej1NdzI4qyA5mz2s1EfVrmh1ot7/C9tc
TFGIfuFWJf+r5NPPMasAEuUhBjHOUCSbfugT8jJNWOSDk7eSptk2XpMkRd9IKho7IA4TGjigSpz/
2oHat/avny46DjxdQfgZVq/lsp9Ot2ZV0zUNJgORYiSdWqUr3Vb44+12rlUaoOFzzEgkuwcz9x32
+hnp1LGjOujuqat5SbUaWNNRtFic02h8v6fgaTjJxn9tep32dIYJn14EQ9yCMqYntM3dC8YYK65n
zDUMwas6FlbXtXhXCJKQtsdsMZ8EBEnPOXv+JoPGR5BXtRsTt1Jtexg5mAzX9PnfYDDzhTgTfppK
/E6wuh4DLBO9z5zMWzaaILL7MDszWsU8QM16VaqRMTR6iwcPAT+LzHlH8Wq4jg8lEpVnNG1VkB4I
Xt6HIjQU/O2OaBc8XCCR/MfsFO5Xc9N0L7xDxHwFJFJFBxHV06pMKOz8UwB/ZhxXA4TNLcUCVHCt
mcYkBCiViYQ8wiVLj/WXAVY3+6AK/W6fP6g57n94Wiu7Nhz5SjgbQNk4Ai1Hb3FrW0OhMJ4EQPsT
Rr9/beHvgtKO9rdnlAkX1qT5MIor4TYnOkIBWMGgd08vRKeiw/Qad4br2QIyOA4e2cZutgpBtByg
cxXnd+BWqLoW/izrTm/hqmGcq8gBlhMYqGXS2Bme2+W2WfdwfXXE0TCDHFJvzH/zTChH3rLVvPZq
UoCoiZlleCNDf+ldJ8VwqiWPCa8OG1APhUhMkep4lRqs9DEr81KtWRzQVBb4DEG90DMOiaNOy4y4
gwuxaz25XnyTGFAw2fb00UbA+xNmxvPZqL+xvtghRyr4kZjQg8qsuGAhZx4dAj2JWwl23AaqrGLv
8aQo4xITc++zkyqsC6XtwdxjIGhdfTJcMRmYBufBSFo+TMO65WZdWOcW30Qb718jvEllHncCBaim
8woys8FkthDEVoswqNUt1vTHvDRIBNt1fsSI/gBuJJS7Q1LY+tJlPe7N1gwHDwp+lveDzgkEXQlc
jQt6BiuEA4Pz0Le/I5chDRNP26eYffPLWaw1U5rQT3vpyUyfNPVoBZMr7x5rf/Nb5arCKd3Zxi7d
9e43UlP5Bbul1cLSCpzYroARg5wYO1Vr81X9f4JQSxeNnIkCpL8v/mSSGc5BDpxpYk0R/hT/Q8Ln
WBgsYY9kLanVhZTeWv3RU5P1ZVT4hS/XBK+XWS6jDLz8blIu7p6sdR7wnR4ggT5B/JTzBvE+D5Tw
I8Z0ND0rAAZhz57tcpxqq5bo84+FPotcQEmFHY5QgXaQoxHTr2gkOOEmzQ+826MUXSfxPdQVx0mP
bC9kA74BDzI6Ex4/n6Vi3zn4YlZ7bpn1mvfBmcXGdAkoPD8h4g1+E31a8hlF3s/f1ZW2Wfj03vWO
JdZrvDqY7Bu6vcNCDV98Ngz5B16gkrFFoo7Iu7o19TotPpM1Yy0DxkKyBpLLJbR1nRBOwJm6yoPF
X94SdZjwKptLq96NBUHVJ40j06fet6pGFlO92m7LgakeONGWOoQ4wv5noWOgSy+xvsyXriaZtmAs
7IW8/qEmKrJ5U9nCaQeYm6ufXa9CYOEhBbS3wMgbQbUL7hnPmNL2pfWGxwXWlieIZMtsaVQQX2Th
4HRCsGxLb8uPZgYBqNUOhSzUpsQ4hLcM9bxAUG16BGhO/gz1D/bY74jfcVg6GJAwyI+vHBw2TMKP
RlPzdsX79uslTfecBWAKknOTHxfu8Sboewj5MelmgZoFlMrWAxGx2b8OyYdfWUdtl55fyRji/J4E
a5Ab3A667C4gUwx/XTOCAO3Mxn2GfP//aiqXCf1mNVCFJmu/FACkSbSbdn3IxnJ7WYzucK+R7zH8
Ry8tlGnt25uVD46ha3XiOzUpXC76o59JyKjBxWNgdOA0dJcX1vTraT0diebCSrnV8K9qPxBUXO/l
ctmY+cG/4SrF8YMoT/FLwMBNxIgbp3bv1eTpiow2MfoKW0OFfSK+ARKr21hmhj/cgzth3jMlvpZg
jo9qGKXcMlaxnIBGZHpsUvTkxKECccVXjZ1HH2H985KfOq/ewZ053GPmFTboZeuoYhy86DxcXmWy
O82KqXxCt0mRQH2g+TBAbnu/rfalzb4iOvO36PyOHa+xqlH0Zhm9ruRE6bWMH3C7Vr31G+XUai0H
Pfr1yuyDvWSjcur0zpMMYbsvAxnwHl3Qjw5HBlDdSg4V4/Ilt3q7U3WBok3zTgSQUppiPiWE9JEA
ScE4HjACy8gAQCMNnRwkMdh4GGE2xT4cQBsGi3Rm9cCMKGiMN7UcLKI0VnQ3oxnuung43OxXn1QV
ssmLjphVJ2+8Z4l3ONRuNL5FYlwmStVC7dwzL4jJGRulwHDva4eB5bu0zaxENnEaZrbT2qsehrGN
fHvvI8bzeDICHh7tSkkXN/v9SSVqbKQgtzhRMX90hN/KEx9Ua2Jrhe853eEOyxQsqcvK40ZWhas3
UtgzFQVyLAE7BJE6tUEGcLSLidrZvkE+58F9S1woH/jMT3gMoWaI4+wGoe0JjejfZbi8rfneTa9G
jOyEdA7/JWShkr9c/A9AW+hQOUVi4dtAalDQiZqWqerQ62HXwkAdMVZk00G5D8xkHYue+2cL5dK4
qQhjVsW20q185NbQCPzmilHZe6D39+1wVk3hnZfIMsSgaTQLT7XqrEWC6qSM0HSHIVMtVWb+qdRD
ofcyB75UZuJDw9qdXX6CX91Bx+jnrUwT15+X3ZCabXPG107hb5V6yq8i/WngyQxPlCx1+2iR2pcO
kkrgUiyZxM24eU6qAI/8clWns4RouwWkpk5myiA/mWNR9g0+6xl7opwVmryqLwFhXbs/bkEe4W1N
yd+DWqN5yNAvPJw8QJa9dU+n8BZUuwDibVPrwEhlNEsRykX3PlZq3OfjnCg4oieMDm/7GLm72b1g
ysITt1ah+QZrA630snzn9T0JtvQHFxFyOWtCd3C2R3gCn4ZUZfqRir5cxO+264nHU1iO9UV3vI2n
ELTez/5UEfMDh5Z780+mhuzUdLGGNGif+ORKtg/LsEb6bjfYuA7kr8Ly27+CYH5FZ/cqRswY34Kq
Dz3gMK6KBv05Bi0lxSRvFX/qzZo75yusW5Avybtt70xr3KDk1YkqexE3m4WyffPnX0wLKhKxaQiR
GSgZ/QOZDj53vAHyzeyQUrzHKfWn1HKxXagKYsm1EoQ/oaugPFTZE5YyuqDBoa0r/ZBD7Dai08am
/dsU4YoLF9YN9QeS7i9ATRhBM6WuAvb60rkP+soXWx9m255zqf+1E3N8d3o8aTEsUhPTiEID67Z8
1R8LAKPBjlVGVgFAuIk41KFzatdZjiPV5pEwBtYXOoSbarOgyd75svBYvmb7+dR0//WZJuPcB9Qh
Pi8KzpLTIb09ZgoWv16BDt4UQ2R6WB0+AlmeNcL9YG/e1Fm2iu6UFqrwR9lWlBSUwiEqH5fQlO+0
pNdUY1KEJjumUQ0QHzLg0a1ISu2CmaueuWJa433ZoM4p3k5LgKOjB9zYEBNEdEcz25RU84Ez/Mx/
TTPkQH57bvQP2ZiTyiJ5Vd3G9cVHLYzDm+aoFM19JiuvUkQqKroqKAbw5yzn3mpIU5UNAIP7zUTP
Jv4KjOpgpX4T1ixgvAtaDkmu+1evnvwGn07zszoNoGBW89A7959TZZv5guy6qQOXph64Udz9xMUV
iUnw2xU/H/PJV4rr73lhemsait4GFW/7wCfB6E69Slfu2LdQ0eKWSkvDnDYc7KXLxATSOF53kJEm
W5/eUnDpA9JmbXP6JBG3b0Z/tBbscwwALMh4/AqxVpvv45FBuBS+JCJJsW7Owc1cTFRL32Wcq/Mg
TlLI5FTyEtvfwF29i4ypPnc9uSrjb9LemDZs/13YT0/Klh506lw0aGjjulBvjKE/ASonG6XzOzft
iik0Ltr5yKgiBHNB5jI6bMJNGCbyNk3Ze35lRixmhb5QUGc/jXFGjrTMwh+gj+MkippZIwD7R4U4
zzOsZS/uQGuKG1XkkojfxRWjJ/NT2puz57nlWVk2lfnCLkUH0sFrEUL6+E1zSoQLScGZ1oY80pzV
5b7ZV53sLW6JSNIVY27t+OxXy7ibeWWuINHdGH18mx3XkLhuXmWaF09ZjwpLzMQaugigJE5BMoes
ycgeonQ7JIWY973P6JTIp/eg91lJIXe12BoMs5KgSkx3NGJ7FPNyv60L4Y+zWWGPXqBZ7fDW6nSr
xjRbH2R/9eDFoB4N4s7rIn1vb45A7QAY2poxf5uOtRr0gGohnnIh0TbrEI4PhD6KPpQNJwZjVvBs
FoV9IK76ZF6v23xxjKAFjF3Zha/aQuCyGEzJNdn8m4XOVlxKvd1wE2oYF8UKdhOhz5p52cxX4JaG
7kvoI4I56f3I1CnHsfn1x12H71lYLWFZPNZCCk3IiZWpErZS9odx/CMnNV4WIgxwyDFqqoeHL+Ux
PjW1Z3Y3u9d8gaYJT5IyyRhaE0ajBluRnwnd8LvZsgdci70ZpmKVawOgw/aNOgD086BtdYtkPPCq
EfdnTtjqFT7sjlR6Hja3TCL2UROr7vKEypJfNhbdl8eoEXMo/ab2ywsFUcCGN4qaG567WToCkccQ
meFsEP/Om73FmU7wzup0842+OhGSNc80GJgLMuhMwXcdsh+lpOEEaMhOKYar1eKDrx5+dLIL79QJ
+FJMUAVA2zQS3qeHgStRZuoLCZQrHr2SmIpJ3jr9BzhialKvDS0AGTox1P6oGzVaXz0tg9azKXKg
HPH+4UBSIZt+twxNhvQ6+HaUe18GkLoRSb127ob4gRn5pk3g746MBZ10XuG8+dQ6TQ7FvJ5jDCPn
geoEckXZA3Uk4928T6peCvbYUcNeAhuTx/wBmW0/5RWF4Op7TGcsU6IWoP4Nct2kMu334ma6VJip
5Cnb1F+Ca6N/gwM12zAsgFqf4R1y1xwmwdwxVJXH8zIxKlbUn9pFgkGMOrywCSWEl2nqQELLe2sy
7BQQSg92lwQa6oJK5MFmOXhJwiZKGlV+vh5KZAoq6Q6aL4L48CMoKphezhSXvBj3xs9r771vOSJP
HTDGJBrR9lkvLbyh0m7kLuTpjp4us0KpxFUnuWQSS4ox7FvjGMxWZ0pfcC2HkxGciUgfEsJn/cjd
IbWKEHJLMwOCGYtW2HrNzNraevbWTJYrKCyufPxgDQZo9ZxGdO5Y5fS0FxiKYsl2FhCxtFRle1fU
79bFFr0Ule5PeMO4ifRaoRerBkYbWqqZ/wlnyR8mKCHC4vpFJbngZ7IV3yOoscM85QJGi6wfBpdA
+ZeTQeV+VeMLqRfcIXH3mWrTUPcjFTrIbzH1TDs+IE7ILjH4a4oHia7Xrj0WYDmdIiwnfH9lCBvP
L/TZhNff4huBulkvjHeLhyQl9BGJqDuDzgL8mqaAX4xTgOWrlYNataZlBEddb8r/i2QJqA4EEkkM
5jr5SzIJyGqr9E+K89duqRD5BwBW4O4rvd6ffRBYX45AgCP8yQxbEwka7+oEivql8ao3QnrRYEcd
lVQS8xu+gvyhFCK0mK0edRHYaZTriC2zBMzF9l0jUe/89E+nQ0PGySm07UBRn4OdA8peGKD7E7sm
x5Pp0swRO85KX5QDJA3vZmGDA4FnSkIS4v1NfiWAwDlRHQKUsWdff+ECZGFKlEaP/ChZhgzL0Upu
RJUNcN8TAiMnMEBfho2gKz6K9TtziqtgXg2FBT0j7mKCBDMYA7FsMyRe5Zs++oOOXuzDzOTJnLhK
xUlOCIxKxHS/3sFagTUmi4A3U+mBFHAiD6WbqZLNtOYxmFfbqo7iXLWEe2LWKjWLPbVVbYVyYIHL
oyak5rR5/6wYUt5mZHmjkCU+6yBK8Wh2f7z64UlS7fI7EZLz8lLC5yjcR4H349R8smwYckK7lZ26
D1fo5ZX/ecJyqxj7s1w4Wgq/U8ygzdbpPKgIQzf2+bTagzt5YJsYZS082BtOzewCwhyCoOIuRQSD
nBa4Ad8N2cNS6XoCzeP9lhy6a6HTsIL7UhYW6kk+mN9SvnqU2cr+RnDj5T8cLTymidR6PziD2Mkj
XFUffJIkD6IvAhv5gHbedL6cAwkb2k3urgxQz6WnkR6RmKjiqKimP5OefNNunV/IT6638u7yThfE
+vdNYCOiNc0UqaV68LoPZd7MLfvebiKhpZLpHUyShjHmrps5cK0rJ1ymWSQl4W+mEEVwwq8RT4RC
g0vw8+Ona1Wz/FXLLFSOEGatmKnOdU+OXxruUokZdRmNo9uYydDpsMPGZu0FQVfspsauhWs+2odN
bm16UxUFd1E54m6tkyTSsRsahdWmoI4VSQTgs5ucw7ASrEoClyHBzAbFUB1Ux6lpfCCJn49k1MDD
I6Lye0wC6EBbza7T2cjDYSM6PkfwyAMGW6tPu9tJNXZoXHdCxyGxMFhWWt2FyLcj35wSKO5qs4fv
S7P2ETmJwGEtHYUeOJo+V7xRXTNFbHALq1goRJtYiiOGlBT4OQmZhiqgRBLl+DyvGGoD1ZFWz9L/
VpOLcCrRN559DyNcT4ODAD7hIqngN9XTzU8CVZyeN2s5ZAEn8dupRHW2vhUA5vtIASyqrHjwJE0+
Upll4y8IJ7hayv3nWfLhgIRTILK3698o3zCqED8dX1LbCY7XA7jymcmtNTUiVsCX08B7NTTEh3Z7
HIR38I9HjrKexD1VCEZRySLKjfxwUBA+Gg+HDy2gSPKIbJCN8qeiqybdFo87hIVRHah9dtGBsLi0
5tHk9h53w99t48bxvUIRriq45NPal7eSDINVm+3PMyi/3yTDea/RhRnDMTcvIvK++6AxwPWGh3Mx
7Rl2bD5CLJlct4CHfAQ3DKCu8xhfE7MJlPV/4dfSCZE74MSBRx5psPCMAPEzzek9/d+3/JrXw3Dy
wsk/oidre7dmglY29XXZ0S2JeWZwQKH9abf4q80+ErEDN+OKrP2xx8ZLJmLOOXOpUsNEgIMKsggI
+47CH6gXtsMav9YEZBFwofTsH5wl3iaVJh5YAhJOH+buujtuEiDbtMH+BV3xWsOjtsRg4eZnXLoy
n/paK+XMRgEdIJpQ9v/X0/ild+//flroejtvc8mOzFdP4WjtrLkeLbV7eKQvrALXsf3t/XFixZP/
HRHsky2gi9SnrcoF5593Xe+8r7MLb7D9tio24f3HkaMkAscckQHjCdsluceLZe8Y/tfQnaUdr3OX
AVFnnU/GK8AOn5tRhyGW7fCP71s6XqMjxhRhpPNOmAoc9dGPHabPYz6C7BK5QdqOefoPR4PVhWiW
sszNXvKbarB6Va+LkORb+zMFgSbhoeSBSZ3KZG+ERq3zBajHyWnlP3zYIkcWKm1gM/iIR80h1xGY
/mkAqs69Xo0IxqPpDE61jGDzEF3fEngGNNgM55+luDjhJuBH4hZNYDNwKuTd20e92TJiI3HYD21G
00r75IDLwYziTtpEH/4su522HQvaj2HZI0BmeoITWjohm9mZ+9o2EySyy8t0MW1dkgS7101tCYVP
6Mkbg2aTfvQA28JWYMY6CPuVDrXeIk8ywr5IG24DCUCSn/JbJrowHNNFfisj9NYbL0TnchPyZyEH
I/c5QDsd5xEnsDauE79AhnmQs3mho3ESxBer66CFGST4yrBNXlMWTUG0oUBVogyjgt/dR2P2r7bI
h0b9LP3IPV1re8iHOeo9LCuJzL8BLMyrn8HPb3eAU7Sg/3cUYHLxW6TL+9wX0Ae8MyNGikrBcJz2
8FarnraXMu2PABtyXWYZ8aYP2/XC0UirRW+zNvy4MutHX/U1eAMVG6tkyIlBNKHFPEursCdYHmol
jDay7UWdo+3W8UA7ECE9IhCNv+Qjk9BV5GTOGtqzlJy8CpUf3iwN4kw+nCc7WHg0RGUPyFzYaCvJ
nH8STtcucMKpPzhhM5S3z7WXfsqbBgE4k8ZZ2FYoDKcre2JmHFv7qchC/pbU5OEREgr7U0Qdvt9R
ykbIH7Ke6Qmt9QJeB+//2Y7YGzF+v9e0PsDfSRV/iZbtpGsDhkcmH4iVBdtqaUDvst13mRIEgtxS
V3DZ61ly29BeR/qtTqzK1I/r5XX4NlxPqvY+EJyyvW/dMyR28MAPMNGH/bnMH9kNg3YT01u2VnhV
uvIfFJWvHYU4uUGkqTm1FBnT7i/R2Mr09h/+W/qDluqomq+zAyQ0gFxjFltMyghftrqBQejyZDr0
UURniwH7YM4a1DRZ8b2rgs6TMXs+uHCXia7y7D3B7sHG3zZ9/fEejkOuMXGbiQ37fWaKa/TYGTnv
3M0lWEZdRvU+iee23PZSQquESaPTI9ZvmmyQhfJ7KAZrSV/5Ouw/BZtQsAdKBNvvFhaheCGq8sFi
x4LfkqEdsPJDuO5gINP4UR9I39/SGJTyZh6IyVASL+WCQRdKY29ELCiTXUFE89sZ1Q2Ikx5vHP9b
8Mt1Ly+YTRpBKtIxfgoTm6x6Fi+w5+m+fihpML0EeahgMfPDV1Ntx+tlZi1/KNblYyp9kDxnAlXm
JAb561bvQtFwJe3I62MfDzKz9rRUE0GZWOh2YtpbCHjKjFMSU7lSxf1qCA0kANfCYuCdqrQNuyWD
gtYBczSbkhjwwHdlz6gHN6L72/kVXfpw7ek6Z17pwHFs+04NHnlo8490JJD4Jqk/uoBLgpXTBzuj
tBbBSUBBDx/DfqCkFWe2qOmtCZPf8iiXff8wMqXui+xWskAeRlw+N9+L0oiz2lJXk2o8vu35RkJL
7nPyyaVwP4F4kiqnqciXfe4q/1jlTR7jDgfUGo2t0jF6mvxr2Igoao4OnGog3NIa3Gpyg5naLDud
F6zoWv2TgaTpYJ4TY4DCR2/ahAPwq5j9BEnSq1W+rVEIt84QGE2vhhEgSHSW5r+794BK7Et2RmzK
3TBxnAWm+PaXUDcPtHQqUhTMfvkLJOFYmKLWrMhKKKjhcqAllAdj6w61HCdSpIIV9Dcqf87+riCT
/9JMvoo8VHFGlkyIoLFTtXREb7Udw/oab9c39RbUMAvYDoASC+oEpl+Eo0UCjIp52kFgyq5bNvkf
b7TNfpku7PTOjjED+9ag8EddZ5gZ62UBbRII/D+2S7Xej1W1cTxqGyHR7pbqTGCvstK1+kKmoxUL
rQVHIfn2Wl6yChHaQ2KcVgruY+2Dl+6x4rVsol5izGpKXLtfALHN1dKQjxwfkeQ9bxuasE5emrcv
ZSP6c7x0sRPpyiB3VvBnGN7oehJNfChKH1wTIkRlenZ6idMvzd8mEr2f269z7EXEQ7t6HgI5gqMk
DilVDbGNN7eSMkFi0HTiIbuqAw9/XJMMdSopeSPoJYYzVd8EqYlEwavru0VWlpjbPglCvQCkFoaZ
iSS4nEV/MWJnvy33wW3asm9DChMeqbyf5KDM7S/61xnwx8Z8n8nu/SsV37L1Mce2nz+oxLQWNORp
x6zMYxmH4HUpiT+m+SKVWUaMPrqWoECLGU9qCrZRaq3fnnZCsLjjfM942MFkawFra3fVf/dmpZci
J8//sxImA91+7y/odHc+ezf04FBSXCDAY1q+UiNW/EHfjDTQGuFCP2V7BabDr00SITBkydGRAF9U
5/FF0yjgd5jRaHZ3ZWgVVJ740xo8Lf0rKOfRJ/llephtzl+ytNfuARzJOOf+YBmTCtMbOcymac6O
LSPng6qOTPlPvV54bKeceh65ymKRCKj1SonQGQKycw7309eZqluETcQKkI2+47nTHeO1E0k2DQ9P
nsx4TqqIWGWYf2vh5nfSGos0QSIYvLI2CTgVLsSGnoSl7pDYHhJiOEBnKQXbjI6u592qznJNQ9FY
3YYAYEzYIA4fqgBd54jWEmV7jmK6YxHLS+kyKdIiAAoaQuhvBoizCl9aZrB+OWYMdktrJ4Jgth/u
OFHvyGqOZuDY3vMu9VJ/hrwTAS1zWOUcHfJVvhXZQHmsYwBmu4FaYkIDPxD60t0udB7rI4MR927P
hYK9rah01mOW3utcDAlH1GzKBmsleNNdvEkX60i5goNBEsrp5mnljt00yL5MXioQUr/p5a2T9Zkm
SFVcyB+Q6A9vhobyphNGetwyC3SnNz0hDFL1Nj9o+2UfkFgi0Cv4YY1Oqd48q/qxsZlnGK6e62NZ
3yjzlPTVwXbFzu2JRZjRMt3G2EN72ZpbnJPV87ASc+xpEPjyCsQbSC6GMRHqxn6EVO3f3zyuhyUP
GPKRirXblXHetfaauTHG4awA6Qw4MR888NTJNJ2Og+2HRv2H+kiXYe7+l8wAXagR/OHFTnGmaNVU
LCLxNXzk1mIVqd/MhWf8VDf6oOmiUOC1oGrJJ4+rNLi11MkE5DywJWwntbJaDEiJicwyphDPSKM9
tTAA4rqvDcPumdIRfvRZT1aQlBs4f7hByIshr7f2XgfoseJwrpp4lScogr29VgxIgC6BPA6ygpMb
MQRmW5dT34ozAs/zdlq+PGboG/pEoubBf8FxJ7hAfmmJPauX7Q2SqASQ52F2cljXXaCPpB6QJvP0
CWqq8SzylwBCgLgiCg/gFN9md6XXIwxyRUL37MLqkIE9KdS04Mu2LZHQSj86P9pLP7QGF9Jx5n+w
Ukq7MmjLaFqCAD2IKre11BUim3LggGlND0hT8jTwNn8CJ0WaYa6cZlxbNd2nicsfPxT5NBzNL/LW
aqcboq2L+WL748jZdyaQPxS5o9RMRYK7D1MTuCBTQNF5j00ELTjPnxX21AwQjy/YkK7E/ZhbCDFu
pZYFZZbgv2PbbuoNWMAts4dSgd85FYEyezWZUZOEHuxhuRH+VmYHg4Mm1SLLc7YP0MSbdPZvPGmb
z8tBc4l1OGhhK7g97QLc6zdx30GAi3UbgJLoVypVESU+Ep7/niU2KGXotaVGbDTNVz+REObFgAMv
HecF4xigRDBwtLF3sh5j7KgY1eYnMSBpD6w9AVQYz3w61BdCOBXMPJ9bR478BFGvlouihi0GXXcs
imrHeKPlkomGYnCxVXFNh9PDXwr/MlxInvNnpRgwrUW2QM4yHfESNAAwxVYJzQoq3kMBLWRMnyQy
vedP9KhXUJliprGZ7Y9Xh3d/fdHIubTo45bWaIGbJCYL2S9Unn5pn3EX0j8XjZ8e9JC1pJAEcTKz
bMVj/a1Yc4x7OfwZAAe6phXTAvKvrfS3aKYSe6Y7kKvnm7s/Vm0NV+IPe86Im3wUeEIQx+/kYEnO
XWkdRZDLAat7SskGKeFg8v15hHsDpMOut+y2kUD+dETzJDCEGExg1uSFrsgAKmJYaaTb4+ssX5wy
JsAT5qXRAG4FVoSFYy3hzbHhQGOKKK1tCB25ylVjbpEwRkMctvSNN+dYOpH+RtVfwGt1bW6yOr6T
Q+0JvU3znnwlSqRBw9udfWokmRLLKfaO9VxK4j67wzuvouzMM7Z7XjqNPkbhTi0wOz6IMmovJHC8
TbWMkLTiJB3/fWPcrK+QI+HLebFgzrxoVoIhV98QjTdaOKzabB/hx6f5/cX5M5eWfzk5cpz53qSG
BtrdSILxcBralvwVUTmgPe65kObrIBJKLyG5tjOolNfXUwXTy+pPAJCHnotGZx/Aj84xOx8d9tI/
r28twv3j8CMDyRkc73lYnGZVnzOe8KTMvH95/pUpHfjd1iv9XKDKw/UM5ccu+/GzBeqv5IkHJ3U2
knc7iHhd4/Sdh1rsW4NvSmQZkmri64DzZTC3GN75mjMLIx7qjCQMP4tQcMu6D1h4JzRAMRHGQI3h
MZqt0iS5OGVqAXa8hYvgUUjKkoVCtPvKlRO/aNSz7rGMvfXn5Fe/IOKgTXFkJcVEMQkKw6pNzQzW
kBMz3d8Bov50w0JPTNRiEFBHauOogBTPKvGI2Ut+uhSdZIfZGabKRb5kOnV7K5JP165ih8pKkqDW
vEn0iQ1uqRSmHIFsK+FFujTwu3kZPrE8imfZQggPrO3ia6tcwjoqH/YT2vG1tUAd8Xetjd+Tup2s
CeeKX45r9G5M0qa6bPYFljDT4wJl4MnlsZs8x2Uq7pM+CwEHChWZM/fk9c9ExlbaADr6rGSAlXTK
u1/sdBPV3knOhTXG3sKDMN4P7zIew4DGvZlCxI8d2JMOFiiodYdA0KIMEFWt64ZCid5Hh7InjqYJ
sn3ClMPz6kipH4mc9l1qZ4ZqXWZjxamXfCrWPvQMBAL8tCDzE7GHv2jWEuCVDDxPX+w1lLVrwTTs
500WsFhanIGPc4Xilu+wufLiutt9mktzyvpzGy1Ah6JduK3xWrTnJCn7psdMAmKsrq3Llh6EmdjG
X8AaemVdVhexkT/YuSwPgIF02PKqwq9xHTErAaJb4Kab1aywHMd7Wm2xCMgAXo++jdsgXZE6jZ3q
XSVpoO4ciBJTJNGnTxSUCVncLhFSFYcW12LJCvfnk43A0xjitiQOwMxrWLdRrSLKx6VwIUrsnl12
AzW8zOkj6eWizupe0pmXQnnFo4AK7wjid7a5zvZPwvrtP1A00K0GgsuAOglwdDdWVFJVKjGiJ+6Z
5JFDXmUIdG/vUqvt1g9qwIUrpFQIZYh9t2DK/7GgRFPO5o5asTkAu3SjlenzwOPzVtYE9e9Iivci
K2sUT+bHIfQcPKRoK6NQ5Qqw3MSDBy1vk6wAx+nFRb4njtgD0dDhB0iTH5HPgtnaspcyr1l0HLCZ
yJ2iEIqAGk/QQ13JSWnCClW/9XPzvyka1HoCK0oWyuEmqAHwR329fEUDXLGaxTGTIqYry+X/yX2s
u8uoXuA+aWAb3p0cXij0GhcJRALx72mdApnvKoDvGleik340WCnAQ8X8BScPFQIkI+0QJjI0gNG4
Ez2sBb988jQzYnvN16uGi+LeMOeEjonnH4++oua1b1R1L4Kd5l6GhKD7HZfuEfV1EEUsXnNW9Nn7
NdSm8hHYSYxiInSFRiDh3/MXkHq232q8+5Hfk+J+ndea+MeI0b/HJF5hjjI0sLBSnhYBTPLnacKm
OxUjSRMANIXALoTcM2CgOtoCg+XgNJ1KZ3aKfpWCx5PPQlwKIxjMJrctwxe5n6yUptV45PG4pgQ5
0eDakwy7J6N47LPbf448/eb2zVdcoRRaqpaBU7iZMimOAe67TIjHSgNKU7xi2CZCzNY1paQkgLdr
OUAZVPwN4P+Dm7Xq7MOah6aC/EJmqSev3y7+rhB97p9xnm2RVOWk5hIFAj/QZLIdNCLGxR8O/LWQ
mR44s64WDuX6i9/kdIF9Ny6Y+/o6hlYTr0fmbBloqLzDvpm7fl1bRxaQ2NLwG0xfvpbkFLDXX3cS
LJ3jJypwmb+rtAO3gEfOjENojitamPykG5Sa3BcxWXOBHDOijKinY6cHUVDiZwehcG2/uKbNpH2K
ZCqV57L9976yEQgF1DSQ/z4opiei3PZa9Nfb24wis0XH5wWJi3e/M9ue2P8guiPvGTy7BqYlHijN
U/CsKZxWAHWbUsgB70yAuYIZBooKl3hEvuqf0ue3J5mfjNJKFsJxaGV1b0dIn8LRBaP+PtIxAAez
ZzeKJuTaQT4Voa7PkhgUiZ7V7EYb+gz7CTd4ToQ14XwzzcCLYzdI0TZzzlQeZwEUqNeapUCF4QZp
Zh4RGYKrkSTTIpSyX5qVbY4N8bQ/hz72M/gEpCgH86v3bq8fvq15d/83yIOfnk4S1+0YxFR2Hqrk
skzUCijUBV0HLilAr1q509IGaqb7imQmw1qok07mCv+DgfceAdBp+pSiZp/mw/dAmkaSPHW1k865
B+O8zqCq//Pe1V09AmKy2WkN9NMO7UE4Wvwcotmd16prvFoews7EEzcLW9NbFkeAYUWMstsRbSJC
QdNIRJx9SkyKh1sVwzgkgD/hWGpJvTJzEkD3Jvd/sCA2DeSSbDZy6oHwp/lB4/4hfijHpU6dydYN
fGipb4hkDyfdFHL3/OnzZOcMIwigTfNkazWJtqKjBEOT2IIT35vlmajP+mSrOh7WZ6uyYOmmMw8O
c+0/bKwXclezandkK9QApYbY68yl/Bw34jLYDO6jNmc0PYb0gvrKhKyvu5pXtnn/L8z07ppNCUP9
NTukg/bchCAFwh0WgNh2MIIDdwlooapN/RzwGXTDlkTGnRNc+af+nB7uBWWdyRYXgofqVfN/VslF
pUkBReURBjnGharvQU9huj9CWWwP3fjxXMlkb/19q1hrIMW4Ub7hnKXkhJeHmjREycWEKXP21ONF
6o2vEfN19H7i02EcLKmjnsJ7CTahrtWmwZEs33ysl9vWi+Q3oivoFMRhW3q2vutvWriElJlTNyzp
v7UVnfezR9qxxeD2TBox3/3B3CM2ufJdrXF73mGn0ShY6lswT1Abj1SmlyFsMYouRC9Zila4UHlo
wD2BGomcnDfbRA1RWV93YqKtpHdQjakbHFlTwdr7CvlA2dCO6cXs+7unxlV2NG9iiMji4mmKnGW8
NxvXbVRyJ/NgQOrt0mf21QjlYR3mB4KOv89eR6E9AGTgmZQRKaFpwJq0wEabkjnZaNUj8oUfZsVy
GQp6P70Q9VQoHzGWcJOa4nZLpiy+shzLsL+wO4TwpV0zv/S8kp314U/YzSxOxxVdA5pQoaJHXtsM
E1K4xHU21QvN+PKIXrDmKEQnhPsaVw9Hu/EdPjfHLtjobKPxbuRAqegHH9qPWYd9n10ntljVgpMH
aWl7qB5D+6jW5tU9H1lkVbAaUX2dszoHpLjOu/7HIW6wa0QtJkpiuX7IXH/AZ6epIze1opUzFPrW
i9gq6fm+2E6kksON4tuykFjx/4fY7mn9C1NsfLIksJ6UcwwqW/puB0mHZH2JaL13rD2SXnsSHm4e
n/uFEcq6G9zU6mFHwyYeo/Oq5d7o19LzcpB/Zyw2ldCbzFI2XDTtY3WbvVqj0+vgMMsfjOlP9eSz
CNIHxccNp56DZWLWoeXsKV9ID2r6PlYLNJWNR3Rd2A5JtfGTYIFYav9AISPFw6uOBpl27lWro7wO
+wzzBd+LLLmV/GuIJXyWH7LBeRxM5WoUi03EH7lZW0tUI1qvwv2gWT5bvWVvQ4NUzM0HnB2+bhGi
EhTs+jutoo4xWrpVaZH9x8Un0Er15S717cq/EmIo7EWF0elTuTN0Rz6qZWEypCFHk4OMO1p/T+BX
y8doXHgYMPR8Ikp5jiOk+kPay7eXtUnzq1r/KiD0tAL9mwfh+EXKOKnPt1VUH0GPUsJ9zcHZqDBE
tXxoOOVmXwF8J3W6TD+PdTiNlqADSFoD48qnUewgZIZklxR4PnyxM4hqsAMy6nzPMyngFLxMfON7
vXzUYypl7V+uM85fTt1g3PMWmYoNIT5yZUdXMPJmrmLzHjez5RkOUproxV131DCEk0rIMaLLJMjA
XS04vjpd21FRboyDMIHAvWCfe2JPQU0Aya0Hm4ROcsObOwKYYqR3W+ifac3AHn7xoiql8OizNfDy
eIAg9kMZBpWvqw9vORVswUh4ddLmoz7dVXc2iXMY/JwqRqDMRgjvN+BPrHcQnHEYtjoWuEbj82fW
/vC5Fo3alEz9kBTwYmMs/kiwdz3H0qrvTCA97jwLsAnBYqtarxW0/1ecrGsHySaoE5uyTrr7VK4n
qtRdKQLjeiBnCs/Rl0c3zQaJGd+nk2l7jizqgNJfu/dgpXZBXd/N9MIfh3LXb1hknPqNzB3Qi3NG
edQHnp6i2vegOPyWpwgJlIW9/EGRdRHxpesRcOgfVgjMmha0lVl7xav0Zb16P4SBMt47AY+yrAgM
BLRyBISaClJPupC9YiB4EnHaIQoO2gjeQEBV/tWvPvN86QRJVUBVzZaSAGohkXLMNTDzVju7OC5A
L7w7BH+81N9HhwKJfgGdnoObQrWSE348huGSBbqt4L9yaOkG9JZFxfEgqWTqpL0e8byCFDVeirw1
KalUSAoNQzcjNQPQ6ALsqQ35rg4gzuCSrovQYgcmj79HoXnFqLA90KS4SkJd5OsWUWzRWzLEO9cU
l+YC1ENHmLoOqmmD8BGeRBRkC37JZUZlWbq97uTDyAg9ZPhApVWPcCXwnYsVyVszzlGIoooDZHld
4S3NAu1LoYWkOBZ8ZXNbcZcv+Gux73EeZ4kCthKt9XJgQf66HVWooGL7zUZezzVCzXLzyrTojkJC
dKgJ7HEYZReIktvjC1b9fBJ6HQKeMN2QUWIGrRm926RIZYyQR3HNIclh2yNw1K0Ipj48VIiyyVTq
V+pAA4YoAGY6sTXTGUEd7EWCmGg347Codps8zJ9W94KTmM8LisKeRoxIU685KTQi6YONpc78sGMi
IvIHQa3x9k4gqVm3ArbYqvpq4bgoUeZd8AGnReAZ/yuS1YTd6AsN6mGA2NCTTQEi5R3F44CYxu9R
ACgSYkDpD5w3gRMd3dAn5rCnZhLa+AQVAey50zqtu1EFNmdyH0oCmLPxcHXs6dvQ3HGeUxop9l7q
TeBrEEx1ZXqEGXnXGn4Cnpik/zcn7Meb04AxhmsV4lm2Qlef7ik1pFLvt8uhS78OCwL7fdRiRpwY
i7km+GVGSUzT2xAhaLF8S3Ks1/ip9Yru/7Y+vjgzeZ7b33k/rihd9kGHc8wltRoy1kA9tCdLSY61
GvgabGAnUd+K/6/aYjN14cq1RHKGDnhyQ67oLKsoMw+hL9s5U0YIN0D6cjamSMV4RMkBmJL1DAmp
Ae100GvZt27hmvCzb0EcceRIgnUQdXef7aK2blX6opygZc+ICXfJhT5llTEgS3hBwnb+hpXsHqle
WO83csgpdU+eSs8B3cyOYqMKkg8oAtFda+hbgzm+UkVWS5FIMHJY4fyZcXTcgRGzT9CAPQfHIqHO
Gmaf4JIBULR8Za7WOjdjoJaVSJJ0l6ufSGCuhJeHJkpA6i/BONfei4nw5UwPqRgdVvnpf4pzcx39
rWZOgzSuyFwM6+1+xfUPEBoivBessMS4A4cJq7nM+tnm7WdC2qLArkYQD+pbq/yHdQN+3lh1BW6a
a9aqdXb55mKKa+gVA9WHtp6zM7mVVesIatjRiTyjPurKIK//98XJs4gk/BFgZGAsXRf0P2/w2hON
P5zYWKWqmICZ8eWRWnPJjKkJ/ctj4VTrCOsndr7C1po0mRXQl7EBP2hIyUOX9jGrqnPUWgrwH5Su
gIb/Qi68nUmxSaZQljAw/khsDqHPZSi7kfrWFGF+WKcLdDBW4pIVnu1oz5I1FtJiIsPu5/AsRrKb
oOpCjwuimlDw6+DV329Ei4w2jqyAJg1w8LEcxBsEgBEehJpzVhcebFNqrQ6oLrFGAsB/PNAnL290
/itaWP5RRFbdBiWAmj6MX/9x4mVV6eT+Cz0IK10v6oMP3+LILlgp3QnXoD8msLehcThTOG8Ho/MS
QCMVwOp1/tJdsSLM9Z6VmJQBCFn1GG1oPaDT/v1su0P2XMZWyvo6YmvKTGghWkSDPra3FBa/bTI7
ZEI9on/fbgnBriW1AvyAPMsrXz+b8PeLl1TkQ4uO7A/dmyVqN0gG9FknTEWHELw7dmjHoms47U2Y
FaSPY5oaAK9XZilzMqE3ywPtFWYsmsPbf5qtCrp70a5kxX7MTorT0SegJ6AAX4sn9PwxzG8nPqRX
X1E9qJzcWMKi4ZJhjJ4G4OXAzikDQsmeTFOSoQ/TmSsQnsZrEm+sSJU8zB+BaaV8gjhINTl3mR1r
7eG0D4ULJHjb+6IVRPXCouRdX8g85t2UnXfdh9ZnKvSE4a1u3lFHEkhSOszunOl3uDeimI5ENdHm
Ea2TTcq5LQ56lBGHsIvP063JBloNCOV+AZ+k0Q3Ffl1nOAXkLnwmM4FrZ2brGSzAOZiSB6aVxcXl
hyREQfRi0mR1dke4GYhb9PYQkBt6Oc6CFBKC7LLgPGcNdntkcAxKP7pknpxulogXv3NtSVrviLlJ
9s540bRCU7gEJ1A2R75n+/0HBV3Y0yLBcnpuyqCNjS/vh+HadTZ5qKwoYQGXYq0IShqz/RcmqAL+
tkv/ncMymD7o9Uf1XmuoOWpaA9e12efD8sNDBH1sxJcniPc8Vzs3Y3/xw1ZJVQz4HZF9bBuuqptH
1LPQ5cZQbm3cpU2AypDAHBD5pZUAEbbE+bmqxNDjMwSg9hGINRQdGT4iWXcOFEcTWrNd3DVoip+e
i2UIN1sv3BbpqAMcnbk9w/o3ZbaDTvxgUhqVlm+Lqcw0cEWO5aa3QMxjcGfTezPuHHJ2ykirUp59
AuIjvBcforTzLfBklWdknvwtGz54D8ILu/IY1et9Kk78ZLANuiA1t88m7JIOF/fNDX2UBVzxzOAh
0bDkvLRsFCH/o25tpVckSlR5J5qiz+VmJ9RmoDTWsHWhtcBRpChLM32D89Bak29f/QddjyJJWbeY
JX40AxTHoXovly6LlDuamtnhHPLM2cyKuWva7xw9/Xgk50KzTVi/vB7jNqD+4Y6HQ1637lrbwq42
5pX2QzunvXbIgeYKAg+nhGmuND6uoWHGF87ArWWU5Yx2bdARNk8nFmmOv7SPzoTGCcjhCOJDAN+l
d2DEjXye0Qw3CDJCT8+6yJS6RAHeL4PrvmCRIQOi1FdR39V/BJZu/yy0Fwtpyzdhsnpr28RVtFug
NhEdSgj1ngcU78SPQYZ59YNtyZugJRvI+LFwd0BzBPZ7E2ScUISF8e+eqXEnOxpYxvUa01RzsBgT
WlTYVABLyCGH93emmfBFaLk5X7x/00CkygfhUSP2jJ1RwXimCMbbHGXdoOnDOu4JKPd9gBjOkm53
vsgld6c8mPmD/tV1cXxLUjxRjUf8tfzl5rU/3cYHaqGGoojbdl3mtmAC7S2V2gA1+ohxTlEHVtSl
WkryNZLriXV8woFEa1gTd1XtwjdfCaaH0W59YflCLa6YaxfujvExyUn3mlKZr0rRymmi+HPYwvtP
nZTsoLs49sAgxWIfHJfJQ9H8WOO4v26SknrfE1H+IwXSMvfBZIGH806L+M4H0wwQC9n1WeVqTt3z
ghNUorMu+tGJJbKNSr+lR+ekpc1eu7kBOdftQrxZsf2XgwFw17K4v2RuZnMzyd3tRYgSRWYo/T18
IqQaoJ4yhqBelCpy4UnldzSDT4se7uHra3xktZwcTj91a37MqYRDfvyLhvfXGfvn0u0sJ/h5HXGh
SW57SSaM5d/2pwYUplh5g2/h9Mvbtl0J4pzPU6peB6ySpAiCGKshks4G22grtMyQrwrFecKrHsNh
FmcLRZvgRu2pckuXJEUhR5VfUeRTfKDTiDQYvhuJw8aVDMJIoj0pZzr/0OGiTsBMvMaxScu9ihhq
p/3vPHPSwU1QwtrGlqO1LUAlrdcplgihPGsG9GuTgLppeN2QjS5Ep2u7BkUhFQk0mOgWhYkCQwNe
p+bFb460uiYyYGtkEC0q39SSLLTcXTyk9ImOJxFn3z5SkNKENWhoHvqnGdBDLtDgOERX+vGsVEnR
MaAyHTFtJv45l1k2QHQmGo6xZvaOdIZm8MlBSI5NTRAtFdrRDrnbR76j+B/39q7TGodofv7OivN/
YeqZQxV0R5VjmTvphR/mrJsQN3G51S9MmulzNKFWyhi335e5w1lcuKcjdVI6kCp6cMqzd+yY2vuj
hWhvJgyjr9C2lp3VaV2SEnSm9fHhihuTqUt9SMj6nIzvZGpUfa2WnWJQBQ5Dt3jXU5kh9QNsOeh5
EXN676ShY9XsUswO/cuZnaso1KESmqiZmYwfb13DOEUlQ0aAAzl10HFPIPZImBOI1OUH7+rx6Dcn
Y8gLoIlvNFs87p1bMskilhiKsaBPdKoOClWqe734PJNPD5Ob3vqQ5e/vc67FNa+GGF4IXFCa68IL
AKnS7DYi1EH8MW1gff/IQcGTFetKTXA+pM0M+GFwwdfTmBYDN6TzOYPoKoO+FEKjTq096sxFWhA/
3oGaDkZfwdRFJxKUHwRd0wc/2VCnlfa+E7dV24d7WOD3K9UF6RA7wUIOQtb/2IIabx2+s9eQbvl1
942NslsV+UI+d4E/pq2V/AplRoivzKtc9Ltwrns0Gti5jNuMB7WBJBHl/MmoFqsSq2jDe+ivJ+27
6aGv8AZ12zi+VzTS9o/f1po5sjSoreqwpTnLYna2u56v2mqGr69cEvxsf6jkfp3kfMMR89j+kuqi
0N8zXpD5/u7F7Kd1rh2iwL77DXypcHG8KPvgsNbxOUZuHi2/n2EmvTm2DHMSfY1uMGEw4jmAT6Xn
sqsQfBS03tPGpY2q0IXco18QSEt4aBC+bZ72T8zeRUBWcPfRgN9SQQjAR4y7uYBgzzYqCBR9hMvP
MUdnpCNBWP4Dh4AiJUlFlIj8lYx2Zn5nRlngpWmQsI+nUFiwvYfHAY8m7BwcjAFEMObq7WDogjkG
WMYisF+rhn3EwDaJRycFY8wxWT6G2eqU+liyzKuImF9qNQfpmQ9XBKSomEpyPi6KleOnqpdt16gg
e1d+dtIiRb+JT5lqTrSPmJ+uQxYUe67nTmkS24nqZxAUOIETTYqlmmCZBuemY5D2Pl0oawD6gSBq
n4O5K995ivCyyxyB6kL+ZjSq73pUskAlv6TfSmQaPLgScs8TxMSx6BBAspQh0WQlpAEFSrEd7dSM
ddYrMUWNfh/qBrvPMbN51v7Lp+CgBkrd72uetHy3SC7/HQVWyJbkqWqW6fJofchOvCylU0DjiraW
b6iKYosJcWNbnD5+KbBS03gLxtZhvACBCJskYeuQlftTJooDfcSxp67PF9iZAb0OfXcuPy+kZftq
KpyrPyS096T3HJNzBMh20FpROogwmAF+0nCuO2MoiSb9L7ysrM7A/i+0IuvKvvXEVkkR2kBwQB+I
LJZpN8/D3M2J43mEQ5xS/8XIYnHZA21cCAk8+w5OYBA+PSsHsqhx9F3hO16jAu0yp3NzFYvlkwCk
0iDACgeSH7xTvKqZKSR7UH6B7gvqp3UiZQdRX3UBN2KEiROQGbKp3tPDUxiRyANJeE5B6lMG8at6
HfeUO/RqDwiIqn/DZNANL1MuDYMClFKasvSFNfpf7pZzEHYGePVIKeIq+bl+VjkemKO26/lQ1pAx
8z3EQf1y4OALK8/4lX6pImq20PZZS4quABxumvUkl0OWju16MaVBU2N3zmuX2Ua7nePgbSQECz5G
f0dk+x57Jh/+Or0GMCWva/WaasfYfiuFnu4jctqWTWlOOWk5eAPqy4RFCAzroakhz2/o2MjxSGLu
mdgnUjJwqm/uIVXsP4TCOcIm65hy7wBeG6MyRWgAiHcvhVKRP6ZAYgr+aj8fUijP/KgQbAuA5oGf
/EA5mSjai6dRrhHrHwmhkBE/lvlPuDzpxpR0ckvNE5Hw9Mf2tFbrAcprOT0A9QThcYiuHgbIHYoa
9LruWDW2MxbSLL7VCoAUXrgX9IXmPGpTpRd3C78EdQ6R2DMeIU/rvVPOOCkeSSg4IWyBUeKBoPui
m1sJs8DCdA/q0Nl6yonq7RaKQKYThpsw8fKim6Zl6AdFeFI0btgXepErGQR6ppwfFiUdQ5mnh6Sr
uGs5okSX4RH+6SQwY0GXNobQi1RzQ3rEFTM3jzwlUCKp0476ZQC1O8rn090g8VrAIB66auchQqQH
/DSf1G+sp7VHu81pJCGDqCcio3UA7eRNfMl5zFFXdl+NDnCGlXm7O7GhzaKqLGlvz+DnjJRjuIxV
VKfSbiCYH0s+15IsgGKbv184PIw+O9iqBLukJrrZLgeVGHEN/KftthmI5le3N+fVtGQNM4qEnGOl
+Jyy5Q6S8jkIyZZkLjbvfPvesbuEVGhlpMjlEckikN4iqSssw+JXt6GgRp1yeP46UmrYlqhV+V4Y
MsmfnUJ6gXc33YSDXm4IgHDagMGubaS13i3pOKfr4jEvQi29P+NQdbJPHdxm91vdVbdixHQ8x/37
/kwK9tlI7VsUoUHjXJKgTeDylV5Dhys2ZA+1ooO5OY3tXesK9YGJOw3FwR/QswjJazPRI+FuKjem
eKquUOdGARaw+OXFQdJVPA4PC+VCwz7JBoDWrAYKfb4tfIJniUOQZV2cfTGGxV4RYYBCL58RPPNW
59O+e6XTLEbKAnTpFOLIyMSJnpNaFD2F2r24D1OR5sfy/2QbkLF110p2TQNcL8v7wK1V/xB6t8PZ
hvU+HbqB4IFk03ep4fa8btcBWX23AX1v4ZxyR+Pq70UKh+jWnDC12VUaKyHjViL+PE2HrJlwy4Mo
PZiqQwPt+v9C/0QzDmmqur0jM6x+kzhd/vXfGIrGiXJTjjGmOjqmO/FZGb2ZLpDuPtBBlVV1KdDl
AJ2Si0vCUkQd6ZChAp/C5OdH/Hp6W+wBd738TXOsSuCFnENpoldyVAcL16iMQP+DayDg4hJ9+Lt4
xAqeYRn4zKFSe50k/kjoUF9sOcM7f0jd6/9c3uxFBCn1l0+IpqWrXCTMnQdoNRrMF1H5WjJi/qdt
cLrn+2tC96sgA9alDJmoImUjZ1+/67VLBrF4KIo7kG4r62HNr6JGJKmHyz/B5WFCYQLj1AMGLNtJ
SX0Ni6Yfd0XgIkb3UHDiDbhnEoU5QyjCrtLGj8lOFdyuN4A/Fs4Ret3suTLrBWXIM77S/jpnSRdp
dX5eEO8aRHEs+/ABq+gQqIYIbPQtPA0lgv3MJZF6iaYzSMRurfdL+uZwA/b1PunR/hHXHvDRIU7S
BtV46lX5/OX8VwbE/tiH6dc3m12T6i1Ep2YJjZgOwJEmZf4PZ2/E7wr/MvNVSFh+YxKeZ3FUCpbB
ELJt47sYXhy8xQLC4d20Y3l3S7QqX+Ghz8dHfCS36sYajJy46+gAAh5lHBlXV6zFfspuyLbSmwMH
ykO2b3Q2xqeZIkP2nZUTzVazn/SWOQHClGqUwfmPAue5nKDg0JmyLI7YOLCVWJ//+IncF2Vwq5pB
rtGXNw16nfKFT3UgHjURRkojqhFPx0M93KPzlFENbwfDTIaHBC6hc4Cs69cpF8YesaruAOmBq+P8
Dc64+chhTbm3W1vFGqbU2lY/K9HWybYtc9RYIlOwyLVUbfiKu8lnU8EBnoPsIQqC6sgTfFUn9U/p
nAM+k8ukjI4azkjWWokea/RcyvftwBSiW8aGM+q0/wOfHILZ1ukg5z8hdK+zv1pdLCXHw8Rrxstl
qlE123AAYpzNFlsVBmW5Y4z7qZoOsNmNTMmp/GUOciV1n6ZIaFL6927yEAYuS7bF+fUfHHdTsJTc
C+30UqjGhyoInY+syT3MTvqru7HuE35LCInxVGX1JiGIDonPXZTOJ+t+67KLqPDNee0YXzwbn/Qd
FmU1bNaqvYMYx1BWY1m1P2i07FzdHLI/8wUIu88YmhIA2DXU4NbjFFvJKE8ldW4sZqI5lZnilYYB
sBBR05NZRD+ALLNtqmxguEzb3rBJBW1ngw1ossbHRU0pNzfb3IgdmgYJTnt5ifi7LrbiZSLwrcGH
s52uzVXkG+3MT/H2Xgvl1a06uZfAEkOALVv49FVlztb98WdxphsO1wN0xCW5eBgp6X65ucg6Z0D1
RQ87CXRKQ3WcU29EaVX85eeJY2zqY0lfXbz8wdug5DuCLBlO4OIjRbUd8vqVbNvIPBbck5j7zLwa
76S13pjz3gajs4Yp8tMOdcU2nr53dXNzVk9OwcNwJNYWPsJcC+qdJnHSc53+SS4AU8n0NuCFC9YM
bUNOmFjdcLqp3V3x5hXDwgHaOa7ttx+pPmjxgY/1VN9nJierBKNZLYhjofLAxlMTuVIx6KaY9xIv
NbiGqGVYFjc0SxhKy5hjGhpvb/bEQU1DSGrmfq8NLtk75vsgg5ag18DVbatSMuSdzLFyVLQmv9Qj
DvMmQs005dBrHebtNbY0/tW9ZOv7e7z/P3rZtUTnEJNse00ykDtfFWco3NJkxc6aP6jxzRIO25GE
AvBXEb2AItPZ7XM8j5Rv7j2QsL0KhYBm/+UY/GWFw3ipQaUoYGoBCnkQeouOBsE0XE+4UExBdJ9R
UhZ+fSW1/5X9S30PpcadoVw4KaHviTFjJay6nEuPLjzHrQe54isb60Yrqm53mY37RoL/YNheWTTi
pkp1hIm7f4JlkaHFj5mSzPBehRTKNQPcJv2zbc+3sMSE+K3hOI1YZZa0whq4Q8cPcZ2R0utrOxQ8
KiMNk8P11/vHRneOO/umoDZ4isFKt+jT+aENIw6flaGnPGLCfFO566061mCJBVle8WXa+POg/ftp
EZZeep2FtB2KrYbngAX90WMG5V6ljT+oqLWlop0j6kBov4IM6NjLXVt4hyjdU+LOi/OIzT4m2yEF
z19sG5rsuVSJQ7MOi0yLaxfgHzvQ5ABPYVVLCF7jJaRCjm5v2bI7JmHPSeCqEMFyA2puWhqLrRob
BOsI45sGp/g6+pvLFqDSyTKAVJ9jqbQPjux1dz63vOuzeedjFHI21K0Hf2Bh6xrCBjnSzl6IlJ1i
nMBWtGUHpIOdF7+JQJrQLkPDNq/nuA1yu+xIYfqnK1qfBETXdP79QqR0wMvEOvnXYvG2DzUqVeUZ
q23FBrOQCm4ONgxkA4EkvYhRbMnS7Jtx+bhglZqSEfO9rAX6/mdQxbcvg0k1/mD2c96j5hOA2oDj
hy0Aqut4cwpDhIF1Vt70Xb3qpEdiXjzv8nFwn96Qka6DhqJWIb24spXL5Cbhg2HVDyfkzF++70Zd
kCj9nfz5/+7j+zQZ007pOupd5Qnm/ErmxM2JfEl1S5BGl+M0qZqPi7FGAK33qDtJUMNFmCV0EkCM
Gt0EHulKgWg6UTw+2PsZgj5gDxTyg0COVvCvQOYUiVRNFza0h7QsfmVB+/mhqIV6Msd13OD5SrWf
zZo2lLEZ5YfnADCAn2qQh2TzuCHZV5uEpXayItNPE4W23IsFvHHwARX7yqOtw+Ue4sPxWg9mcAhW
8ZRIMEcc+WNrnQpXeohV4tRQXYv5upJe+I/QTZTmdq3dV8HU6sn1UCg63nZ/cRepNrfZ6PH37WLM
DAkjKxgkaXL5iBHI56x0yi80t2SXKu5OSjNycF09dkYW2Wsq5WiOwqFGBasxGBmjOF9qPhZDJCvm
xyaJBPofC3DTjrut7phxs3hJEsg5ap86uacE5sqo9cFFyaroMucZi4ZY+ZSqVWet2ywfxqb1n4UI
M5y4/ZianJOAJviuysSnD0R5eawWiNMbHsNDJwrDvoBdpJZDTDM5ugqJzffM2eIDig1MeJEMRR5m
dXnuxp1qXM7blV6+ymUvYgEPcNozUSDs5O62wroFecgwQ6HgoOb9EAp2c2UBq1NZv6/mG0zLUogK
w+9TBxndUk6FAPiRJwRGPATrSZqhVPDHZtoO7smNQER8D5GVANGh4ATsWQeDPFWfqur6rvXPNYo2
YWKfKgDIwq1GDgIHw3SFVrTUtnolIHgsJDjxSyQu1YiGSojf18G0SrE6p8OQ5eCNmVCra97GzXzS
WfFre/O7NZoYJtwuLTH88xF/UEvxZMZeBahRSE+ZUpXZEU9G5fxk06mxV0ecUw+Rod6m6KMqtYEn
gu5HvU7oSOebdTol8Sl7xUwAwkYh8MxdDjYO9MissBdm/yNCR3kkCMA8VB8sCdTd3HgqZWhbgxeJ
y6VSOIcbz1kD+S60PPVOZvlosijGSAJMLz2hRCE/dZ+1ICI6YDC37MggTMjHZsNMH1GXZX41Iy7F
BsS1s4WiUtE3r94ZeRnkwk+6SDyLFRfxJnPhqvkjTYhjuKRlHtT1zcorehvA08KUTSC45dvvaleM
tPi4Ow3eaDPvKXzfVEkPRxuxd3vxm/0f8A3ZCbG/itGxAx6sO2+nZY5GYJnDHtHXjLIORwp5/YBn
JNGHRDBOq1Y1KQcMFgKze+Lq/tpvobn7vTG13VO9Cw7iz+VZ2ip+UVAa2divm5VwgqOMi02tuqTW
KS43UZmw4C2uBwFZu3hmN/Mr093kOCDC3EmYs/OLaghHIHjWpZd9n3rVy7jSZbAcvzgRPbGe0f0j
5caviz9VlJf+598fIwB4zuLSzRPVKlCX/pTUlk1UUHaIK3Uw2TG26eAMETzPNEO/oqYBoPujEXZ9
Sb5Aa+V0DGdhs4ohJdeOwAxBsuW8eW44jNXMh4oyZC0THobdohkQKywYbpC6pptcIy4662JLw8rV
vtjWHzvXEx1Ut0tKFz2I7b+xGv7OM8gwVZoT+6X4sTNQnxzdgQDPZZZ9jbsUgcQp5HUeTCl/UxYD
XoshIQpMPQr8yu4UWIYTihGPFuLTmfIYSnm9MyFZP3kgoWVMnjiYjTw6zrw7xCKNCcoiW+HYiUFv
m+jGjH2B4kcPxGEQ5l4Ozom0PCVoHXI6flh+x14KrRPZiGwJnPwZ52S0byzWu1z9r56Wflcob3kE
NqkWHYvhlDzAaWtHBD9WB49KG/NIGk7GTxZQ3FWB/mM1+seJ9vCJGS60aUYt+HYnZDq29ESLNru8
oNmPz+kcmYuxE/iiGaYRLRTEJSdPArrbntZRrP9nvbvqZKGfstHCvQVbw3pP0y+XSvyIDl5tT0Ef
R16ZhhY5kHCus0JLpcQDOQy+wJrqSPV98n2xABejvGdcfD53h1ExnyDSKtFn5bYC1ld7u43TByu6
D7y6FXcmENjSzJmqSqrn/5X35Omsu10SiuFNsv/cG7ZYsQUG/i4Sm4mC4VCG9/sJaJW1dcClHLyx
jGjhKKmNj0GZ3BDls7aYb+J6KJeled3TQVYPbiJ03K4oH/bb/kJvsthnFUH0+jiqbDLilOv9qDwk
ukUANV6J7Xac6xtPs0UUvvT4kH5q4Cw5WcqlQFpDa+vbXMCnN04RUz/THPJfgnw/JKPMRMhfdpA0
2PO80nVh7sngGj37ucm0GZrqs4oQBzB4GlBdBpW3rUKYbyPV/rzVkRdoNrd08ev/U1VraOnv/DK7
gRwrbIF3GX53R/ySfShEaQQU9KwmrpMpfh68xFub1+Pfjae82P3N2rEEqcI6FRGyGMFpNkNI9wOq
e/QV1GsMw0LLpa7tLhp7hLHgaWgVSP3AV3IAHamqqs4+DVR5K/2vrF7pcjXQ+QODlpRS3jftvREw
fmk3Gz6MA6h2jKXsLMFm8fZqn+byj8L5b9Rg6++Bzs3pqH8t4mjZRuqVTgjT9BU08qieYjhh+0io
4nyBoB0PCNBiw2/TcpOF9878llxzBfIXvDJG3Jh8OZsGIvl6enWe+AMTELgRtWm5Wwqg3KLPfiFI
QLLs3zus+3QffiW/VRwev5hNBvucOxQzSNAm09U0+5CWTemmTeUHSXcfuvbbkUmD5niGjAnN71wM
WEXaKAu+vB9m5Zdvm5BqUwzfdqb6tNYTuTck9uNlR7upAPFgAfYHAF9PCxRYjmMF+HLqOn3lztYm
mrQlrL6vziQx3VXhYspHtDghEao8+wDnLme1/jtlUg6VwrQMopAEXwKM2rWUojSyLHdNjfcET0bg
6GRKIICfOmZdn39ZtmuyopbOA8BFRGWeOUk+TDT2kxT7QBG2Lspy2XJr8Sk8yJ18SF1H4En2t2Lg
bTmJgwE9aaM7wrTk19OqWejrVwKbZW2Jq84A+4H12zaxy/rdvFXFzEtLEbCTah9lJCN01SHPKfqh
QVRJZ/6xrYaBY/1zh4e80I7wrS3MTd5B7PZ9BO00jUJqz6zThw8a39xpLQMlcjD4cUzdMI88SNVT
NYNFt0mNEChld8Ji5jSWAvpYt4NkqxoB9k+JXqKct3a2KSQ5CrnHqM9+CYTtZYP+aaGYiYDD+Tn7
Ue0SKhBREhLCo1vAIqQ9cfXcgGUN1JfT6pm3bsncCQ6wfCpMUvo/aWdKGrYCtjEaVs3B9MTMgP1f
W7L/oFKx+FmKE8eZ2E/8caVEJtcgc+dh85kq0nzKfXRPhC5fqIYY6kjYTDAz4HGyCyhnqfsqWJRo
t6uJ4X9IdpsF691Hczj4enr+aWMJjqNjlXuCNXCGfMsckrZd+ItjJTwwiv5dYutJ3crCwdf0YuoK
6wUfiqdrEst1iYzoaQqmR67wXYgsmBXV8EsHr4ncUS42ZYtfSRtWGAFq1RHQ7+87aJfzSycfKNwq
dIxQHgg/2C91NDlKyhr/iV4ruYxSczc2g1c2mf4cmTQcSeILyaCJBPOftkHNpDi8Ys0TeOmWFMzy
5Q7hIKwt47tTpIlxQqObGjFhw+K9vO/YIj4OCgpiJ4WQ9K2Om6FvfgIJkb4nLOQtuuSKwX0wYiGS
RkbIekg1fG/Qb0ZLKp630a3shmg5vEjOi64BsoixTV4YCqHe5x2VDrj6fzeTyrecrVYQzzs2Ypa4
bGqcaG3ufrooUJGMP0XngBgNsGpMQKMMDNPmBfrK2X1OT4XJK0qkQJU+6o4mKPJt0mC7pI+UaQFG
5GbMyRlqGgb7hdi6l5CnIubHmQ3zBnkRPpE5cOCp0Gn7z64hNQRAcJQrKllB5iCqqHLq7HPD/JjR
NybXaZVeyPlU9FIGoLqsrEDTKJTmY2jku5pndWdQ5GBdbgAwM412g0okpJBJIs0PUUZ3l5Ko92H9
kIdeldrNfd3eD/epBIvDXueH+xiYXJHLBs+POhpYX/5fur3DtEQoNoy5fGkRV/mo9qYqpH+Wlo5z
ys/j25n+vdKl3QFM5u/5g+72z9fBT20he3zJFtbTEkDm14ACPMqhCUCaWOFF7yMocb7vTaDOmawh
QXVCu4bO6sc84wVNCKexRbJ+xH2q4rxp1N1Ed2cQSIQvBI9fSO3rIKFgvYm6WSNGq95JLrmtoqzO
w2drRg65hb3aGmlCQO9mFA+JU+JNqnlWg0lIrUGr4prEzFTfkIeZq7p/90DARgT8bEFfnCprDygE
oKJZwAkQYDSBA6XQqjIx5sERqrPXoHCz3Gb1wBt0dgEoYe6zZ6RmEsqCl5SmVR/GzbhMEG7GdkC6
ZX/MNp8gMeY2gcZ+JBTtZdlTJM8Dq3SHfOv9PT8Vdv5uXQjFimAXS1jzjBt/VbeOrUppuw1PTJyW
veL1078iYnLFi5zaPIqQP76H3fGADFOT+WmSzGFD9vOQc30esUXvlousmcflGBOGeJcgXIsom/jQ
78Dz8BuwyWpngqqDh6bsjll38rU2SGloUKWiGZEPN78bs4z6MteYHuwUZ8s7KGCifJPTE5bLn0Me
HB5l/kzEdfWBdn5t4BsNMqcHYb2BJAGkXvXcpBXBPrWcK1ASv7FyDrPWtXyx7/uu3UZhrcAf65X0
6sU3eUlxImTa+wGShCSdLzm+vDTGf+pdtCdUobXv3GblfasgoEwkiRmJz+EDuPjAo4LFZojLDDfe
+1hwloIvgv9SC/gYE1hnp3AyrbNx5KkLqHEshblhMgkQg/0k060syRGTcj8yfb+fXjurOob7xFqk
Cu8hz/g6uJ+gVWsDWZ53zFvbgYjRJ4xyn7i6Spt6vkZs1qm3newPIGX9mYHcI+6pWqI926GrJmGM
0avkKJeUo379foOKOkIYIBn/AHo5/kGBxcFgEUVDXbFHHzFCyClESaEeLKF3AKiKk15WO0R5us27
6hl2zyaqf3drTPYFLtv3F9Q4/njbcpXwJZ2x1z1L0nYRZ90xT+Ul84n/x5oOWS91ceubS9yXI6Cx
cnRaxF75tRhoihb3UvNOYq9E6XxmgH+JCYXKbxMWV3C45ocRpNtd7dFoPTYgjdXi6Mr3ls5llILb
H73v690cF+hJbnbGE8P9j7i+77c2JjqjB5jASauF96e9cCRviRfty+OAdv/mGu7FsH59Vrxb7QCO
Y5IpzOErSsIIasBZyGBTrl14R/AmZ7BBA7TKZ8NiYuNYdDg6XE3LPIwhRR34HPSLGEgsfDWFT4sY
fbh18NHAeByatfLKsLGrRRcR8DTf1QN5zfmsReQCuLXsGXGqdaEhNgT/r0cceBjjvmwLU5jNNvl3
BLcCukUzKmQTnQCnmJVlwVp/jDCv8HVpCP+LesMX0JHqg9JdJh8M/WXHAwtP+5PYgFZe3LXNPWQm
iNWJZQoOkslm5cgb3aEHDco0BDxhHEUtOuiWDOJF3KC0jtP4+F6IFo70VP05iA/6nLOZ4qIDMgmT
p38XKtP71+hOQmX5zgRzKoonIFN+/nxd9qO0jnainQZwm8PoHNaJtSe5RudKoPUeGp4k+Y2Kb2E+
yelxfr0WvWstE2tzuHVYTXqXwVg3b59Pxepok8gNhp5MVRZI5iXeeoIjP3v7UnBo3DVVymvude3M
HrzPid2EPqTBpKy7qdJQHSDhcewZqc8hWmA3zq10qaARBe+FB9nyOmRvhs1eApoEamX+Y9kVA+50
/uIFAsifFbbotx5GpAF/x5BvsO95wrZZhOwhi+IXV+SzdYQy5wmbTTpzkTer2XFzQol0jh/gOHAY
4srWuL+FhK7h0esQ8ivfPpy9dhV62IAsxSGGBVGkc+pmaWycfsSbWp1mG1EHU4QHACsam9SyRy1e
4m3zj3987VeIH3RC0wyc5lzWef+cmzEUl7Q0TPm2Np6YurSgMTMHdS4dRxgBE3ttm+5qe1fGYVem
ulpJrlL/4RP4OZPiI6iVxQGYwkNIDIqGdrVyyBtoDKARSa5ujVbbR6qFHcd3tTMWqiFsYVdwIYYq
tkqiP5c3ILfr6FHt6N1ERsLXHh2aPMkBaztHllVmanMXMWSVXea/WZgU0C900DlXYcNpjnkK4VPv
fR8wFWuEcSEmvRs1coR2MP23uQHVap7l3dHwpc1ZUQDfayoGG3cyTbNrPKx7bqJWKyFu6EiAde9i
Wlp7ptD6prn4jJcI38V8S7ITuGxubwlQH66R6DGGcdgzEVlgwMyRyT6uIrXaPDcv782g2n+1RVm4
HnA/a85gHLbq5BsYf54ghtnlkll9e4AKFzLyjbmkrDAF0HR2dR/5UghmBE8REr0bHR183kxUJg/g
DW3DK4IOiVtfpeWpASCuKxl1OXrCnlVuohS31QjWuvtKYBRNgMdNQCS+klZG8k8cAb0YFHIuSIL6
u4h/1l8wWNALou29GNH2f89nhrsq9pUBLwaeqIecV12WMPX9BeRKbjS5v5Ah6AfWxvFey97eWuV8
B+BXvQTHp5zz+7+59VswdpmEsIAKRbszDXIlNt3j+gVIldW+BtIaKGbvHQfUOy64rnDrBMg2bRoq
RHwlQQJ5+egV47mEqEr2V8lIa6/FN5hDZwOg3REOWOxUuDWrXhfqgTKd5JIPxJwcDFaDSV2qxcb+
ZYkbZUhd2xiTH41CSwbG6vPPtgXGnXk1YURHaJYtGzMoZj+7CyB2WkImP5q9zJhEo7ogim0GwrKX
vZ1FtRcIDiDKTFnXiw1wo20cbj/1Pah8xxJqgCwItkEgQxDdqJ38HNgG+1YX0exFuul8e9PQliT+
c/1QZOl6s7ypujrSlErP+HIY4PbhIQJE7SS0ovW22uo0mlKHPnvIh03EUnS9gertPG3vh/vPNLGz
WHHqAR42GC8zPeDVDnVlzmdQRUsLv+gLfNB602TvHd65BeIxyg+pJaEhsbcMUztaLCpkf4Yb3Bl9
ZmiquI46yZSGITm1GF0dkxDI8Wul1oqliduc41qjzf/9kf2/TpkLMP6O2F4EwFGgzVxPZZXwJXwr
c6wP+yiQX0hjF6CXNZg8zVPVV9hdoqoUanDpYTNfI3YFuDvnCQB+XLnxXLUN3K47FWGJB8chrLh1
+CqBPHZeSMAHACEkLvYHdSifUFWy5q9mmSTP7y21X1uJjYVFvASglrB3XqnZVlyG0CN2fMa/Xdnz
dXb8zIzCTo2aPIyDQIGDG3xaq6/s+ya/CQaOcLRzg7ivjwpev8sX9jkTV6j8MV90//4IDvqOD8wz
xHc1stzNAMV5pgCGn5SXBsg7Z6rEE8GJSJAy7UN/aND+2kdQtXahXp0Jfki3qyHkRt0AgACOHe2D
7hgpEkQunBDe7nXdsFfdTs9aTiH8nojijl+DZZcIgmITGYvabhJLy1+emEzMTREukq2h8uJIAa3k
otf1Lp17Q6m+fsyuzspeY5P1LcjUfOpDdMZ9FvSi57248SCvLlZfZ0Xu6mtfsLkLV4m+9kX6+bAu
DoGFjI5pvJIyoPtgPIJS3ioppWuQRLqAw09WSTJqcncmqtdZKMEF3RKjtJY6KALs0TZJpI/sqs7o
gtzpgatdoAFAslqQEWDGZZqws6eUWQMSXqchk7G3N+Xa4hNBAXMa5/6zXMrRB7kSlMyI90oBksgC
5f0HcV6UFVagMKGFA55wSeZdWiQX3VRdcBPZjbWBP6p3tl5BvMTl9uaXRdeZlucrbPc/hHIsc0BM
Z2Aza/mo5q+eGS1KWZLL+Mbs/H/WV9pA0YBAvX/qrD3xG3vAReHgY4Hi+EcWgxZsyp1Fc6bbm12G
Ff/X3aixy6vBurEx+9ip4msRocCUD/PJzb9a/4bCfXZQb642vbnMY/zDlceCYPhTBu7FXFVdu5yA
seKHR3a0rpJev3orDvk967byDXUVu15xNbA2DlPcv/nsGZYr6zGob/x1N0PD1rWwWj7VrxE4MGvY
v4taS7tYryBzBP80agHkOoTBjlNUYNx8aE6TgDAuRY+hOYazpmLl0KmPTSeHF9Gx4ZrdikCctlak
PuUMgTax7CkZm3/SyIiKGr7yG0bJvu9wknDHbUBGJhbqD0aU1mfs7JVsIrun0t6JwFq6gGaptDdR
2Vn379xBb1EkdX2ZK4OVtuzHvDQWaGTh5tTFWYcDN5OvfsZrPV2xpwJukSc+hNtjKSyV8Q1Fb4M/
fHmch6yKPwzcb3LTRIxA4P1JcRfqWDoQYQ8oYpCdiHys+xLP+tngZLX+NFl+ASMyYXoj0nhmDPnP
03BokCbBjF+H1I0s6x1uqzCm8SXHPZ6CUNdOo/BhNC7z7MKtsSpQyDKdySNZpHy+4TFm/70VWR/o
htUSF7HOmlZIlewLe1FbKvv1sFGS3Hp4lOS7BD8KGTadJ9mtq7ZalVSLyAWunRj5is0AvZJ/+IPD
7PtfZEnP2ZJjLmKrpDr7iTvUM0vlAHoGlsfrWYYn7L1oSb7opCoDMdqFwY7VqKMz013Oo/oAHP6y
5Yy55kdyIv4GrTWmk5KGVbg5yZUcGxsxR1SPvivO0uti6ioWMF7zTtISuv83/q38iYGQmCfjTca4
YJCt6JQouGYMwyDFN0R8m2ftV4kd8PpmHStO0FhGdu6/eVtTBi9OIfnO2d6COegN4/Xr9No4g5aQ
19es/zAsSv32sRFpxVrNNTj/vqk143JIiXwq9YEnoViq8NDbGN+vRBS2tel9a7hpeygKIB7m/glr
JLS1yHAmLXfdW9zWbk93bFh8Vrw4WDsX+rGsX0mM7pdF9MUK6p3oamIm571rXCfEtQZqUiya4Ssr
TyQyRv0Fun8AT30qgWyvfeyU+wfnjGpj1RJ0AEwLFuiEljEvRD9Wf6q1DbBwFX63DJPHIsZItgaT
dppdU9YHFSBnv5y02wRxbCJ9pDk20PC48hrHsoK1AV5uKkahslFmYqwWNKVl00sENlRE2yZjKgBL
a2WO9S1OZPL0gUU/TQOtyzFLwNVsP9JbcRIHZMumGCCRA2hCZj9SlGH0WmOF7t3sqGoL0a5oM6at
VoLjqoGu/oGxThpS7U8TAmUcci2/1peuj10KdUl6s+5Dkeznfv3PddifmGijO/aePkfqCMXsOHts
Tq5CIXe/S+1CUy3CICl37DwVgCA3elpiIGoXs0/bn6vvy8vNnZYaSABvLBWMQA/D1+qcqPXlV2mR
IeBpbS19sQ+0NLoGE1PAg0Tdkv7qwG6x96CO+tgImqjPxjSQgsXHeCVqka8sysrrhjd+apIlJflT
4rw3XNZlw0eRwHoWM6Iv8CdwjIPYkOEQGdZ+Hlv4ENla9utGvN/Wf91WJTLu6yRf49shaLrNBGq+
8LBQOi9siXXC2sMTHf+4nIJMW3JAISfvXbyreqLL2XyBQ2dGjMspzWcIP9qddAw3LeKsa6RzAsZx
kzOLLhuig1v/272S/M3BCzxYkoOBa3x6ctuoSIDKxTzg1Dj8zpKmCXQTnYsAXsVfohDOVjPOxM+q
xAamzyCpFNRHxMe2mTO5jtqIqoCYMKPSzhejaR/b+LukBAjMalM80w1S9IgYvWMrWdgI5GcukSqR
pgbPUv9IZb3Blm2bPqXHdXj2TJFfv3NvgLEHv89Sk8cQYcCbUyNefy4/9GwbVb2kzn3t9rMNYUes
+M2QYKKx7wut44C05cqUkwUt7IS6a0k6edaexIQ8XvUwokqJzWKOXUN8YzsX28WIAm5TRDOw3Y0x
/tYyXv4sVLh6W1ds8VBei/SCsWksuy1xgy0SKrh6eCa32BF8eqBqIQ/7heT+IfcpEYKIMz6/7wyy
FOxEDwSIql7fKSS9S6FZUqZhIs0HGUutlMjeZR7HwrjJg+ZMRFyMN1qDToCc4hvgXC7EG8ltKVrP
s7AXBvBgKTDqUaOylhcri/ru3Hw24zheUEWvzrR8iHi2tCfn6lzJ3qLaXjuamBYtdwrZgJ8VCHF/
WTlqmU304APq1+icVMbvSVAgP0MvAe2ydhbAC+OonJNbopn9UiuW/raSjIK6uB41sVR2nU23ZH7x
t3qCKtnHXoq92vjb9R6Vb8/esYaOgYXtH1F2fQXfyu1tANCeooFjMQpxXu7ndsQhuoBxpLhTJRsU
V4pVnjkaJEU2yJ0tVSEWcRrd4Xh28cT0b1DeS0jCTaQd9N2fK+Qsn1GBEKuyjdD8QXiCYgy+jdi9
npxEPLmL9CLRN5CF3QTZCykEzty3GLyOMCCWMT89WCYnaV4u4Z20duXk8u65eR3oP1Xdj2Z2hKru
mrFSS556bVznBqGc4VREuHSN9u5T8+ZyKRlO5avDWHcI5y286JZBTeyiX38OJWkyxmIwrQMj62OU
eXqiYryoyw/0oq0dtDolgba6/zk20ZSLkgeWmVA2z4GAq8truEfOV+5r9FZCzzGRiAYzumNKmfpv
To0lMf9EOE2RrErDeDwZN+mOfMJU41UGLTdeh0MnH94xti0RGKVieUxii7bFABWokGrr1oRmsSx1
GMledmlcCDI/YayTg+MHFXG4aNCpcphnNJaDnh4mS5XcRZYFfmMWaUU6CjEDSS6TvNjsRTrsyQh0
sfUBV9fseTEJyEEhTvfVGRb8onQp8j1L4FUwuUCA+mm745vpyDT8j2VhmQJ4b22wb9ibt8W/c7EW
qVDO+dD7JDRNcggjY0vmYvS8IhjDDyN2DlStWp7LYm321GV57ywB/ZEpDn+mK+6I2THOflOYb1Hj
JaBA3q73bfn2ZBImy9NmsEmVarRArunz8fLYBqd+A/QA0+AkvsAFteRpl0vrnSMIhsf3a36eYRvl
ZWBCT3alDlx+z5i/2Ohg5x0RFSuwCjXctg1YSJTJoQNz2GGkf4h0vsiUOl6KIrZ6FwPrx6nLhKpF
tw0NRDemx7pzRsoV+mZoSIMi3cRhDdb8dvn70D0cgiGg9VtJKW9oL3WCTgrOvv25EOoOO0dcxm0R
JwsIvT6NTdlqpT+7YV9tcRCQ/nOzpqJXPLJHY1a1oLdj+RKx/uK5wuBqMa4GySxdN6PeSQ4Oz+B3
8mkLymsfDMd6K2AggOuvXK7d6SvUKdjJlxUhYazsoeFykdw7yWDJ3NU2U6u8fch74nm+2tkHFlNY
py6NAUcKQ3P10YMrKOjN4+Qksib3pNavsDpiu/HVucIf9E/hvD3ANSmxNFR/YUklMUbVbWZjfPRN
CAXF5JGDCWcm4XqSZZYtFx5C3/VsN2+EpZXlryB5kU/pBaEUDpjN1QdLkAXBBhEQyXhs/2kbpJsS
qEC09//Na8MKA6nqLVAqGsC4ZW8S/nj1wPlWYVGuOmVp+MerkEx+Sk+1A58/8CVsvCRMQ4Tvc1M2
J02CZExHWbev1jLBpJucFUCGhCMqUQgX4rjZTfpUSjAlbK2FUSZFRkhfNhE8a2Fs6Kwnwb0VAp8N
b2htXehuw766Atc2no82axxso99aUptcBRiBkjijEMdrDgrcKOvdWmklL1S2Gg0+PN48ZMG+/g8n
gFZGbGNdDAkxvYMOSDfFd/exM/f2sxzEtwtBfMTNTz1EGFyzQZa08hzOfAceWvSM3RuGWtlUUuJD
LWblg9lGYM7wk0lcGL5D5s5Be3LbG50PgUEYyuO7I8B46Tw4JKVIpeUuhMxEyetyWlPww15NADxI
8pHywH1d73QakVNCv8/Y0WDGsoLhDmAkCtLiDEkyEeyl9SKCGfEk8NvR/hE5kiMPBTWP1TcCNvB5
itqyjyQ2vuM9wohG5CbvZZ3rQbpi/4LackGHjk6mLkb0q9uYKnSW1Q9YD7klOAfMSzNWJr9mtNoJ
0aFvd0QtKyrdPvL3dnEX/SUS4phPHs+U2CaLm7deX5pmcNxEdc0UGbDWLdBPqKJR8IdLixQvSDh9
2JwOBgv228Dq8iKQAf6gwqQ+ktIVRMr5xQZGhWFLH7KRJzj0l/PWq1ViE1VAga8ztdiUsFjfljBB
FhC0WOHa4CihwWmV+eG+vJLu0nPDVYrDsIBYb+F/7xBfaAKmZJN4nG6lgSFBVzfp761n6SHQRy6A
/axZ/EBypj5WNbEoJ1jQdffRdvhwWf1Rw45J2+gaj9pVXfO29z/I8WlyGOKzhivSTjXJYuDrXoU/
I4t2naf+D6bn06TjQm8aHdBrWmfuqJcElf9ibFtUGbDPnFe6udYn52SxMBGwdi7xZsZqeDtH7xUe
VrKwKERfl4D22lN/CjahqIuhlTe31y0VQao4KcryYLSakbD5ILlpyI7QoemmxpGFbS0PQXxf9qa3
s8h5XgT6mxQta58nAtsNRAQkhURU/7ZqEdjoQ5WxGsroNL1kge+a7ZaNZAgNd3d+qfsuTp3fd1FQ
H7PbxaM0OhDCcalSQ/c21MN6iXnVJBx3TvLliEXbIXDQFWOd8/zqe9HA1YZKQwHeHr8kJj0z0jph
peUQjBPdtH3GaLuygHGVHINFE/ChRJp1Mwc11tR/ERg9p0NByoBr8RMfWIGM3AMq9c0QHxdS4LZ2
ynMw3Ydz/0VLCMTnC9HkezcfytCCnMYBXalyC8it+DK3EDA50zFvRfJEF0yNWmOzF7fHEYLdSDIq
q4ZRyYR86BydOKx/IqDX+VCgVAC+Dn6wqA0CVvez+Ayyj9F1Abm6T6sRGbVmApBHA23hJKlsbuQ6
wewCzxXSjugWL6BlCLgClTvhKLi9KjXAOcXmQbaeYhNjjfdfq+uy9rr3kB/X6rrxcCRGIr7RCav+
PXhIzn4fjP93ccg4rVmhUTuvuCpmvELoFD2IxrFbSAe4aKg02tyE6OjuWzixv6WeknpWlcG3o+/T
QFk648A/Dy/vYJZ5FAJ53W672xfWDcpJx0QC5mBX/qc4vMuxOchvp60klKYqh2Gvhu41BRpj1xlE
vbkrZqSHBRqswi9oJ+BA8SB1aKRaeNlFLDcjxBgB8ksdzssTCmoULIoKXDjKbRPvr/o7hjuyypgl
e/MciBkV+ru0+yVmKGXZYhEeCz1p9xQ0D6YQq3E8mmpqduQmJ6480ryygopc/zMnzSgP4cyUwAbw
M3TmYysHbKLSp0RBhpH30QhKvVkolASe0QDsLSKpzirzjzmYkjC0AJURZEe+zMF/dcmvsBdha3Nm
KqmmH6v5jMMfyREfESX0wBrpZyKHZRUtu3b6PzbOX6S9M/HGL2ob82EurVlCQ2h/YE/3cdp8S5YT
prXf9roD9orIa3Adlsel4+uI1NrEoY9PIq4CWKUFk4IH1JJ6ims+tFYQroPIpyIKCqFm7fJ7uILs
VEPbnlio//Cp6Bl5/7Jw+RexNwRFtdDjTVcMgRAzlw7AoI3w37i4oI8nBjLQipmjWXNCn0K1H3Od
ze+P6Jwl6cJDKZDrNYWynFvWtQXCX4KjuEuSJFcadijNLnmJzbwZbZWqsTUMCEDTMkH2vjougVx3
VKKXSQk8yaUQppPsJpTK3WYJvlqsj54gs4wdCP+SHmpUVJ2oGq1S2eqO5IcHfenllyw8v0Y1Inya
M3ZChVTO03KEmsEr9t+GONInfpuSuZBjDFelO7KIpCNtdNBJajcJ5yJ7PMwm+GJ0Pik42oLOGRWF
lHMOsYF/FLsL3OyOyUbGJVt7jUU14Kyzgj5FhrvLNyWGK4umwUlANpLooRi+ZcgfiRun3EdetBZF
JTj/OpCwOhQKrzyIEx+NndWgN9DGXP52Kkr+9bxUPcuXbErLhOJYzv15ohywqROG3IkXFjSi5/Ok
IDTd+l68wqN+iDfXanUcoz3qSGz/kUqu3FG3Jt5zbfrjaXC2pnnYQBJ6fJrIzkhiRdcUfTU1NOZk
hycXK0p1UgeGsYypeNQc2W9IKBUhNzRHcGe6jLs6DCkzHriCvJlzXcU9ID63rKIA/hpBMkCpDYdE
akbCcfc1xS6FzI+FNv4ezbQYzEVL4zNRkslh0K3WwR0c6bV4emqzi/telcFACIahJLvP4dsCrpuS
lipvwATJzsO642CujGyF1FSckYaqLzfZFmbDuFoHAvlfnV2VVzI9t+SXbClCUWKNHxDJKOoKt7oh
2ZRflXiPFLkJDnrD7CYUWY8npc/13k9ZV1EhA9jW41ehtqeOnFK56eMOCYA380PV/AQWuwA/+QgA
C6600LFx9J5Ocp/8vEUZzkH/LA7ZpWWXA6CC2+K6Pqca6Vn3Gdp5b3RkEHf1D7CdjYEIcvjl26v7
RC8UfNQJw0ge044SMyGG54wqtYe0FDewCLkoUeY+vO15myjdB+1lDvdcYQT5Sg26zQBVgqFlBxwo
GxzV5tX4xhxNtYesf+L3R0ldcNPPkPmamASx7aD86OGKKFhqLTx5gn0KRoPc7b0tibwcZ1KBU+8d
v0AWKDzSsrP75h9p4dfH4O1mfq2LcmSgsd2HdLcfbGAQLQwMqt3fNEKrIKG20k+z8Yu201stR/iT
TCg+NguAGt/UOknAPz/Lj1yNqUDOKUjI0FqOa5EpKqTpw7+Dxv51pi9UCiUaMsz3oTvrg0tqLfqU
8lMmeQkogQk3ICr9KdY9cKK3goGGdvOUVjkWNG2a4azKbWjDX6CL7kRg7tCsqpGeaN4jWVn65KrH
BcSLacTcGzpz5oiY9lrtiFJ6Ram5MU0GBXQ/WUyv2tsZYkgDn6y9EJ3Am+dkcgQfoaR7OINTmOYo
P0ph3yorxHqcC4K3uM4ANwT3fdmZMIAviMKJehTFvcRFtxLQbgOxtpjf9u9i3JWa8GHcj1mUKz4t
V7Hjb29MzeMSS9t4IQ6FfOqNB+yuPoTO7vFC+o9sB04DI8L0IWIZVmHpMuYILypEObLbEtafyoek
V8Cq8toLp9oULItWz7qQu5IbLAApkwLJLS2/5az8QuQtngd+U1WNEvUA067W28xImOZEgSB5+mDB
fx/UpYtng/vmF4sd5sRmvrqk5yE2EojVlCtp2J1QFykQOXmS2830tG46byDnbVQXacD27gp6xmTZ
Avo6YvjUQ1MPD0pBZRx31KXq4ioCuExmE1gn1z9lwbB8fMuoWsJ3iFo5FYU8UkXXb0G5eZwG6r5G
fvnW3BV9cwplT+2vKsxaJEQWzhjTMJVJ4Peh7TU8JzpgVBM/OGOp7fNP9Rcr+Um/UpxI/bHLFQ7F
mNLbYfBCUPgQsSx8iUK2Vc5OgZEFHENIsDJmkVQq0CYhpdiOKRYBv9Fw2xpfyoF+PlmmBEXjQU4H
CDEQfsK64BHyWb+Ew5AmQGEPfHFAJm6Y0ezsUAJKxZJy9CgqxQTUSxiyhhG2x8bno1f9O0+UJIWz
tNbBjMH+AwHRSJ4hMTgtCEOJci93S7ZnVGY3Rs1+PEDbzszvbPDCWauoFh9xlUZQw7W5DuzE/jP+
yLs6C2ochnu5NMTj9UZZa5FCDFHJGZfkCuWMMCWPgvjtPtrTbNoG7kcrWR9sKLAGJRHeMHo6VNj3
GxjtrfYQ14HxaaWhlSoJQj9sArOW39Lr+ogGHQ48AQRP4lohcQxo8uXceNB0LSobixUS59eYV8WA
uCEGzIQprnvN0F7MnJz8xmCvpiF2Po+j73PD1UFpOeqOGdgENlxBdLSiuVfmL3YmUqQ/M1Eos7Ny
ByPCGDxLq1y/zEXVdG/fQMeXGJRAI6STuawa0r5u1e7wc7eEAZ7L/O4eCqKGdpdACFrFQTEbxij9
XFPU5hfmEbVa0NQEOEMJMaD/CEFsoGUKV/VY4u7O9LDUmNIXa4ljlf068I11gZNTj23nEWxb6YSZ
7I26WR8xFUxHZXiX+1mcCMg0gNeAg5+Az1MNo9pzemR9JeYDKRpHbUNVfDxi8jSRd/yZmh6UsKgV
Ln2VHCfUJfayeArj8tBNoZ8qTDyUBSbkcJfpVSoEnfkDPKgIWGagVJSR3X62VQUMBJTFNJdp2Mvs
yKqeRiNlmTaa9rR0/k8g9cp3FpLRFK9SaxM4RVLNJfGVLnFi50iSMFlOrLKlMaK7LQFCS8fy0rju
BfVVkLket4SUC8k4zsX0H1pik1oapbgWnHOPlgYP7kdGveMzfe2f/MA15vQjBDrymhQSyPGDRviQ
WAeM1HCkdCSkInJEgVQpXT9G5GPBF34+vOw77Jni1GwXxrurgs4Hd03y1E8nCrJh7zchUJCWHjne
j6SmBv5hF1Nfd8cmNO20HLWYxt7WjrqmXtSlyU0vYVbatZMlsllqflRllZiAnV2+lbLHsKLV5Wur
2zUhHT3jHpLddqtIWiX7bPEO+VwJVEi9dttV+CxHDG+G65+l2YjNJoNXIybOYZHSl2UurJr+NX99
PAJDwcui/PkJF06VZBu/yoKjwcpps0Wu/uprMKGS50ccfVsAnTkvmKU8iKgHIBED2EH3zYAR5B+s
HRe9oO4kvw8n8wTl27ehBxGc3CcMtstCAhLqoFjG56uYMyEZ343NyfVp0RSYMCkbu1cB4VgOxjLb
RwjfzDOHz6ofuR75yLMtQkqHg4mbYOIrY2tOkYO+3PQsWtmJ7tzhEwdqJ8vCyJvXyzi5zaZvPRcm
U3IaIHUkjkhNGl4R2AtDCkDi3VdqjZ2UaNvQRHrxCbNVqKisKMFk5GC6TMqOvLIOo+oveRmaeuRc
8tZk3VBQzcHmEVaJbCe6oBgQZsfpQvUpRP+GPeGk5w3+1vP+n1xYNdcKPCZdFG/RS4EllzfS52es
Ms8UZAOyI+MrKQNVFfGvzkGU41CCAn3+Ouz7m4cXR9EZzFjnjsODMTDh4Cj5EbZoJg0pejzCsQfW
Ptd6l3EJpFr7DsiIo0xJNAfBKXCPBh3bJZoLTPiWcFbBZeRlB7oZ5voCwTC8bN3kW1cui8/Pj4Qz
zlqkd2AMkKoro7tijMMLpqLeUkZkgHgNAgN1eBqJXEh/hK7631KitpvtcgT6BFW+hqvc/LR7AK0n
eDsm1oLQ/A3L04o1VE3671aMZneNPet3fPvDwvidd6dLc1xc8GaDyjvLnEnUjTbBzLxT7dNsbcUT
N+rBqWQ61kRO5wW0sb2sjo+yVKSkWYa7HNXNpnB4RZAPzAdBL5/IhlV4ZrAKrUQNvjTxluQ+wkLK
91CeJBW99okNpYuo5ktnC3KANkTq6YJG0hw6C8Op50nHn38+XSoFOzz+LNDi7v8+lidY/FLqQQxK
X68J4FDRoICwTWlZTUjt9tPvJt1zza/0+cedI8DTAfz6BTzYVGMRIhQMCcuZnKWGoR/W7nr7SnLU
k8BIKrVuXrxy0py0s5P+udYPXAEO7I+4eyaKI8bA8L6CibkIeY9U48nv0RPM3G/Tir2K2RrszBTX
E1MuVJw0rxLq0/VGHlS8f61+HhA9t1pIj3rVrPWBq6GhG+NceJNo48HUKndCztXVYkatIJ7zHXUV
/0Yw2/Im5KWuEw8yP7sIDA0FG8QodXpL0c5KCM+7We80ab+7ebHnnJTSpoWfdq2RPlD21MCbsH1v
tFB9THiAo/jH0GBkVt0EV/TRXcDOQmsMl87sxIyScwXMPVicArqKoJ3c5fg2/HZzXy3LAtpR17rz
ifbvQpNY19C+JDEJQBtBy40BDR1BI2vPKKVtIpvmbLqzU3xVOOpck+YDEthMg5pjvnfYM23sH+6s
tAA4No4CEpKFZMKKf+ZAT053Orm3U+zVqka7FpSKMv/qys1t+uZ1GkqRRBf2tZWQyRZ6ZaeIasFy
nCL4W6sJgRgeQ5N8+nTpxX6ltGADfFs4deddL7J3j9BHrCLCK4eRrjcUFGXAmWm3tMZroy6NtQQP
LKELh3oNpeaSRU62BXYzrD7DJ93q2vyFNrgd0E3ACCgb1e+W3mKICCSlJT9XzPVdXsMGFrbWpnwY
3VmD0Eq2ptBp5CfjFXdXZZ2+e+cQ4QhyJz7cOtgdLnEsnC85YM5pL0icd0PPkm54NWQSTy6+OTHp
5ObaBy8HUbfHINVo/K4r6GquZWN+L/q1/PctdE9fUnG5FDZaj+xbFvaVRf7TIPbxAc5pHkdJ2/yX
axBujrncIieqgOnQw1JUhg9+WdFgBtl4jrNmX7IIhVzbqkoky2nOeNtRF659XC2esqSUSqN5N46a
dZkeh+sElS7sOsNFFNq+gVCADu46U6lXPaWmaAbgWTCahzaCX0orAYlVmwI8W9Cn5iOOaQrH+OOH
yzjkAjLzBldfBqKSPfGXVYr+WrnfE9kWl7UZf+paNrKcd14DgWDHoX11i7xNSjVcLhvkkqpCOvZ9
oHQ4y+sEI8wIII1tpD77CsaamfZ0R2leyJdyrFVGVRpJtaMth1fo3UQfCPypNXt/UdWl4RltKvAJ
EIR6Ks/rNG11jpurwZT4yalsyPzEu8SSGNqMZbV+Fenvsm9+gQGmH4W4BOh8zfo4gv+2Fc8GW7zQ
8MCQtvO41rlnQdFWt8JzU7XsDWIMIZ9kYI2tKey0tfdAow2mkBYYK/3Pz/wLHvx7Ym+fG/eePHIq
HM6cRiE+XFGcYcS+S02Nphcw17tmEDnbsaMVwAJ7EtTq4fgh2j6V/NL80pECJyzvzP0JvTwZbIo8
HJDNSaU/0+TyfuL7L3TiMbY1ChdvYlPb7oX6gcLAA06oNtdrAF2u1e8RnBLiMz4lFakrSQYh4YVq
0wrYCt4pN/1GReaNXu/nspXbYhqCC+oBWMbgpUCuJ/8IlyVkoG2L+i6Bz51zOjs0ziXYaAkc4q97
Gi4xi0QWSWY63ZHER4mkO3dag/jZ0ScHss7SG7/BvLdVHiELboaE8BFDz9aa+uftohf6X4vRhoXX
wdG+psM9FQYrbQT2vf1A8aofmA4g0woSFbTUt4efZOX2W9ly5do6qWRqXG60eT+GoPfHNYO3i9rk
EEEOyN4v9N6MLicJBbuZZK/1Qm8s+Z4mirnCHy75Rvd/JxXlaEMWUSz/oPLOav7BK1Kk+9si5ywr
eDWbj9QXNDQrlm1j+fWvixigQOciyaQg0xtvG9ARsGTSEGmKtV9PG1PUSEhUpGSrsyt925QBILDO
0tJgWt9HabXgz0BxW0LKhqm5W14QES4kLAeu2Z4gOANOD1UoWzlnjsQUIwH9QIXziGA/thDaxfTX
B/gNPabUVMq2FAwo6srQitYBVR4J95akz+QOLL4zDaPCSkcRvfl1FDwFcep/+VgLlJy71vnTdMW7
Wqg8rOwyfEcYCD9t5T/mh73YhUH29mvlzfYbfPejf9+Fj16ZWNBsvIiW4pwQu5ZjoWnfDXcZyzDV
HxAWm6JwmAVnRNjqpe4oQWPmFC7S73rro/FMB5YNgOC77JyaFHffTWBmEecQaaKjPQWHs4EWjMjJ
G4hLz0f9OrH3tWJkLOGIZBfa0qdVVQMFPbPtO4W0iI3AnN6ckbpHe/lu4B7PJIGZ85hpCYgrkBPQ
QYdyj5oMwENmp/PsBU/YQpOdhqjE56fFGo3PVYLDpEJgTUo8xhhL2PbkEdRt7E+ZzPIyqgwv29Pl
4FXSlAj9Q10nSsZtPebQ/PH/irrXcKiKMIle/OhyGzkGLoYJyH78bGkOGNqSGT3GF+GZh7X5f7rY
4EMQBTZQk++xTbKu+i5MN2k7Vu4yo6o8VBGkKHzf9LS2u4nKSWQd4z9laPrqGiAJ596zRF6XBEZs
qNQfMxOoem55LMTHKWfLCFsvfEctgmlgK6JvvdHYiAFkNGfJj+pCUZ4VqQSQAajAMI0JM35UaFjs
cIXLy4v8z+fVDFRPpL9aaIW+UKPLBLBohLd4UPDkpEw3KDFgoVS/BU1idYZGz600uByMnfGFDKgp
WXZnXzuc6S5/cRoIZC/FEZ3xdAulpRGbUtEwhVAkCijq7NKmPMHWx3Q9JMFI/K2mSYAZ8zZwO9QI
o7mRRHV2SXAZ4kcU4BnPKyBQ8I/C2L2RQSLbE2qwj45DRcW8KvfwUNy/anHlDKbTz3WH1xaP+y3q
4Bq1dUUHDpvxj5mue7BsDzDjMXQ1IX2Vyxa2WnUJf2ihYmC1gDAqCHigcL73Tl9KSpX1n5jJEnRp
skqtv8H1ZpnpE/0Nwtt0mAUfXl6Cgyq+4/+xyghk3peOzBfFDrUdiXyMTC0uF7MbLmP9L/ylf+tP
+MGqNxcyL6G/36Q8aH68GC6szMgcAQKIH+wLoKdSc5jOqqTU4qDdjs5fCsP25t1gQQkxVSSbNM6U
FEZNvViZDXIFnotdwiHBArLj7JahmlsyWmhT4hBnU3aHzimmwpMWh0pZbCMJPI6dbHV0HSI3C79F
Y4ILfURu34qGuTV840lnGs5mEzGp7GrNV1rvItqB5laNTSnjTZBS2wwKkn3j3Z6pfuN6mxOCdabB
xOKOlvJsdjMNOU8mUMv/9h7s8f9XfyDHp0T4W8v4NWMv8emKZTNwZvza38idBbiW9SQZDKbUzDej
lfAftuC6czASzMaLSMGLB6IE+J+d1ugOF+Kzfy0epjgJsjEk/uaXTH9sjEbYZdJp28R9DspzT2DA
sTCCCn9VlzpTATdHc6SjuR6lA7t+4Dczk452G+EOKeUfgpeUUsEuhU0rvxjMMEn+DbsXQrvIbAmD
tYeUtYeJ8Y0DWIxQ4dpQbOUtX/VV+XdmR/hxy628/7XIWkTcU9CwwWZ2XIMyjbjBk4sPJYh6OYZy
9JtT65Icttgv7sNKxQJO8lNGS2vXFCpHGV8yPSTWK15mkKWHxPFh8Zkf0laGiZix8HZQvjc//JDh
yq0LVjaC3+in5/vNkJTEyQyZBNBz9XpmpFCzVumvfSoC5M0WEsMZ+Hl0kH3ehDeccp9w+BmD67AD
L+u5RrR3Gzh+R4e2t3fhB9UeOrBJXoPPqGL0WLKbvuWahnnboMXzdWvEEiVHzjqsrxjorbXnD+Sy
bTUz6GmO4hkZo7WZ6TmteAcCDyIDo79J8ikME6BrDNOGL2imP1FC68n0tgYggHp143rHVi3udr7D
WYk3uVJ0KXjkdRrUQ2ako9HHzZVFPQqJXZDGrkbFJm16kM8QRQl3DGTNEVKdTtSFQd6A1jBD6VYh
qLV5Il6TadV0VL6obSW9lkC0heK7QJ6531G0SDS7OlNWbze+tM1fqsLx1opI/M1BBLAsJsLmDRZO
xJoQJrlzISb9OnaVJkI1HktUAUk6LAdCkSKzFbjMB6xciL1uT3IwW8jEUcK58VuYJoaJn6j/L409
D5MDfEhaQiW2v3v4gg8IV5n1rBfhZjdLw3cjYvVnBh7hHtMxxIdC7bprO3eCFgVsjPxx6LNiCE+K
umXSoBPvB+v0V8mOKs8ck4y63K+gC8BoQ/kxLehCGHm77RgKxiY+1FCf5fgtlORPIhKdMlMu9ncq
3r33G47UtUHbateEiI/7QdLksbI/J/MJLT/wlBsmVw7x0hdcJPIyOW3jgqKngLP3bjdzKmoZCxOW
ICzRSzMREG59PGzBvyFGbLA8SXcFyhZ71g/wwjnM9jWHngToA3EZAfXTiOLHUSZD9pLeuZwFfhdt
Bn35snXIZxnzVMWHKihbkSG9CoXP+7PUTNO1+XqV09vdeVvoDJhSKxfUB28a53tUhG7cvJG2E2Br
z46nORgp+ChlcAx/w4kNrtSI5qIDPMh24OnYuKkaogcJRloMuYPC0aJS0NNmSo9jAEgL5PP2SNCv
+/vb6qxOoQG6aKbtTjxtWaKl1hVYi6rF3Lo7PTPhQ1ZZMI0NiFga/ddOMwLvOS/JNTxfKoj/dsxz
Z+gvp8kZVEhM14uJGja6q/1iuOGS2LDRtLytlfqs5pkHy44Rpyo/ZEW+sXFjAsdn/cpUiy6hW8+9
1VON7gnic6PLFmYLQZTWOD8oeVV355YRWGjHFiV03gWFo4g7DGd2VjbejyjlhXE6ErfhTIAB94fE
AzxM3x1f7AOTRmBn6IPrEnBs0gc/39/4kE2riZNVQlH6LQHnRPFfA/iqeoqp9FFNmtYKu6QAp17h
w3LVYz8tqsmnzq0GEFSdkAxrxMhgD7KJQIPF/Mylz3iI69dYritOtfY7WDiY1TWya2SoH/SECfjN
Q/ZZClAxjv5PayoLyDtifQTyQSM7kHNA1KoEiDnrOYViL12e8RCiSEVf8fVSQYhZ3Xq2vx4heGc+
zjG5hiRQWEhW/RUtcgsAi+dMDvYH+nhJYqAi31qsei5kk52RyWcPQYYY9XfdILMyLmzxJ6ZWJn62
L8mIH4Fz5jw/qHGMqb6402XumlQlx1L8w+s0LuXAtQj2X4I97t72cO35qVRxxIxQAIHRSVsrIyJJ
JqKoDjIGVXQ5Sl632GBGoZU/mvjBiX+F0RrpYTPJE5JC9BGbgCWQ0/c2YpmijzpbzEBWSaqcfx+2
ukSM0JOw4qGPIOe68mG8pU3A4nWKDclewxOr8qan/T11xsHxbkovjHxb6GB7S9xrDP1/gq+qBy/4
6tlnN35OuF1j552DnbeJym8TCdnetjO2CNdvbsJ34MPOsuTDWmj8pv+Vu4vw7lVqh3cCI7UrkmMJ
cH7V4CAHh1YLviwYcXFLFjTnFc6vwIRdCW7ZGcHrD7NXGStjGBzSsaUwHtSr4M+j5mEgXfJzXEm9
Cc0prSXvv/xGHx9sJJ88LxA+i3UILkQNR+9JR6DoPKt4A0y0lJWmWo0mLj3lFLtQHQjm1isfPut6
qKUnYCQfP16bRDM2Nt+T5fl0fxl0XfUIodJWjWyxhXpsU9cm7Z0hSwZuk75xe8A9m9NsjldZ1kjo
htQ6o0mr1jtrlaNtxHgQEVFxHCory+5z/I/08ig/uhjMoHG1RboxM6Ma9xTMYjF2UYASQuVu+AAV
7Iw/2G4mbcb+xUpw7LodZfYhl3xpYpYTfdGsZ5hmqaLh2miFfL1vVuARou/tHByfXuxVcYS96Rm4
mmzycJ1VUR66UZdVMo71+sA9MCGsonteszjRdad3CWfJd8wbCJEkcCpdZ56cpWA4NgJppmWueMOF
vk2uBC0YMvfdug7wDYqv82pvDK7IqEg5nt5u/j0O73sUiUdiIspj6sw/FtoQwCUpRlxZXJq4Mj1b
BzC7Waa28ek1MRcbQ3HTwswLp+9ElRcJWjo9za5xhiR9SjAPS4goqwMnF0pdsvzMPXPXXTTydWgC
rGrsRSeVJZ3sPLVStc/vjBaKC9MXTpGzeoDppy7cQDFudY0YvlowKwb5vMmW8MT1RHJykx+kMcg/
uBm/GZf/ilkRrXkZhUcwrt+C3OTLoAJyKmTUHAb3b/Z6FNcNDRsUlgdqhRF/FtVhuD2m1gksr0mA
Pq2AC0Sq/iZ7IaksMeTCwb6xYLRMnKWwjAI6mPse750PitHVobCMXpVn4Bw9NOUahc2jzRz+bA2W
AdHIvWgn+EqcOfQpbyAso0Z01IKKHeyPyHTfpaf0h7XUpIbjShwRMWuYqgRqp5D6VIS9QVt2TWQW
g7fQgAT2vsMQo00Cq+tiKBuxcwz05n9d5ZSViO4uI6+l0LkczYSM1Nauy7giL7f20DDi0sO92dqG
N0eGI21KQrW74Sl1iLVDRMJa5uNO3UxbKIkxfJcJhT9fBQM+5lKvjL9E3khZQmjhm/ZWTVIqqSA3
0uPu92W64dJcAyIFknVgqNv928v0TpO0t9a9/hcVFdq2RPA7PUFtESgimH+j0c9ZzunhHwL9Qkvg
n6mZZ4kYtM2f8jgklJ2ErjoKPiv0ohPGTjISXIsyFrf4YseArH+9/eTPi6uCh4AsJ45W6upfNvM5
4YdQPGAO38suDBYr8GGEnzEvkBDytntuVxek+lw0dFEnF8/8cT3EUwl171qs+DhjHbf0IXC3Oudd
LTciUk54Y58wkf0uCe9ASNrsNaW0fOTZVUX5/HKORGIb/A2xYVplzfeThHsI/R4nZKMgTw0JfqVQ
MybP5yXxhjC4EL8IKELDwP2X5x+mof8ReeRJ2LAwSwsZf+FsrzQZ9sWmKdm+eXoERkbyEiufalb5
E63g7NRezmMwJzC2EhPiRGQwd7hYb2JtY6Ghli5YTliqdJ3rmMYOLdJUyo8EGi2JgtjDyhjOiH9L
QH2vHNh1hplxPtLyv0S16Fw6I3nrfzZ4kf3nBFFp1UtnGhZmziYzkWQR3bSnxQFRiExhfJMvDoOe
5KVPHgZ0qbsiSb+1N6bvnCJiE4CW0sl/BuyKQUc8pruaMMTdGmoIAQ+8kn8h14z/5csGSW7adRAk
ut1CtEVer1NiJobYCEqz3/abWtcUl5p6Gz748T4dXUl9+eli9oGAZJcCz1yfc/WN0o0xewwyJ5H8
sFzj/n1oGyOgheMY9KvWIcl72iu/dAx///FPW/j3s+c4COQ9VniKP+TwKY4PtLPzgV5lt/HK6T4h
k2Gn9RZfGox6/WAmcKZc8TSz3zjgwrWb1x90qb3hqegBgH/4yBW78wZdpM8GYyx2VFTTQsQU74N2
uHnvLCSpkZDEKyy3hDwyzxa6BXjlla5bgZcrvoLdnk9tcQqYz5SvOuWYUukKtFnOZQj4y/lqKNtK
J8n/cMzARIlUCvgRRUuSfy9Tf2sHRB+qf5VUvPQQkz9B3iNfUeY7r66CB5gkaWk0r2m2xUNx1D8B
UCCERzFU8+ylXXLsozRA52UorprLiDcNNMqSDfyg7LpGIggPYoFkKQHt4fHBlrJEniHwjt8zbBFW
N1if7oaDKAk22oowSTWIL2cjlhBWByl/Ht1mH8PJ9Zt+3QErsR1xy/dZi92BnD5zUzAQ9yu8OA+R
OY+V4wJqVI7o+3Nd432zXI42fGtbdmHWy5Md+H2KjYOt6B4JhhQHBvsnco/tqGAhw4Nx3y2Jx2AX
Jmq4psJkMj6fjCGkJe5OOEveF9Kg4UeBpd+1eYrXpgyqgDSWBztMzZcaqGB5AlHcFE0xM75705Wv
dMaj4ZQOLGzzPcoug3SzYWfYb6Kzlq0MZ1x2o8pmLY1eYMGtdsVA2IA9DUIbI6QEy5wuc9pB4fYq
3LBz68GlByaD2ECdfAVoyWZjBYrt3eMwR4zSyXas8b77gTL+Uga1nX7okVGJbgwKO1YwhV1ekbg8
A5DjE0Tnvui8NbLvkc+PynOhD/NJB9IFjmaavm65GwesU9ZCjHD+62bbGLNyn/C0w3uovVh9vUCk
PekiszkWX40TilGAHfqU6rjfG9wG08b5Poymy0AhEJ0/haU41+d+hY9CANgquQQdUsBW4Kv4CjNp
AX3PdbOp/E97CIrk2rFirZ9a6E+lKYWw+zJjDxrMIjNPN1aOA+iJgHLfDO43xi6AFVbt9y8bNAHC
5D0rmCa2QoDDYaO1T4mmqZUVPbjxN6plIkO9ljYKH4uNu21G/b5IOQCJSRzuPsAhgo1a2/jQdDtP
t6EuxT+3f9Gwkk8rdbf69AkpX86dzM4aG4tvu1WrZo4G9PJxBaIxGUVaOJcOvDx/oJkVMgo0UIn2
D6c4nCvatIXxj06n6L9bTd6zfN+h5/aXRfkbP7+8JBJCiq6zaNzMT9fTnqJU2/7CPylS7cjuskwN
EDC2NZcHGd8VevySggwVpX+2LGj0BrM+v8TP9zVqrBfKxgrs+LhEQv32NwXLsoeRGV3R5VPUseH7
A/Fz1TKJWw8yKVI2tMZvsD6gMnRd47YNV5VVPVU1EaZ69dvQOeW4N/UMijFhtSsI7Sjnpu2IEmgN
BVpwjUTUZF2GLrI5NNGo23oZ/8Xop3suUmy56M9byilPXQIQZHtSFsoBc2YIwQBrhZ/V0WCqaoal
iE51BvQUrYbqZ2PYvmSLheUlW6JEc2XWsjU5ZNyUBIH7Pm4TjwX+3r1xO1GPIooetlxgcWAoFoIl
xrt5y/uER0xpTVk6IcbuL+Ms5JlzcJiIq7a0XXGoSnxt6PyvNNRwI1UI711s3XWvnZSHovRkrwF1
VKmG/5KxL2PYMCpwSBM5ysAVulfZolzl1HCgf3nnEQRCrMmIW/dSaSTUn5DHW5Pt17Kv16Xk+mdp
4gxFxPl5h8lTkw0yhkwRTovmdS2NYcrzLPBTSnd8029V7HAPKGUk+Pb2zSTfKJYxALe31ANAp3d6
9sGQwp9TIZys872UHA9xinAp5o/S1vkvqsFbujcDxOoj/qtsndtJWOhYx+UA2mx5/8WrHyXn3VU+
wuJJD0v65qtT+qDAaVE/8csNKLs4t9EH2fkAlEkcudy0Vnd1wthnOuxfMamliixvDNEyZ8XLp3ej
z7fUkJuA9shy4H7SaQhEwiiMrOENQI+jS81QxiqLSTp2QWdEZXsttLCoEwqgVbuwzGSqQrpzvqtO
JhSDh0b+7rqq7s/mSdDoAFc4P9muBhZfFH4QZ6iBbmtObgBAoL686I3273g/JwNo+0+Sm0LSsNkX
g48WoDdAwgSDYNbt3XZgxv0J+okx0avszu6LsySalbcPVjqsTySq39a6qHPF8NKLrEFJD77i7yFG
g476MkcEM073oFlTGLKFfq21zILr4oNfm7v7D/1MkXzrTAJtpr1h4Sye4Bi3mG6RfKBLALTgUOBT
9IKTs0/gkucY4GaQ0SMmvuf2hQXoBHsrrhpEZu5oMGirKC9/LixhdQ1hWY/2QZCFfLidp1/M3nFu
TG6OX6ZKaCgxCQPxYIH4NDArSI+YDaPpADrIOjGsty2ITKCBRbc/YzqJ1pDHbb4ahlo0OQiJ+7Sw
ISpbdh13uwvlmcWv7fyYG13loV613E1N2hy21or1n9LcIwlfyoQl6cm1BeyRuPmjsgm/LTzFhVIv
Qf+qfjn9DHl9ydOjwJnTI7Lw6tNxc7vzC/xbiECI1r2UFnjdf+WSGpthJx9QpzPua+N1gHqepXN5
TJLuZ2uLghCgOZ5kNwzVRalYZRdqaTxMJCoDa8bLi/jDos56X7XN0g4E4uheVb4Sbhfpv2E/6zwQ
mUNP5ZWR5UmRfoNnIos+/hna/39QgcfSQOHSyKWmzztiiRteyC7bWnrkPEPYgebOi9IygHaM5GMd
iMz1lW576KvlZsc+ukEzqd/e+DcctWzPve1AI+gJk6Tg4qzC0j4PwGjv7EN+EFePo085D1VUwg6H
m41qR/TgKgRe4nXCyeRzmrHwowm1hPMucOZq6owZMKK+NwYXuxULv6IZ1jheGaiP+1DrOxQQaQD3
rN6LwWoEfROyiDoVxHYOyJWDbqh9PBB/gj9MbyNN9lXb4HItx20eBcFi9Z4+s2pUkdIYUgBTjTXD
IqWHOF/swLjqEMW+ikXC9xaff9DLhLrjPzhqsAgJ0dybPyAezrlPBJIAdJ+29kwwmNRqfJWHTo52
O6sWD5mK1aqu6j+YagEBEk5tHtQp04vH0jigVlUDa/2rki6SXaEBBK5rFaHupG/OceOtlDZIZgrg
UkYkBvkMPGAVkzgoum/dpW8NRIfsKelNDYcJqyOcUguFyoqjmgxquRGQx1uJEEz1dfJVhhhKksKh
qw89WaqkH1WQ0lsjzJj8wiyrxqdtCW0g082u+P9BiyqzHOPquLBXzmxnh+hw358SKDXMdwOmViVf
Cy8t7ewIVTmRMpHDuZ1f+s4zBxjR7R6CsTQA3bSiGNCzrbmCi3R/A02G1vzIKF1bDP43RFc5gcEV
6GR48J6pjFEggMfu9gydbqx2rFSe+6QLhhehvmOSO+Rfr/gquZJqqgj/0935mPy0qYo+I5/RAq4Z
Jtv8+G0hf/lMSvaBQeYQi3ZyqEivKvgxVXCXFPwP1Lj7RyviC8XHCW51tAL8iftmzOcdr4dkLyfI
YCw0qL1Tjo7i9ptDPRBsHLSNPiBkaSjhAhPgrIDXwgKct2amdYRpxKhpRG36O1rfmqa2ZB09n5hp
IpIoruPyV/v44lsUXgCNa4XqZK92VbaSbYetueUFyICBQ8dqkTJ3Z0yCv4rg+5lKnNwoOv/D+KdK
L+5YSgaV736dgNCkHfsEvDvwo9B4vG9nw2VIEPL2S8aR/OgncxKVCEjcAtDbavTecTVqQ+FwLz/g
Vd3QmcCv86efLkOqAIZb5iwa38neF2juckq3Nkas1tbwITNrmmgbjhBKjhpWKd0cgYtJ7cvltKI7
pZavxrBCt460TssS346XcErfV5gQ+oCxJUMAkOoBC0DLh+GqKvoJw6dyMefFaeEecZStMXmrBHp+
bqMEfB6vy6U4qFr/SEgr7lvpktfiV10WnOqrVQ114+lhDKvF/zKDuiMkUe/+Aoco08W7Io3c1O9J
jfyVyQi4PYS7U0gJ35KhMGpj8Jn1wgg/vXmbs3qTQbKRLp7K2VmMIvhF9Qgs6DwsTiefA7ii+APc
tER+FDyCchy8gc1KKV1yUofBMtqrgzzDvsjjW7lJyH/aDzyPF5qMOMwq5j0MkPZFDPXqS4XN+1G/
b9T61PSK15zrZWnpi/yiUUz9u2yMUrBiOKYCasx5FfDKlxdJv4GxDnGChodKz/DFuLNl14Iv6Egk
lWXOFdc5W7rBw4bDAJHJm9h+cWT0g0yCcOGLAEZbsAYC1sBx3no7gg/T7hZN6KkgdXjjYi7H+zC/
9WSUXW8l+jedIXgM7niu9ftamZCfZ1LYIv3wE70zndIQayvJjTpGwEahp1g+HbAt1QVY0o6/Vefs
3Cp6in5guGcWDyO5RAAQL766tZ0dv5sbYxICbmc0w8uV0vPLmyc9+lS37VyuewzPjzXH+4BteFDH
VMCmRf7zgGzVw0N4q9XuwxTqAP7j2Gg2xolpJyVjRyZVwzo5ApV6Mcilkw9ZuMFF2cRlcnn8rwtj
gW74SUo4x73IBwyUnohb3+JCU3GcuniSZEYkfyziu9V93+cH+EptYOz0mxKBl9W6Gz88aBlQzo1B
NyN/gInGCJU+2FqEeIRG3PQ2P0t/VMjTveHJS2Q4ecldYABy9dymuHCxExcvMHtq0bVCrjlkMYhe
ntWz5H3mtHJy98sJ7z/hShEq86MmlDMACkTB2fri+274egAZfBQmeOK6fqUYsodBdXezPkrraCRw
mCH+p4gFHhTrC6JZOU243CiIi17d8dYBN7+5UYG9F5PKOLvGl1xYgL3p4onNe3RrBvFgOBJEaQgC
pRmErjsBR21OPlWBuiIkjtPIVqxPL9dLQp1Kg2SkK6SLmUNx/2ftit/fBUw1loHMD0H6YHgO4x22
VqNHjQkPbQxnecysLwKyugM2ji/gM2sPncosE9nwSqIFPOUDpeN0kEuph6PCPW1BQnhH38LPjVe3
TnQ1lPoyE5PATzEgeCRXzFCnjDXycR0XQEgFQUE0NyU4ZesGL7+jQZl8UW6tz7yJZJVSFjidvYiE
U1vzW0GlRTISZLN6WCzO63ojDUWM3XNhlkHzki7ocKHfTji3aIDvBQiKw0jok15lPXAPtPKm2Lnb
YzH9aLTSYNKg/nV2MnPYOiK7zZoyt8f5naV0+8tfzBC+c+U9g7gijVYKgeMNXbUSNYUc1B88Gt9g
Rrt/LHl77ga2jv3xBDOBQhu4J/mG3i83C5ye1XiXFi5JN12GDqZsmOsAdg03YdtOsyfHmAedoW9j
38S15XmLDq/3CZyreRDyDR/boSqgF04z5rNibgwX+gzVypH3vA6+udU625KjdUPfd/oaIsVvciu0
j5G+wUt73jDPrdzHzDsLnuf2xP//pXMHRn+Zacb0t/FMvUvDMs5pGEmzHc/y96U2xAIhW48GSDha
MKigh58AmLqA1Mvjp9BCNKDoNL/gVg4wWHaQx6MANVYHM+6NgYwd3I0OU7pBTAJaXTrLHmY0H4Tf
eIpV6g85Nk9fcPvwR+PC+UsW3wAPmEuAt76zujsk1+3vf90ap/mmdp4D4yn21/EKC1wSdNLUXxBy
xRQn/UnLQcmvCiZDR+T4/dyy8qL1gytiDjurtbrNNh64o/1aIMzSvvuV0k+obatyn3YsrD73A+r/
suhIDdRMh7FIvgNjs4smT7lfijBIIc1mm/X0WNqteyWPXCDc6TZznOxLBexmuq6IcxKgUSLcA0sC
C3sry6bEgDsjy1O7ZPKpuo3aCqwjZV4hI5TqZ7GmRpFETaMIz1OxEH5WJ2bKH/hKYzWl2/AAnTSW
fI2lShUBu505xek0hiMf/eAFNSScmh7XXSlQzShKFVmvC/xM0BU3nC/AIDpWZEkIwTIdy/lK1N97
xEkwL4DwPj7kHfEQWhe6bZs8thdrTnabKpdvgPFW0TQL/7veYN5Kii236CnnYg/fszNgQK5w5Q2f
BtBTQxHuZsGuu4b/qEmDar1fUCRiuikENbVFnKtm6UkRhv1HJTsfbSwaVQYMxAyuDvB0maIH5Yq5
IqrtRTxzUoM/WWYp83x5NTCq6nr00lyuJPmUUWhRWYsXMWgC6WB3rlEcZCGvdsWtE2Yd3TlmiUtu
Q3CuhqJ5uMxTKF2Pt6ppidgA2TheMBG8R+tvxU4gIOPSSEx2BDx3vIaYuR0svVePrWimFOycpGPm
IicALqKBHUAyM8aJRFUYsmlHcmgJreYm+iSumcudhX6V7x/KhSx8RSzgdJ34DW9E3zVFcPiE0XZC
8/OG/rMR8WgJOaTKHbmEM5uIqleDhLg48K/sWkDxLdK3e1JjE4IUSpxt0veSjDXhnv58tBbmxXEc
3+CprKW8XzjzPnmxaT6iaU2DSqL34B4k4T99gm+fOhh0YtDkpZiLtv5vfj7G8FG7H9iYBtxNcRFC
FA45sThrWd0uM3VD/90bE06OxbAHEbmP75zmEG4S7Mi2TPpZQXi0qa0gTa6KAcQKTK6NInwSSHrp
iEoUz1aiViVnTdrHWd7q6GUnqIrByb1pRu4k29g8mwVdQ/aiO6kyPOjGgAHjA+5V79pYvaivfhMN
IpkBdQjk2m1SLgl2GhYwfIcFsr0LApRVbwCLQs7tjHh5v8JhJwLv4VQA2NaP3JfPT7GoAWS7qjBw
8vD2OX9hzbie0pchrEI/DsQR6gLUJD5qYgjtpllPDLVDS0axK36Lb69G8wkQ5e8Q1j8YIB0HdZwy
w4P4UzjyIEsE24TaLwZOVbydI1R6qHaApjWSLEhpZtfm/3U8Lxw1t9uOMEZagYOl/1A3GhWZyrqo
ERyRiOtbdfhSoOFZyC0wD286+r+Y/I63oniDaurUUZZOhk7HxJxgn075xiC2hYrtz3k362lAHfa8
XjCKJXSjP38/NSZcjDDnZ27wtXWb4Re5mVJMF3rt6Xiso5tUwjZKTLAMUuyEeQatgSqu+xUtZDjI
iADXaYI7Zyzm78wojBIC8yWFvSq4Vei6IuY2eVdoVSmaqBRR8lZcyEvedwT+BBIB/sjA8g/yZ37Y
6hf65Rs2Z5OdL3PUUNXHurRNUST4PeLUfoISy/08sveOFeCGt+xws2Elxa4NxJjfgaH4Wae7tLQA
ky9XzLUCA2Z/asZ7xqtIALZrpjM3fW+IvXGrolJBdjDuOdvIE19pkLg1tTE0GqwBhc4/uEefr/7k
5LWtrGRvmbGE6Khs87G0RJa3z9agIpObYIGcEKrYf8jx1vo6j0fpHkuBuFPic1WTpfRly8ujejhE
uScu7fbGdKD4usEkL7vDq1Y+YkeqsOGDDunPdLS3l9+0QD7luOqh6oziI6yZZAYfBZ5yQDIYKFt2
d3R6H4HE24gV8xq+mDcBL73JJnwURsUA1zuW9LCD4ZISfDUVGyrgM4i2N/lC5h30atwzyF6R1TvS
D64IXlQj51uW4GfcO2pwMvSijSwtUjVcD8+v4WOCvrQbVzZd8ZwXScIsvC8mZFEwBCjkqGiW7cU/
T8ilhK6Wj13fcJfVdKDAiLI4KNxWldzzdrS7/pbj+OEHTyQ5PV1YXo+lku+6aw3aHTOvxnTyyluY
oNPh0WOrwWJObSazKfOsThR5GZV8mkGQzIN5KTGrqsHkSVNChl9IAKceEr8l0AHxFZ49/BDUNgM7
BM8w0d0Yk/nayh/FONiSswHhOsqNGEIhjQKZFT9+lIfYyMVE0Y2hCvYUKQSyM4NeYgW0RSJD1/rp
opkvx4Tx2SRSMjWwsSISsTI6tpr/ks0LxrWNyx0Daw+VwTJ51UDtRyyHPmoIF3rhrxlDWhOq5oc6
aX+2V6jZh20G6dvn/YmmMU8A11ppKflhdSHfJ9dCzYilZerxmNuvrTSmZafxHSmZMeRyADAoe6fZ
5+S+gyxOBlKGQYm7ZGQVYB2CIz6AbCKLye/lyRULSkwxvL/lsYu5GhCnff06Pjz4/qfyAfvdpokY
jZo3TMNS0D5HKJIETpYbOaZvHOrb1GjEfAbmBOfDiAlNtHA3WNd1ng0fCNQQF87NWVTum2zLOMQY
W2FN+EwmGOzM5RLS4B57UxNZ24L8kEVGVVbJC+Sd7Aa7W90P/dpWU4g386JnDpHh0ll/zllsqf2D
vt7bqduagSaTlEHWiV/moZH0L6Aj5AFxcxa5pibCQKqeH9v+cLTDCkWTffRcNv2xPscHsBL7Gf5m
oJpMnXJykDdqJ9R/afXBol8Tf0mPw/yxfXwAEQt0pgRX8l5fcbrBl3Z6Zpp1R7Dosse1VyNtetPr
v/oaNgyla/GRMwdHWSOfotOFaTJS0Aa1qPxJC4+kBXyOYwVa53dNpFQP1u/20EoXAVSRoPWNwJkD
urqDumAbkPAU0CNdNtATxfKPXWYt5Ei4mE19MxwIsYd4Q0npJ/IoN0cFTVeKjz60MgRGUkDc17bt
54McKcHa2KKwqRWfM7z8RnbdwZPAsf/gAuHE7wQqXmevFc22iH89TBqsLcyJkAzP9O2HdqzKH3Ig
Gi2xNAa3CUCUBzN8uLC45AP8FgVq5wG3WIBvJDPaP0A4QfIYjwlrUTMgm9CjsCrBUMfvPQBb+PP9
GTRszy/m5kjeasgcuAiBmIyrlkxxPPJcua1BGJ5NgWjrMDEzbj0VnOZwumArIFD9DrCjxzTifnKF
CU0oeYDrxSB5roYG64gz/MEvvNNR1biRx/vr/GeKTLOVfwlBWEV86bjYhKzli9i6WgAyBgZ4kMAG
KzV5HRq7/G3ZbdRroyTF5x2ed+YEJvAwlOCwDWeW2mcQM51L7HrHFR2mwf50uGeQNrcDUJwGqTuG
dWcbb3BpC5JJ/X1wyuDh64KnVsO/cfKCKeAB8qDHODcXftnEB+C1IUh0q8PSfy3Vrz80ziCmS2r2
wM0zZSGu+FwTp/S4FB9IP29GrluMElTFJhS6zps/1Zn+sknDkjs4aJzccwbtucA9KuoMtGagEBJv
nfoI93BSRBLQllP9AzlOAmh4278BULuCitdDWRFT1VwxnI/QG2i5RXnNUPnzb3cjvG2FyYkTQb1a
HRjirFZjFlP8ZhqmFCAkJxieC1CrcalNPfPbgmCJ6c53MHaW55j6XOVNYqBrPte6pIvUS5SU8ib5
wfGv95B06DIm2bxG3NWdLuQJQ4wWyvOvZeon4mcyqhZQVTELu8qyFenJNosCnSK9xhxxCdqhICi8
HyA35NnO8ot32EvoHvQCfvRqd3QBHfPtf91aMNauQAE/28wgWzIbVbQMEjLhETTM4dM0v0MikjId
vqfEVFqQiVYI6ptBDeFcBTAQX9yTBtvt+l2B11O5Vmr8cxZdNkokVGAIbbwrowIjDsosrv7rIZK4
7S8s8ln69tHazQQDL99U+hI/gpSjJh5b+GHcUDyJI8VchnDBpnERqLQsUoliI/lM7uznC53gOMxU
nWzJ9A5yRDtgUWviO4l2M6VQrL6iKhtzUwn+4H15QKn8od2KGKjlLlBrYsaMBLPVvHMnI9wcdcWK
m+Lpstkz+lnCZ5yd4W82uvSTcf74Cgm26qruBmRn1ppCHI41b3ED8PnxP4Ji7MT59GKfxla1pSDi
pV60Z9Du3dYAEJvYXT5b4OSdWXA+NkOvg0RCPfdQV3IdxAwWRbXUzJQ4EJ89zAvX9GxY2S6N70Fe
Zvqzo2TdkGBe8ZVbLC0XHFK2ppB3T/Vy9iFQD+6nn3337BpGqWdVVBH9W02Rzu4UCx2Mu5mw5XSL
zlZlQasuIV6XjLDuSDuK04TbK8cplPEDRefsIUuWpdrvGVEnTDXOxUsd+8onVA947OlQa52413OZ
m+OpOQMDMP6eiwq/U3oL0tO6PmaBbuHvapbs2ghGTRtqR8iRhKC/brVx5wnlyZ7kxj+Pm1JLx4eu
bZRC5wJM+C0GOwqwctOqj7qfH6YiH9bHHvOd/t9JOXd2ge/7RloaGz0yNzIUcNsO91VO1XpdgJwn
g1SG6VGV85p7xau4CgGwN+j99C14YUtpHYpiLeD+9eOlu4Qw7QqX6p+nHBgYWt/T0iI3AVALVXlj
B+ljYVgrBmRULCxBTAnr3NavpH11I1mrZcwc9iQYfB3A2c0mMg9X63I99GJj35nvyG3YFIjE9/tu
Y8hY3Zt48BO/QU9nZ9CTj1bO8lMLCH4k47W4sZjowRhAbwkeGDlCrzd57sHQ5vAMxl4VIzji4+Mh
a2aF7WhmeKkGUUL0FJ3omJM09DVfuQul4MHIpLyVLPFfgo1C/1tryXUWhLn/JDOj+Qkgf4XiExxq
tWXSl8abcakHIvvKf/JAAfSoYfNoOwXe3ptv4hvJytqvp1r51RbNb5EPs2ji2YrOizr9CrqEXE0L
4kE1nxFCXALe9aEwpFvzx7BkjKgT03RH63jjVGhUyR/O7o/TBkTpNOK1Mdv1RQV95CsevxzEgFtm
qFFUBd2DP4lh9eF0Nve0nM8/k21mX/93nBy/iRQvxRp0EQ6xZevEMg8lmUnk4hwLL4NWZ6WOCDQw
eDqbAjIV+biodMo0+3YRQPFfKdWYJi+ZwJZwXksnTY+BjJVomf41JXKoxFRl5bo6y5fsBJqAs0wn
lFcNY1swKSxtfIvbmWA1fklsz6SdVAZ9vyLnp4hBXfQF8R1uj9fKw6HZ2Sea9ZiP7owCVcc4M16v
yVtoI8mpxwecJEQAHWcs9ucASPB30+u7snzeAr/4F+Z3P6jf6HOanzBZAV5mwmB4FLK/6+i+goco
hVnfQ/234cc4bV2IxT2AonRj0JG/Vgqh7Y05rPuWvC7Zz6cofLlQteBcWRzPEX42sSFnphcUUZiA
EeFc5O+BOv/fUjzwgNfIFhaaXZ2lojAhn3uCT8d359CPA02fVYoJJYIehypPUZqEvDBK6TCopuPM
DUfOKD8syohKFD9spUoGoSdhOHbiV4ajuA7G9ldkhYKsSn5pxD5fmpXBHp2mzgg8+pAjsG+X9xAY
4A3MtATWZfdpWDu9NeR8jAcMorqqHlmsRG2wvv0z+iGXCrdS3j8hV8e2a7M/KMr0zumZIMTFD9hg
jChhVHw6JB82+bfpZeYb4NDTwW5cf7fQu7PIE5g4vpyhiscTq2iq7dSSj8lqZ49/QgsQiVW3HfuG
bm2foPzjw8RxCDJutYcLHtis/5+2oDJin3fyeYaIJXPCZ27TjRTZ0zcuuSyUedXjdouUdZmmKAA9
BKL5+iebKzvatYwbsnE4bVoLNykpjNLrAQ26vR1eMBAIfSehYLHtAZ/WkAMNl5djCU/6RRKtPOtn
9B+6Qaer3STxUqs47Jjxmwekz1wAaDpnCNeeyyTQfLbswzLyZcFoaUAQ5dP0pz3j4mo1Fqw+Qylw
hu/wrr4FQH14krrOH8T/4iueCiuXAscXvW5Q45xxCwz+sso5Ju4h6k1e/2SbfSjloa12x6ZD8p5G
m+oGjyWbC6vBVaIB7T5I/rb9bwgqJkM9s7RCw1QbXSAbukMCG+fQZKc0g9BRA8e7G5we33QGbfxn
/ZuT5nFGdSv6FNr5apqUooCYPzRYQa+IxFuIBJ2W/q89q0AIv+EHmbAMSns696rZmRhFkQUzNgqa
KnHNXtAul2PkYpoRUEN/bM4S+t24PphkqIPgss6M24PU6+juvxq+VheWjxyPBM4HYIZMMlo2gpqT
6O2UWMMVUm/zsdI7HcOsT0glJe3PQmdTejqLJim3CXAwhIzTAsauPipxiq7jRpBzia1LyWEcslnZ
GPQlIjbwokCYz9vlgMUXW21FuNpvWsZnDUk4UZDNJ5EbSMId62J1tcj/oSiv5R66fGrftRYDYOYU
lbsmjQIoze2A+hFZEbvCzKpD1lh4VmITCK+kl7xs9QJlyiOnFOw6+gFCYWbDVpvvIZkLSIvOdW23
956Yrs2ddkADWZJlJg+424oq37VvLn2Bjbu7uj0VCKS6tuvpcSTKNvaGQ/ruRp3rdsZFXyzIYxYi
ee9r25VvDiyjg94uubzcJxulmVNlMIMaSe2a5Xx817aMgUnEupBPEstx61fsHPu0bbypgpJwao7V
IKjgqrXgkPRbUAwT+zvdLrMhIE72RXMGaadilRsq9w41RU60XROatKdit84oMuEdVGH5uz1vloP5
Ellpvl/5Bp3CiM/yENvmzGLov+8KAwzcJTqHQ4hG17vey8mY0HImNH8xSyRnuynwkGQSNetHWxEL
q93wCEslqndgJ9ngAX3Tj8NbtlAYN3pi/fXKVR26J/Ko2Fx4DuPM/V56X8J6bsiyLo6tvDLcAVLP
3xHMHFEG9sy+ihQfmLuqELqEoJz5vuUvt0+9APyuuhhSxNG+HbSxDIFHsWNFj0k5RA2R5i2sN3Kc
U9qu1UYWTMP8O2J5qYYWqU9n3IfSw55tyA/sQWyY39+CzCisqlZPe4Wq3MUsDvda6eYW6Wv1xwbf
zuTMcroiR0+IeltUhP6/4JfuEgChjfnCLD/V4ypr06fF0O2pPTmgfPU4Frg9ilw1XIgUNScm8lDq
cwg1uJ6ACESGxmCMyUbEsk/KvYm72jCwXT3gJySnXOy1BH8qHAndUWyph5439xOzR3fyGJEg3Wgn
fPl72c0kDgDglVo5z4BZl20Mj0vHE8ADG+qMEpGP15MlPQV0gq0+CY3DvnO6uMNeB4QgHa+XeN/V
YDs9Yw3J/SrlgDdE0UhHPJID8dTs1Fsu+UvwQaZG7azZjUdhJPqy3Dp64WL6+bqvF80+YjSzJfwi
V8O6H7xuK3c7QJkEZlo459sQuFTl6qxHaYWQPCatHXAsn59/aiDasRjNHC2Acs/9crj+2TRY7+Al
vTYOMIuIkn+IzmVU4V3xQS1Xv+kJDvmwETLkxbOa9Ur0dNL/O9wbUMaeYGbvfo3TnLF3AAUEdhDk
QVdR7AQigtBmZkYQjLqjcyxPNK/UC8Ycj5LWu/L8fJpqxCU6L/B66J2TkPln+xTMji0WReokiS4t
egKjsfuVuFjvChuPUXUib2WvRtLbcAuULA+Tp+Yw9MKBSqbV9xmU+ZYj4k7ASi7ovZGtjrnqveir
1EUxIFMseIoWmDmM5eKhCJJep2y6Uy9Xdavc/a4UXLJwdUduJH+xtFvWnWmur/jD3DdaM0glfQtf
lkUYqsYc0ADMcZt180nWfq6QIY8eF9wD9u/2D40taA1bdWdG/+HU61i6mGTsDNjHgYPck9OxjByI
clYQjTv57IOlEfHq5AvuxVM9uOFekH5sDeija73mOahV4T8mtA09gFoJ7JM9ImBPyNpS9ZfytbN5
77UvxxRwnXkEI5lalUhQFt9fYIk9m8NewGuF5t8Vyp/Y3HDB5nRcNZ+pMkolpJ6c8nqsq3Y4JT7R
vChwdLUe0gpfxrs8/5fwEblTgZYV+WQ7KVPUX7iDBG7yUv5BQ16pydRDLxYqzCKu5gw9jTdMipD0
SHdoW5cnau3mfHGnXXKTJmzfO9APaG6pj1gdXnvje3ZHBsjZ+y2zAPnQtEdOmjQXHd01e2lx4m3L
r/FeHnk9u5xpAk7b7/vVyB3poRBeJ10fiwKWutQdc2E7NKfD4V1L1Zzy55xWxo6hJ/ZiP+AmZHmC
7rRWufK/PFSUUVo+g8Lcfhq06sYjdc2LhHgptUrA3A1zUM343DpKgIliAWOTd///+xKmxux+CTLy
b/7SqhApq65jZ/wAeQdvrWlC4XaiA3Fa4qd7+5CUk45EhN8dAjZkBRzBEA7DcCjmaCkTYl+GHp22
Q1iIE5SGqa10DDtZHdIktd2ZqukLFlEkJhVk09MYUmwblUgyfsrBVGBP9co6WgArJANdVUdmCfmo
u9G3DYVUwNCnvgbsVUnRhXruQziQeVHn4l39IEUDJ/21BshQ28D3vxDjAHIaEK7iMxT3LwlUVpjn
3/aRTmc08XXU7iA9n09JndM9t8jUSI+mlXB0cSWx0WqweIIa348kGCzKhDjoYfWBJIkjRhJ7rul8
5rSDDegntIjg/BUUsIpmJWHIvdsGSU61oFdTD4vyHdWU2OujFw0nQzdeuKYFa16Zh/i/EXgguw2d
UGZhis8xGYva74ha7Fs7Q/hU/NY5QyV8UqYhg8anmmR4LHwChuDZCvVSBY8nXkY4sjhvagsSr5tK
MW5bfl3F8mJWlksimN/Di0dNFn59WLF2UAzw0SLWHPmYNB2WKIHQrRHoF6fmudYmW+H1TlnxzrNG
dnBr+DkSjYRSQlt7UTnpQ+Ikvk0tQkkVGhSn28qHrDQrAdbdcdFw//6+9TKxgCcPt+oWa+NIP5sv
jFPCbnfWjVhtD5vRXXGq+Safprdc28ifL3xQVX/4PLsUSeXsXW8e9XvbyOCKdbknTHPbRIM0UL/O
/wzIZo81yJ7eXmN8FCOquTV3lxmSgBzdA0tY6kf1Tf9Jog20ujaGINKP6VPB44OpXdlp/EqpgL7r
i6EeA/UVzoosyXYu9A+NMDH8oW0pOv09Gt8sAsE50Q1kPlatooIOfcDDv1YJqs3BZYmllhlxdmC3
CghhOQnTmSITErdxusldwD1fp4chkuHswbyAzbd1o2jWYrzuFqNl4CyML15jMx3OPR9cFgbqvMeZ
e19F47VJ19m+QEu5ofqAR8LK6o9nlZ9gphbuBM1hiPQEuQBhP7nN0RMYtWhUU1/jW0wZfURS8TRP
nmev69MFMfMkJF4lhGSo/MHdVkz2bR0dur4pd1SURwri6WSfcz4RCgqyMD5k++KbIMPY6Lp/q3vf
a190yerGiJY6copk8Laebdkzw+Tp0fHpSLlXzoigAlDTll63lGVzbDFFSgeDiuHv3VD9cqBykp48
npD5tppLFU8I0hwKsOQk9VTJf1JHCiLPxyIbQPBS6gg/3/g8X+e87yUw9u97B3YIxFX+Lbpf+kYP
pFi/HiQ0Z+ubM8U1GH8S6kvVDbf6W8ZE2NTYOjjyDFG7zMo/mUqOQQHfy88Tbzf2JjNYqIfWk1Ek
ZRdl8K7a6pGXBUuzkuNQbjbM8AW73AKO5TPurtavIvo/NNHJ5+21iWR5fKXNh9id3dNC8asNDPuA
Bprs36TK5N8khkErb1g8jg/+K4qF3TtLON6Wzk/njwUzPjQcY8UMcOGRvQcrS1c4eSQWCemKtOF8
7kC05iQhk3GPqozZoqDFemDGOdTM4RmQk84Jt5m5E63Dekrx9E5Nvsit2u+4dMveTWvW0xKWYfIc
hkliq4Bl0qt/HSPZL3oslfRsHzV+Y38DOfrBno8MAu53PVpO+Y4xS6029yaafpNKLgNu4TgPCpN1
TAVHKP0OtQMBS03TWTPnVdgFZIPILzEElcqAPXkj0VdtB+D/XQ5z7Ir58hrrbDJOE/mWUujmClok
N2UsA84vaAaIcCzs3HdtqsQc8A72rXbAaUgDd/NsC6kahPHbl+2wnjYHMgUryF4hkedRC9BgundI
Z+sFptaTrRA4SrGmBe4uEQjl4EtCVPQ173fn/gV97w+jQZkBTuzxLaAGIyLSL21pFa4KJd1NFlpv
RZGe2RUQBdhAHKgxMdI9Yw1msIA+EViFPQE0PQmJK0n/41M1tze98xawxOfmM7WuGCCIHXlDvj7X
V+JDXkUEIUKGlQQzcruy3jiutTXShUME1wVkQsypOAuk7vzFN84GAEVMXPeuJwjwFgFloinMRPvD
bi0eVd7+ax9rslIbBZAUH1KvvLOqXkvCOlDJIU71WNGBWe5nzv1Vm7TZNHDeUyHASjcr461gYQKa
nArXHK07eE4E/D3MtmxLtL8r11X9Mpg4v8pgiFDb/1toWWn6NPAIp5gsp5ufOgEU4SRGefT6oMuI
Msee2gDDKWxCKDE6q8c/zdQEgG7GtXR9NNnXG588xjx+m/7cth3wOr7j1k2YCl8zNcAG3w95iF/x
M0b/nex/yGvXNJGahlssggptmcWZsnIuwGL1SPZQNTMr9tTq/YMGk+OZWZ7ELVtM6Y3TjQtfTIQ0
zfNvupDaAOu79pztvmpbvM6PxHFsQmt8daDXWSNpXPv/lWeRd8WYl8u+hCb3rzcQJi7pAp/Et7SA
BkilZaGb2Z3akL0NzQy/nFOEv8ouUj/4xUkjkW00PENkGnN/4QPmolnTJIiZMw/nFoFnwm+jZnCU
pcG9P+tOu86DhLbMPUbfsMcxrOFo3octh9+tAwMADe936SmTVsr8o4zv3UAq3OglobuVrd+6t5oD
pbieYE49oeO5jGOTcx+8KnNAo80pK9Fg0VSQGuzdcBsifvcKJKTGXPCXVIwStCXFLFhZTX0vbdVO
hhxolLCyfSobso81PrwinolK3RAdqvXL0JS5r47SusXwE+v5vkkrZcrdAkmVckw8nEasU/9iUaQl
XnTQfJH1Ao+baIge8xOdG+/Px2AhOtdPTT9zENBKq0/3KJEpqFBH/Hz9fO0ZpztwmAfkPFYJ4bCF
XWZVdxYXMd6xRdPp7MshDqMwKB9fvdSzWPqfLsbZ9X4boMsGkH60eMjlBlEpaeEkNWfY4mb0DYxg
pBZwzRtWbuZGVLw3/whmnIsF9Q0l8y3BAbQBv9s6voXOFUASb7oHRogu9QkPORxtiREE61kBnilU
zwCu15i6fc2vFpDNdbYkxdV5sVqTCSYnoMTYmU3Xqbex7wi/NeGpaxZStR1cnjdWdQe6NuGrSVrM
nsFlsSJE8V+0qCqJvkipZOPE2wMQB6nmD4G6blNrNFMrEdNrU4ehSgHwOiBw0HugKlJ5G9o/eMHB
Ru+p25PDAOzxqBd04/8UkhlzFVGvwJE1olesdWTWTCVsqjwf3dnK/7HtKOKuFi6A0niX+KgR4UAj
9dvUEqgJgYQgSsdZgw0XyfSHdF+jUL0vIXT/4fUvZ6/oJUV13qYZZJplUbB0fUBeAiLQCPA5Tbr8
tIn4x3uopgxef2QjvEjWZOleMsyKflLHfuFOBv6nof8ZpBhWdpJj680AqUxrp0oJLUUDyPeIEURk
fgnlDsqvMBXOiEaOQSNBtpULWfz5pYTbBUVA94DqECuUe6ssJOMIyf+iewOm1pkU1f2uWtNWlnhS
DjynVWrFpZ5iFIXHwtp8QjhIce0nN993Rm8nkEicvmqU6UZwZsQhAXtAhtvKt6JRYVXLZgRp371r
ErDhCfagqZgnTamJV01n9npLr2rXivg34eDBkBgnSwOp+0PvI8Hm21sCyt5eOUJj4MsyHlfjpg/4
ZyYF91Fzig/G6EE2hI4bjwE+nni3aVlxJo/1dsuZOCXge5fxANejtvsZkFNRUfSkwjRAD0NpB88z
/cxvVihjP9t7l3ABKVw4mH9EEP0Yl5O6mYkgFRw5jHcaW4pickj2nMCtlBJ9lSQJrvg5XF5oA0dy
tP2Fyq9O17wElpKKPY2VKptExuzr8O7zrNir1yTF133s7m9ueWCerBaGm5T8IMPDHc0IwSaGMoKm
YHP9LTo5cL9gEpm6JEwRK3wJq64L5LsSY2JR2Hs9H60/9MfXGPj5p474ouO/eWhP/tpR46wddSjb
MXxOKAjYqhM3Va2dLNDDrcSuJz36Fm1BI4zEv9PGLNrjG+HU2EOm0eU7Q1UGo+W8n0Y2Z3y9sRC3
p2wwe+b+HswwHcBNnCzgZveURAQaVUuM8ClMdsA0/JEO/xiTsKVHtWuQf9+AWCQaqVRixUn2moQi
0tD3dGynp5n11qpSYAsi5L7r51J9oajPeVIuRhZUKzqihGrdjJGdmrE0bfZuRir4bxR1ViFXCO7+
qfOMSj4drkfUldrs9RJ8KR+Rmyp0CmQX86Y4/2LVYgGXeAw6ZVmdYWG4m0WZEWYQP4D3Ok53+5qp
4ok7kypL6G7xDIpVlHTGI8XcGajNxNU9bqxAMSPyCd4EdZX+KZ5li8SwoNuRZ67iiawFIxPryUdR
UGvRIXnQDUewNHsFRXqHuC0XPRCcgaLGaF5EAM4jkM1W3DAdmC5k7RDEGqgsGicljE01x5VNkBsV
egbDknMTO7ASj4bvwfdFtIuwlpeocyJhHgsrFbwbzJtmkp9CCYmVMwCrOI6024xSzyq/GAEXis7R
PRdhkjey4sZkR09fit9EL6e24yDqaXK7jvtNuCTOzLMeWQX+xxvYZe1sAl97Y4DMzA+v70G/gm+g
FWKnOkf0B0ttLPfDDnniJwsd3/sH2B1uMe17m6hdj3o2PzK+Ugy22D2QQ7jhQWgnwqhx9uHCCzCM
mKXpQxx5WHQYqgo+HOIJh/PHuRHPy0XAuURwKG+MyoxDYT6Xa87yZtvScugpApHN+oQgiD3o4EJy
bqS/NSXFBzdxukaMtRYfi5mxXjaD9Q4XDYJSnuVxdb3r3J7rxN5mD9oIMSanNUeE9KVGfm/EZL+u
Rwa4znMc3GLjy58HihovIwQvGw0bmoxt8Y1eiVWZSKgv9CKx5yq96hiI50wD3u5yFkGV2f6Ya0IC
VOKVWPaCg99iEYHwKm6ziBuLJRvAlyIASvjwMdGkBXo9G1SROR79xjgqwrAatG82czebsDxZRmA9
kZPoDBSHChIosxF4vfdw8CkXj5kGQxy2AJvT7wP98H7bEdgy+EvlxJ+ZnfNjTRszkTY9t9h7vCYY
52L1082dcpbvYJbWBM7YYK7b6Mafw/rmif4BQReaX2F7BxGvidyXE61i5AgSYWrjBEPwemnUhXOd
+ZdWCb77kTU+IRRghs9TrBJzEHrxgMfeyEXGzQGyd75fLnJ30x6mGTNrebapl6Rp1NMu40VRI2Gm
w/YJNnYJGQpYphqLucfE+GaercRaUBSWN7scLTkjx+zFAeAa3nz6pdTmIBDP8O/ik+yibU3RBP2L
MyLUa9s9QUSBXVDyszXJquy6NHXsuoaYCLZgnr0yKD+CElIJmQ4KsfLY1AtfFhVDtbLScTzWSZaC
/p+IoP+hzeC7CWmTkJJtKtZGOQ5qJPF7f5Scs/PGm6yaEynm8F4sku/QNupcLliCRYuOi36q/bKX
8FBoD/uJNoOJDgwZwHte7DiI3neZMwjIrnxekFkeE/aGXeVZa6LlmPHzsuxCvrTrau/8OJvmku+W
QAkD6B5MmTGUfVZeLYO0Fa4RmROjmvfR+5RIGDgWDdnUmxEnjQJSJH6JcVwbau+OWqWOX2ImgaOx
gKxyZuYUYFJ+3KyBCIQCBkBd/Uaeip5o6heTewekPGi1QuWCJbW/mLTzJtrE/f3LW4H/woCqeouT
r3swdfzPoHI4tGs4YF4x8d4DvR7ypHqq9/zHrDf3F4vJg1ohZHW8752mAr479Qhv9Z4Ec7SwmtBJ
61pD5fUd2tFgw1mYPfXASBGTXjYokFJLJwgiAS6RHYo+7ZovUniqkC8CwCTBwxcySd6G2QPd1APq
WlICJrU20MnzXK0UzDdkXM6NiRA+y+TOEKlxakd22K0ilWDFStIElnUc+svCb367lwF0msNuQboi
bcOk+kF94UQqH3OaLW3JRRMz/hrK82eutgj+t8epxBtV5Ykn5tL96eNoDgQEuzPI4CwV5wPNiX2f
cYI1BVlSjC5jUvwddEVT7b4sfY34AC+Asi0Up8HLB+kgZrNdMn9lJAl5pk6vdAjlLC1HP4vbDyEs
G05+TPdLm6vjZPJsOD7d+Ag5zjZ2dvTkPVimbA0OsW1JEeXE8Mom8xWdtTEH8AYy1ov9wJa6MGBC
T6fTP7EglCryInNl11h917k7q83hCQlinacY8g7Fedfbk2GcbbYi00T9exql6Kpjr3xx3jiwyn7k
wdCOVSIuA8vqC4DnBAiksQREQlvrhdbgvXChXJBMGb1S/QnXdWm+jvo1OQphJWxmDySgFGcLhDJx
QxnfgNoTK3VGsDgxLzHRD0CsLV+PIh/H7i/A4npVNhnJUeBBQwJrVAcTUJprqDbQd+gxPdLuX6Gf
sv9aEI8bEaa+0eDsUugikif+uEl4dAngAWtVgspCTkiaUejUe8ox3/oBaLFTBxtP9k4zC41dbO23
v8VGb4o1hnUsixBUecgVb42yKgvGvO7BywcCNMeySf21DoL8f37UIZcKkhqcu7ygX8Pbnqzvol+S
jkJBdmnZf6XqEU4jPZGs0WUfWY4RnrXODU5VjwIZo1Gbw5O00OPg6j2bwCSl4qugaKYNukirZz0E
yBG9j8KTeTA44SbJOSzc/GZ/999L2vGuQCjOcoTX4LVSNH3lNZEJO5yKm7PdBd0CdJGUqSkI2mNd
pNU9Gcwe7kTajwnz6gVIFAqCRWOFoOIRXloy47fhOdjZC8+UYCPnGUYKT0QmavY0FusqJZWHdSTv
rD4yQa1dyLibUd6URTDTEkZunfiozgXWM0xl0qxlHUSgxbozo9VW6nfsQx8N6P2GGc5yZtd4axL+
2gF0hbuBj83iVMwem1LKKFhHYF2OI6K2Pk+UWrXN+ipulBbxyOtokFAuO2iDfwKj8rrv+QPfRYih
I10Sjl6OU/MtnkUplrQG6qz3KBOVdX0YShcRdQQUfysxB6eEq41qPErCT9QmW15O+jK39NHTNyDu
XdJp5Tn7rXeb949jhXuHWP9J2JaJHycRU1D/7XNxVd6sYhe6s4/qilmr97Fi5Nrfow/U29j53Ayk
GSfQlKEeqqq0xkISVesltOZWFOQmbPCSqe3htqf+Ah85f+cCv+5cCmfi6h3kCITI9q/Mt+Hz622z
nxPhxONms7OZBcG2F5WjIapmsJ0xLdXOhDfdeVY/OtvVHR5uFVlp/RpwUZxgaFw/VZAoNABKmSGW
C9b++BG7BrOKL/K6Ic5noMHn4GZFYybJNE5rzcxsaKii4dEnnYLiCcKBTtea96yD/occSfoUpRdt
iJc+yDmyaGkrPwvfyckry/A+VT4KsDVOxiT7RyRFFSsPIW56dA5ANkqdZ/upznDCu7Jtw8YRlDov
yWW9QjxHCX9s2/sI7T9VaPE4M8uWQSMAyr2iYuYeHrJt5mpd6QnNjJEGD4q6q7l012dpaOaP3iGC
Fl6ADwpKffvpCtWr/TEgcvJd+S1Cd78KM7zo37ZrdLZJBmQTCgtfXJSJ5OzMjOfQpt2fSsunt70H
eXSeLmE07ORBO3MpQsK9ocNg8WPxDBt5UIcDsge0hr4TET7Lg5EJC3nqJUp3kUlLLs+pDqbdSF2P
iLoxg8dkGp6z/jLeg1UfJS742eC2q21QI3yHkI3HX/G6axxtd4ZIJ/k8V+MLer7EAYp2E9wVBfkv
QYN41h4moFTsuG328EzoEwqlw0rIQhGmpRFLCiSZJGBrWtLCLO+GtthozZGYZf2y0xZM4T6qoKht
s0R6Pmsj6ePTQH46Mzjn37iGtip55Amw+C/eTSusuR1ootu+qfkfwb1PAUmT314fEUsLKovY/MIO
PINWefgwDcLa9ociLP7AHMECAjTtl+XjE4kXNCFQAXes/uEJNFf5gGAi0hFRDJLs8VlIdJxlPCLv
mqm+aoVS0SKqjucwxCJ7M0j5X8/ngOl77CVRV2EdZ7oosdtJccp6ir/rjg4l0M8oxfVSK6y9bZFD
G3hq1GgcwvNCyRVTdQrqj3JaQM6VRRvoO8VtporE2VS9RvQXL22Ktev5//tTl/vTAW0dD5cVCg1W
g7Z0lOjcOly50Hx1VF1v8sDxECtC5UorT/er4DicIPYxVy3oKGf10ybv0/mcKlxBnXCTQRnmyHNS
C3hir4QdLlPFxpVfDkAxo7YI0wD70xsUDIK//aPCEn19LKDDF9PlSIoBFTu20CGLkqy9U3vcUFvK
MtE/Zy6GcT7jUm/8pYQ+I+BAE0JLYORcni+NhIIv35tsCoBRztnPw59VEZEENq41yRHm+FS0raz8
Fa5mcHjFZEv73OEy90vbcYTL5GNiWBPoaVoMFG9mPkjvYVMI+9Qm9oz9tsyZPO+xuCpavobCsT5U
MbjGoaogxCIzPZUonPIxUUye7Y2xCGJICM9keqMH1qOV6iSA8iiYLVqyOtX0olqgdQIdCrTkrW1A
Ukkak1BnMP26uYVh4uEEajOIAbLk3oafIhzLyhkrnwks/PG7buzH71BBuzbA4ilIkpMo43FDW+NH
TAcaJDCEy5oX8jRVUcxHlRWYb2Ef3J3CEXEVDzS+Woqw7RRx4WWxKny4gq+BtwlgAvPZwXthtRjX
iS5op3a+f8WqS/rhGdFde8Hi/4UrcNJmF3jhaR38HwGxweem9FpfF9id5525m3p0GwWD0cLrtkOh
CZcdCw9mL24pvGeTSzW2bd6MEtIn5+qlNZjhk5+8NPKzKRWfdKLBPTtbn4KCdIcXXNaywmHEhSVO
FoKCsRSGbp0g54yt6UEac1An9wmbPzs5Yh1tdKUrvifs7L/kavIj3tQOuQSgaVCs8DkiJj5PGARz
A730acuZKmS45uT9sOADT1xYftG2o+EuAKGijDjdU5PN2k8RbDOP4zIF1APqkbhaXcbgN3TyWRCJ
m3ALjbtsXM4p2HLvgdWKN1tyq1MIL5cALj5IT3b8+lPjx0W6RY+WmGcmQi2PW8Ut7dMTuafRfb5Z
v/zJof1Z8tpdze64ujRiTKkBx3/H7/BVzg+PEjoW73Wfyv07mkzQRal7X/JYDRV6nAn5Ii2KdTmb
FyhWccsaSHQTU92S5Fxvk3uWzrfNKQ9umqY+BkcEnqL0IX0S0SBatkCWwRZcHpiIKuP7zDDfACgY
oeb+jMG96L00i5smE61RPDmUmS5IxW01oVB6LWTAwxnvhg2o1Yp1IWlXNKm0aaLDx1pTYKH0Jqhy
yt/OA3KBaDZiLaLb2u6LmR2Yuxq3WzNnTT+ep2W52Zy5yqMDHHj+p3V5OGxsDQYwejAeqhkQx1Xz
h4js/qHJv7Gj76SpXHYuSZcmbACASrltpkyATq4RJnUwDECej1Ffxy3jnFSK+SzbOtOwrzFtp0Ng
jhLfLmxQEc63wVYnS6zcOZeue5vAte3FUUV2GvDoAKyMAITTMFYwsNWUigAkXKyRduPCYvzz8wdH
WNQj2RPXeZfMFLyz4m/H5W11idSoNLFHuZOTRMho5Z67AAsZw+nrxxk+hrUYg0uqn7F7e+MMjVsg
UoTydOCSKLaTIZ38tnno0mRmnS28bMgZ7WjuQK5zsbaBXRSBwFvYJ4/4B0psNYSKWGQzqb6L6j4j
Ttcta50uT/S5QExhzIq1PF9LEIVN8xtHCOSrY2lAzMdoBcq1c1efrQCp3bbEb4IQMo7CnfUqCHKA
5HFVEr4ECbHJnM21mVlaIf3n6rMVT/TY+T+KYY7GALTN9hRDeuIxP8YfsWGz8coGg1VuNEOXnIyI
+7dsUH7tkbEfnE1iYs98hd0exl/lFaMHZvzP5Eov0NFbrJnIdsPUXDGkD74Xx0QfFh5w242+Jlxg
Ocg8DFElp9TGftgr06BYqnw4OxK2KjeHWMu70pRJplgoWEs0OaIrWaPTIuLuLkoJ2zOIOr7o+rxy
ZSyuXvtGXUhkQZqjhCG5AUs42oZmlyDe7wcyB4T/gz0VNQAqsVkg3pOB/tS1M1CizkDrN2097C0L
+JghRUadXQf09Ifg452FqvGH95m+IA9gYrsdYwwNBP91x5owVJpSaBistwAOWyOm8GOcVmI8fCQP
JamjxFnC197kXmJGStUsj652C2fl6PVd74kfthRS30eVqCgKbAYOMWQc5wZGUTqE6CDgS9kodZAf
2NFC04e2TURlXqQN1t6TICdEhASWU4N8/pCnQDoAL+CC5vYlrow7Iha6y7V6+/H8oadmlt/AVbPQ
0MkIcVSETufyTVO6t7NV8lmca0TYqRReV55pzDRKdXBiljKaBdD8CWnmBdO1FJc+rlpwab1P7Jx4
O+O2geldhMLx3hliVLW0JpqYXYlf7Yjfr+7nQykL2iuSZb97BWGe7kT5ZzemIqEm/ajOMm75dW0T
UxIY0Yse8AJCCTQh4DXWdvunP4pzElKK7FX1Xr0SZOEsdlWPYEAsy9kAAHKTvabFZM+0OKWr1fYM
0R+CSMswz+U0cqhOuG3K6faZf2nddhMzfH5u8K/tgN+S3fKERZlUIx85l6+KEDze9oeEjmEEBfSY
jdD2O2Xr05qWZ3E0JdtAHsg4DYaRqjULa4UDxmzMhBHy4S4wFyyQQXEekjeHn2eYxHcvOFsdEoFS
2mrCVgoD45TmBCKWeRLGOFO9mOubDn44GYlYTZ5yB2efhOWolQhmHFiHB8JbVS4chGHfAG6rjeTm
0kcjbVUQkIQ8kwcTJaNxoXMViS9jNwkzvaMyVglYpWXV7QI+bdRUQx6KimP0bzaSrKlKhygDWF7J
B4jargew+siggSofXKeFwJqYcYMsvS8DaDMyx217wXxBnYNXK0nohumwL2Gc5S98qHEa3cndQDFR
ZRw/3w5gKa/AIsnZnEhHy7RH/QBPgAjAOFrucNtKfsDAzm69kT7YZU2hoBYjf12yA1Gq43W/DyVi
oL3zCgctJ5mi8+SLeyKGrNxFxK/0rsHghBMlRV9tGLCw+exmSZrp0i7b0j3dhRj1cSpvFamoswFq
JaxSjePz2T51SbwynDAHb3FHbsPZG32r6W8/Cbb8Cx+bKOhUvWFNqyv9QdNKNQ5UDcUUzvD2f5Th
hvutJxFCYV7n/ia5h88WGlaigGbX4AC0VaYv0bSqVt5abrPUdHFSP5RqAyOeXXLjkrmH1AIAg04E
wzvqgpKdEs/q/LCwKfY1rmeRW0fVesRflVd5xLnRf8LlbuSYu8TwkiIGO2NCXU6dqjTOKjWH0BbH
8eSMBGCZqr1VDOZ2lZzqPlMxAJSMlHqFH65O7SyMnpZfWO2nowUkNRL9jT7myuoP57h7FtAThyGM
SUMSqpCvdZfmBDWQUTIVPJoPKEhyR/g+tkAqC8KHSd7RUEQMSwdy4umEQVy8IOE7+uSCw/ddmF3i
NYMF79cOQXOYV3TOmBYqY2rh3k4YVo7SPC6h3rD/8c6ZEDeGXMuScRCSLBwoW3KZxaFZa0XqU9wM
AamtWPci/as6UAQJpLf9g7g6SvDZDP3v7IOpQhhHK+hMgsLLjvgZdhWH/kmiwzNk80mROlVxpjr/
jqecIF4kq4AoqGr/E0sBkA56iiOBFbWsKZwLV+9kO+1B8TbdTY3ILjPb5pKBHwSQ/dtD72CXG75r
Y0m7u+ZAYoJBcDsfWm3+xd/8O9syI+Zm1eAjv/5P2O/QAzW7u1Apu1q6VHQiBnsseb1p8/Rs2KbM
or3vNwoKq0e+XX/ZqEwwID/KYBc6w+aTCCaWYc5eroJ4lMMu/6ZWc8ASzNpS9M+8kAtBEnRQMAN2
LBtKCX+7PI6Dpfq468tCGHo2iQxC8u/HXLwIwh9d9GMcomjHwXCqcFIkxem19eiULNLh9+NbqX4c
/sOaNCmp+B4XeO9NaL99barDE8HbAmJbJSKtfilgfm3M6F/38vOQ/QnjG3DvL1A+Q+KAtUNW9HcP
DFVnzQxiPOK6QR3OOlre6YrUqB6f4mp+8uR+iJYbYdHN3xXlAU+f5ufCFetvrnxashOJq9N+y9jb
/FIXYK/6nLXu5IrfoQVrGIgLhXJVnM9K1yWr58wdp9Vb0mdACZFuCE28k2n6x97Yzyml+iLNhf54
RGOAz6+/9Z5SZSbRvQuC5ZTTTakB56Pz64cz7b6JoA1Ppd0wuPVyUPIQo+wn6tTW+aCiD24PPrn4
Y1xn4gyzxwQK7LjnBCsd54dSgyVfaTy6TP9Vpmj2lK+YoKYB3uHTZ+oYduWEfoXbQNPUFciAy2Jw
SbtlqMZIKt4BLWUO5f/o89SF4bV6a1LG9OilWdEyx29xbPfvj/hh3pPXyBPnVNmzxk/do+CA03/1
kgJX+8vdeKxps5OiWPqkY7ffydu/hUrmPpXTyrRVJng77zo6QYX9ODlJhbHn/4Zp0OwdGdaSXrzL
+72AkTaMsDNqELoQbusyQssoZNk7bXtRQeEilr+7uxEZ7+CU3RGGsNmtcOjFApDofU0VMCZX37V2
OPNEGXHr8jAdHQVnJ7iCkIZI1AHAhc9llTAh/CwcVgUMj9YlxuGLeGfSOgoy/QYfo4FekH5TWgXi
NGvnP4AOocBoUrti65+rdJtBf9VeylStC++dXc+NKwk4IY/EYx2GOzkOyl/SjCvf5Um87hfBuHZJ
fmb7ubYK5SLDsKOCqqizlL1pAOElA9A1rqlNflKKyKbYVFUJsyJ70/mAB9WKNJDCWqTjsUX/ZhN3
K2Gp3tvq0tm3tm9ClHoQ8DGHIy6iS+srSxld0AzIkSpMKxGH6SWunmKaECab1DgwBLfai/i03yJY
tV9YipqVh53IYc3nj9W/0K6awrefjNUEJb0SojDF6c/uvsYK/6Cm4vT4ndewLD820DLipdxddDPM
q1UR0iCGoEpT2EaxRa0nXRZN2TDplr7Yaqi9MLsK8suHzUY5MJXNdEhI54tyAR4fReoARtHYDVsL
LLkM+TPNrcgVT1O6HTcVmxashNQMgvTfcGP8pLT67KNSpCatckI78vULA0iKzSb3Kjc48IIFBrA6
il1JBJTI4k1RAf24oADFDqefLh1Jmll++pdxb7XmxRgbwfKnvOZaVHb/J+3FIbfEmdpbwIOuTEMx
1qNgFnrEW4x9lrgizBzgyduHmblkwTh3+M5VUM9S95ua/o5GlHfs8Mvenh+q66HNf8/hGzkHl4sv
3sb4lQebVisa+1uah0ZTW0NBy8NF8B3imZM2exT2uxCa8rPn7hXGsrGi3L+DXa+SBmMs/rZ2+Hea
Mk9Da/Hq6SdV3LZ+b4ecgou0hsQ28z38idmcbsD3DLu8HBvdx3R6vWQZ3OfieRGlaOSnG43ihQYF
XiqOJChHP6NpQUeSXwzsfmJcufGijoCm+RzOu2XlHcCA/7fe4AQt6TRtW92orrG3waWVZ50J7BsX
CDMgKCqhpKeoOXks/EBZHy987NC/XczEUEo5u0XyU1X3SQf3x6s1dHaHAMCtzjPuHB9/R4Ypm5AC
xVsbAsbzXTcM2zAbGfCjAmED/Nl3Y5HOrW27ZRZ1TJA9ScV14cYgf31JVZxtT06aC+crNuxpgm6D
VMkhEW5A6KdCzIkVM9ZObz3qGrAjmktqXw67Wu0IWvRjwYESmQIxRjs6zZiBAe08KYNn3VhK48OK
/nwnGsRrIhE+5HR0SiOgKU4MZCj1r2e+jbd+zi/Wwx5dqezIcvYSvP9qteG1yN/rso/rWUvJ3tz8
nCdx/bzZPCA7tgP2r7h6eurkl3EMFtv/vx5+fo/lFhL+EsysH9xBm9SMUBuqM8tloa+ppLnWDjk7
2bDQREC3ms1xHUvBHwszyde60ud4wHcQgB7XO1v0q26n4HUcwIud3NdLXfTLh5ovFQXp2aHM770T
foLVc2xqAa3Id98MASfVRKIiw0iBJpILUXYDpjQOg1IQc7WUVOa/xfvi3OHR0PbqVf9tSN3h7CdG
4ReIe7Wd7PcrEx9F8gZZpiba+5l896L8qTperkddxeh+tCrWBIg/6yNCxSxA5VNYSViZT5QjZ43w
D5sF/NxU+oGXGhFskpm1qBfHIEZLCtcWt9EjivMAKk9meydk4dGPGAO6clRlBXMJSthWbkU1asJ9
UqJb/TdhiXN9yigCggeU4AGdgpKjFC+JmJyYB7sssn1tUuqYYMLM2AJ4uahVm8kwOcSXCmeTAfzB
lyH3N5VV51PPGvsoKUpr5IJtVCZqoorknR/OdYYMqOAe6AZIB9tj45amLrSBDvqSvE6h+UxcJ3gg
EkXxuJw9alngQRnKtqHQ/3V0J60YXRTf53T1auZFBWa/jaxNGYL9FVoQ4+OiIFEROwYMUJSPZtp3
KwzEyZmDx6Zlo1zyZ+GqjSScIbCuQ/QmeygkL3cZBKh99UmyDhiNMsBxlMu5KIQSfk8Ld7qBsm3Y
lScwpDx0bzh/pQzkTs8SESXKrz/izkX+tVK/SiQCEDCpQ2Jr/zvSbdE52HwGHVHkCb0Ou+HfkfuL
BDoTTKlexZyXe1if66mMRZzUbHgHwMNR7nR5FD72/MpM2ZBXSMJhpntVxUe2ygq38iK6FLRWLbYq
N6kf9OMfSrxSA1CKmEGEPR4LCL4oHBSGOYvccdHrWQkks7q4k3UdNnl6ZoJPD5Ztqi0fLukmjzi+
+l9C/XqxSTjUr4feoWZI/zgDLVz2QlKNV/45NTsCCdJs9eaV1EkUICvgPe2EqCf0MRes3AarmCXn
zxzJe0kiU0r7yk+DqorXX/b6IsOCOS3PhC8Sy8sS7iWmXYJB7qv0RyIbqQ5RkqANCguvpWd4VNB/
AWUdkcb6O8ppxwJjCj7PagKH5/mMyZrIFBmIi4LCbZ/7abyeJzDG4ue2Iigh2KYvAiLduco7fRYu
BxEU4mlIH8kVOqeR7vzViSADPyJogNHGBCLhXCNRcd4ff5EGdo3OIK5ZKz1c5FMpmMOHjQ5mg81J
vifxO610NRDabtYs0zmdyua23vyDcj03oAmHeIvFaNPazqwt8mF/U1iLBqyMim97dYvI9L6zDDD9
ctbwW8LViXRzXce4gvihahW6Fj/SQ+YbBL8AOeV10QwOqDzYc/SZK1JBbxTXuD/6O6SQWXRHQ3+4
dOilvAymql5iWPObTapCG8zpxAGNY1f5xw+kt07/vidR1WtzEskGtNsyqtCr/w5okHPBYVHv61i7
eDJWBNrV24W0Opk3MdivBDHAr2YxMh/QuofAbJqtWSaqFP56H3mHtli4bGyE2KN6KQJt8Xxoosyp
Zv8e/UBlpLy1NVGORisEk9yJRBjsX9jqAbnBivTH1GM9YQSQvdy2VH5kdpc88wlAwJwzHSzejotT
KrRZNDQ8WNpkxtAtmEXRBHegqpXAXY2T1biVqeUlpCWPijO6h0Umn/1WsYEp8VyTL6r27SIag7F5
BiZN2n4GfSxuTEsw+ds0NN2qKqJ5M20i5Nk6WeIkmPteVaaX5SpB41yXWUyK9RNVEszk4R3pJRjW
sr1llyhRJZ/IdNXK/hhLsMRxeHJD5LfUeFqgk6I+oqokyYufhbMpK0MkcFi+e0KexMBDTOBxS9Mp
vUVbu6Ba0ABYhFWw+8tU8KZ+aWvvEYBzZUwl9ggu7WdKY4HatybTakk6WuHNR4WdcVeHOoL8Lr0O
+6YuD+Qp3mDrO06Ihy3qPMno3idudT4iY7Bgr391dq7nMh7q5qpLwchynI1zISWeOqvdH0Gcb3qf
aN72kjEe2v3jwFH39LUCzs822MH4AHwC+zG4ktR6i2bA/mAdIF7jFyz+l8rg9WNalgLjVOWgQ1dZ
8+tYr7yiI4DdzSqKb2j/H/5ddcf/q2bVde0sAacwCXDqk9wABngo0GVKxchGGb6Q/UuKirra4O47
rgyGyNmNcxu+Z16/XzxoC/+nP56+mu31WxCGVJVqPTFHHo3rGM3fMt4mlRE8nO1HI2nptDLGWKft
1JGnJcMmi795SlWICYBw+9w0pHNfqgPbMHAqCTHGme9kMs09AB7AJ25LZsqUaq9K4VgHwe0w8usk
q65oFbP/fey6dA/s0VKStNphvIesy1MBqZiKoHdgMYcIsQrznuPUjm5UeVVcki2YDgADNiyl4Zha
ZyzxB/VR7H6egClf+gTmyU2xnh+Yt0nl6HVaWtfKHbGB0WbInjlCq0wpJBgGSjQCFTyjz4mMBLxp
T1XkMXcH+gpduMDkJwOnN+3c7x/1ov75yHq22F/ia2VQq8oQaPJU4JVd37lMyRP3WQBovJcKg3A0
5toBSlzMbmmZX+j7DJv1hkWt9Vwam91glWmv5KfREhNB3EjWfBvZacog5KV1nRO+Xifj/wLzvcxd
Oz96p5HxxKluCzVQhLoXEkHpisgKDlAob5DW87izNb2WqoQxYTBJt3ogXtPdQ+7TSn62oEL5BBfb
N+0gYeYsOTOXkenIwCA94+afzZ7/2iWx44L5DC/bqRDq0wXkBmg+8MOPJFm1dcP+YW50i+dM3Q/L
gnRC2WoI2wwfdiiNObA1bPBYsxWJ0j8yrqy1nWRyS9CT252cmYUJ1s1mgsYGfi/mOs48qS2a/TG9
rNgrUZdQcTZB1mLu8i4E6L/gRKBL4BkvK6vkOHVMPlEl1BLvkPRS8mJiSz0mUz37Tld37ha5uqwx
MC+UhkGJNfVoeaRgm2lFtZtN97R8cFIinbgwsC0D9FKCzqWlMWzUIQeiXuFGZeRK3MyMJvdm3ga9
pOyQj1wTDoP9PMrcQMGwWKdVXpKyskEPIUzti6coNdiMELeGGT2hXR4R7mIG2Mb0uhqaeCNR4Lth
+kAdxmkkjVVhIB04zR+gXCEQuCDkyIBtFiC2pjnW6TXsASqhHkBhimvzpF4OG3ReamMH44EhjhOv
7B51G+9Nin5aSCQi62AFdQCzDfwj2CJUTcsp8xcGB675ANHh8vDrVHiTqJ7brTbywtlIP/WGbpYp
lYz61tB5avYieF+eS0+vkSeWo8DHF0sv8+U2IDvvM8eXZXeYtka00bseWiKxnJeRw4mfD0EWiEXG
6IdYDwX2ImcMsgmb7TM6cMstLgBYeWKn/V2w+NaOJZP7stqcs8c1jJn9SZycTXXHkcHsx8WC+0Lz
tvGRlPdRYoNzuO9y6xxVft17iRs+XpnqKuC89b8zMDWbjprWpI+el5gjVuj3PDr4UD5S6WRzNRoC
CEJ+FBnw6HhGUwaeVkjw6GHwidjJw2Kj3WWP93CGTIPkDx1pjgtHdI3T7RNfFTvpLzJU6ajKNu5P
6u3BsMHgEadvxp7LXdL0isNmAjp1N5RQadogva/2E9//ouEeNqRiYtkpqOmH66a0wZAlaKPZh4fP
wA033tVjUTqs7tB97SUe91QYtk/Ims9zpVIQcWKOWfo64I18lNaJ9jf2wfcjkleDxPnReb/xetnr
72a0lvUakN+k5nTEtYKBZdDfXcA1qACR5LmgnwH/BklqOdpR5JAFhnPhEI2JW1sG7b/8xFLHvNQk
cHsyBmNGPlWfszvNLcSr8+VD7sgzARdHgbY1RnfdHUL8e/kOwnoVTtFl9DIXVjrf8TXCesSWXv/N
nBhDAglFtxNa/EJ3h+nIjshv0m2PLmTYLNRsKCpyJFr9XPTgF6AYr1Eesyi2MSD84iUxhuJQ6cO6
UzVp13WvOHnqcFrF2q5hHESsH37ugqzeMZM61BwTTELO9GF3qV0qRJsijyoaNbu0OyRXeco6Wolm
NN1cN5nNEUgs//g4IHnWYiKcAewFFjq2PP0RyDceGiZAn1wYbz0hFmrjyaoiGBnqEvqnASq5v0Yb
CznFC2gchDnCH0dDgIn61ktTl3nxUFv6CsA2lrqhzghsVuiaGRSNK8T+kO13TSBTXMqnlDeN+Mhp
bM4kukrqc61nvu2dQVBL0M1syRswPHdv1CLQMyNu63Jv+UqsctoZBtequo51UdIqyNJu30eKuywY
NG5ZO0szxZeNpAAph3V06ZmWXbI+wjlwu5KF8+f7IAw/qQcHiGf3txxtuTo4TGbim1lVRZXb+331
zxdr5HPgpUHXZLI1nE9TufJlw7Owz29xEUuTQvbRHKNeOnQSPPxFp3MeHgk+8d80Wkuinqf3vjnz
G8R+nXk8WnFVQ2Odmz7JVMR6yNGYRsnmpdzHcg9b3ceaQyUMqxrlDaGJLbLezZIO1Q1oYmQk+uM8
7ICS+oO1SGGoq8T0dOKwXgdwh+oGxZFLMLVksjNko6gdRU2iHzaCMMdps7PHAMzD9rXoIYBmQzwq
/cMJsh6+KBeLlx739Ln1vDECL6PXg5aeIXdXhWtgFAaqm5ICBbfALWy9264P+ZFM6WcX+cxHTicL
S7qHI4Ihfx+xliyc1YMe5Gqui574NBLRXomJKqrOgdlN0TiWKfTDgwyVZAQtqLZOzg8cSOmO8VbH
lpC2E3cr2OLuynsx4lhtapGivunCn2vMcjNOHHxn+fNFx80hvECDWFRvBWuHauF97PGcwvrzDW+J
o4HXeY285EUEc1W89B9NiAcSKR8fW3+Wa1iNvGd6W4nHXaMpND2wX3mDN4xoLPAOMzPZ7zERpez9
y+dIHmfYwp6AHfgaQkq1vSRYyHXL5t8MebehuLcE2fO4GBmEwvQPx7c39Wac/sjrzSn1R/1nlNKP
Db01hG7bR5uLe5EXm5SsNdLdvrL4ONERQavINa68eqi1Q3Qjh9x0oxvzdPUqx9RNi0t+1bz1J5QZ
AJPLuIv9DMCaiPj7QgWTYsImwElWvOdQNCgd2dvbeDytbmJbtMzGPtBwdfa2H92cmJhgUXWOm0PQ
G8PJVXymOSd7vDHEkC4uMdBhAArxgh/vvX/VeMLQWPf+nh8GJTVY6n0IWaqPyxCh6eqMbAGMvsKD
q3jv890Dx2jDj0KLVZBZRdUSDCmJlHQcuMRb7IDf5L7hWoDN5h1qKgVsmQLm2TnhaU48Hx/N5Zkd
KV5EEV0AHmbMNCkBw8PW7TgQr/V7/UCvHvJxnuxFyPwDvKzaTBfQq2raQbnLf7BOK4HGtETLPl4t
GAtZh3kOABmTgsgi8p673YfZDhItYQWAWipm2PE3goUOciPint7uO4PhQwsdw9i8qzvFDg1lVGzC
Nf4rfHllufL7kCSmJSPEnx813c9hZsZh/CR0SIicvatyPr5aOjZTcpsoC8SuGYQs/LYorP7ujvaG
rOnYQ3Q3KgkMKGWVV/kcklWz2wziO+ZG3Xte65z1yoxXv9K9a+hIkUM//nanuJ+Mjq/CkCRl944W
6mLoREf/txS0gtTg8jpsRyFQ1worfmsWLEJbSXEgvRh4/81lCfmf9ZsxL2cT9AFo8kkMbQNAqnf0
BpbpQxYe1Ux+SxwdTpwrWzLH2Q82+lxQhMcM4WsTKnj0X2ZB4KWLZxEeuGqXQTNJxVzula5HitUh
J+xGP08il41M5/03G5Ea32yXf00suT2Mho//L2ZaJDGg6LlQqb3YyRymolKBcfoX1Gqdn+T2NS0i
7Uwc40ODry5+zqLzgU4CxG3ejGzLXvCXZC30hotmj86XLVs15qH3Q5Y8DiWnC/jufe0v7vpn5bxC
4zYOKEvtfs3glYGmpomT4SLeMga4dpvC8BDvADAtKBKZW/EO5dSx/+PGB303wvZLD6WO+aS27Dgb
QVN2LCkawxoejPUnB+iD8Kmhf3hMu6c7jxukaVhx++qtlv6BoA1vHNATJcMpPbBhL7FVgRQFHm7t
zUClDoAufQbAXx/9DfPlD5ItbU8a0kd+eBaNEp2V8AQ6E5f8uJwyMNAeMllCqKC47lCgP6QicWwZ
zNcE6MIR1F3Ps+pBTqnOCRwDTwLt8XlVvKdyr1unI3gLe7IX0XrZFsuSXyRgY4Qd4cTzhAlVPue6
z5z42f21DoW0Pgisbk+olC7n5FkAA4FxiVQJDk62AtnglVKzKN1riHsbk7tmzySaZ+Xs9QUwWx7j
3ASP2X2s/OtLlo5WR8IiwsYY7xnQUI51VGM98uJYyNRC+DcYHl4UykGyCikOKu12gEtBsCpND4/y
TrPpVJCgfN+1CFRTUBGbnXDIQd/moLp0jLNpzGAZelBWVpeQttr3oanpfftNaEyU4WPdTSbTUK9V
eIHqistrMJDZQirqtKuOJOW8Ghnr2GVBPDHRnNUEhjZfK+1TAwxop/G1zsEVPwiAYtAU2BH2r5ZO
xy4MpACEcfcW1jCXz2+4/xiTh2ztqDog9Iv5wyQx/AdTff7qoFkmpO0XNxIymXmtToZph8GquEkI
9pkif//fwftdqH9ZcdrlhOsE5rSB6aKnqZFmFwtiFYPFtsWtn1ki/2Kf32cqdXvR2JlIcaRt3zY7
j/XFYXUocDJulMoZvEyT1zE54qfS8iLeg0NX4SAYXOn59XAlIE8JXcCLVJ1tmQ/h+zv1R1dlTiXk
oTe/nv8GsaJ5I9OHZHF5C3L3xj3MrGGc8BlKt7OBmB0SekEKpuZvulyKPYVOPs6HCPCHQLlVc8ku
dFv7h9C91DiTPzTuBM2O+8zSBlJS1CsTt1fC3eiNd4uNmBYFGsF7oOBH3x8qqS4mpogqQnoPHyb9
ABYM3+KQzvrfIxpkhZheoa1/12txWCZr2Wz1s1ZiFRcCthY6IxwJfzqb6NczgItLMrfViCB1Qzwa
lGptN6c/Y6afk5KHPjvsSMT+QJe5CmJhqErJQmkSQZ4VIy/tWvDS8nggG0D8aXQrgCCTJw1bZuOr
qjobiJjMyEf4FQE0N9I3g1+Nrsyuy5DXdNgj231Z0A9G3suRMrL7aKnwEDxK1LAl+0MFZHl2WZSn
Hcncu25onu89LdAHh36ZKhpsJn5Mlbm9SJEUrk03AlGfi/VhFEI0rsTW8HGLj9eNEqQR+cid2H0I
TjFCrH29MNGw3bo6TSak3MGP8pQZ/87BYri0pKtU156V89db0Aze5bmKqen+oFwVlODptjpIPOfn
6G1VVyqTpgpP6XEOxrFjqAy5HYn1eLAY2us0wZ6H+XZ3YqV3cqERksGs4w6xLQLtUgcL25ZYWMkp
v/AQgTFanK+XshWSsVkSb3Pydq5DNw5Da44H+nr6NFlaS8hdZDYsK1E6Y6EQO2X/soRxiEMq/ROe
FwNA7AfhzSmvGack7mEMLUnBQpPSzvzYyvODHpQbDkBuAFbn3bQkOxPz80QU0lwUzmBzz2kIdhrI
aRlBHvzAJiZ1LIhrQHaMtTUInzNg6W+1lXoHQDT4aRK5fMi29ot+cLnzGCi/2V3joiQNkZS6x4jE
aHlPubep4PId+r7ZVZabLcC4kM9M53Wui0D+DFdtTtZ6IsE/LOLB7Jz13uEhUS1el0hhrS4Z/tO2
6/LbVMaVeKMMcxHTz45DfAaAAAgXWwXuKT+TsS09s3GoYXsFHKlBudgSPN3y+sc+OAUJ1edQVfsK
AFhduwekH2cLNS5BF5uY7JW9MY6vdqs7BfoSKgqDwcSMncmDJUxbn0LLuEfhh0or+stFFS8IQy2+
4R1tTtjLT4CN7f6b+i0LRGlp+Zf/T0YYqhwTA+AkK7JEszPQFkudA+2b+QDiSHg/nIIJDGIXwHFa
PtrAfAuzGEOTbfDMxb5CYcaS6OSASfuujYrL76sgIS2BUZY8DFmua7MtUaOK9xvcudqM5G7h2eA1
vlXsONo9n0NhLWbJJd7lMQ7ZOvN+csDV8nseRlicuUfRV++E9BBUbXqrBq4qdRtuEovLN4y89XSZ
6HhIPReRSYv8tWzPKmr2V6M37cuGiAXyongUR6iOz08Vr3Cqwk6k2wlyVRsmw8dkCCKbtumLrkes
lvrtGkeXNYnDxPzieyTI3i6l7H6mDgz/DTwpmqrhNLsgi5yjQHQUczJxzQhdRqvPo6EwHv6s6Rtd
twpV0KHJS6xWkA+fmXdZ5p0NMMLDC4I/uoTVuqwYfn87d9UU2CB20clQS/VSQaUwP8bWP+lDpiWi
iycPF3relGiU0dllJSIBAQJ0o2q41bk/C7wV8k3CdEhrbz5GyZqKhOAlS0MH6l9PTdD4fh2lJSay
2KTlujQcighy5rlVAkGXFQMbHzWpQFyzVjU5KgC0f8sCc2vWGBJXfbuC6RBzUoyTT2L9TMNU8hu3
7HKZOPqwxX+gL5kfPS++6dv46orhC9PuSFokbAoNlCkCmC8xYe5HubXMXA0KApZiaLNUlJNCxFux
gPeoqvGYS0/9NnejqhpzZjVVg7bOVXH849qWhiJl43DRC3c2N6rw6MnwNx52Dneu7k0lxakTRsTE
ZX0jGxoRETU/faoxoe/8fPubc0rNgBSFY8OEOn95mbYOVQyM5RGt8R/zdhvDqEUjr+cqc1wxSXUt
ZVYwqFKDtBmiTtNDy/vrOtt56hyCIeo+JfQPY2pS7Jd4EGC2+WGqEPRv0GYo49t3eo5qNgMMuKEg
+hdG5P/QRNh9nQ8aAjBucflMHq8mxRlrwbWABcrLd7lQKX4Zf/9D7zoEqnZ32XzyN6o35GbEnoQq
/3aM7TSDHPS9/97FSOIoeYlq3H94ZvXc4d+7fLZ9P8UqAH1fQcM22XcYO2UxS9Chjx6dKYiKLmI6
mxrctK2T2TxzVu1lzaGxvXrj5sOe0gj9vLOFUP6pOtONRAJ4Wz9FxJBSlvRTCu/9QIsJXNHDMEIw
2Rtl8126cn0CReJQ2hnd9JbituGtrEk6SwCSuA4ll+ISnK9xXquGC4KGyJAWfy35V7sbyOphPlmx
3UjzOjqsNYqIj2SOXQyLRz8PEQBaOsjhlm4zg7kXXEkv0nvQedMh2skKHOHGZY/tVIg3yKBaRvXn
0gQKH5PnoZIc0EE0HYpSKYNECkpCeD6NNd85E+GdbZ8jN/81Tg4zweoEAhK7yI6ArnkqJcz/77Eb
cQ8hGIMsED0jjXpE3yv6fUeA/bb+hDRuJNIFxVQgXnPleiS5qx2JNMROtgFDjfaUQqHB3ZRNyugw
8YW4bBwiwFjWk+a+X7yZ5yHneVn2xRJFpMRuIzS9j4iVFx4JVnUoO37mGK1iNlol7obvWPkIeN1p
YVQyszRdC9yTgGusdBGreASQI+iFGG6p/gjVsqGCATsTtBAqjVYasgAiz+fslXQeLobj+AvPOgB0
oPIqFi7poIzYEosfqTZnrR9pZ3+ODQxM48Rv8eJJAC9gsTdEZ3FQNfhyCrleolRk1euvZ/2l6och
of2x3axLM8v59x2e/wD7e2vQnKH/YbdsL+lBqNBbErxYm5UEqeDBig3ibAHswWRyIyrbaghM5ZMn
Bsif5w2ifm4bUtE96gUpEeGoDTKftOU8DSCG3Z1JHLkV6mcU1hO86USrembim0HERCLjt+sGGjyN
eS7fZIthMQdWz8RQlIs7DyQdK6QFZxoBxfR0NAjQYdiYJ0e+P1Pd/pjG6IaOo1nri3+5uTrrY0kC
gfdvMQtZ3MBVCLGeW2Mt+hxBq+R9LxhiXPe73whuqDMj3FT8ZBvWOoXggw2zv6aoK4XW4TSWD9X0
3w2nD0vKIgseS5+ty1cMWreA10hDGvuNLmQs0tURgl7QccUfK0mXyxcJt5fGtYvch7ZrYnLnOopo
AgwmplT1SPwUcc+h3u3iFxI56Sys28itZm2XcfcxNZ38Kefi5/4oDm6kUCiM8yY2cRx2cQue5EUo
VZXfziS4BogNUSeVnUzdVovTlAufTTAbs48XvZbshGvZWoMRocA1n4PykINXHjzjGdXlDXpaldkM
YXV+dIrJ6FGf+JFTUkTC6qD+kSWnGUx6Ht62gBvBtgc7wGxGwVdZh2vJlrpqKapr12ih5jwdZRnx
I7WeFzdiT7o6nvK1z7Y0COsjylpFdC1ZRkuebvZdiQB+Eix/5GJ20FmTCGSC/BWR7ADJSSbemAF5
ptpVuSHy5kOrej7piiw0lVKmh1L2ARcvbR3QHpde67JIEOQX2KIxR532iO0oWdCq1NoSNvNKziTk
U37aaXu2shLxQgyf9Q22vncoS3VHr5VNGaQAbGPPljWaKHQ61zDz9yPmc5DOeXjaoZPmUgLY17Z0
lgzknnVeV/0ZjUlBCCE6am2nQGVfrExkKMkd0Y7/feIc3m4YzwqEHV9MaKv6UIQQ7YBL0vLkRUBK
jjjDF9M8dAj8apgQYprTJOz7yuI3pc0cEV2pOXOYKVusUdqIKqO+cAn+39aklAOeRDXUsCXlafOL
rlu1AmEy7sKJEGdgO1TsC8OrcdBPhwcwT9DQL9pIKt0SaISc+4ClMMBC1JOYEWa78dcovyAfS6/0
AkWTpky8HMl0mGaCc/LhOta/rUi/I4LOoVrrBydKDKgGi70V/YmVo/YM1y8+tdo9lf6JvwCXrMPn
Z5KMgtWs6f774gSi66vHZllVTHTghlcks3Ba1chLZO7vfc53J0tKNq0h6Nj+vR1UFTyMsJLTN3Qe
amN2sS/ZXnYwszs6KwqB2ZtkHzuyhUSYlmFXbvcAGKYurV6t3sFQzL0WvPIWIk8I2x9Nb4fwJ9mi
d2nM6euFOeNTTzUpZia1n5gFAvE1qqZA9ipU+xC8rTkJHrK6xA2hTpGcJXdgO7YtcRjyoh6/V8Jd
JF0u4NKQnhkE5qWSNJS/UGjHcgX8xuAXg5cICNUkJtcojzQ9iSZP3wsmDF+J4wRNhVydiafhnWoi
oRTaPDG/Ra4ippI7gesvpnjMC8yxFs/Bu7RxbPPZCsN6VEyYUclNIZdHAadvHshPBkiGspY/j7Mc
ILwimbtYrTCdPzXuQyq/vKvpU0SmwxF/3MAmHBJj/QkUeuYDrcC6Q+hqbzGsefecOPomHTOYyA1U
81ZmjTaJNnw6/FfXkHYcZSgXT0tq/NvvQAs5rfvQ4x1hwKAYQo6S4k4oO5lGJq4n4sI1bdthHI1U
NGD5Ef68fiy69JEX2Fyqg0M6Yr4YibV/uTnI1ITcazhj3v7WztovQuYTCBMJwESRjYkf8zhhmluh
eeAcc6uMo2APGumPoZQNetCmtA/fpu4hGirf4vrHL8+TpWjemidByQQvP0pAoxGTc+QAMULc0hz6
S0N5pRmq77Rou2TbRq4L0Mf5cilmJLeQ9MNiCnRXrCL098xF+OfBc/nJtOgZXIS13PiojP86C6Vu
AVuytj3+kLl6lUVpfnOxsB5V0JeEvYX2fKV7yjN75fwLGCnHS20Dw69n0S6G8Y642Odo3wCepycd
t+vx05vfQt7MJO9YDZBJcZIRV7yuAxYs16UuC8Rudham7vkXQBEBIc+Pk3HefPTDfxAdx4izz79S
D4e3QYPzVmLOxchAFTnZGJIJGlkfbYWPedzfPywSmHFRoFbS5Y8qOK6kmaYoVJoItDQ+dLe9jO/a
IJmbWukWbZMrq4ZZrS3uXhifGYqEHrTUHKqBIyLnXkAw2SCr0YrBGIbOZ786KRFhXVGPIWOFKosD
F6TYS7T+yLyEgSWsS20pCrowxk1sjR10TsXFYBJRY7SDSoxhfGzXon/CEGSK9zh5DsRTFYG26Abs
DJAOd8kuYSMMu/DSPP+C0HTGTu7meoKVFjGIFzzpdoCGT7qObBp6QpLGBTvni88jd9J+iQg+Efxz
B+WwEDkLbsiU8jdeB/FZX0WPyDeKaIeFVDDg8/dnDPlhKa8bsh6Zb40w9JOs/MzaI7PdvEYhnuMJ
wEWMK19jTvXnpG6iQN7SkohYy4+hjzZn/DAqSQ83sTsOxH/kqioA/DfOjHZanWXtLil1c6Eln6qq
oOwW0o5bNvBV4IhMQ935iNkSzUwqi+VTnCTtjapknEZx3xH1StRaxOId5bSqhswZh1iuDGI9US6g
WOJ5IKJxmx1scdWBdCsSyiDAC+H2qUZpCBBBnVdU5rRXmQWRh0TPAYgPlzMB34rCrST3NfSdWudQ
oq1F8tag4vRfd0IUsqZvDV15DPCEXoVU/T7Et54F5am+7wCLQIV5JFZx+KH0UmB5ZxiJTGd+i7tQ
N3BtHplkOW8YfZGf9FpEZc4HO7yGs4UHTIS5yYZtxUUG/hL495RCYuvB/Fj9FEiXGFtMKFiNOMvn
eqeRub8lwtWcrO8Nt+aHTUa/9vAmN4IUpfZSr6RHnxwL0Hilbtr4RxlmFZK9oobag2l8t5P3GcC4
N1vD0llj7R6uyvxoKUviVYS7DVghCmJfPpVLrSa9SDK8PYVwwNNVVeNqMDKLDdCG7qAHAFMuTNQI
bBgKzTj3JVfnRTbtYVZKVMDtLX0qxF5xFp6Nxo8eIleCQADJkNQ0hKywwYlBJlBG5uxM/tTq/k9B
ndSoil7MFVK66HmGb6PvhrzO/c3tycKpZoAQzl6BGrr05jszRfLqgs+w2NwL+OimUc8djzaxozIh
Tw3F4nNUGK3p6OS2cdYEbuSavnR0FhFy/E7LAXyaiJVBv6mZToXaRCknJZoIRATwVRLqG/VhTddv
zfeSlDAC9pbl+MOESVxSdfZthMVQAy9chX7KStwnDUtNx/DWQJK4llaZjjK8Sy18QbLdFLl1Nw60
5Uad3bXYYT1Ip4CMcbEsnhdE2Tyq5JttZwSLGZ/QRHM0i9IU5EGqtr3/AtMtnEykPZhpXfJt8OKL
eG7ZjEHfJLg8K7WUDYvKSt1xkOsEGn6koxPVB8UaCEw+kK2Pv5Sl2cpPvmpqZmtZdrFdIJNIubZi
WWr53U9riwY0DV3agR+CglLc3dh//rUuM1jIz6WqBJmE12601UH5SWRPLuaqNhD299JGgh59KcGw
ctqfOJ6sYYTpd5R1AZnK/s6MvUsWs0FBoQd7FRsx1vuvEjdqX71ztPhi+Drh2WK68vuqjd7CavmB
Y5ZDRkchoPAU1NUqhQpaFdImszkZY5fY3bHGlakTwJ7S8YFw1/GdjcNxnJJEwSWtdAVVDjAuD5Fz
WAk/pygwAQQJU8Ghtgazlc5SFGG/EVzFV8a5TtuowbwxqZ5mVS7pMfcIrXw5DBaBBCitylqkwlky
Ao0aJhFjmDQNbeo1UZ0+lxnTfzuez6Ao5hnlT0x2bvOdYawMhbKdqJ1LiOtFV5MLK5y4RLr8LXiJ
8MPPVrjlbERXuLKAt7nelHkbhb1OFSxs4HCh759SukyBcK484lUjqIPp5a3oBwnRDvMeYKIAe78i
5+8qCLFAhInYpNtLwiHFVzf16YPAlT/navX14eRo3F6PNnNc5TkqCe6eTmrMZBOYTjFo2DBbXDc+
IllXku9JPaCJTIzly1d3FBzrzEXGRd+uynR8ojHp5xw8pWEHP7dfzCoDd7fz34xM1K04CmL8sLIh
uYGwCn0+dPChm/8EjlLjsZ/x89nEx/BbENWMoh4jMZvXK0R5O7QYG87J1EDDIfZJ9v1krlbuWJ53
hineAbtYCuFplCtz/yCUDYhQjXsk7j28DichRXtzLLt72XL6QGnMeY//kuDVjct4s74ABgdolHys
kh7mg8i8Y1yhP90sRKZWraiYmzZqa/WjdR7k2bUFWN3T0CJz+v6WFZTKRuK3U1xCwSkLB8gC1/kQ
/fuGFDOxwGzVll/yuUOOE/cclcouJkPzkoAZKY1gtqTQLdeYZOL1pommxJFkXNgvLR0uz0X5f1Ce
GO37WydoyoAzEhCGVI7mCm8CT/l2xcl1+INrincqzqf1YAlojNKJ2aogsy7qEtclTIKzIvDCkvl/
BsxIf/g3tRx8QPFXHZk6dAJh/FzipsWM2nNjdpd8aQZ2ci3kggeD1iEZoo+p0Usri9AtV/P7c829
KeKGrm4ayEsqT3+yJqroGJz82zaL1ZAQdi4JVmdYPaHzSvC/zwfqRhMAxYIroxBhGKnvoWlNO6EM
HccmtrdEJd0v+2rYakXwyBW5QB82LNMK6oq6DyGhdDi+lDVWojtV+ciWPeW0Qc65vReASkTLLMxs
ptp0nn+9DKD2z0Z2UetezMloSQRDTFZas/6hlTBRB+mHAmMsHadGf5TtQBNLiPIVc3IgWVuuuJWa
lvY3Mihcz5SPJTOvNoq4sGnQfrqbC1nd1p+PSUKA4PPcgTjN1WA9qy6J+5Qb3S3SgPUCsHCRP+5o
R8E7xstJ356CtqVfBfD0pMI9LxubNUC3/vYrwFllDvpPlH5CTcKgiIUG9vfGk7qX2QC8wwtGjXay
0VCfEXvCBZEB7YZ6al2lcF18qKq4/Kh2SS39zMzQSV9xApulZGyhO5zPSIo2QZpGjZeju4w/ppCV
t3JveXvCzfsb6B28eJ2f3A75fTK7IDI6X65JAzyS8q6HoQKwMdcKD1QpN2UO9U5PUGTYFlnXLjbC
v2HPEYk3xX5St3+vHZ+LbWzIKRKWDcDN/RbotngvaXx30CKl8DivYRPBb6efXgGpmBarTBBbt/pg
b02kGHhrlKUucxvVc+DqDH0AhHWcAz1tzzpIi587Xy4JRN2pLx2t5gJiJfAc8m5WrV+KSQSVXOEo
LQded+Xu2sIgysqIxIkUtRKcc3uA3bh4+qG2RbMSAQtv1BvDeoXkn0G/DTHIxBthps5lSFwVLyhL
jYBJvtlIbHdUUKcgMkPdFVoz5TOedm3SiGTQ7c2pSSg1kAHguKWviSiBrrYcuFyNcsKvG0EPQNHz
axEkwX+GyGSpOSQPXGsaBuL6Non5wN0waiRv3X82vNXojouhCQ8q7fRJ69jOrwIbYkhuXwKX2Joo
Osj/P4dg+K5lK6fHgqGFL6SmLMrZGfsQ9f/WfQ1NkgmlLggArtcrN40yQprvcPSA4Fa4AZIFueVf
5r6L9Mv3MxR66Sf8i4pdkfyHs6ilHIlGgtxNgipwpuWoo5JcjaLYVgCYGABnNXkDoZup+ZuGV9gm
aYtzVmycWCWi4+8AI9DCqs14mWsvj92yk2zDkxyIPLuRLJByd/um5nPM9UA1sFipZwMYwTvZO6EJ
aKxyKvBR1qDjMPn7EDfHycuWy+vo3F103U2+PAkdaEaSwBy7U93Ij31048aODuTzeTXAN7rhJMv6
QdeETCxeSZ2rHmZhFRnE9O/S3hA3om5so0XiFmowHZaqzFj7xXkDZaFCinq6DDyK3lApaMM2vVxt
d7j0GUitVCh+gFP1fZ7v4dp5r2heyFF96VPKKKoylTpiQjNTy8UPZ67NTJrb76xy+aiS8BlJSJYi
rDk831sBIuAoBhmmb8W4mNCZkAcqTJGlYnzAKzaENHH/nuFI7WTS+hgd7Pehyj6O0WNQjwEFpeGt
QTr5T7u/YSoLp7rZ5O/K/ZBT9YoB0rkBYs0HjJQXoc3VwKndkVVBBfhefI7fdd1HCRR+J1BOcWU+
4mKsIi2/7vuUMhcS9OVM4WAG5iahtl9FJKof4e9Qy4qCD5vBsM6n1zb9Yuza3aUE9jhxRhjcEKF2
W4xxEQgqpoa32H8p8FBMddado/61rjHzvP7TePVDSI2OuES4Y6nLjiggbYKtle/nJ3IILPLhy2gU
RAsh0a/B8qd3vAz1UR1OtamZNNnuXCvMLyigaX3vTJzOLFfm2Gt3j2PxvprwZI9KahtUN3hbEH69
4pp+Yh3jgHFJ+8UrjjwO1bn2tO2Hb+s0mlfKdRnNEPYwJnzjRWTdlHaEHzwiMtE6EVp2r46xBrce
yiTpx8ktMAqfV6AHHuzqy9KPfSqOY+eMf/YC/99wS1ZvFi2sLOYW0OzoYPySkFU+frVHxnpxKOg/
eSsgBalzP11Y4F1u7jOAgdBL0QKNK3bqjoNazpyXFVRQPRV9oqyQ2loBaaueNJWsNQ8TMIZQsiD7
UF1S0Q+r2KrTIz2N2qfaNRQXm/p5QRZAr2SnzBX1B2BKkU0Qkk0ES6kA51PoPj4ySZHNhF6bI4Os
fn8Lp8BMKiPYcuDHuh/4IQNfVuUn365MUgtClLwBmeup0TkXX3NDAL425AQL9CBIo4Fjm4K4JDP9
IWTtNh0V/WmFK6EW/gsrh9XLgP/F5ny2iAn7lKTTYmH+Bzi0OaVnSp33SvKiyuYJ7TZrq4b2dfmF
O128fCyyGzjpe0oQ2oSD/+WdA/0EkQkvX/o77Iw8sCtI12ZJ7ogKVy/L/FbGvG2K6BEqsiNC4xZ3
TAKu7gtc85vEJAoWLjgIXy/ccfT3KA9wcJkb45eLYMYDpvYGChST923ZAQwSo2OXCYj3toTMgR0m
6q9NCvaQg65dXas3VCq2MpKCMM8IoR1kWdcJlGLXHgtfCK4PaeiTAI/hxJbNkFAUkoCAYIkxysq2
KyP9wgBrRp6pJKHRAnwnlxRMaNgdRXsK/NIaH71uqhFi3Wm99E2zFRPdUOFujsxjW47WV+xpCjNk
ZuSIuavUlryklVP1d14Q6fOIZfuRD2K6OO6MCJJPk5LC3CaPwLJ8uS1pKno2nZ9RyYbyvi5ODf9E
LIh1CuyV/fDDIcecJqGafQLVf8fLRzRrnNQWlULGoxmvz3JXwVqM42MG3md2/TpD5xYltfoiAAhT
QqYZvYDr/DkWvwGZVI98HYMyTpUo8Bfsnf6IJD4CqauZlD/Ans+ILhlz4ytm9D0gAgzS8lAWXcNb
DMOU9gWvHRJ0E3F8Wqj9nUyiu/a0kxUE9f71PkOATTfDDCfDjFPhZL9PcFfde2xivsivHO4I2ZJI
CsTxSnMq9IBH/3tmDi9/l4ad8auaFfu4sjKFIt7Vq/3aNMarf0oLa8paxBf6R2pVRkNZ7zKQ2ndK
UXp2jYeOT7G6Lkt27cAtfokdh47PiGpqtsNG8EebVdLaVN2WjodHSxhkjMYdddr3069f3oNhIeOa
LlCx01AD0y5o9+HpJgNtRSCOZZqC/I1RRBtzTFWXRN49qNuKFnHHmtQwdO05XaDMrRLcI5TRyRBX
ln6u7GGK1l0x5ps3Jqa78Su3kcdvUX2SM/z2ju7frV6Ijm9WuxZjrlPayghWYZsA82YcusoMn1I6
UyVMmVDIqusBgIdop5mF+/h4Kaqq4br5NbM1HAA2FAZwjbeUMYaqkJHdjtF8M/voLZAv+IWVQP/K
9d3JT4bVINW20v9awyBhUN4/gH9nVVV1beQyOFRvQlJ7Om/Jwxm9rfBqlA8EmbUSqkfvclWYxS6k
+T1T4m+K9VswLTItW3OhLWWqUGnV8uXf/bpq3hllIAnxmMoatnq9Rd0XjzqvjRqF4mXQpb35BzHl
tJpZj7rg+cILic/HLj+FxCZY3RGdm3jy0iiLz/U7ZRrndNK9VrSaIF5bCobxyeFmEsU7f2IhELVN
p0y2s/K8GrOVJQX3YiZvgiYtcPEBKjpPLnr4tZp5fyIZdQBSKrQESnGyGjiPYHJ9+5lTkNwwZa7R
m10mNmJUEX0J34JB2OWNvSjqWZ6QC5wiNwGqi8nJrNBSP1LTfm/IbfPrlLLgJXG3kG08QfQaFhq5
Z8b+ri5hQKBP8sYTMOqFFesxLS+06T2Bl/F8yCkzZ60RCdhoNN5EV2zXjbBCDjszoz2qUMVPA/97
ps6y1xrzWmejErUthuFXeoq3tjXNjUbyFv6B2fUL3/728dmrpKP5vlF93hVwy1ernqWriaiOrG/W
W7tBPfS7ASs6MFzlifwjjmVY9ektPoDKzByzRgHStZj244DWaUdNB4mBtGnNGalWJVQXrk0uiqg6
5Mj1TDqFkckW0CcTgWM54eCjavsP08ngkUJ66EONLI7Q0OehLtqf3LRTxFRws/aaW/m83il5TYkp
g1iZmguG1qCa5VHs09+F9Vjz8pB/HEIQztevdnpqMN0LjnPO6VQAGmrYCT1QHqzrsWR2KrVuNiIW
ObPAmWfMbjFJ6zgcIWFBEQuOlrVR7kLd2eRg8nKELwgUp90jRCMiRtReF9BNaTwyGbDzyYZUqsZK
wc7WCP3OXgsZJj4GvEhZlohn7M1IOlInmkKDVby6KGmw4IR3ZAoqcvUlAgQyD9ROQle+NXDQbibB
w85+GKDufyrPMzB5+FtXYLj6UsEhr5GyWF9v51sYN8dYI51rHC8oTz6iOpAgVkQ27Ps6+aN5WhPu
7ni+Sq+AKpTyD+wVmgx2ws2pryOCNBmkFwMV+4AuLsu9aIVNr6gFTkPkiS9n7+ryc/QdVXSkv2Sy
eNZIelEriqXqJ6W0ZOO1hCqORkESLb7mD3zs9JDPZ/daWKHFBRtJMty75Pj6QAe0Tz7UnBCpILj+
vZ31YDERBkpYo5wpKxNTGOc7qQvn0t4aGn5E2YTat7iFsdf28PMQKRLcHzZD2cBFcvlucxYndxRL
5E2g5zUHXTSzua0vyBjUkMmt44qn3yUMsz4zId5R24YFxXuoRMisPi6zv7JdPiesgPwOEGXSCiXl
gv9S4YSZCwWflY3OCGcLhVBPHtfVrdIGDFjeVQmjoiW6M2D3fFvqEePN90RBjORq4PI2F4ejS2q9
vZ026GknzDJ0LyI6jbT5OkjOE2kYFk77vnO1KG0eVsMhE8UfkQ4oDzxuOEykIW5vS+ZBp5G2G4cK
si7R9zlq9eedZTPLO4pDDbTmLgCdYIN//SN9Dfg9ql4N6ukArbGe+LWHZeIHyAEn1m9G4JFSl4f4
51RQymOBcUeWFnyE96U0TDtwMohqX1N2VJlAs6nvIaNn5JsIz2fO52huV+Cfa4Llt1UDDU8jjXIY
Ubm7wv2/FR12wVWhst1TTXBQt4cfLsyHuXS9yCUmBPVJBUg5ObWvc/gFaOOBvF/ZrR+jTw7EfRGT
7h59EFEghYEywh4/7x1ifdp3P1J3H2sWtJtHd/9Fj8CWns3/f0E5fO2pvf5IaRRcAxiCmYUvA0Pv
ydJT0u5wXsctiYMF/SjRpB2NS52PAIm4dEtHn7a0cBpCtROjr5jqNXxCVQAL4bVOVtk/aRNZ9Kkv
xa8nWtVYqVnGHqSY44X+Ou0rovLEhFPhwYXjzl3LmcP6wQQcvSHyIhUpIMJaodq/9+93RZsjN2P3
WzeIMCgZbQOyuXpwWZ9/lRCdIXBTDTpVV+Qj+VgcLYBi7dvcAkWaBrNPlDQ7/mOct4IC8KqfRp7l
kes19w7LLUzyBS2+HH51ENnQC5hXVjutzVVVjeOmdsJBxsqQZzB+dlRt9mSfUeWHSXzGkDIIQ7Wn
lA92dW9qJPKmHxhypUIIpRDTdDjAjfVk/K+CAYdku2M6kCdzr03YSfVMdRa7qKoXlfrqqL8QrF0h
NLGCtXPjS4ObV+cXo2Ylc2yqSlMpcS/UAYDOoscj/LVC6LZ9aXmzfubxst89+UTCY6udnMEqZnnN
ZAPKl7pSox2YjL2ulQOuG5F3qy7MO+SFcuNhQVnXOlbKfypsyn7NucUf/M2fUsEk/UPEdjjfCHcx
fvzKvVwaXAqwoqw7o8De1AiDFgBUqbjzhLAuJhw2CqdSL+XMZFNBKMNF+4hBGxo/nIueRxDnGjFQ
8Fbwq7wwHoy7aY93zphn6WuS8e0+kcvg95Wcz2ktHxfhvXrMU8Q0fKlPDPjFDErvD6Qgp8NfIyT1
vow3BiekfLC2AySkSEW0ecQJUNr1GM5YsfaQevxnGfn3lokDAQ+8qIviYI6GAVD2G3Or/PhY+33d
Tas7NBgXg1AvdFgJufVJH78lxyJadNIVa/8nxqcdD8RYMwgzhjnw8uj84Rjm3aTTWqVh25Uhszty
S20XGpCokXPqo90WfExU4gEL+7KXJCFnPPGHqYm/A3tBq7OYEkWbOEO911HBOvkkwFl0WOxnpS9Y
BDhp9K5Rc35SM6cap5wdsk5s1Gc3GjkCNDp2KSvolSGGkh7wer/IrcjQHT6AAMAI4I7V3q2A36XF
Ceu4Dt7C+JCSiqY+xgImloPaXqoSpZwfuKJb4y7zsx23IOmXsYUTQiA7tPRgLhIXopW+lZMQvLaW
D/YKq2P/yTLbAS9PL7lUR64+qxN/PZBwuzThW1drI8hS7u51ox78Aq6LnLsJ1hLfwYz3a2IzHruE
yRAnUmTc8birGPvZkZa3sPBgr14SP/K2YUONezeyKK7gRyNuXjlClpKgbgNpnPtZ+P6LoDmxS/7J
33c+q2hiqQL+hSbj/QzeaVG5uaYARbodigojUH2ZuYoGlS8vh+GLqY+d1sh5g3Wgs9+iErFqaBdY
EX7eNNuy9hM/RXsy5fksT58owKcZzMnsyFUkBu068goB4VlX6YY0RvXwmXnHq5YFkTY7oaMTWCXu
LunYtCMIlUYBLV3DBr4cYGwJpjtyJN+Z9lBr11vFP9w88olI9TuqTIXQYrA6/YaQfXbVgRuqNgfP
YvIAQDbvQyflqnDwY5HhW4kRqT1Sa7rNfEB5VGBViTQAAu2hHwjFiNw88SItIpPLdSzBzlAmkCUi
7psOcgxdepk8rsV8/6WbteEksBHLKEe0aX9RX0pkflcoAfnjiiEG0wCKRmsmTIKTaSQH9pT/mW4w
CkiQd7YgqyFMonZvWNBoIWZxl/Wd1K2iuBD36baGfHVWJw1QLgAj9mI/qxfY+M+FmDc7g9Jz6skM
kI3Ua66PNY3en0isNgD+d+sCCWYgY5lRarq/d2THNHUggbKXhXTW0Awyg0rG7fyNf+h1nVDC8Q3o
IVrc/8XfIWjn6vVacV0e13RjMaqWMkFCuSY0v3Xcc/MPpQ8TzhK3Usv/eEN/w6g89vL6oHnrAQRw
LDL9LBq6V2lbJw2Lvou1uzJMdejxWynDrfueZq2P87u49vy5F6slwbEQAxved9+u55WJVxlaKkWI
xiRDlgrNgj4uqEkFKcnZB8/FVlRTpWJ3Ajtktx5dxLZpRCN//CnTaem3JOkxB//3udKQaaq/RT8P
8BKyB1T8U+czdjLfEF5wuW/QLCSfwCIewVMdVizAQTgBZHVAyqxYbH5ejt5sccfRd98uUjCjMoeJ
yWI3fEU29sWyMaWosS0zmDNkqEJSZGEGZ0H2a0Lpt594O6qdDaMxXwkkRpKDq8b3zBaWLqECf//d
el+sqN+CTGSwTKeHq5g3ev8lqh7mI+WKdY+H8jHULqX2AbN8ieVd1vdKkrFrkH05WrjoE9p+vzbK
+9Nbmu4bwk/7tR4XGyN3NJGepgkhQR42iGdEn01j6eDk4wOi+mJz1/qnyYHkeRhf9RST6na+gzuw
MdQO+3payvn+4VQKITXSNJrxmix4zwEB2pbfWH5cJx4qQe5QKJp2rJRM4f1omGjctgrwIAYL7ha2
m2NghhErZAsez2Rh+V1/pgASxA/urfyGa7hY0aBumQxZKiGT2bHVF6Wq6OFw4IWCuE+cFiHUksTA
dgdX6gwgg3DClPoJkcZLGO+/kq7JpwBDVABaEP+0tcIgMHO9KG9v+k+sjfHLrX+zd0t4bmEsw8/3
/BQ4AAu4RzHtw473FjjR1PM3RNb3Ri+G1t4fgm9l3+rXvbO65ZbCNyTiBkusFdmjblcOGJQrd9Ld
2Z00q3aN9WJoNTkwMvM2t4x2RiqGCAMz/F0tz2OQEKgG4i/z+Jg4lI7gZlp3aw2HSu5GRU0btDKl
DH3/klNyGI9Xd5pfeSoJH8tHIJFxPxA1NVEiu5qMe7yk9GxeSoLCFUr34aLus9Fcw0Mg9YulX/Sn
QE1RpnaoOo7Ws+JVAagrS6pvFz2MvPm1C4cmlLzTdUu+ETmbnjeyQIfCONM47zvn8kBt9RjmisWQ
4X7ctcHLM3dnpejoo6o+JhhRuZo1fiRl4VkoC/+TfrqmojFFp/M6Ap5ulP9P2aKvWDsmMhwGDVem
yQhbUFxsOX1yqkddghKbKU686S4+uEkeoR/thgOvuZTFk7R8dsrxDfVeTexjguu8bZlaZ7xPPSb2
FXePW25zqWt7fgxuAOvmed7zNGKetoNeMEYJHCzIq+NTB8WK6m34MrAsokHU9BIng838XkhI8BG+
1/4Oxu4A/L8C10aWlX/UQi/vkesj/NZIBTegN5VK7QOxjEbpoKV/h3yQFrDj1YuhO8CFIEJ0g8PI
wzrE3hrRd6AHESf7C1PDMkjVRUnz5nO15LXPWxNcfC7fVBsPQlOGOM0kZFGiArk2ARrV9ffeICRV
W/suJlWKR6o6U4jZCMa2lrpp0wEcrKOWoNzQAlCRi4S56UnPBjbX5xMTaGhnbsnm6DXD+Orlfhia
WI3NIqhiHLtCqkZ6iNyCsuezeBWVibrh691aiwKTcRU7Y524LBm98jPkIiaOv7qQOPxVggF42gJa
25ApLsQVp37gU9fCNjvGrDuCg24YAVblUYjy6Ez7646AwT5mYwyqyV9xbyDOg2bsdWfC8eaZ4Und
ZCcssEm3+E4aBppvjqQX1hFXLkmskL2vwi570wdtbQFw1Fj5XHsYkgZxSkXy37qcNeFL0Rf782vh
iD9xaHZCINxcVr37m+R4OsQTGpg755gWuLrermjhdshIyalXuYV099Y8KPj4EGVUB8lJkpOnx9c6
srDUV7d7l5S0+Nqd0ublDZFzNzxKZ7E/0O/mZXPhCSmjCKZxx0/nMlD0Xi7HE+5xodpaVv95RZLV
FNxiH89ocnmQaGdT5p9yBzqB6Pdq74bUx8RU8zJtPbwPuRI42GlqjfQ5vDySaZRWn03oIGPrDJ+5
/s/QH4kpBkklRh73oF/pm/WulhooKpwSPzHlp1tC3U3G9plI46Ai/u3KzxgPWDCoUkJzwnLUlOkF
oAK6p5yARiAc5fNb4HrZ3DVoszYW+P2NfGwI18U1pHB8sNtG+h0dBs0Hch+mRqDw7ZhcW0Mowj7l
hDrOpx0wwFp/jgBcVldMmRdW6BtYAyKx6lquxn+69SLaj4F7lVgZiyrixLJnBPTTRyx/ifBvBJKW
MHR72AoP5j5HDIwB5aLP3AjACkWwWkmvEv6IEDFzUq20SfWNkMmogdRixuqtBbGP1ELPcVmhQLTu
e7qyluYQqLLr47EK7UxEJLnbIltE7VYce+8iVq5tkcIiNOsbKi9hxG1gM4NaTphoXRk/tyJM06gc
HCorxRDnuOtZ6fMc3iigvPbd+FBRGEs3P0aFCL+dc8w5HVMVKwza3KGdbdfm4bitIKHP4VJUE826
oInD2MYvAygJseik2OZ6AJ1mumAD4V3yidQK23zubXLivvGenLeKnrM/HFRWhnsj0RkoOVhSz9G2
EnLVrlExnsgdny2Ix3WFxJH1uJHvMs5FcmVUvvtFINLTnFPqOez30/n+dXSxFkqSHYTWecJg96r1
Vh2Bt8rcNmS1byb1gMjjOOEz8LHaW0mN8h4VVzh/T0BNes2aMbRg6hl1+2NhgtIT0iXO4gKNeZSF
5IV+h/CXAEbTk/43iQEr286C6WnSD6ItES9rn8F1RwKs+pd4indpdZmOI4ldmo3UNZSUcm5W+2Zq
bq43lII3i6WZ7q6XJY6nWpRtQfm13UAZ8mMzo/l6z6NnIXCPhHngtPnbeLys1E4W7yz02qwNNN9U
lxWMmKLzClTWwEvtwt6D67RpEYDbE/+qcQDXAccQWnP6Bmkp7jnY6a8KKnn9huiviebPPZRlDuLK
fvlgLfK+jXf9eqUYuoXpZKVbMxIyGuOhh93VsTywiHDDBGG/4N+em0RmgxcpXU2FNIXaoVTIUXo1
iN8+XTnrUfVhQ1+EALygo0Ysj3jEWbq7De2iSv0SvfZU2bIAqSD+kGoqsyOvYMrk4/94uurUwWul
kmJPb1YKhV1N79fHuozAZAUQ1DzRXhZQCdLxAxbbjSESO1sXpArMMhaRJiAIXdHJrm6BLXEXLrGR
VWcBmCU7lM2tUfF4/sXG4mlCXvQ9jVm0+EyUyzfHKliH4OVjczkrlFVPaKgC87tdA8cNrMkrpEtF
un6UtrvX04w85QH/r6d4gCwhc4W57cfHTtCCKOKkpSQkWcCKXr5t+++3lyjL9IUjygSW7PxEWTmi
xLk+0G9xyfKxm9p7BHdaZmozqbSCt4u11jXnq/AMPDZLb45D83clthWpkq1xllrFPqw/IcU17zTl
9WYum1z4ILuBou+LmlNGSryZWhCFuabpH0iO9UoQBeiTrHlT4ONbab+hRcF5G3qc+b2X3vK1GloC
TcCQGv3cWFjSP1hj7g2cHkV51OQ4VEzFmshXMD/xcLlvvQB92GqqxrbUUc4O56e1ZJ4rgOL8gSO9
I3scV1/6zWGGxOQGy06R9FoOJXFuVjSJ2DUGN3xe6MslcXQ/EqsuQRzKBIp7IIJcsuNS1tAof7sE
bqDgwYaRLlW+akVvZUkMG0vl3XIMceoNrVWRX6AGHo7I/0UBSXuopsiSd31u2uJ10sx+QNmfQWoD
ipvME9DbO4NXD5EENHgA2ydnMzGR10EyGufd56hbhPHe1FHy8k7h6zGLIosxs+YNC2kAc3iJ29Ay
8QfXKTDUHINedmbp7hgEFmIkvH/zZtRTiRbFHloSH96Whnt7ML4sjMI3At8dG7CoEbMrjgcOVTH9
tCU/cyIrtDsWWurT6kzLqLa7bKdZppuwqDH8hu0v0xhlBGGoMjuo5z9vqqaX12W/pX7eoX6876I0
XW3iDDT2AfnU4OJOFRfnu5hD9UV8fmcwtMnQmq0JGqjEWwrSB2Ih7rHwF4qcIMQ5iG9nFSKlg5KI
86VscoJxMPznwIS/ja0iwjSK22tgJD7krOd/n31cTGFR5FfbpKLX2RkxWCqvYTESLItkSqGIYXw6
vHrBcguxewDWej2Gvqqozv6zvvRU2niQn5iVcpz9xnjPVtXVgqJI29g5DTH4TpdEYkHZgMS+5PWy
5w/4RYBLI3q0/6d3h3cv7+QsSy2aOeI1T8sTc1IYglvreuc0os31l0ftoPTmCjhvvykx7XH6woUa
FN7uakmBZvXWk2PmG4dr1jpePb2JyzCkQHDcn+W0J+wjbF1+FkMu09jnkADFvDY3H28Tcdmcw8hf
surijpi+v9Fz70PR24AVkPp3tOsNqt6sXx1dW9BbnZY8+PV7rKFw+Htc330OJEeTNhuT8ssBhCrE
6Aq2qeuyLu/6MsFx4mpjD8oKD4NyWWtRFqhIEfLcsRGGQYTEGWPturGxBMjAWnbB5YL2tybvCDTL
ayUhOoff12MIfypq8Y/pKJnTSW7f8NpTsw3VqrSFQPkD8qyCqiwr1SQf6zuX5ng9/nj+qK6iqWpz
tP9QfXt4cY/wMwOq1yBU7P1rH5kzdpHIej2IF+JiECyDabp0mLDQFqU5nxBtRfvv4q32KwHaQcNC
id8HTLA4jbuBeUcEpiEn4qPbJ+5lDaWYfxH8aR2R5BVAWUWZERwmaweoHp9odlEcnoeVKpOt4Std
yY+BhmGjQ0lQNNCHGH5vRx891xs2lCfh1mSGrBKhwd9tEDsuw0VcbyzpNlJgDq/d8emLscEShFnJ
zPMU/Qj7FDiu+VuRhQb1atjVgxzBPa0nlnF3DCqcH58MdHAOvqedQH92Pjtnw4o1rhFw2l37SHeW
w4Eyrvi2G8diowhKMxwp1oy8rmTU7wquNIX10P9KEmNkGxJSh0USEMQDjvv1uKv83IMcjdJp3Sek
aBFwjtONFcmQF8hwZ6rZx8HU0TAS0M9nIhGj5rKWNOfD7H1j52NlgUSG2fl2m5kR6b+yyW2q6yiO
Qa1v+2XGJ227djajfG6Ky1UqpTneIbK70D9Bvsz6CjfmqWJi7AONoSbeiUISViBY9SPpD1l2PQ/B
k12QtvL11A/BUCyDEJsOaREJo1Wu3B6bmOFCG04Rd0i9+l+arMhfY6bY9orFjsbYbfE5Ec5ghtEX
Sr7IaB3cVX3sNdxkU21q7fOLfLhZi93728kkPTkruzQEo3+z7hdDE9dXO1aNPlVeXfhl+rfe7aYO
SETSvBXwl9/LKXmSwxcED3l51uKFAEpHq155TT++adbyTUvODX1VxTwb2CkrUhbnrVUrALSpCJUm
nhf5uPWtVzbWxuAmKN89mf0kFrGMa7EnL/hQ7CknNsmvmureGoENgSWlmO8VYxEeJ536sxdrk6fI
lihxzyKvwHt5TUfci+QzmFbVoLvhwEuBhDL1ZrNhFzcc6tlvoOhnuksvnuJ0QPe/I4wtkb+jPcEJ
EQED5pYYlNVQS7Ib1eQ67a2wFx2fHaM+2UbiCdLtLEk4cf45/kogG3ZMgHr9Qfc90fXIWVDqsijp
AvRUO+P8+cn2+fl/USV9KzrcVua6vtRDRiUs+ihjnTZPoI//9W3sE7Aiu0Y+eSu5tJ/qvgP7Km50
MJUWt3b0jzRnvF1AupJOP6x0jsv+K3JiKy+xnK2naa33Ay394mqXt4rGH+kXeV4GzxC+J/z/9TOW
WHXfiTPhR9B3SuIAhVcrd9zbjhaKoFGduxyeH26XTQuOjGRj1RX+TCHcH9Q+bxCUQhRfQSJYTHBf
PIxe5/eHuK31Li/nwmHbq+bcPAVMAb2M54vvbkckO2AYfRKIyqBKa07kzwxgRNbLRIof4qZsLhn0
4qKfEhe1uXfmDMsbg//8OISkXUQNsTzc0qSA//vVslFslV+THsizL7etIow8MySbQtdyZxss4aWH
hMyTVw1Vftav7VHq+YaGyUuAui5kl184z31aAeVDMCmTG+Yu5NmZH3zh07LnRDsa21n3OpZdquIY
+jWXHtDjUFOFB+cokvYLR7ShEPKRyCZp86zErg9DLDn5YiyFLIJRkVhIBO9eiXYHrIAqsoNW2EFp
G6quD+hyz2vzBW44oikfaPwD5pOkMfld4bXbIqtr/XmaCkCLHPoS7QGevMBZkxD1QGUIMr8917eu
HBRQQtKrR5iraNz4q/DuVz5QVQWkWzckuZC9T6kulOJwn8Zc5e2TRm3mVwkKUL7l+e1Yy0d9iSLA
8vvkUud9Ax9OxHOUGhm4yuvbGLU4e8Mg9LDlR68EPi3pkwMvQABitQXfMNuNgue+asawfTEE6TLl
xZ32YBqJCPQwfNo9QYvE36dsPEL27xmBDOxTE2XtwZ7m6iM2RJxcYaygnwuN6X4cfV+ytt9kAgo7
nj1OpjEfl+EkunkpmQ0Q0RjmiiEUVOaPYE8c3N8MkQDuDSkXVP9lbzO4HmUh8aTJ9WONr+zLtQp3
NSkwEVo482S6zEdKLcKYR4qZhJ5f8dqjZ7mBTJfLRjRFPA+d3JWr3YVDc8iJyRQxHwX+02ZVV9t6
I0Y6prghcFPWvVgIQzzI11Plh/niVYIVNRdLcM4zLLCuIodkDqcUslYJS6zYN9EBpkMRoWE7c63g
1dDhNSF3xk+H26LUZqRgrXYxo3ZNA708I8CdZBTn1Et+HVL5NJIPNCmu08kfydRY8/B7s12iiE5D
zYFEOxfm3lh+xzV3OxlSjk+8ku/R1f3izA83llNWpOMG52xPiUudLqdZZR5shL/Wi2NwtI4wttCu
0IWpxzczbl3i3Db7qipc5/azsQ3y48fQvYnPOfx5Sjri9JSQ59q7czmcV+gquqSfmkOOKIJ/zfkK
L0hAMzk1eJV9EJv6F8xwywWAp8k3jdvRvRhwaJQ3r0ibTL3h6TQ8uz2ASYl73KexkuKsjxRH9Hk+
/bWA7jgHcjiQ79/688l2fNI9ulRjKyDbvINJmseClRE7ZVBTyFO+jXcTYguTvrgrmFuZX9NOKCzK
ZXWpdRTH1gaPBsKkREhyxZNmanKBNqjgBSvbAnYCnBeRqke0vjzG0MplEnX2bcC2ExuGQlyVFraq
jvOa1QPqt/vJZQ3QMV7YVMPu9OZh20TnCruLdxmCp3gn8fzohRwBukkdyOqiGQb2STD5msGY8qyC
nDd5KEI3FOav4os5A3+Xvcy/9+P4O6BWw1SE0ox1IW/rF1IWtE5WOkwi+ZWgsUuCb7AUXqUmGc+G
8ZqZAFvZwney+cKP01AQui21eJCP537WGVFReZpvMAhTI43MPEC2PaeqAqnBwvfL1ClQ9C9Wh75Y
bAM7eUrDWlWRMoc2uY51O7YweBooTkrqfRatA8P20LrBlQfO41M6a6g3x+ocVBdsctEXsc1f9QdC
Vh9DknK59RqO2peNGOtffquBeqTAeVGLB6RZB1GG0M7C4jqKh027MhYb+Q9BWe6erFTdSNB+0fGT
u15SdQKmof+4qhfMbIdpQySVe7xO5vPE/4yyYLNHAn8mbN/xEBuT6mO68DVCSuW+C66ZkL6BJJ2s
Yjv3X9r0x68iFYUsVSYOavv2YyxS6PUJfkMKdMY+pUV4124hn6FgGliCRj7uH0MSd3EAG/7w1yez
7yQeKlkdBZWDEZxnLQGnyFZHHFnuE+Vn2zA3y3vI59Y/G8MJCzUQrPKGkV9wZlhO/C6PKADBBY2W
PItwTdwtNbxAgRfBA2fcg/r8EGKdHj7ZrxcHYRcLJuTnIFLKUGUXtYeTfZUTkWg101Fco43d/WFt
uGqsFAhg3DkXV6DfXtILtrdYOgUroC4N530Cehjkwdp95Jott2PeDIDYAu3Opb40eQWU8SvM3QZz
0YbLK8DLj0op0uf+JAwjifCeyeNNkG5BFNTZUH/Bjm6Z/8U6k8XlwJaslbbtTM/qXfgSSHNzMaXe
VqDQbAWGTvZ96DTBw/u/3Qvq/L2fqUZIDGSVMtxLL5EIqLfKgOCDrENbFV7UAgBig3LPyBGr6h4O
/nuGhG7cMJ20AJykeXWgCrtvWxkfuAkzNDN36gxB5OAH+CbSnoW8ib/4lU0i0HD3Y0w13oq3aR90
iKTn89Z4+Em8AUlX036/Auk/hWEbdyC06xlPCBq1zlgGR/amFJs1SvdhDLlXN7YUaI8VWe9SF7zP
Oa0uw10widAkR/ps9OpCq+T5EylMcKtlazeWHTi0j2eM6yNibH4wE4t91GiOizdNauE7+qGxPGCe
goa/hXIn+pT7xX6Bn3jX794GOoPYwJnOw/xl3ydjn/SHJmszCiFxfKIG4Vs7D82slYIlTG1C3h5K
h2N+CxgCjmdonfdy+pXtBTJWXWqkQuGS5Es0eQHV3YY4kcJRt+tBsjebvo1RNu5FVQf343snekfq
qbifPOJwPZb6pLZ1KS3wlxN/zXQXT2PQfl45Wbv+pNmWjAyDy8sT3sL9ppbVGJtXh3pGC0KLdcaP
EhYakk9ySsFp1MeeT2k9YWaipBdebP+VQZqNLa/VvkDS3RSL4XQQC7NLi4TRbCg9wdEYHeNYJQwa
RhftgrejR9J2RCrJvRpr8nQ8wiHvgSMiByheuTZzpo7Q3ynPSolAo2rrwn0tuXK20eoaCIZr1yIl
o922whhonM9lzp7Imn0f9uoJvY+2fIMFU154MMZDH+1njPiKfKzfaPrXST0Z6P00PdQkPFRxUO9V
fgv4vNF/eb6kfhHTqHIUSesfa3U5lUsp04nRMCFCsjSRxfk3+EAl4pIsWRhdDpYdjTpMFmV9z/6E
0cOekLeOi8Yk0X5Sw/UKsDgjzoIvVEk54JtXCVU4sXl7Ot53ZPhn5Eid5lNDcUV6H7ZxfPRFvD1R
UgL9NjmIu2v12YmPh8iYjNZxc/awtvuGszsmwuFxKq52wbGoZbEsXflJK/lcqHNcirGpQNXxT+ih
SsHj82B4InJIq46xKwVG0cmp+wuEOX3yl/k/cSNZYfot0YfhY4f/AvFqEZzm6PcDxAI9ajkwEMj6
53HcxuYJVLsAjut+8BXogwnHsop04JQmQrI4QcN3WOo9HtFOdyNaclDvxG3S74zGP8ah0U14AvrP
gClqenyr/NIbdvOiV+dpgERjCTO2KMudcM8X5oRcw2pGxZZabw1l0TYkDcEDlc4hKg3I+aJC5MU4
92Lr6U01/UvWsQd2wP0jyPTg0LJ66BX4J21jMCVVE2eHHaCFzM8qMetMJgFwBIw2tIll0v3CSNq5
r8xD7tbOwtcS+LUVlXfeot4CA2Hr48AH6cENh/btoLbzYPr7mnpulRkEbdFmDDhAe8ngfYUiAC2x
f/GPffNrKxdvk5B5usIzbTfjTxt9IhILXpvNIHMcxYaqC2XBCCzH5spYv6Ie0ItTCQZIlkJsiPXe
3wf4os3UcbVeWcHCb4ggEoULNbZUN0lIG4eOK0IbBGWgyZi9CxzVOkFaqA//aZOIJ/Mjo7L6ctqz
wWH7z5dpojwXhdQ/rXAhP9ZZH0eSHTx/+H8p1ryS8x/dPSA5ljR5v5bQIr3nDinmCriwTyqU+sNI
xBkYvXVhF5cbTtYjHc1GeDqxXI62fYyVTARvg1jJrr1PpYtGAGiIa6tqbN43O0s2oJTKHo2zXZMI
95b7C3zBDuIBF5JCeuTD59ObdKfRprcoAhWOViwvcxt64AIgpJUvTmqQcjwV2xOGq6G5uILM+uJt
bHqIp+MROcMp6P8s1j0xcWNP9t0IHF4PBqBsYq4wqOhR/hZrdwu94QwBmF1sS21igZ4jOxRPAtbu
gkwjlVdm37lyFswtvU31pjN7HrGN8KZDPXRpzPxeG0DhSFxjDrgoFFZbJJYWMy2E3KdC1/iyws/a
7e6UAbfelr/ZlHNSNgLgV6NEdBsfFKcxLA+xTV/AHPrQwcmpsM6puZn5CRd5aUcQwdw/xrBFgXbe
XDcUv4LoG/32vicQwgodfpjaKe/Nb3SfJpKcogAvSxiMzuOaR5xgLHKE7UO5okouugWoYyu7gSeG
Vz8SmPKlcqk8Yx4/MSysvOQm8K+h41UiXv+V7q6hB6HrB+Re5ZOV5Jf8Aae3fdVlhMyEDwr5o4kG
xldDKK+UwGT9u8t9UqICD2Je8+hcBfKmtolGss2Cgj9/jVsLd4SN6Hi8AZ9KIFFcdypjJA8WTsn6
P5dyfLPw/jZGALw4x/i0K5Yd9AQVypLcRgB1MWFAG6b6Ix8JZsbVo+ewYcYh0Tv8TnfKHhjSHtWC
hlHej8Zud+oSkFulfCnEFrtPIlUjQkjOEClKKi4+P43fSx+j9S3i6lR+XDg7mApXWaM0nWui/Gkl
JeS9j8aHWLnKYjTS/GgaUdq7GpukxS62XuF/ujfx/XtR1dCu0qzddzZdCsucVmiJzpCW5xou8RVa
4X6Gclt0CK9TcFMoVIHMkl9aYxdRXI7R71h9u3wdZ3PMNG3JHXvr4gQrM9fvGiEcXhE2LQttNQvk
yyGZMq34tG/BTCySOLqemcIyotGupHJiDHbw2I6Zritvm5uunA+rsf4qfCJm3EJm/MCE0pz3FTgy
xPTau5T4doDiAwCpITCkChcsoUu2CQ6jGX+HueVKFNuXwB6UtXI7/Kcn1lVEHtiisSbdoxl75uGP
YrIj+DXXvU3yDUvfDi+mBsCb8sf7AjnJVHHApctcm/XbayKvX0vB9VkDO+ZaYUnCSf9cLk0kj6wd
sTmIVJVsy6IA3Oo0u4xxD9LnJ897iM4jhJG3c2bYl+YedWFmUsNn04OlEx0Q56Q5zZ09GhHP8573
Dri6dlVWqCq4uUrN3e2eQWvt3YMiyROMJgqPhAk6vWSwFb+ZEQrYTJG/e/mRiSu1VuqeeaLZCrq2
VMw7Iq+4Y5XVY7h+ka6feGJAddqbsfCL5OKweqC7LEeQWP/I3uOzWLeLysrxEQyLfLuw+rpykD4c
hghkRzVHgIcj0VwaAP1kmOXnjwhs09Ne+DagGHCLP64MRQbh2hbMAdXcYJk+IdcpDNTe5JxEKgAr
p+OT2ZIT8zzksy8B76ezAu8HvxKxXA/FXJfutSCRULBSHT50w/lu03Kl8D0jP1PHhztjJXDn4x9e
+YwgnToaWKV646xpAclaJlyIJGDeIgCpYfaLm5fhgmWhoio5j1zTrcVvWZ9Cm9zR+iZtTfkj2tST
t8IUuDC5o48BBt63UfbUoq9Rw2nncNxmZ9eyCfFXgZU8wefL35uEUfUK+Y3Vbb1MCsbNrjlxoSA9
wyJURHBkNLvFPbo4JfTS1FsC0dN12FBHJ/z6IRHNB5k3Qun1AX2PkWrCDwTeBNXcBePQp5BUIfd7
SF2/kyYxGefQ8Mm/iTKCADSuLMSRRjO+KgXU3bUoGyTKVgJX3/nclCMgUpkYlGmV0oRSB+W04Dt7
LXAaEEVCsLr+JNAn3z60AsuXM50Eot5Swi9fHXxyUxTbbFlv9TkUrSekNiImYbowNU38OnS+/2Uw
r+nh8MUwkK2iLatOoul0PcUdrqSp92zHT397/JDR+7cfnQSqOo5LsLSpRogK7PI8Nhc/H2eOofXy
vavsuKXMTZAcs+SdSKA7TcFppOFlqMkrO3EX3V4TF2TVaG6KWtEJf9QUZs3bPg8qk6w5adGAZ/NI
WIIWo9pRXnDht/FUQPaZ6u0tT0yLVEmdOYTGZ4GQDVTxGx701LBN8XlyLzGvFGfmxPyK6ywBmj6r
82vpIMGkm+YQ6TyIjpfO9ZiL2ywdvqN0JmeThUj7wd11db2UphMGTPv+PxZCTMcPx3i8Uan5NGdD
HOV6uEutpI+Ap97aYh+s5KukQPb9/ypvKVmQmpkbDwSLOItci9QIc1ItqYJzdTvgMxrm9roW9MgA
Zhk+pcUxvX0d/+IJbled8P+K8lk3HXhhaVJ78JvllnhyEFh4x0k+dtSNsPmAOfh22HRL79sRS2av
kCR4d4JU8pAMZHfVuyDA2AY3zTGGbV1OewuunOCLVOJFKlNXuA6jmWpTnQXWT/MwHdBMCGxNrApZ
+x4yihYoo9uhIoKn+FG+0JV6ljkSkh3vsNUuUK8MGefWvAPX61NolLwsVf3BnbE2i8vQMJ4PkA9Z
51LjQ31TwBzQun7cB9uJu2YZa3zy9mOlb9Fgs0D4AXiE7rDD6NbM2Z6N8+HuF2NZBTj457n1EOAP
5zwYgzLmG5tmBo/0junGgYK9LG3zwSslEYlQ1ioBNn0vRP2ypSJS4Tw3jNdQeuNLFDzSMlLDklus
4hmZqwqC9AaZ6DeyhdKKRELE7iJfrdESLvAvyybjE6SkEtQRE5kZpxnXksQBZLYrYjfq4iSylGHR
rYm6v2iu5Ncc8SN7jEbI7dZLRgRxLCiCTLcnJe/fvK4A2jq8pLbIxm8PtBYlM1gm8bfw+j50+gXg
94DljyYFoy14U8nqs4mmM925nE24OGOORC7XqRwIrWHw2NDMdAV+O4mxc+NqYpfixEXtCHtVtUn5
qmgsjfCMcVxXH9jQL1jSxjEu4gmFLSD1VAgTzJZEIzpnpq7woNusdlD/f2uAbFnsKRxgbWYF5YcR
7PViA3hOuan53DrAH2FyJL1pux3fm09nEEXpUDmxXciSf/4/tQcJ7rzCSMGnrvPaNaKx3cKCwTIc
rnhxfnmBSeyZNMTK1KYUpmaCider/fTC71kTfCMWwRtULuIj0B2yEZmrNK9pJD3VJe/u+USoZUSm
CFJN+5tMae26Eyhy/Q9/ol/Za+An21eEtymomRJXOwKiBS+Mw5v9LJgZl/EFDa1onzf1serglCPK
MXUCL4X9O9ZgTLn4lujLlXkC1VjHeU0WSJ/HppdQ2rppM3NRGHG//8VtIBw37E7MwcMwOTpJzdNS
Da7kdJq7rQdWvpmyzrjQ8fmTwVIE8ywnl8a5Hb+WXWbTrCP3WI61QbLN4g/xXkUETNvWiowq+6k2
f1hcqnk3rRUcpCe0s6uvTUZNcN2VWYdFuj42KcsxvCK1spSmPa3TKBwDqOhFeIucwsM5UtwuRKib
knxDRefSoxCglBl70hrIMDd5TMGxTCP4BSwfRBkzHFOKgm/lSOM3AugaUdRHQPR9yRgg1oHlIX+0
9MCfuqitDt9gKj2Xq2CTNUZkg874ZDd7iFoZZUvafom0YNEKovkk+C4jjPmfQhJeMr7dw2OHT31r
oHTy/aHSloOCJPdZOolMoOKKKVnYHd1G9f7t90TCpDCl3/V3xsFAR+J5mSekH6aAdIwHZfkurtvI
niOCayRe8IDcOtOd+peB+5V9FEyYs4o0+NOHHpj9ftpSZgoL+tdm1Rl7m+zGK6NcHU1hqFX5Frkl
oB+RoPOxECtsuPKo3aD3/od+rqTH26WkzONS5+L0ZMNPzsyI5slhfTNIgpsa5Ula3+CRY8NyVO7G
sHc/6EheFQ7Cx2XXwG4wlf7PWTL5J6T8wZ3IPuwbHpEmBB7cO18E7ZWFQwToSzlJLKWuzrYZUOxO
6Hz2/KeV8J6Extv78aJAPkbaVh/4UoLDVcG5dhHAurNbItFcxkZCsU4KFnII9h29mOkgyGOTFCr6
mE1pLfb7TCWoY/HHW7Jr8S6OYi5+C1HNPJDc9Z7gumyk6A3VHrVpEI2COxsnfZNZXiO3vhYo+4yE
vLmARgrNqCCtKAnAlsecET/K8QU9CDNJoQ4Q32v32sGENObTbjmNn+LxUoQ4NbwhrHUFvPj3+jEp
iHweexQzeUYfXcmYtEV/hqQf/M3rbyWgAcplutzgKJx5QrnAVubuDIZbidDSoo2N145S8AEExCRO
lyAtexktXKXHIJ06NkmQribd8U6m27yvJB3W5169hwo2kQocMJK7fl40ynloji/OMJCcC2eXH5fe
Sm0B3jMLwwo66h6UQhkyfIw5fj3GQGjbddwucRSxU8lYYgKkpIHYZsdm+ZsqJQgoEDhLpscpxpFF
XQ5PvVDThaK8FbCpTGvj9QKR08DvQDHziNIKD2mPVvx5+IpL3y7GRVsvx5tQPDmAsWVK1wT9KDdL
zm0wbxuvQ2CrkqONifTzWSH755Gz/ibN4uGguyWh99sjz7zH83Gs9zHEcugdSFvZAkNUfdsM8Wya
L+OBgxXBXOJA+DHGFtXo07EazwNaGO/2WSYHHHZ1XjU7eBlga3GNoCQTfriOqIg18KcRvc51jIUN
emC3b0ALF2umbhE911eUxIPtWWBf+PnIznoevmZr3sPSEOY4wta1wPJc0RmKlVrx4OCY/4HP3L6t
jcUU/sqP0R55/DrvSOgvQZl53JEeIQVUoV1Y6Gc6mqc9jDR2X4j8pHP4A60ldLhL0ZXkSPB5MU9L
R/3MsF/iLu6Am4F8HuRjAY8k8Er12rtCOVlBUopuoZFR+/QvzCdkVo9RdmoYupypbgppaGcdFzLr
6+SeX1qOvBnlIPDx+Ye4IF6kWhxhXILrcD4XsnuPr7R/4Z3wZX27r7Ij3ITu5DQ2Pnrj7bq1PBOD
IMZOVo1/BHrAoX2f9/uVtbDRVjp3JQhLiD0e80i8ff5ScGCKuqWnJ9/BZybCqpaZAaqST0SFL9vU
2xPc1M2gAnpyZ6SbkDif1ejnr5nEHzGNgyPGmZGLVHntEw4awfWk9ugcfCzluCRUD1G5iPWCl6pP
HrTkt84fmgrsLVzEX9sRg5Bth6PsfYzIwFBpDX5a0e+md5KSO4xRAcOLcn19aCvCKjQSVTaTehkf
5M3Kd/3Wz4xAl78ufwZ+4bF4yVBlL5EN1HTufu9pjZ8ASjTwjpELvRq6E9qN7VjMPEacvIOGRDoN
tWXDhoznBugNTVX3NMWjgVHbinyUHPe1+DQBBcAjOnfT7H3NicGJgjiasdH1oigBbxAEd00doJuV
z6RI2y3MfJV8J7OlnGrGCcqE0bT1Ry0GKL2BfCVcdaIduRk85PoQOMEZSi/0Uf1YzwUkgGoOHaok
CNJmfKIuKs5wciSaeoE2qFI/H9fYppRKAWVaPFEsdIcAPu3f9swtwOgtjZQtPAmADQecpKsVAzXD
kfTAGRa0nGgYAGU+aWh7RBOo6PLnjbKIKEWFQaMqOcI5ebH8BFoacABNJb3heJue3/apBQ3wA6cN
5DPjA0yLymdnJl9hPw19Wlq7AOFbipNE8e54Dk1pFcH/oYwci+T+FdiVpPwKwF1/UccrMiaPYU9i
VQNsJuVzSxQStyuxofgppyYq2YExaAUVPS32eNGXsNyYuHhvPIXh3J3dDsGrif/qPCX/JDbYUO/9
GZM1QuH67hNSsvHQcnL5OrxEzFI0mA0G8jeLSfoF/pv+ennWn7OJjuCeBX20Gq4wZyQ0tPNpjbia
FVSp20pBRTbAqeTMNxLTdysPD3RCzfAZj5MZzh9cSsb98Qbwl6w61i4MLoa4Z0N0pMZeX4HjDlmY
LlUtjSAXkSLGv8nyHHVISHpveNY+eP3Njg2ZgfcR3nhaQN/Sjt/B1B/O7oGsKlu1QGi6upx15Vlw
1JJhIQz1iHFnUdQD4sB7IwmUQ1k5XLlOMzj8Y9IndHCuYfFDZsraWiZjl6XX1MYmPJCu1XMuqt2m
4wgpDcbTY93/xmd/YQodUwtfWeMFE/0bCxJZQAYNL/XQRO0dF3nQ995m4oj5mnSa8Bn//fW0BXsc
BUa1BUruJEJU+ThV1ZiszejUPJebebWT3EnB4HX6uD0paGVWjpUmh1y6HsMbX6gXxiYXqf+VlaB5
VcF26jc1i0Ja1+iqf5EvHkhzINkVD2/Qfh85Oju5dGYhsFTV6BqQkVIZswFo/D3LnEbcYlBrtPFd
aBVk5sUZuRTktSmKZ+wXH0/yegH8QpNctk+0U6ct1hhreBHCEBWm/ARIhxJCvfWzHTf+Vo0QT3xv
rdFcKqWECoxAqdyfLtWmDQIxXplmPHRYJDdsZTTp27jl+z6ksyB0FyEZG5XAa7NyTJ4tqRMbOWLQ
AqYFnS/k6bTBNOIZcb2E/uOZ3Gf74jqODaBGQR8hCAGTFq1seT+2yvJR1K03wyGei1hWTwzGsXIU
/Gm0311Ay1s02pxmMcn7zxuTpmeWyMFMf1tLxJ/iykU8lCeizRkPxBJIToGBFouTssbKCBem1vIf
VqPjfC7Htpc41sE6JkuIevgn03sWvgaMnQ5rtz/Ey0z6Hst6znvHKQV27aidRAW6EnUC37oOOkz0
AFV+GnwmI+EwyNPvG1eJe28gCO31mIfBzoOiL/ro160sFWLixN9XiYvhDpJHiZOJWHnd6MjGpyDC
vsNgjAgAZtIOInuA1JSlNSa7SfAkAgi5JYLy5ul3Cpcblos7KTWXDje8o41DufP4UIiPg8yRAtqs
UL17LgTLPaicNNYjq8prGZGoiKSnPh1JGPYU5ovFTJIegLpHkprm+HaAy5lgQ5kWn3/ykqMqJl0j
YeH1EsqlvJCiHdpMZSh9dbWuGLLie7GuTvIMZK8vk4X7lshcvm1mbYWLK5xgQF30rj4iIvk2Pcpi
Fvsa5ZDxHnIA7HL2iePhosXFNKX0sFI9uMpuw25z6cVubeS7sZ69T9tez4vVletYgzD52kQYHdOa
WOVosIqdWl4+ybzcw71kLSWlV/9NDI1kTzVxCELU9G+Gu38zjYLboolDtGIFFPAVRK3CtqxOD8r7
t/3SnJ38dugl/IFvWoHMUqUFYAFSNiMBRaNSrHSlE6SepkmuJ24mjInPnxOE9x5i3bZma9ehTeO3
CMUpExehsZv/qUQuYKzNeuGPozif8Hdt1P3aNu6MjW+UFu5Ok5TL75eKIZ5agPYW/Eu/1i48AGfF
4z6GQAG5mS7ZN+dh/OHTYDyoV1/oW178BM/reckjQYz6qrhcI+a5Yp3AA/pQ11QwLe2nlmZfKXWm
y76sLs8GP+A9m8ChGABJzdHEWcQcJ8PhYyzD3JYsR6CXAKis0rRTq9WNw5/JyB97ipZW1a/eKtel
jgaBpqSJO0WxL608/16VYFem6QJn9bVhuVDu1OCBKLHdHoBM9ML4D3uwgTB0xXH78hlfKiFnrjnW
34bG5exvuwCKTowdIm+d2U1rsaXCaLt2BwzbRdkJrkANfp84cqREeSferGbHsaxDGvAHStJ2sUIq
oB3uereFg7LJAVOSVqYr+cfZ6vMAW94VQ/O56aX89+EzSbiHdApDvMu635W7fCidarbW5GiAaLa2
ni9C788cECKB3wE82hA9amvw+MkbiW5l/EzKaPfC2pWFOWAI5OjzaAlROeYIf4tdfdHvcXWIN+90
TQpdFf3YFwvAhBJmljWCUrKmcshIYnta7xUG95HkTtGZOCTmbv+SdP8HxzCZcLAPFM2+jO/O+Jdd
Di+0EYziKSmBPqBu/6/nwqxCibQopGmZ60PvD6yV/dgqSXuifzIp82zLlU5wqn5woMXYLdbKIsqq
ZRmKnsZpnkF3R+jN4V63kRRk9d/nALTd0ExXFNY8Yy2M6v1gG8wxTeQN3tvhzN6cqmmYB4PhdULx
uMh9KJo6M9U3hWinj/Fn5TS7wUdtyHJ5Dmh4kkW7k6qgGgQKrp4q1AjKaSYTg0az+RrUOuCtRs1u
Q1Pwaz8UW3JOl0ww+rxAR5nNkFBJ2vfjrIi9Y/htdGEdp9ewn5MIwITR1z+2Wa5gX8gKkO0sb4C2
DH1wxDs23R1FHnxf24BBzBIqpTDwvPdv47H9ZXa7ziXx7Kn2gLPJuSZm/drPCZFqSLtDKe6lBN8b
rzA47qYq4615dt9q8Afq1sI3aliTZbWbUoa0yaV+1b+XOotjk5POZfC5VI1NYB4gQplVfAwwvJ+2
pyISEifmBiF2GwXVAmqsiFFUkWMnIz+bmdz67+KEj+P/JBPA0wbKZSGP85s+Ys7hh+BmZ9peSyTC
Yd467OwIM13aPv+2Qc0JAVmU77uZ0aE3CZDiVBM8qHGZDlSD1CV29jMVSih3FinPqxQES8Ml+yLj
vC2fea6BXXCJGxeurL0gA7i5TIkS7WCLin13ESt+oxWuJQMTlwHZIWR5SP8ksgcE8zJ5kRCUr/sH
eI3ISVcgLYs4LyfTY9ITtgkcgubITAyE0HBnWS0BE1QNj56mtSdtNrH3izqNf86O+9IpEgsVVKpy
orvcruQ4fU7vJnhSunadJQRYnHG+skaawiu7NIVAkmfKwLHXwM62tnT6soJ8YoggD7AJ/7BubmFf
RcOtcBsi2IPr76GDHq/7s2dPfNaQgagSgKBuh41EatQCV6CEyL3srGrv0ycztMGGjzYEEtUIJeQU
Px98Oeq+4rOvapaiFQRdh62jvM+/veqMf7HagWXWIDLxOmqLb/vN9geDG9vExvKfvMifgDW9NajF
35wqsw9FMuW+0dGDBOJ9FRVfWNl0ml6c9usZ+1uwvto7DyEDl2yW66gARj45KLQyUx1x02DrFbjr
4BSFb57j3xI7kve9m+aRUye/wcUflEMcjjhQPOboxnPpeVLrV20I1vCw1opilPaSDdBq9mS0wCmq
D1gRYzZOx0Crn14xVOKoEkmXBceAqNtiBbrsBGum39+PjdA78hdhorLNy3rFdgYDbqfkDuXds9Jg
9w07uh0lseVsP4+QGZo4GuIJyxXcfRqRfDzGgKrcQwFNzcLxQ9hbFriFooe3TnD2NbF6xV2LvMau
YU0ZTYVB9XQ/Ws3g6WbXRjKM9FGkjq2vcNa7PCEPc77ofRqk2IjYNNKI/tbLnpwxezJPaIeHSDpq
GR2TWxbSIg8iuEBbLmOxrFsIFBk2Ba21CiDw37c53uhDu8ubOuoAk/OJG5fC3RTbd2/7XzFGGNss
DtR/lHAfx2Eo0ORXWfypY+iUW/AYuVAP17l+g9rviFrek2amkRrC6760/uLbimtqIjWDtNfAsy0k
fdY5L6GWswmI5r1+SLhmzxR8z6JFVww31jK0H80iAeas6stBPtan+AS79nGnV12cPePUp6I32cVR
DTSqT5fZ+/GnJFgbXgwLx42mWGMao8Rb+95M+/KZtwDjlYn2RCafeCLTNfvARuHQLKJLkicSYRNk
a08CHvI5HGoCW75QDaU6+bXjVyNZCkIriqw3vmnekF1Jcv2ExodJ7+jt4YiR2fWS1FDRTDV5UBxt
Faj3cA2R7cpFCS1419fmVm/dHWHKYzSzyNMSYIfL3CBZ2ea+o/qln6lwUOCT1KgIU7z5zx/m0hF0
uwH2X3c5J0XAv9x2h9vfnSH7yA+n3wLeKcyWzYNQUk9uKqpfYJ3YFF0W4V6/BSjzLFQVY8RZKY8l
6B2UWulOv8lKuPvJJ+cma3MIF0A1Wv9ajXmUf42Vz3snumnB/wTD+nGP2Ci8j5whyKndijsos0by
hjCiEmjWReML+kcIHT4mLw0DHd4vP0PRSD5eyGm6gKuvEGJwYrYbYyEQzDH46ewVgmRTLYOTl99i
mvibwRXzk5PUAXkgIvICNLPPWyUlBxNrZu11sVyLR5iJ8Vxh+D7e0QyYuh1r9Bpp8eqlaJUgHhlK
aQYnhHyAU0PSib6EC8tfyQMRWkPJt3DoDzUV9ikU0xM1MbL8rLwPpKKBytJRzOBk5Px7YNG8nPql
15+DQnYu71sjEc8kx6pvS5RI6lNbE00GXS4Kyf5/Zq3jo7buLxrfs15KJO0QopsXw1OLxy7CKHDj
hs8Wakbw6XYudLFA4WyLyLvb15X4fS9XgtZP5xf/j6rtOFHbhZOsZbzjyH48ZF8RmfxpeqpBeSE3
NMtUO+uoxRpVviTdUc/mSWJStuX7ntpTlp/JW+N8WIIvfHj/IudIO11LKB+21PXDUYH7gRfti6aR
m+mo3DlUMcTl+ph5dVPP5W1v6+QAumfsb63fXpVrQ7Mk8UEUb2HImMHvdBsu0i/JM4MubGtE30MU
8w0JRFwq0eQmC1DGpgJ+hH0WdHpeJS7zUGJ06GwtSA4d0H759uC2SkvE99W1M64DuViRy1EVFGez
kH/gUFJ3RyfQvyCBAW4/s8r1JPYuKoLzhgzRKi8udaJQwbNNPZYcta8z2GfqEz9kHCQohFpzcHIO
233GxRFJzQrLAl0ruNYVss5aoV8/rdWmX1oHpNN/fJJagmRDNChvS2OplQeToOD5Zr034rlrIkKR
QNk3RPOuTVDY3HUM+hUOWb6YqponPq7XoEMZz0cwLk8ym7Rrpyk+REwzr5Z4SQYhZxwzgdYn809S
wUrYHNsz6xEnfy0CU2C9beOPtfhwSBbqJGA8hyQwXabVbpRr8Hkp/SCDMsS3vahuwQNKvjaKfCV5
qQP3aW5SkPjasxP8lWVB/S1Sm65V+6XCmTjrYoM07YA0VsBnwF3HzQxWttJ1FS/fbR092Be0y2Wt
h/q5NeSH9BFqQvvUqpminpErtrqBYNU1bHjHsMrxg4zI9uWj8w4YTeUhNFaE4kxOzVohKsxY7hZz
dxaHY95qt1yXOeYbEZF7/ogmXbLfV09k6a1Kn/vFamlz/n/OWBmv9kKlGw2H8gZIVK4yo+MNH+XZ
S5l7ZP5ac+J1fmoCHVLVpYvrBcrZC1tWswU5aEQbnHl6LNjrrfZohuSvaLf0z5bCIxyP0QKxnNss
DqKHxLwE1oPGql0OqteqYogRfp5efyvOuRxmVcJPwo0R4vOpMq6yCeLTwo7FwLMZorNSXWeuAyKT
CMTAyykBAN6Vh+jWeJgOupDIicJ33fHmrQb6LpvXqIhxCqKhgwRozGH40OgvrvSgabOBzOO5a/eP
S0CXC0l07p4ruOYm8eY4Tepg3Jaojbs8T6Q352b64yIf0RudTPejVgtNYAIA6DohXU3PwYJk6Gxw
3CHSyqV7hlpK6TfHKyZywEnlLdFRWOZ+ZYt04JNKNk4f4ipt3goyWbmrW1cgynYHZpYpsWkaQRAi
/WT7j1fIw5q4w/QKVesbL6DL36mKFdPAWEZQeIQlvERF5Vy4erAeV26hxKZAIB+s8OcVnN1MHirA
+ETvEa8g+Cx5BYu+/6GOpYSwwJ6dtHg2CjA9v00pOVDWPrhWk9fBe3QWPTLFy+HJWEwWxmsctX0e
hOdncdA/GBnVV5sj+ThjQJdvFcjzMn3y7ujYj3ikFg6BMA2xWEJT/8LpZltrKEQufPezgbHcYlg1
8orWSfmChSHGDZdiMszDRB9t6UldW36+1g0UsXjVncbYYTNwjyvKyAfRLXDr9Lb2mE2j+H+9nN9v
KTwOXj3o2NRAAw93b6+63QAtnK1+JNizoIxmat1IoWDTyyQz2C9LUjCaGVIRbmQvvoQu+IP/FxSA
lp4hHWznCRZ7/stY+NAqQkZDyPcoHgN0r7a4LGdZow8qJsa7KMediYg9UxM3nZ6y+vDmPduF9hZu
vjC9LZ/PnmoSYtDdRIM9UjSq+H5tQ54FCLJmUIJoLfwyIpTNcJIHLvwFy2ljnOCjLdS8+5TbFqhm
wlj9qKQjDV2rNB7Jye0cndf6fy7l70KX1E9zqRX8P/JiDV98j+xlD7Ci1DnToQm2jBW8Bc1JHzOP
wi1PAorLe4a2YdqB3/40iUGBMKX+nzeaprZCpiQLnXoWByOrK1BqWC+e2fW4QItcdhK9JLa8VTZY
SuP2hrBc9d1j9K2BHZInuXHZFGdzAThVGP8nrvlGgTL46j0AKdKHe/dvTRCwO13P4Ep/mZUsHIy6
DPtCB3EXqlL76pV6VkE3/yJD5MSxDYfXoYg3YNeYO3A/HHhUmTa+JY5JXqZr09zCf/VjQJpYX3Bn
qxbmJYBJkbeZP/dty78lcxnTPJ0s05RJNBY5J3BD/UD12XchFH8GSc3m7JyVvKCKrMGjbw02Ms8r
k54eQrT8/OSRs1ymK23IPWcAE+6+KSKe6Ffc6YpcFjcsQuS6Oi8sN6ziLW+SlhUkhsHgN5kZ0NXQ
8HXKhvYtkiJuujejituSnLAOADOBAuEpItgxEivyfKJT/tXCarVXUfIGKSyCzEJNycXZ7KzJvSI/
OVSPtWbO7egZLM1j0Ty5ApUA4wjl+6H8caYGDcfAtFxC7gZcQcGlikxiEgdtIh14gj8oVXiJDikq
CT+APQWd98KjwqD63YkYms3eNtV3aX3264EP8R+9uELjo0B1Kz4PUOUcEXU+7MiXT6BvseHEi1Ea
HLSCRX3I8a8V9YGs9KpH4u1Tz6Mr1dvoHZk4lRRlx97QduQfuphoonWR/tvW/GAUdWjGgn2MW8p7
+pBIms9v8lyeXa2XeSXKWOUr76yn24h+f2R3UOlz+V3ZHoRyq1iNW+1ZhJY9/cRTQyLi7cOW/ln3
WAFysiMJKBTQ2XyOiv+9dOhJ6KmXqONH17S0jFKA6QJSOOapotCoirNByd4SKjs/aLjQcEayl2Oy
y/psRyv2DxgrYtXyRn17T+B6HiWqqctrt5D91JwBmxR8pz6Fhqaxdav1CNnmc8D1Ko++QYocAqHG
kUd2jl/Lxn5wmHWAzCAnc+E54qvkAK1DeVOoQTJniMNKT98fNeW4Mby1/jTct8MM73tkKTa6qngJ
7J81CcdxeBUfx4iZfk4ls9KvksMa6uXY9FN24IyQUjS0lgaNmlzZjploRYyJmYkZHnXLQsdI02h2
XiEuc0yRK+peR6mPrJmEqrlXOEh3RfmP6ChWgDnaLURP6fsAW2xY+ZpV45Peo30aKNVP1+wFXBio
yuyo/nBBIc2gIi1bYanS4HDZibXHmPxay0fG2k9UkRvvJlYKP0GTgJSA8rKqYLUpRFpPLSaleXQP
palH8t9nKIoKFdzYWfA6btcvw2nqHoBO4AUlQOa5e/zFh4BbW2NpndKlMSxpEyiHGYdueh0LroED
gbeYI/Zdmfj572WTGBvIlXhx1/se9XJO6dANUVRwV+j6/WHKlDsx8Q84uMTgYTjDkDCaHC53EclV
i3fK1okiXKVow2sxa3gCivqndniY5aESYjiL++vc5IRv1gwGWOOKpzZWmWzIpJ7z5A33AsXSjlMg
uLcobK+G8quV55DY+dRJPYQE17N2ICe2j/zR3eZ2U3HnB4vCpW7IO/KgFnNkWpEDDKsW2k4me4lK
k79LPxCXmme8RO2XdvWluvwaCVJyZIAu05WTZJf3Xw1PC64EAJCAMTlbXiDYgwAL9npiCyMCGFKp
JT9S7U8dvf19NEKkP+jHfkHoRSRB34tzvybuP2bb74XMsPiPSgLBAG3fiQqY7a5wD06Jc9nlwbKI
NFetW2eDcJGhBYKmVYwM9Fs5n2M9c2fuJzsLtJgif7qh0wDYl6Q0/bic5EouexoifYVlThOfNBtR
f2Bg8qQQi22k0q526H/L2H603Z3Yu74dNnyNxK8dPtupwlwsQ6lRxS0bUqw2JKqnwlakjae/HxWm
/7ORBz762NaJnZpIFqKp7U733b+ntfJsphUBo/9LfS7Zdm/dm8iWkHmRQWp9Y1cZDjJtTyq5U6gw
qzPIAi705A2+4tLbza/MpYH+pQttiRNpcwk4Dx+shxsdogUBfDL898qOK9/mfwvgrTOmYP+4PW9A
h+vKCXGa1d379TQOytFR7/FeQpn5qH8O5JcQoeshZpCeQDVX91w6p6TY1geovUJRdqFXqSHwMJ5R
iGrXjVt/njgiI0qRJ3kwprkPHbNG/O62AcdEZ9Jis31lQurRwubksNskNwClWXJy8LcWAo1Z/tp+
m9HF18ysPIIGp/Ikve0TjeuIWVa8BusKVGmMDo1b4sV+g4RCHbPTabM47Rzd/VnoSZ1cjI6/KXlo
8M0yPK8WTqdr0gBKmRG+qSmT0bCekzMeaanF5rhu8G2K1mc3s37ghxZJTHfouJgXBtkuLnsNGH8t
UlCHruNzpeadZ4nX11y6KRxAA7P0imzbNiaugPdu1InSrgrR84kE4iSWB4nMdHgV0WuEs/Fknvwy
Up5xIiKOqXqfKhRHO7rH1GqlhLtxIPp21jv87bPaZBEGEPZEh/Pi3KnfJwsyYpmceBY1EMW/1bY2
mxPiN3aDDH5hhYTOE1VOLk2stBkCnEiHZaANZXnuWzOYB28hRvvo3nvI8eFhK+t6gl76T/aGKuC+
TgMUcKv0E+Uhk9/fCcaAdwSK77BRdRbqNJI6KuM85BkVEd70RFFtlmPK7OqJx3EEEtHHM5T/fWVt
wEwL591RaCP328Hc2Xfl5DazvMqYQ6ZRVVHpkceYoIb29kN/RKXdUQO1E+hnAglmkB99dr4xCTit
2+HHgqOCOTuRxqyLl5tRh8WN9Es6gS4/QUIl9YRVfDlS/pnrt5Zvw7ZIM7+P3ydcQg4F+ZRafuwH
IKT0T137lkGFgwxyqgR1m5nt7JmFRjJDDP5NorKp0FKBbhEirnYhH/ICryRVzNfDYuszqbmu8ZkF
1nU9ry+YNNqOEZovjrLE4rRiERWXr/sKd+jAjGmcyp5RWSHwQOIuKQWbWmbrGKfxY7nIcITgxEXU
Tjnh7pRg5sMc/8VdlcT0OLyrXpk6rAV7IibgfDedRkx8edpLb5H5Gzj37VgxcRK+5GH7UqGB3ifl
CkFiTpdrAWsyd1/SgkHKj9mgv9lGe3HsbwmZdmIkl8jp8LX9kua2DiPw2pvsT/LdJDBj0KsU1r62
m2O0OB6Fi+aXhZ8ch/yqpAdNQe9yQ69tk2qeNIng0POg43/qHhugkT1oNi4e1i3V1btyDjjPHuF2
ossCPkn1kLLD4r/DaHOgKxUxJFUTBZtlUrSClhKc5Zo7lQWukaJcimNuJbVV4wxMq2cRp97iNfsM
Q1jWcfHiKj1B6sWdUZ89blYuuK48GjkKrM+o4TRBefcPxgu7b27Aurf5NYx4UE+BDIhswIa6z6l1
+at5RyG/mC2QdD9r7ZVW1fesSMsWhtLLAqqdm98t0vWSdeH1eotvdD9ZgeoBUWR/PZbyFL+dsMiK
/0w8bPdOYSnyqDSKD6zKm/+2pDz3i3s/tOdsMk3Sjfc7DUnbivBhuzgp+Mbj2DMtRRdVW/f4tJuF
FPQsbwAOrdobdTcTFbHTzsS2rJuyEklSYAbnJcdvHzXmu6UP6dHFgc5i1jMQWylTspiXlDyc3R8D
c3w8VqN8YhFGyetZH8dkvXRIcFlyZpqLNBqe4k57mCZdWy4R5V1RGfZhsGOhmTHhKnk+i376L/ki
prETNw4N+7xfSs4tGrScLZOsNTTIVR1iICK22jeve8q8Nl7KTbf6ZcIXo6WnR0vZJGqPhFsMbJk1
ewTD4n/moA+zz6wdmCiVAtBygpwo1Il8IIHWZw0QcmF341xS8WiHJgZSIL5BJewOQwlP9FU4jULL
OeE9yMh4ir3+7v6pvWQYRRepQeC36qN9eI59uqkzoWqOI0tdXul90UCVlr1S5QGS77UwefLwhZwY
//uPWu7UYflofoXeWwgcL6UaMwB/gLcQL8WezRsTmv9sWu3DtT8I4Xyfr3ISsCEvp4251MoS5zY9
BliQ6Jh1/Lh9uZW502LGpE6WzrkHx1vVKQUxG3AyBHFS3r8Vty8IEbRwM3hSuY+8Mmf5BhsBbymC
Mi6ZQcThZo8+1zQ4bwNgQb7iYwZRMiYFa44TvAf84jtsGB/N8WldFaid2gchLzmlwnwg758/cDDK
+lNSqKa5VGS8IG0ucGBWpTHkHK5LagjLMFPQYvNQJpuCSuAtmd1fEqb9q3A6wLxaORduOvzaPPM1
3RfqQKYdDHCUfFpXGUmL8asX7s5ISrmvsWdnAce5ic3fl/miTXpCcBrJnx3PPiOaH408g2kPWjrq
XOG+3nRfjWz3jtx3nhRxDeCu5D+LXJeW8OsR6wYZUtkMp46xgY3laHxSQrfG81+76YVknPBpSPij
i28GUkQ3boL39e+sIcIWDz/bUNzQZWYhwoKaIYgksATSY4+daoqhzzANj1E0BFQAfINjF+RhPHfm
fQlQ93o4oK9Yyimg0+5eCtRmRZ6fwmk+lDskKciuEYw6pQejwadZfdg4jGYPz2yymLXc5RV1d7P2
fQ+xcBA2nY//1PDjOo956iUqYp9oKiWUoLerlLd4PdzV/BpgkeSpJcRDnSvnR56GC/WIC2evnsu5
+mpOFRj6+fGUwNLgO1YLsl5O12YPd6p/GDRT+rT9NWsa3ouc37JDrWi1sSJpxbkbcvOuSjwoaITz
Kx1DJBJgFO4FdkJICj8b5S4jokhvsb8ypFCrAdeytcMbLAGO5KbN489x1IXxkWPZ0mMlFxEBn1Di
6V5SrNwOlbEytp5mUnpra0MpviwlOKkBh/zb0PBNGVIPLIDbdLpQx5CEAnWLQOz/WQIrf93JtWLX
Tq0eeJco15g89520tBXe9GPI39JvoamSlQM3mfcxJaTKDAowUhSgPyQ3PWEUYeRRPra4ZccRgOf7
AKhI9xxNKsBuqPxlTIDfQzPgSMPvMORp41rXJDiCIwVx7NrKCSg2z/QNUqsTRp9jkASHs95ghVW+
/OgXBftMDjXKAxiwFt8MW4eqmvtL3EAa2pT38qQrkNq+ukUd857cP553Z+/+4TjyCe8X/DuImnhH
1lthBwqUgPg5bkpCV6H9oSQZIvT0fDUQ+kzALjEfgLppNG7I0ABBLBIXaW4oWZuutmcf/HmdFg5U
0T+CqRKmpGSubGTieOFZIsjqqaCpQqLjqyltiZZOEN5OHLw0BcWKqfvGb+5S6Px4oS7VEnm3t27Z
4Wafa1xyzZQ61lUK9MKhhrhrGdBQ0osyI13KuYbxSabig5XzH3Ki09sv5t9tUyMWRZhcc84ye+ve
WucTFs/cjDdS+u/+LAZH0EDfiBDVgUQVyg5WdPnRR4q+lH+ODVlP1K/G7vga8hfymcfdP6OTiKl3
J1+XP13Cjzv9xHlpuYTTbt07U3+jfLvn0qGUcGVbp3zEKJ25PjxnXssO1yLfTKf0pS+GnOhbI69F
hPdNpu57wWBOjBQH0iENDnemqvY9wGzxqB74d3kMNkidUa21fZMH75eXPoScu3nxoIsCYeIC65HU
A0dUVME2eJCfU0DcN8yUhxSyZv1iWJcMC7MzAiRcX6DGk38MbftwHTttFvuLmk0k59CpxE0MPFAA
FdFvB63IOdE9g+WW4R8k6hLshmaxIzWpURJby2DLpDUv195VkKlVw7kY/TI3r/hpxqS04cG9j99u
WoTQsWLDKF0xPgyZCptu0BYjMPnaHEjXuS7auoexot+BvaRg4QhZTe0IlPARPGZJF7sx5FHIzFpJ
JOKRj/nx37v5DS9vQY7n9BXgPG5jLU4KMp1j/mLcv38kjf24s34YPhvSc6gDkfjviysW+p5h4DHH
Oxc8AO9H5HFJPB5E4ZNo/zPRkR4KD/sw3SMzrHuLcp+ewzcj42Uij3/3SsNj8pvRCtjlbIuJmCVm
t3rFeaCMcVQpKNWb5VIjVPTupaemSjyQfTnb+BtvJD4ELN3umx1SHuBBQkdLPMOJknFsMkVEH40s
sZtia/rHGyn3Z6yhd1RtX+A0PaQYpvRXsffuNFlbgQB30jzwXUYPbSapMhJ+iLqSdur6RoG+T+Hk
XhbsIatnPOQ3vLxb6O1e0NZxwUcSjdKj/py34wWrkRK111H2Ra63nJ6U87SqULAr8wiNKL9Q8hQd
8WPxo8AuWoImGxYeJPJZd/6TQekZ0MwxYf09t0s+vQ0bl1P5GNA7gyCth74Xkv97CQXicf6iZCu2
Piv3/6gAuAfvbXfMvlNmMeUvvMXeo2UVUIO12mOEPPACKvY5IBsan4fugs3AmievTdTHpHwnnoIl
ADL8ku6JSCvJE7/sT5TDGt70iLmiGrdrR+SbwxqIvwUv9JdSNccHIASrSAeGcy2cJHlkmbEaCzsi
s1p7Qx8cPEGXUB840Ui7UgFSZ2459vL/8VnVX/yTi0S2caXLik/opMjB4rBkxT9nQf6EcNXJp0pX
pnuWGsUwT7M9sZRWHnHOhjU6EY0983MqXfVByxZJJBM44Uk8hQ/JOwXPps73Ew5PzfWAyzPkae2E
zhzSPsrnMCC4MWgq1Dh+GxASlpc45Cg8d2lcfXN0hUmbUOHkhcWqLZx9sEKAgO11q+ko++w41SoR
6PgqOyI1Cp+FYQUkZU82TExToWILqoaU9EGDIsjB1jK8ro26Q7rvZbx0ZCrBF+jL5QeiTkuNCe9t
hJogL2vCtmlyw+Fs7+ebsTqJ7P2T3Krc2SeJOQtqdu+XMaTStGREndX352t/AFZVRTstuPSd3yl7
PAQn4jZuFt7p4DVJLxlXo6qll/RCti/a9v6mjN6IvY6wAomcg4xhkMuTOdYOBAkxMKOnqvWGwwWN
pm9TQ/QPDrLPdjaDn44srE8LDouwyCZcucUoHylUmcMLw6yEL6ppn7GutD+aQvTiHVrDTTN177MI
wTaSXV67TBpSb51wM70saO4v8/mu8Vz/fNNN3zJ/fxYayAFBN2QN3O3rQksGeG/XdopWM9/vGVrH
jKZWgz5PfviAY2XU9rHVwZD4LkPWsDbV54P6C5U9R/q/8Ry7ADiJ/Lw3i9F0FYFdWZblEybTRvHS
ZUij7Szp8/c3ZqIZTLPm/G223kfKNUA6msqEaS3dbY4xISkuktaskb1Up4POVOBe1FMHYU2N7+3z
7cyFZeYBGEs91vT707lnuJngD8WLjb63lUsiL/1zlHQOGa+aHpprgm7rNcoI4kIEI3YGikiseNNs
ZjX9GV63lwpwXm9m5XSpUy7W/dphSSXlVAH+pBz+ttxbLE/y/Jf4bMDt64VofyLM45xe9lG7TBx6
kftpXSGsaItMUwy3/gOAHUb75mgtPCnPoj9ABZ5T5LFM/M4FgO9rKyCa0ZjXTX9C+sNWosc0uQEI
3SXYyg5VydvtQzwbuUxgSiZ/lj5+dg255geF4wq9PrHUZUS7zG0ibr09KPVzC4y80Q90wI2d5fl8
ZItpeueL4uVRtdYO+LY2A1n79GD4sCo0HPIqC3rjJX+7Rf28lI+Tzn1/rEo7h3Xu6h5uOm1AN10v
1WU7SpgXorUpmmo0go2fa7K+AOAszqS2LkPH8QyT2OEikKGrjENA2mHUM5A9FrILd+IrMnFYHzmC
Sdfk0W6gkIztq4f6YuzBEx02DX6OiHgU0T3yCaGrWclq/NQy5vs+n4F2Jkmc7F5z4eA0rOM8oSTo
PuIq5M8OfxTx1Iyqd/apbM8hNtX+Z+zcvCjL4HwBSHDR4RH6ISk1Qy+Pcf+BRTvYG2PWmbLcMvtL
x16Woy8juKAQJWA1nsxlXdsqW1Qn6fFOIh/ZEWF6qEInZOLiHaXPsOfu3TssGHZYUM6sKlHUOsaD
0uuALVCgl/A+23x6tSIyNI7fqViuCCOyq1WzvwSiZuqR6Wc8iq80tjt6wGqzGCZIpRda4BUGLzwC
MghdvSvrNnpOrFhGBi6Xg83kTvBlQtoc+cBk80ESApMDAYQS65OGx+jicQ2mxnyBl3u/KUZjS4Bi
uTX0J7btC+xTy6Diz5LhRICgrFytbQPzubuZZhVuA6afWMaYGCzuGwKG4++J2npB85/NUIpLvzxu
iYdW33rsUfw3FgmK/O+ROyesn7zl6IkzHdAjZBFktmdhPx3PSFJviRx/uyTwowGbDX9sgNOGuxXh
NGo9hrsstErh1LHc3KzN5NuOdr0r4OYtb1Ad2ZUZ8DGUIwQad6QfYhWKVHYac+YWFjl/+Ji8LEFi
4bIo9QtGvu3eSLyif/ALckjf1yW6HMovqfCeW0PTJu9FuExMk3WqwAaHIgmvLfpBZtwdMtx91GO+
kbyL38f3FAwARD0TzjzscODFlSwOUF8vdMCI+b9Fp58CiKFwBfdS1TvaZ3sx0+7HNE7UybGXRrqY
l1ZtMek8DTg2G7sNtAStZO3Cd/IUZ6qSZzpMi1VVVLWycL9rP8d6nUueiDviLXGWk9s0VTZduwnW
PjaYRtDrgFGRSRqd5BrYDilIPsMmFgmKdr6wtU4jH5GnfJ7BVbVWW4N4HAd4pa/v+s5HcBNXFDrT
HPye0K2bQNF6Q1m9m/RXex7/U0Aq3k/OuoKCmou4zPxrhN6lxYk1ZvQOJi7JeHhF1PFFE1ZbmUFQ
RAxJGsRFUYXmzBMwdd2RF0KBJf+5UWJZqLCMbfuBwQFrDxnCHEu1BdDzFNOed85HvWHLwIyD6VYY
/HqdGI4QVnguYey1ABsh3YwFHjk4V4ku0xL7mcE5wR74KsKkKUFGPP34ELICIKeUUPlbbAjbw/0n
QPAIzW5wPxvZXbWKTylwC6jsUNviO91IvQVVYe0YXSVXNm6lxNPUCKvrwOXLBYPGpoQxDvJDRq/e
DEvpS9cWyYfBNpCtUOjOjAoMW4avq9VlBZcX3OI1rxAca0NolitTkR+2LU/3ZW9GeV3cu8rf2Cl8
GHmTjlbgy4gAlZ9ARoa/vrqMRQc1GZCJLXz+ugkYO7oJyFrFannN3GjFmUafRAM2+f/7qaL2KFa/
whk+GtAktsjE1OfLMdaJS0B5OAqWnmM93v3U9Ga3SKTKGmnY/kbua2WEmfYg3bsof011F9l/00XV
iHhjjRyJJ/cCZzt6ZVxZ7pg5AkCdcfHepL7lfpF6KpMCYwl+B7jyjsQUujcPY8pqWJhRIkMNcWJo
Izlby1BC5R/aYXUjuLX8neIZJ7Q1hHLH8m9gVF15MYKtPssAYBvVI43UIfyUZVCvRlDeWQGgC/Dt
OkPwKT48wIBbSjAJcW5EflCTjswPJ5AEfxAhj62XqEymrYWqjsNbv/moWOhElrkLUGUzYAEjuJST
Vvh0OiJrnlCs7Scac349xxY0ABpaC3ei2LKdtJ00L5+JGUmLYe7jVlUXGC2t8hBf1OskiTajduZN
jppsV+L/qYWzUZ0qPCtHZsz8ajd7H7RmlNxr6ghtRFIz4WXghNKZyVykVasPsLclPhaJhnR8JbVv
BHqtO/D2kEtoXYzPRtOGKXo8qh2kO40CZ7dunSs1dxAYtxssaJidFk30csCPx3PzTQObKwOFwofa
ltXGbPUQN/WDZZOkNnbsI4xKfD0ayUKU0qdUpnGFjWZTchOUzkbusq2LXkHoQP41Bx+FYbQiDuav
s08o34U0siRbY79nGKAsUY7OjaaHtyDJeRRy0uYHk9gwy+HBtuuPOD/+4t27JVEzMt+qFXJOaFSi
2y26bbCTnBMia0ZOcGflZkrCpi6PfoOaQFh4S9rKZTfkYYsTSM152XnUZwu7AjRf03TWHOILjdE7
Y2XZwZx2YHLYztR4rh7ykL+R/SBSt1K3KF9zH83tWzjeTU8a4o9FJOg1oW/Zz1HBgssLy5q+ui6K
ErboE0ACJ95GfnEKQEu519skOOLSjsSDwW9LR4XxygR2Om0ZNPv/YNd8/5zSSuH1ML2SKeKYv8nU
W3Z7fBmbRUuZmiq5mLwrBbaVcvFasMAYON9gSeFqL0xBLqA1nqqUzCF9SsY5tci9+IUYV2HKJs75
kKJ1JYteDElJHIpK2TPIYZtEVK/sxPdojSrYy99boDncpzb+vHMpM11C83xX5vlCljlyrLqI1duH
k9eg7VV0iYVDy2CDw63UGxG3R1VxETExG2WxnqcMkCiI37N76VdfpSPjzBUO/ZHaKpu5apOVLcJe
uWCQP9e9bkfTYjhUy3RDXycNJw//9oAsOZ68K0aUIFNNtEsp3UeplnibCVrFfbFdeqFY0+x8YeUw
pAG7YynqaLbbulaRGvZZXFnUYIQu6pAebJEzxfh0oQjuY973xyAvIXWH3LZjwMzExz77olqtSPwc
8kl81HUTXrVMq7XPhW8qgbsYTUUtEuhLDtU58RRueXBt8ejNs+d1i2DAJEr89Y6BOCAPWBvx3XHk
Ar1F9rjlzVCQOcxSnMnMUC4gUTZjn31kcRxM92Tx0gEjD+OqHgO0X7lDlBpYRiq+lZ1d4Zmlf8zI
FAyAph1/PXAU+jv1Xk8L2TN0fdxgp+p/d4swVp8B0Ue3H2nbWOyNFUKuE+5HMv0qMvLjsms8B0ja
mdpmGxFN2Ik0wWn2eIcMPwKbcDp07q3AqLww/P0fJ3/Ap254plr3vw9J/U5nK8Pd9drxPS6DTat1
HS+Dr5fK2/Cnh+psRmw5/72wAaqXYRs91kvBY7RJJFt780zazoEoU4wERlmAZn0WrFsQ6AHVqQp4
KDUIAy/WA7KVPvbJsj/KjXmDiGy9eKVtOxgTxzrMOLp3o/hSViiCG2vVLi0srE4t7AlNo2/TugWd
MQK7dpxVH9jNzUlhNhuqyIiDP9e7on33sOH1tVJC/Ndv2T1Q9fp8w8MxfDkjkS9RjcWCf8QKw/IB
wUF1BT3WWivEWlIxvWhiPLJBKbcxkpnx133y0fHcClnORhj58ZKscbiP3SUAwtG3ZvGHs+Kn/zTU
iiBkkNRzJbnRAUxJ15pDsuYZhOm6ECJ7roL/SBguR+tuovDQJ95j4BQ3Fh3u1h/+L4aL04F9JS87
CMvA39jb//n4+Le5S5MfpvI+/kh1hSjQ6obzeemEUxpCwd+iuab6L0OMFdKDJAIPneP09g8WpIut
nxclkTNeMNlMT8iNFvLiLvEnepbM4aJryt7CjsXcs9V8ATRKI90jsqcDRKuYZuFyS9g9Vc9+a+Ev
Cii1MDp2DBOdDCYBABc0BUUYcrn84+KDK2t1GZZooaK5m8S+HL4/P2WfA4esOc/t1ThEOrh9D/Bw
+bGDP/+jVxJsRP/btWkWK0WpYLo7PvRtKJSDFIPuzDT72v9JE5XFLTnPzrZLHna+/cMo1pgLTZyR
JoYJydZurk7TuU14qC/IkJlAjanUnscs80uGoxfraxkJgKbPqeeHTw97gM2GO9reZHYNHq6+j4ZJ
HV70N87yeX76fSbXHt5HPH20qKPMAAHpxOoHdm8EN1dRANAWKEbOh/Qmz+YDC5cGkTWF7OZnVtpL
HzOzaXBtiQHVd6Pwe21esK+ky5NZktmQJCJ+jAHt/CWmH/fStv0cqHk3Zovp3vX/Dd7AGpYCZCWL
iXw4xJ1XlnfVqf0THL1RdmO29JnOrshWByN11hz1eHnJWRoLkuUd+AIpmbAYCYYZBChXFk1aAEwi
hWiEaWLNNC8cpZjI1uu8AhG2bbtqDLTmc8oBSBl0Hy4GDLewdx4XaF5ChTIB3+i14GFqaiQN5RcH
qcNBcRaIyuS0juc73kwgOGQcypXmJICejKDVy+WZgHe7U2R3WXOB/EJjzAr66QQS0pgUtdkhgg94
dOdHmNZBvdE4lDkyNvg3vnX3d2rmtYzJKJEnwLhftEczyS8c7ynp8EqyTgmibVT9dZy3Y/9cvxjS
t5apJ2TzC4EXpRCMqQtgPehFu9Wj208xBxoM41uQgWZ8/snuBtgCea5IY331HL/fFJz77NKNUA1o
LGqB6HLOIUtJqgHRYvmhXY5DjaOJWOH859cw11UfDZgzaV9InSW2caDGEqe1w7EkYpiY7sbNC0OT
kOuWka+JrDoidFR8XToA5A49KUZ2EJzEyvCdN29Lnz52xWFHnFxJEm341oVtA2VTArzlOYmwAwhw
L/fmZU75E/Sceb6WmrXxkT635N1f1FtVJm3GScPUW4aT6z9p/EOG9R3hj435wWKLf433Gb+yy7/T
muDyVFQCL7ccLiNyTcwic9cDWfCPnph4hJrUYUSKZkjo94F3qWiZJGGkMEvRZvRu276aFDyODSqz
wUQmmIeL4pMW9wHCQgU9pEhMZkIJsE/rSvM78cW25HftQ/dSr80vwLGvqbtAzYzzVrJ1Ogk/XM0E
6TvB6b1jI2Es4ea1F+tRfQDYQG7sT40ftHAA/9b3/N7YwHID2BFRNowAZsquo0PMXSBYBhmabvPU
gZ8TWTuHn1vpZExxL8bspiDh3OR5VxyTUEYWf0Dn/AONaQyNDouKglZ2LdW4G5esBtIlQ/sWrPDq
xrWzJ5Emz3ZmpwIbJgWV9gNRVfVBb/OJ8RtO4WnFexwzvdeaV2N7xapwi4KUPbr1XZtcd8a7bd76
uLw1w+xg0/qTSuPE6NX6HaGgSh6YKy9bv4BmMYX/AL29L8/o3ewDeklnjeGMzwaqcnSj3Bvr/9cH
LWtaUmKcCU/UbVx1ZPGamXAcU8i8DFFbRTi1v2LQPHD/oyi9GbO5rClUkvMicPR8GIfmfY1f1WTf
vA2NBPfusHxp6PtZy15LmmlGAfSO4VwxJPNuQbIKnNqmDGHGHlFQ6+C88uXQZzO5s3wStn12b4eM
zZXLT2acyo6EZ7mf7AlOnjONDcj+iP//oLwa1h5k40AGeXHH6Zbdi9v/9pAh6cNqZblBFq/meoAw
JgHAhEkb/1BVobGbBQ8gnJqZ9U2D6jpDugy0znJvs5s2k6rzyy12rpG3CNpH0SdGHxBkFXHDfKO9
dlzlWZC6hGiXVQotRKfiQNodhKYwTsiiBQCG3wdzN/20PLAjRLQHx0ACRL6OZdxUkAbEO3Rvmzc6
oZJEgaYuAWqj95cOJ8uahR4zTULdldLZ3NdgmRKAUCYyXZbKFCIqi5DJfqAezjqEFLUKBgJwnX7W
PKr7ki4RbTKv8y+I3jWVz2CogAiJqZ+TO1sHIeQqE088+e2RIy+FKxTEO+oerjZSrWlsc1tnzlGf
tTfNgiOYalVuMx14QNPY1UEbqKEDRClfnPG0Q/aeQYQaVzoThPJCzLOaI4NdIC5ev2/9HlGszsV1
B378Kxad3H64sqX/p1PFha86pjE+SMhenfUnbcBpIgMkFZTd9IlY4HdF0Er/hZibShJZIvMosnhN
2wfYbcNXMTaZJDpzDJB1jUxWNVbbi35DAxjES0utltVDgffQxY30Ro1VRGmIS5MVdZ8g5HN2TkSP
uLEUSjYjhPHFxbSf3mSUYxKqYkK8AgXS5W8zMHMioELPnwktjZfC7PNRxX07+BP0kdlldgJ8uH/q
B7YOVcLreltt5+lBXBnS19YBDbKwR4qNTSSpZV7hV9W3ZaG1VhaI1UF1On1GWa9rT0wIRnzI6hTd
u8BrD3J7klinZVqMw87f0mcek7ifd/2CmOCzQYsiPPk3ZQbb4gA0BoS+adO+3n2SQ1fjPyJQTRJ7
AAXq6/RhN8x46yy4hfnk3nalOTGTg3wGBf8ZzFnGna4Vp84mcszBkWmZa5Rt89LGsqofZY0nhJce
ZPtnpmxkrio1ogoqCDg81eUzCdI3ntlXjuiySf91ZC99R5n+7DN1lGsAlf3KUQ8QqDQaC3ksl3Oh
IyFa3+3V7kOjwrgozM5VXVGjvZgZf2fM+LZU2k6s6Rh3d/yqXLdnBdDEIouYME3qBWQGffxfn9fO
0wjxqs03I/+bcy2JoBB3wbJxsLbIqAUYg4nRWwcLMDQCpAIC6l1gECVoQh3DH92kwcFBczU3Y8l+
TOupXTeci+Nh4zUvlzazZlq69SqiwUmaxkq8F7jSISBZ0HXf0iVIDSHvwYJjLhZYS5DpKJNFNhic
Vaa7gdNs/qGpyqD0E93Z0k5sKTY7zw20kNkW6WgqearOkqcKJEbbMb7itA7RyXBR5aoS8kMr8/Nq
MeeNhSxeUS8Z3rAxzzPKaLCQPWxIE3SHnvKWIbkwngvNzKwrHNg5kL3mZaf/GKTKs4sx8uhZZ5ys
e8w0XgPMUoEGWifoSk670etjWv0WytIus8FPvEdsknrVUcWRxmKgvyfNukVyrj61FaIEVXqVJV25
G1RybrvHrUHXmZZ9y7CqQQrAsyWRzO5nwMUV9wHFxtjAPTMer//ae7gg0y6WJ2D6JJTTxRXcNbyo
OqNaw00jW3u4vwKytkFBTxIn51khL+Nx8kO7dORYjVgTJRjUg18VIQqsefh2IwQfqSf4KAeTVWm/
3CWVS3beh6QIG19Xm1YUmF70x1WYhIdngPGn/62C9zA5RRXF2owoYwzr/eqe/sCYGFLNtR3nDx2w
2+aLkYI1PhHdHG0+Xzf4iBmzr3qLpCsw9IPlwMJ2fl2LocbnfAIkjl3aVzYbI/h+OIae5lTtNSeW
5KyBp6Bs8PZfiPK+nyKqHMkoZrSDGPA4euFnROvncWSuqNK7abz2P8wNtNEJoQGCw2SRzZ5HAwxK
GUO+WvZGA7iD3t5theJxHv1WU4n0scj6afEhmGyL/SQvI6C1e8a5TmGX1f5zoJ93ODSHOSGNBgn2
caUQ9VR263+BQ5aW+GT3BuPstleVpJ4gvo6QwVxh1Ycbr7F7kDgJbnA93V/DSUz/nFwLhqngiSnY
xAYTMYmv/4dqImoxPYQcvziXKFyxjVVod5m4ed54QtQQUhvYHH8dg3Yt4GnctTyu2jF3M1Uqe5Ff
OzgSjwcK1OCy1HnGtdUfA1EqdtIWyP9ycNxhiTOBcIpQt/kyzmS7BIPYDVlwPvDD3WKx/SE0pM01
KbKN3LW/vj33Ldr51RrzAfuhfkJDwCw+njsIvy5KqaidoXtawKFdB/IS1QDReb1uUooYYtanoe3U
J/uCTjNxoPu/gyNkzKsP/Od8MAsNI3CoWZGzotJ7JcKdgu/al3zm86GXz3+pERKSM8pKgHeXdTOC
7mY0nQHza0HzzDpbtP03qZRydMX/wocuD8g2/99V4dP09rmHAQxZfYhXif/HHYqO9L1l85OJ3yF+
JyXvENA6Cf6q1JJyBTgIsmZg6bFi+WaviUsLtJtQ/eWf8MZbdBnK3XuUEmM2H+eqFgoEUj0W35sH
9nttPi17K0mvukKopir+LB12/LGzDilWOB7ITfYfDcPXRrt+srV9IBnGJZDFNLltelGCcuqWRjYU
kmtvnekqfsf82FB/rpsOl4LcZEeOR4KveSNpgymcADVHcjknflZBVqJDRIYte8Z2jScxI7SJne4Q
jfjaHuDDDNnhcmTV0S3mrnVeFwxc3wt2l+TBF9/fQYhXw9gIarp5rITsQzGq1O92Mcg2qgRb0AUy
r/7AlZO75rq4DCMegcrTe5ZesEyLWjsFDWMQEvsqlOHp21PF6lokYfJwbmOChiGanF3tv2ESDjSw
UYwBcV7QszyMFMmJoE0eBkeexnU7fO786MDNMQ6VhIefb2hHC8fzghKK1yuYg4ciguIy7DORAcDR
qN1uqpJDFCHU9hNYVd94ibA1qyRNOMbVThZ7AOhmh9M4COAFb4b8qBFQN1bBfKfMuRCwff0j1VDa
R0NCF9B7IqtlqtEVOTyi950X9wW1GwWun9fVzHKbI2YN8cLIK/nvPyHGJF+w9cC0+m/KO5dJdUoN
URE17jwgaLomyoCpgaSHQanIg3R/zkfRpMuv4lYAI0cJN6j7/HaWdeRQDXYiI8A/Pz/a50D+ybtL
3Czg3rZwR1hq2tKvUjtJ2SZGEe+Hz6JIOjwFoP5sgXqXWw8+lR5oBOWq+kzlzDPAcExyI0FUbsjw
1ILUH+gptskbYd7odpOEwFxyAUt+uEJKxuRsAbu3y0t2+Poymtg8o3yvlxl2s6OiUThifxCJl7he
xjWoksMFKKxZ2s0PsjnA/PwtCwtgmaBIDKG4/pOGrDpuOY/DU44KH76KgTNHCQmr4YRjZttAcfeY
E0dlV+pk/Sdsp+/Jfhiuvl/Mkf0WjXdYNsSuR/ay0pq6loNDp0GEb+Ya/+osbcZAdM8hiRe4ABEg
6vc0l07JKA4SKSIY3lh0XXcDmtn6QVvAN7r1HKuEbPQ2daJ1vn4dbNOqXyL6860t7AnhDNVgW90n
+QaSX6IWaRkItRP+z8FG5ffM75hzb2x3u9wN0Dpvr9iPZxW+N5lVBFrzAqwVyzjR3+5FgA0WA7R9
Ouy2IsntKSOBfAd5fqi5vbUgPe0XzgiMEaBEHbBrYtHvh5CLz7wxVPHXab0DWT24NHOj/iMkcJrG
ARb1jzVSba9gZ1i4ayDw66dcc5owFUCB16uHaMh4hh5JRQHZY9Yl1+FVZ2OCEZvi1+dSI0kUedRG
jZ2poyymvxG81OP4i8WOSilQ8IF88SUSalbx9nVwNToLIxP+t/7yD/xxcC8FZl7kdxGVgrqFHYQZ
PBthG+SMsA8nd3hGISo3ay2m574/qRMVflK28eI1DAJ/d/x1UqQO/jip82237uhpZ492rhs6Xmo7
3UmgeqPtaUDjf+ipO45e0YhNxstFXIz8/BNhwV/6OmnVOjTx1UmDcbAFlq0DYJ8JxmU7hAIl4Fck
/Vveu4l8wexOluB0k1aUULDEmhCipj4QZM1bvbnUNQu6yvvQEiO8XZ4qLRUiO1DGEL63X1zOmgKn
el7Gxb2ei2zFdjMYuRkTxNZ5TV8COgOCUQuHcap2QV/qyXK1yn5lQzjl7lp89lsePYBpS3+uIk6X
5XimjTdvTQAwzm8hINyx7Ng6rjBlO78DaYA25vdVX66+GDCLr0nB5HtTgaeEHvtv35gZVdZgi8Po
MPY8IjxqgFdaL7eANzWIhx6XObZMY4wRWTSmpGHBI/UXejkLcQy1NVv55/JfNLLEvZiErlOpbhYB
iq5bdL8F+w4K5z325qdhignVXm2Dgj7yDrhe4Z63O9dn5V/wue6+KOwsL6s634dSezX/7BCvd3EG
UgvmRSCIkq9xCb9RS4gf4t/pfdEJOs5AXYarD24zQywqmdb76Xa2fjwIFfcCTmSacw5mf8BSdcFZ
z1edoTvkTpK+NuRA7UeA++/XjBXrpoHo2PY92NS8M4RldXg5Muv3dSaDPhlrDJbVSLy3/7XJORve
upDxC+7oe/8MnTzofm3owNOt0Dk6PltILaYSL12hQiuTc3GWbvIk7HCIolRd6aAV/mn0rlECTL0t
XZPimkq2UzBimZzhHUjgmMtR9c4pGN5W+38AoP4fyzTwr6aI09OB+CvjEQfcheH0xr2c0LAnBN4S
f7iv2cSxPbnvcy0JAGcPcKCRdtPNCStwSmg+V4gV/kLiKZUBE0spKjqYYvB8z36VzGWYGOKT5RZv
15OaSelLWsd2X9hRdwjsimzJmn4Kt/za7MZlUNhKvjP9bQZwBVKRF9x8LXbjz7243WCWQz7DxQ1j
Hri2zuEKsoI64J4jRZCyX8U/Pc8rZdDIUE+0jAbqd25+POw/XvzvDFpIYVtX4NjJtKqsCauORBkX
gNmKSBLlKbAwxZp4kbyJcZXXvwU2enFuMajOVxXJz8Uj7f84rzbT7ttQ9gHub28lHwZoLJtf/5CF
qFr4vk+yv5r3IS7BkkxZWnzahHxB9tKHggtSmu3QJkbh2ACukjJGk1O30W+tGTXvBK3Yd+CHnney
9UDaozZrhr1dSLbfzRho/v475XjJfle4qxx76nICgg1LZofOsizNHC1HNAQBV5OwpJD0YdeVlI4o
qTWUY8Z5JDMPHXkZ7C3WpMx15OJ4OUU88Jm37CpcBuZLQ0ZgJ8Xpf2rBqeeRLcP3/5Ix3zdH4Lbk
ZUmHBNTbDgE3+eJma7Dl15BBOiJNJojkLubtj64dDVbP5JhnoIRAzcCMPg5VotopMapS/CmDSLjz
KQbR88fY4BIk5cqhBWHMw7Fuew86bdB0QA0x2CE3arJjgfenbSZHwFvuym56a4oXmXCJtQtxfosV
5+YEwyjZMLNYaLNGMLGxGQ/zGaFR4MYJxeVBZfMFjVPlLoCCZehDYozmpk3NgFDYgpw4uRF+Wb0e
nebiUS4W9k2TP6WCiScPxFTr29Mi0wyr4kpo7G6cG8R3QOa73r0ICtymEt+F2wCnzUmo5oPht3eD
bvZ9FbjG92Gnf4965R4Lmw6EIppjxqwOdkdgfQkzdjqiMeYJ9zeygobCyNHFhUCto3M3FUUl3Clq
ftBb6Y3n5tXhX+sEjC03SpGZOAAdd/sVKbA4nzXJe+yt3uL55QuLMKZfiEEHGnuELWaNb8Iz4A+n
Jip5yUnFaZxI9OpJhAV5wlA2XOGU9Fm5L5ySC8cLG6N4tkPjBwt86p/iF5VZRuMRYhlQgQTtMRNp
t4C1Hy867TkphXCaxnYOj/EsNHLEi1eFSqyH4jh/bA1wR0IdSUrPIqflc3Dza/KLOqi6i3s7m7WJ
v2PgV10RxgcTw8EhZImQc6YkaDoSpP2rsIKE1Ov0SulJQzZZRKsFKt34mukjlrBtUWuqG2hr72Nr
9FBkki8TSlcGMKtQdpa+6fzxWRvA/8DpNyVOnaPaYVebtQifZx6F9bZagXalObLJ3k8a6GwW1hjK
BoboFaJyH1gQlIbRKnwdN7ZosWtrKrXmszmIYl/UvZGUV5b2/e9tTNhCdFHoGHWUHtq9+zYQsZal
PDn8fpVfFBmH+OfZAZHiYI3eCp77njbhjeOkXe6xDG4/h3onmkKPiSdzRshylkg0zaGZMERNGlCj
aQ8EAULBvqQ3qy49rtPgUvO6oGeVer0sv7qSCelsS1e1kVGz1ff0bK3TofroT+umBMsA+5E6VOd5
Kioeo37MUtQcsZsY40jwlQOAZ+YkF6Vnn+MxPsh8wToDqQlCNWb1CrOVhTog1A8UvWRwFaieaYKo
gQhat/O7nnggrzfCDsN0Ohd+vOEfo3Dy6fzOdOzd9Dh1zdJxPy7klcXFXQmQghpvdr+/51bFjQEf
68/eCtB5nbaFjWElOrueCqrKRRx3bMGTiDQC8zKxMQPNcItJ1ZWSIYGDgon80a6cSJKiAaGxPySw
nKgGQdSh3porTgF3FJtrVW0BN9WK/s9NdLRQikG953uwKyoe94AP75CuzjIn/f3eRcTt5xkZbI44
gcILwHWW2AUGCxkA8KdSKqfeah7Cc/32uMqbKc2fSTZ+nO7wJNBkEUYR3yxutoCiE5AjDj8EQ5ja
TD64sZNWLdAWxHpk1hqQkoOQvoDanRttXh4/I7eh68ZDBB2Ej2F8WY8HwDq3yUMSmWa6jjtLMFwR
BVM/KbQCiYPH3jd6c/cCAnnLOJ6/bEGVRX+SvbKD2YtREmqB2IorxXdMfO8alMOMYo/HEsZoQHNV
/I5gsLyfuB+JF0v8eGvtO3B56ZvnOjmsb1guKeYOSzhOzbhOhkUw9489UHzGXTjVyc5+nlD/N3yi
9i45FR4Li8gxysawy4EN+9myGQm4C0+bbv3xwrA/zZi3cjPADNJ9H3inp2LlZjn1rXru2zH1YFbg
iaoa5Tqf53ISJbvE06mBy5U/pJh8HdUXsTVu7zvIpfVGwo31H8CUrQqrNkFGYj17mMEoT+Mz9yPH
W13Zhaa65PnFkhTOg+2FKkmpMh6aOrW3A7LkVJRa4Dk5SX12OGDdbLfk6O/fXIt9aOWpcH1FsMJN
X6mO9EOZttdUzOM6PtBaYgMcxKDCVJH09BQImQJRCqtJwLbIgBt6vc3nCJFYRhpiNs8QdiDeWbrk
rfrSENOxxVfsqXd0Pmudldonr686C5VbquS7lz6E33F/nKb99urEjxqnvPW/IFtIEz3VPj6hPPUA
mPEPCmWcBxj6sASGRuUt22GpDkF1RnCZivZlRAfFTmpOZCMJ/zg1X+Ao7IWDQcA9Qc0AoYTJTvEN
9XV0WVh0e0vHimsnwIK3cK5TtMOxFFJq+VJHuxSITQbDJ6nYFIKWM+7lHGU/91Gwcmgdhx86Wt1P
ifTin86H/ss23NWbBbPJlmwb43Fzo4/x4YR5/L2Razi+5hWckxnTfzf+L6CHJ732IrrJffM40AW/
KBFEgJQKrGVmvqTcB/DO/evBHrj0s7ZlZi6x3PGMRtUu4p6R5KJfq6/4vd+rAcyy/AuRKhMDqLfG
FFhVG5fmsaZc3CGoffWHSNsEQ9pcZ/djxDmm1gJ/c40jCcWVmI3cDCELxezYH35SYbTJk8amR5hP
lEbbjGnYMlOxgp5BOrx0+j35G5wtoBHDV7lvpFwuY7yR6B6kXMmtcBD0Mq+pRZK/uAAJ59PKFixl
0QZdZ86KsOvPjj9cohJ5eEGqHR3HVlt3zfQoWJ1pfxH7gG4VaY7H22mYOJElsopb9E81JQZSsyV+
OaraGloS8yo2MUdJ/ZvlJURzOmOfeWp4Cl9OMtcyqGJgiiKjo3fT+ClLlt831zKHYZfyGmZ2WB8p
ra/mygBvDRPUWosx4wZtcP0A1BkBdSmuVJnfZZ23xpXKLF8QWHdr01WcC1H5AbFJ6YVLklsV+cfC
qIjVXWCQnoNQtJBg4FlfbMg4KhwTpxmhgSXdwjcI1XUkOoCro45bIvRJksIgiriE+cxIBPIHp+3n
QXeuXPBF4yEzLSxX5z67ARJNG/zmfijlAn0uLQmqW4RngUl0gT3azgexiySpvPvDZybgAs2Y9sEL
/GzilWWDJ5huDcV9URcyOqCr9AxoNGROYwOdO3RLR4CO7SbJrD3MwpKjtlIMiYhv3nJGCMfjbTUp
dHa6P+MUVPmc3wKTv3LUkr63+0BSks4jiTyxCI/CzkiasWsI+C5+PLrp/ZeCb04Ly0oOKZl7IDQd
xhrAF0RWxqhNV2ABGmNp4doOdZnYsOuQmmeNgR4rawMYVcXYk3+xxQA6uEb9p+7250Hetan2w68W
Jt2W8ZuCQnVF0RF9hwyejkft/1LKmw8MqFBu100H3Ok0qN7bAF0//QU353EbQvt6yIoBDgbE5AQL
U0SwuSeDDNx21s3bR4ZsXJpmYLZS8FmXzWa88gB2vt5twcQXhIVRhqqNqTYH2qGSU+Nu11NT/ZeB
EGAWfb3KwNfdT2SgxMsTt26EBVC13sMXY5X7/8x/yMC1BmBYfrMolAMP8Nx/U5b3UE5vtUST2TSh
uKkr5efazWHCv72Csesr/64IhLsBoqBB/rxHahBzrEQilwzn0ujMXzWhR7HNpaMn6xbTA7ty27lG
2CzcXwFdBfI+sifhXHCSDiuzALq6GW6mwJ1lCH78mrZ3NBv8x3lCTdd/HVs4vT6gpJFEdETf89Uu
EJ30RLcicvqnAh3zNbtceBwmxl6+c1Zt4UoWFagKJiWWwQ0bLn/indmOzdVz0Srz7n1ZDW3xADIY
cbmFfL8LTr3AV9tc+D3PIY2zLpGBTPNi5yzLs92nEOPVdLRP8EnkSM7EtmLRrElnDva+ItrlozAU
0KMTZfAkpXelMvVCJUwlxzsVpr9YNRrGsYIdkR41L8DTOTt4O46vI+AdaZugdAjQW7xKbjPkvORD
8lXi0BEcXYwlgLtUy390qtwAzOlJ98Vl3lcAUlGMLv8oP9B35R2h4l6OJH6O8vZWAACilCfe3Y6H
YQJXJV35ix3lQvrh9SVH69dEPqOKJlw3LprEOhreJN4Oh0td/QtuPzwBEiYpwPFNfxf3gk81Ij5k
hPDEwznUuw80rz7JqR5TbnDr2GvN6H86G1p/NpxMezZIxS4OlYh3Z0FNRCLP59wkjQvWkrlDhpT8
rylA74I9OcnBgiuxHxT5+kUmk0vOIjbiHyGS/IJUWeQMeCYljq5NREMcCfQ9e9DGc8WCQ1ytBQvK
P58pOluely1KLHEzen1+mjqUlnk/Jrqn58y4G6kDusosVrZH0WNOFPuVrQDeyDssZDOKb4LJrRR3
/cW7mwy5CSRY+bCm1etI19+B3SWHbaQINTWk7kP+B8p1XEQweyvJJgTCDJzy6/V5CLwwCudTryIE
8xdPX418SINv0TK9njH7faPpaIC038pR4JnbpkhSSyV3LGvODBNNglYGRk1tOP66ZfVU9P0Kxqeb
P9j2NiRtKr3tkJzkFeoCATs+xlesihIE4GliQFrOOlnaKZqU7EDAiZprdBCmwjFSkOSfBG8ZBP7Y
w+k1JHMu+P1nnb9/659iu2DStJ7dAi2eNtYkQFLKaC2nSNqDK75O204/hnFn9GxXJHHRVNCtWDOx
GpIq8EQj15A+kmeGfWdIZIqeK4R/Fy1kasDRY2jUYF2g8wF2wetl2DKe5ZolM0xKrLDAwu1wjTLg
v1Vo+CcNnwCRofCb38WCK2FHyA0TQCK8g8U8kSZ6bGkkHF6p1Z7DQjqFXJ9dLEkFTsi0SfHG/W+n
ZqM+NEr5UKInKwOhihIBxQ8/7Ef1pTS46x6p2xQFLDOrADRrQVEsOqA93YCZ09+ymBhtCv9aj7f4
8ON1d9e4g8v4/RF6up+ROwxw9S8zciEa/wDk3QLdU2o1qWq6vHcKOMukqW/FWUsQGm4ZJIn+MEF8
8eD77nk4F1Uf+Hrj166M8gi4XocR71LeEJwBtaV2rfPUyY9uCenQ0ndwZrGt6GZfzeGrs/ZBZIxA
j4co/Bdn9f89e3Y1cBHu9dnfwzfoJMCbiTvTX52SdMDxByBGn3CM5zmhbGeyHpgyo/oNtKptgDNZ
wKgq1Z018ClZSxKQxyBhjxfniWfWGlIzAKK0MMRgyqLxGsH4liQnva2DRbiGS98MmB7ubqTL/yM7
NoFrGyFklVWSwXRbXImmjOflmIvEGxZPYDlmXBq9vL/ov6CKhjW7V3cIFSzsfkPuVns9NcS9JCJj
2ed8A01csr+mBs7IxTMWX4kxQIvqpxNlVXay05GMRLzfZkzkc7jrB3CbpPtoWHuoKVI67woGOU3r
VyP0Mf1bEEVj6zXu2apFjz9RfQQUZmdLlfU8eZe0/F/9YrjBF1lXYf5YfUuiVv/cChIxmn+TGUha
djabxS5ySoCbyCqOsgk5p61bwYQ+n3cYYN8QhxXUSKspa4wXqCOn8dy7/O7bbjrAWyTgfEL59dRT
i7IYD5FQOP3M8iTzfhrWsWPWxiqCT13MYoqTEDqVdFwV3ubeQ8nZF2jYovLMQI4P9HD7ITr3Yw8n
xFMNmQdrEBKtPzZ5Z+IDK1iJmidBBHhUKMprwsl+1fS+QgCQWdbx5HDkKDIzptKeda0MOc9lpAWX
Sx6senL9TNvhKSKsrSRkouphZYjWE4AjtwODg5QAuT8BKCjhzN9T2xQEWU+1znWySQGnxrPXPK/7
mUPP1nGS07yfP2Xaon+T2dy9xgwlTptPU98C7bGXEDnKuvQeRyyFxZTlpoy6Hz1mFhy6k9VO3aeg
4Re72vQVyryFkQZ2WYnDb5af525KXe9b7d3w1WMFWYd7AkQxqlacIZwoA8L4PX4LXVssy4rL1kiv
uxdcWmPjd/e0seSVMxmUt7PT0A7gBUpI7eTH/DdrydnLGImVYzr/3xvQ/TDrlNI/Fyso2MNo8jT7
Ah4BLlW+Y/J/43/2w37mgi1gZAvPG55sFtINRSF1Uu6ZDPuZyuMTZNQ1IL9XwrNAAdX3H9H2QvgW
yzEMipSRLiXyRuIBjIHe31MbzYsaRVq0SnF7tnAOtqaJ3chq6uMV2p/m7uf6znBugljA8KYGiLPZ
OW6YXDVn7LxL4wiX6e0qjNPrWZpSepBTGCLWRq8ZXeS44PtgX/68hF8FNUR+3O7banZClye3pcQr
x4hs/+EUYcGe0kK1Ed/QHAcg1dAtsWjt5DhXAgEcCTvjnzcKvXiSgUXiCtlKyi60LMo7V5oXS7DF
bhNlT6W37OYnnUEThpAoZu2IPY4/xoXTZNiNPlGRndB4Nu8wmIzYTRdE5zAEQAxUJ5W4/lQMzZmA
vEDgZAmH8SyTOmemGfZQGQ9aDpEa5G8Exkgdsf0hlZUWXhx64xGnvUrYeNAAkEShuQN9nHIyq7y6
pI/8NJPo0UKdtfsW1C/k1erPr7zQAnW/YrUKDGYfWYiAJ4IktGUVLigBHj/9T5PhJpfEbVv6qkxR
BEPgk6+eFq5AWXcizlSNtkBoOvYv0ci5gi3AnnnWcR5aYIPHKgw6dWKR9w3DxNg20cGdmAaUMgJX
DMO8SX/8n5LvkXyvfajtGYIgM/x06MBycP7gNwYiZBq/SvVgH0vxn4I8dNp6NGx0L+FSXelAcZbr
MCyeZ5H0F/HMbhNlwKnJIqDiMleAHi5SynYOH+HJZJX7m5xSqv1HKdJdSLMFDEbTRcdFHBzv9VWK
7HSovvTaqMRxb9xzfjVJLuLo2LV4pgzqjHIFbNSyTIlk4u5ww7TtYZcxCXx+JAprTpng0K7vQuzm
0nRA9A8hjmzYydU8t7P0Mfm2h49dDuEVEqZIxuw769OFS3U4gsRDCslUSDjkp8rwXXBhEOB89SwV
auFwVr134SzZdSGbAX3vfu9Gdda4vzhOE2EDNi6qYRei0jtk1m/lZ2FPA7Sp75lOo3zWoNBMkBYr
CrGtll/PZJ29EhzvUh9wuat1dahbNsRbhDGk9QQJEAMrw9o7z3AGmUOm65yGaoMmiLH8jvxFI0bz
YSR8vXCwiXNQ/nwI3gs60xOGvI40k0wQQ/Fk4yTKYM49/6KcQvlx0MyMdaGEy8cxOBrn7lQpxzNy
yRyAf8v+qbL5m9Q26tMqhHk8LKj2J/sNg98Wu5xjFQACHoOQ0jrApOrTbHeC8FFeHKpm3O45io93
pnK0l7BGJFaOWHj+2j3tRH5biSCcu9Yp7teFDrR2ZBQ/LOwGZumCcfYysThPGbzINkWyHcaXWgwC
UMvoyIQyhWZ7gv/3qP0nhrkm+kHQQ3jhj6tmdqbYJRrmyHXonzxTYSZFcQ/mnpeElaHGFjhVpaNW
MOKZmbSc4kcZoncRaeSM+KCy8FLE1GSsNrOkXgRv6sD0vjh75hS2OCDD5ltMCzPn6An2AHNTpuaN
XSkuKMHg6EJlhv1yQjd5bX8PYLs3B0xeNLY4NQnK+a1M0HlZGzKEyfbTM0hDoYLhHYGDqykC8ZbF
I+m8iiqriPflkJs67R4Bu6ypKTCbX2bYqrXmGF/nebx9T2jl6LCFtLUGu0c5JVFqOunlhgGu69yB
zKE1NQDNJwJvGyhiKJs0BaNeexwKCPLOLnbe19G9lYqqVsQAscel/zU0qDynxpYIFg6lAXQnbbn9
eQTrTbt/esKl4EtcwaC4xyTCsozx/KU0Z+k5ZhU1u14u8moSFe8ey1wKblJiE8pvPgKQ4//zNMX7
FxbEeJWo5lZMK3g9j0BvTytctcckH3w+6Pw5pbt0DqK7GIfK2t01Fy1+lkKfMxWbnVt2XoX9/1qa
S5Y983+ATGWLbzmvYGMg5rpO1pQn/2ynu6kexRWc7B3vj3NQRasDVXUOsySDO3qXwttToo0dpAPZ
HhpkUtb6BF7HGlBzIEdWy9yQkNJ2LX1AmERDpim38cE1ZA2XgSw5u+EwmiI55ska4JhIjkMXdBG3
GLiln7EtwNgk+Ek8aHlCaT5WWn04l9dMYyuyBx8QJGaBNXoP28kv1H234Zmqngn8uVp9PBt6LSCj
xgGUrjslxl5URVkiWE/JOkrUJgSlrSAPdDzzcX9Q2WYgTfhvRc0TKwnhtWMxsYW9EJjTicqEMcnl
QRBdXzmkWq6rDrmM7Mzxqi8Uvk1ueh7smXrLD4zwaY6asPs8zW6QJ+6ga2vN+Hx1PRN9Kj9JSreo
boxFZkVdwjoI737J5581hX5miZdcbcsEeM+RLyDrlTkP3OMSwWWSa4iD8BrW3Iayvvxb2C0dfTMi
GpHlyL+FUsl+cZXAFwA4K6OwEbB6V3nwttSjnMVLp0touH+mUHudhdgimYaEt+Y6g3Ifps5xR+vX
wXp7pky2B1UWoMipjfMU5ceqtJtr919NJkZPPhLC2yPygyzOCBG1wTOWx2EWxzPYp/1GOToEYkDH
i1Efoh4atX0o1szdQ830OFx4JWSJQP9akHsGvORqUgiYsYbCalVdxuDK9MDD1hXdq6/bWxFNcjRP
abdiPYghoZ5PZjgpEZNbe/UluLvnQQnbo8BPyNUfSRlduBjuD1UUp0RQu+nFjybQjnQgrC+lC7aB
tdfwsLyEwc19j4X40BVIVLUb0+dGOwq9NflkSf8av94IQWu7scPC2gRRnbTZyIeLGfMqfWzVIBOa
1NpV56o4XfakJnVJDTL6NZEGhcLdzkZfXnCxaBP+gPXJ4zXBdlqYmgqFPexVfcrKqywGQyu0INIp
8G/vhPFKNOmzDk6OJMCX452qMQV8iIr7KqENlik3P1He3IU01Sh6316DQiwvSEkisbdFSCXX1vTQ
u2PEwENXOj8D3sQANcyIB/KXnAFZM1eBwlsm/CtvKRjk1HGMZ40o5t1mKMXp/mlQTxxOvqiVxpEe
L76NqSPz0H+4tyOZ5mpnzYPIIPDs5jvD77kjI/gSHh5aYVP/6xoki59e+shtCZ+Dm2V/9Ahjr6Wp
Ym4zkJkj/tObKBG9S+2ae69yS6h09dA05ztykAUXc5hbS4uw8oZ4xDTZUa+/2uBkeMSN7sTD/9Ds
Q00JAAqOwqKxMeMVaF5vx2+w+ppG99huxeW2/GLO0C2DrqjeHaq2C/xAWg7wC79G20Tjj08gAv+e
cPvRa4H0lAN/X1huxs0CcBXYw+NJw+ipg+ZmsA7Q8s/AQcUHy/9PfaT3eOaGN5TmbGpT6jaB4UBL
zEovysUVfiMUCMzxoBjVyUqBKFbYPIKKJrIUj5xASh+w/5BHBlqjZ39h4IzMMGPNixMec6viGAdd
d+6+fcfZxeKY2G0WNzBiYmHmJI6F2os9YxXnx8DJtr4rUHXmZuDPVyD2JTtwRewC4Rd+/P2o+rK+
NPX0u2qQrUxZnSSxDE8nUir75v0Rdi6lYcnX/kVvQ62xQZY+W+EXmnbM5ZJ0yADBvKULmovwdU4D
63hF/OwV5W+LNg/ZZBR9fdkUAxpAHvvn8+F/wClLsKEVycByLrN1b0gx6Fd1sdv6DiB0QiYIX7FI
iTO/me4/332QjIWsN/4ybrI+oNrsfPmC19dgryeVVgsSetitroKeehYgL26Z4bQd23AtH8y0y3Im
esmdRh97ObsQCdIz0ZEPiM5PAmS9yQrzVTevQvmh7iqEtYfT0B8rR15nGwrFO/hJTHEiO+q0j53K
8GS6NoHJHbm+Pkp/1xvf/UaZXI2pn2i7R1DzG5fwe3YDFYjMWR2qGEDAudK503rlK/PHAZjVRjJm
yZdCQ3lU2xwgKnj8lonVKGIArvWGSwqHf8dQL22AVCTImYNR30x8v88DXgyLK2WWezpC2O6oGW+h
qtE7meFG9BOBazAEHMF/eM3SabQ5EZpKqYHcCsgba/a0aDT2H6jhsEWDIpfWLytHyVCLuereaLXM
9CSooSTyzkyENx/8fhyPoEVaJo1UegeqCqoUxMpMkYvkB0MqOnXHpbVqmYmCYsSRoL7KkXtKb8hE
b++FtYjrIz9Ur03deO2OnvVSe2tTXebBKB3s8pCIxzqqi1AVcJEZIjFaOALOmZH1u1nS2fmlFgOF
x/b+Ls8oXy2tE3rVa08XXPw5x5xCW/XzoQc5owFUG7PE0EWZKt7ZQEUHBoZatCI1bbE7bhyz2L/P
+E7nJgnivjxXXXaYLzq5nrdNG+lQVI+W/Ao9nAVDtfBqUWTBewRR4IaI/xh4vrF8wfQlks1+3wvj
LeZiZ0S1y7Qzp7rkSx6IKwe5SDKfZ3zuvp3uP0r1Gw4VunXkbRwr0y0Pedpn1hp+0C9vBaDJDoWk
K/9jCcBLxZp9uVzqI4ak7ivgGMoPm+85NQ10rAUSASINHhbwQCmVjcjRcQtE8vE3U1tepwAawW9y
KW1l1okojX9A7obcN3Omhzuw08zavsAe9VEwhSXelz8anxvul6KPL4aNeSEBRwBKA7OAE+wH/P/+
3252q70yaAyLo6dmokeiqVyJoygjoCaXQlFpUsDDSzbGAvvg5kb/1Tf13eSesZgGlYu8J4NaAoSv
drmAKoJbxdNaBm/ysgFlTp2PRHcEVnFbSUEnfq+5qRlXyeftAWMku1G1D81R8mEQEnsRW8fQeqM0
TCovcVurqmT9NZL31g2yJVs2q/zK1Yv5i6SEQFkghnvIqIIEdYzXqvtNJkzkdLcKT5MhEgF+zHTH
kaeKMc4Y3lXT0oKZsJywofL90lKkD5yQGQ+lRobr0Mm2pyFmRFTsbTaPZJK/kOmdBXQb6pbF2I2T
2ZzIL8WBRn8GM3+M1dUXHMAd8U/qdUWdt5IupJOaE81V/gb3sijKOQ0sblwJAArR8xDlLITZKaOg
8lUU9XK2j1pT8kJx8OCAaeYCoryi/XglT7nyABwGc/iRoNcLgHJlZRdei3KBroMNDC/KHXGw6TH7
qKLZhIIoH5EFbk8gGXPiiSaVIasUvr8dpYKYAgouweZ+myxm8H2QkIC6k84TVu41A/mo2kOmmuDd
p7v9Z0s48w4s3ftGlFBx8EYEfXGCwqmynutW0K9ZOZF5StX6jJko2rIzOBnJcGG+zc+whwmnP0QJ
7g8e9qFlvjPL1IaVpkwpJH2e6JaI9i8D7WHhbQGs6CXSPZu3iLaiR1Ls7K6QYAGe8O8Fr9VkeLkE
oGNYyDhAI5vxtz0Vl72pjsihMg1RgKGf3Z8Rt53WG+p18lz1+gnoqN8OGUFFh1WY+NBlpwwuEWEc
YzKy5EGEk2tf+hxVJdIVPkNkL9hl9z27rhJxhlmHwZUHgs/tqJu+wd3i9p7CCzqDWUSaHrHVte1w
gkEYpwXvniSL/yAS0G2u1x0GoLuMYK/uJCMH5cTvx7uKeckJVHW4pFgJbAvqNJBl8cM5arP//Mya
ep/fy9tqwrOwvpvYBRyGxK0xDadU3OaX06YvoD2GKUll4DU09wJj65ZsFqapRjw1MHWBZg7ga7fS
nfgnRvb+doTDcWBJVrKmjDnQNNB0AiuvhSUom6G0UwaSwuaHTigREKBvj0zc0GL0uTu29p72FYYL
nauXhNq7CXWSD8dh08LT3YFP8RePatVMef5FeeHGSfX0Wp6753+FX0zQobdUbZfMcpO18WwYAKLA
SUrjqEtM7XyjG2ZUY40N2AbrAwY/F6g/vjbyybpDSl89SSLsMg0KTVSdAnfVBuZdKOQKv0DnRoam
B5fAhQ1m35PDZ+m/18WeoT3sx826TL2iIq+j+BWBbb0fJSKUXxUNIK8OItaRFjsQw3cSU5SjAata
MAgACjO30h8Au9xhFLWlFTRiSim512fhNv/xFEXmLZmhWrNOerL/jt4Vqh4srCysEBpKLhs3XN4d
sdAdTvF/gjL7iY3ShhxWJ/KB8TiEwaS4gyyR9arNylvIxhBy73MLQ1zB3Uf59qRfPqkN8vwxJOlv
T8m8xPP6ZJUjQRNlGrrr4ukP8r2nxgjtzdgUU+wWPfLgfQUIQrUiLBr/cq4G44vbeUuRX9/wbT6q
Gdqd3K2nWrhqFmevCQAq/A2et9RyxzXx9xNUw0PJqSOC2o5JyYbYXv1knjLURSKxHI2eNVLc0kK7
Q9W/RJ+Wcc0gJpJ5AMOvz759QwB75lleRZ/QJ52bVEh/60E45RPNi3Vg4l0XRTDV0APaOgTOmCkD
2o17CqFbLveNG/20I8PDetVULFRBRLJb5ogXRs8e2ph+nn37/DjfkQljQHFliT4uYeLY793UiE8r
zHvIBVbjNAdiycIV/pX8NNSdZ5HldOCk+s+/mRHcodAR293UvC+oszRwCOBeN5xIanoos3jGMnPF
vFfmiXcYvUFkXKbvOjRXNAxZPMBPmJq2O+Vsc/rypYP9LS3jXjz3357yQ1e61yF2+1YKvVtTrX4S
KT/PwDQ18Wv8vyyTqhbW40+MNDqRf7VXsWNIfTtYIC339dzAVmD0Ix5iIGQ+t6RVzp4DpyLLrxzq
11L4YZ/hErBuFyiCD3P2QycbwQuBjR4IF+1V4p6b12jUFPsM83ooTfHFieJfeB4n5Fforj4Tw62n
EeN6zJFTJVjvKzD8xSxekCPKhffZ9iFPbLtwvQu8pDPpgiEWghl398VuHhz7g/UUQlNG709ug+IV
/HqLWk3HFC0O3Y2rcaXXzeZULkCaK/aeOfJGwxtNXIRRnYX7qCYCQUorTSQnKIxMyBP92+bt1/U4
CJ2YSUKSupqtCjW62afsxnM8uwOOivWCqfRrdHSa4RHfLYZ3E6ACgKDs+9py/z8LakR2iObpQVm0
F3hz633TiKFZF+nsd1A4XcPKwcNcd17g/fjYXNtLtA77JHy8a6iPQo0pKxv0VrAYvR60GpqUglbQ
LoyrP+BLU9wZag6WWrQWCs/9yyCEvKecfzyxLLxgLKnKT7Tt7ax4Oq48tpHMCUONpeIgs8oduZPu
aHzAKySrKasD7FELoaNmQa9ycKHGQhdHNDuLQXXaV1AWVri8MolDfbE+yUTyDBU6z7L16NQ+mZe2
DcDtIaRafkT63liQf4l1Mgy4NONNt1ez8QNdzSLW+1Ukk6MZ4nobTxWG1yIdCUS3hwn5ivIIy/vZ
41+zkzttMnny3FDEO6TcZWUyU6X/DUkGyDRUfMEPkGT7+ykX9FjrvDh9L1Tgy9bfTmf5vWFcjgGm
zHaCGD36yIInueCO+V0QehtU1bgOV4qsSi7/KLpBVhi0NZFwma2PUHPdItJVr/37nat6VKsR1QJF
7xiNocQcqmUWTr7Ops7orcC0hymI6YCFR/BjGFn4yVRMgw3mDB1nN1a5SQsG+gTjiim0uYZYT9YL
9H0mAj4p6Xtyty8bwwlx6XyR+xg52J2FgJ9UkmccD0OHOpuDzVn310ksJFqxS7vNSWEN1ctt+tq+
3fU8kmPVOaPSKYaKLwXdndJWAOO/M+KLlBMPntyrmxUjLqEhRvuxOlWoRWN8FXtcpdlptdffJz+Q
9NNxRxiROyFJs+iV5+X0O4kcGkBIBiDDJHTqRVhbaNpyeub6blEZecSoMwD1CqCHGNdJvNS5amd+
dDN9U15W62PU3fmvDXTtDAgkHawzisRe0xNV+3EQH8HjxhgpCVw4Cm3+3PimAzy+zMTz0J08nK53
CRDVz70VVmUbo83wQ5lH65prMAadE6odRhoA9+xI1bh6i6gxA82Mq2QhXsofgLHMI4WjDKvjoF4O
dcAkXQvHApOuVteXxMzWHkMHOFjfkljmx4R+6j1ABohtujL6kYPx9Bq3/z0ALKjCbQv6I5EUo7tu
1794ebAVV6aLTHTiHnytFiKCXjrzPyssk7rbqYsVltZvRvg8xkyqoGpFDRM07jWEWqOt7QghpeYN
/6GehXRoEWUHiUxWA0jIIGkFYkQqO75U7h83tf+MRRjO3zBTRmP5kT6oKG6wnLR0khirooaGSozI
1a51hZxdxKnt3BhLAFEwDIdcHSF7l0/UCVRleXQhJgWahK6rKfjzAe+wpAWfFixHOKC5iVM9uCzz
uAWRNBHdW8lfR8HruyNTB/QiMSU0aINiquiTl3uWJC428mqastBoSlIra/dkjmSJ3HOe3A4VBlX4
shzYtRKojL0HXjKUTWDHB1Y0NPytc5BHBd8O23nMzFmJUQINmJ60XnZ5y+7ka82k80LUnH0SqW0b
LKfBW93E3Sxt7kfpUIJaN1fWjHhkY8iSnydwgmFdnG6ggJffO+kRU2AIfx5l1mePM7lBS2zSDLu6
Q37FGQCzVT8Rspt9FI7wFOsYbS3e0N4z0EDK29jFpm8Ewtk7h72Bjze0KdzRXj6Y856aiSJKP6zK
5S26GVhRooo7x6jPpEwCs4if0Fjp2t+MTopvpJO62lsTSpeWr/z+50TbJNEx9RKfyp2UyIaTNCvO
cHnnilrpQP4kOiQVkzAm5VID7FzG2bWw4hxPxDYG/u51o+/n4odKA174iVG4aSJ+SZjOewF1lJ9Q
GFRHd4gGmXFctkAV0+7IQmbD2ec0PATvV1uyB3pWv1jy1WGzIWrCYnJzbwHzqhQ2SoafPTEAopA+
rxcSZa+Lu/pJWZqxWLjxItUdasbHsjDovXfyVRk8nbJSBMqQI4yxAFZg6MT2WqzbNWEWwkaO5YOJ
zV7ZD859GCYIDmLlt7lZGr5uE8P6MNIdB+fX6nRKVLhiw6+c8KPCvGZ7KQl7rjAh8AuZ3acoL8xy
Eay8dOrehzIOFx4ovtHUfY63IfzOPU0uOlamCsoq885gEnQibR65hPGce8cy/ET5SL9JmiDOC5zr
Sfp+SDoNKWMFGT9D7jBQdLmmTrPZ4M+EuoUnDm0ZVsR6NjU6AhcNvQH/XRws045JxhIQfkpCrBOC
/AspQ3ikOiXeY88g/qST3ddGIuB/ECaryeMdp4SCovxvqbhKLybfR9Fy9tzrLxgC3zmGaRL4qMEI
2CaY+dLHnDlbvbtLVfHuNnpyZSA9WvJdgHv4g1NlEBo32wVcjrGjkke23lfu/BfUSD2DiY5aqj6Y
c0bKLt6e1+HOPPgh8+cVCoRsky9lb+WlmheKWAqw655cqXMnO5LCmJH9KAoD+yTOneb/0/1QAvSx
3k3erpSHIv7oXOxJmOqM+MOqN9fmflh1ukZigD0Fru18vTmzj3zZODud+LHHA4XXX1iGR9YvNtYF
KkdonKfTYmtcTNC3vJ9tY9vret0adS/XQ8MGUFnvSEwCGXiluHHvVXk9GtPODSi0orK673DP3XXD
4EFvk6YMKJxT6tAiqi3buinEqAJS1UK5XY+kBraARoEmv1Dif0wn/NJJbrtcJJOLsCRkeFY0sNVI
e8ktwEHqmFl+4DTTYXbqdxe1tAt1g7ie91/NvPC4YsrZl/ftOjE6YMiSxkY60U50/rWYwXPbMepG
qofb70LAc2W5cCJ0se72fos+QWbv3odXXC4C3EbJsehABJDo1hOEt1elp8KqDnmWMjL2uMhiJHDV
WNCRnJVikpL5GjmOgB6A+x/q5LPpveYJMyf0D04to8cwg7Iec6aDUTWhjC6jxpRxxUzr3CoGUFWP
5sWkzNEmIFr1fKic+HswB74ow7UcY0B2QSr5GKlfo+TP7DJGUAWT5oPrUUOzQLct6swJlC8OTrzf
oOORZ1d5LKz1cleqf1Akr3pGdftQH1A1+I1s5m5lppRDrhvs5AkEtjFUuB5HjvLCkwPlteIFwvvO
KLn10UMtVtjp210niNdcdr0nufF3m7Ti6Na9AePoh/peqXgVHdf1Z+5zdKUOmdtR+dp7TRZbvpAS
eKFxuGsYw+QQ22uikXPoIWOkBQ4yraVo66MHSjTtbKB6uCH0Nm6cbDnT3tGm4XM700cw5dF2zaSz
dJGJM/2gn9JAKuz5TSqQUag1goAI0YcQCflgmyCnuhSSFdrPjUiz4NlDM/Gi7D7MSwIQ8R5lb2Eo
NIXK2P7El1Ue0YDP8d+D7UcEXCGy2WpsywQOoLJg2e8eDGwA1M0KUHQ4Dlw/WVh62AXA1JNNr9Ra
EwouusC3v7wCA2Lo9mr0tlSEFt5vENLyhb2lLjRH7TqrYl6XK2f2WQS7A2+97bz5GD+tQ2cqFWRW
Nuz2VUm8X/9x0hFV8mNHzcfDSqK1/TmzCJnGL9Zc36WuzRqfYVOLnCwnBdiKCg8G5/o+oEMpXv4o
i1DK32DECV1TKvQV+jTUFRQw9M+DDRUKZ3c+sb2HjP3pRjZCOApDtWlllzG9lRY3C6MBeCszSCRj
cqpXwXXufT3LDzZZWJ+2zaaFwv38XIfsNLgQ1TDy34xojRRpRx08Zun2UJYBDoMBj8ONOzYSLIo3
WP4STU4MPzq57sqYqh8nVh7ehHkp58YLvjZM3RpFQ3OBP6PtYeD1PZTzT37ChR72TbM24x2oCom+
e3zTyRzqzrvIHWN0rWJ6inLqD8SQeafsLrp/9zRKPZKkVkktan76LXQbBko/chZqbTAYCaNUIVR+
PTcQbp62q/y+HnDCboErOxmgyz2XQ67osbrbihGawFdc3OoAuxPGOXsIaiV4tY/azEPRgeRSTUZt
zFEqzaawZ8Bt/pPhHZdJrlx0vQqXvQGxEK27Sr3yEqz+AuuqqQUNsJ8l8Vxu0oZ4WFnbyRWzAEGa
ZpaT1fp9H84FrkvH7QI41cksP+pRSQ1bE/YVuZ79S9UlxDsPS0qDK8FCYVQGRBkqlWQU/Wh6Tua5
TQJRB6rEUUpFiIIu9zcsS3UwPgas0f9BylQpczz9Kt/IUWjOEuxEYOoK0urQh32emjlel0H8RjMw
+h7vngteqQTJJF3teoA/x1fxvGYtZw2tS6E00RZMAKM5uGY9zgsxp32PV7XgaEgGTUUuBcf+aPJT
inFG7xIEbH9ttTlLk/ea2f/pbu4vrj0suoiidfZ1CVDdoiIgIx5d+1QbcDLfqsaF+MT1vTr2UXUl
vu1ufHlbCWP45hrHUjkx5K4xN6Hx2UPzUXSyi1tbVwHux+GanpWzJoZmEsYtGq0gAcTuU9jZkmZZ
HKOM/KoJ/eIv34h7BsXY0+2fBrp5cuGv+7emekmMv6DWHnINaNiuxyIPBgJ4i7u6wz4MGbnbqR5v
M7tYdkVJv53vAf/bDJ7qZuy0K9t7WYYi+FUlTedCTtB5Epm306gkh4r2ZIwsCB90XXnWXPXqkSWd
8KJsRzNhhSlbLAM9WzpnWI1XyVmOKWX6iITvX9el7m7T1elyo1CUR8fPJ0jh2pGuvlrEx8muhoCB
2pyzFCdFKEweEJzzao+t7bP2wB8Eup7/0F3P76dmOzpdaMyW1LMgHTeJJlABsd1NznZ2KB/eXh92
e0ZiR12gDOfRJVpoAOpVpu2vRV9aXpLB6CLU8/qp4MkI7wGLLqKS1wPdt0j6qvwS2MKN9tC/1gc0
NIp2cMNz/wOxCtxNwZNqTb9myz9DmKnF2hksX9E6PB70coKAu/OgF6rOPBTAaudFLjHdGBRuya8h
m+KKQ73/HQ9NzW/7GfPDkzIZMlC3aTHA1ZsLFiWf6UK5VjV3bt8pwZH4RPGP30pzmbMS2Hth3wKp
W3ruijXgF6j4CHzt8WWMA73hEgKcdcbBL3XKXen/AAQSxSx5Q3BVrq2ehKbnYmDLGQ2r8YTqRT5A
WSAem4E8yJw99HgOnAorTytJaIpA91IdfUBitsiVKlQeMeht1YkMmq5GKXAYCJx6CbixLFj5tH5x
zREED1eK6+yYR1+/hU4uy54SGGeMpShP2QNWieR70z2o28oyCQ+cmMXtOvkxIUSTHYwlROJZoDl9
xIpb3U/INwIIM6L6RSwHCN+Kfy1oXR5EMgYGHkY3gVzA0xSorQydfHuB8oEP/rr8Fafv7L00XfYT
+nSP/YjhmiaNv4fcAPDMAUIu1q7hM9AVjTEiaOGmvB9IyeHmZ6EstPJsePikpR43z50lw6oUZYuc
pR/riATRm93BJauYrmvbExdZjkseEIqqay6j6KUAbjY+rZrrY33hayIf4npEVFDdwAhBf0OfO3nq
N166f7wNEb1RC2x+V9x1uHQXW3fjf2WHKX0tjXzXM3BRUMNCL9m9KN1KKz6WTbc0pa3q1un47R+L
o9i1mquyko6Q3PVnTBQjB/MorcorsrUyoK49w3M7Pi38swVfamU/iUDx8tQ8NClg8yXn5qSbCWGC
2YA8RFAxsqon7r8dSIram6cg5T5RB5aiuRQUqI3TUhXtSGomm57XAwGQ1Uxx5chF07X4EqsRXWuI
YCyoyB4IGDCm9oCAxYnJUx4xc1f3GUmQ6J3k3RFeuheUNtlE5WjHxX/yQtz+TWz9g/hJG5tsUhW7
iYmidv8Oaww3luJ7+fzVyzA60KdmY8AXUFsJPpjRM4O9qB+ctxcZANXVK4+ILZx1dknQmHCpjcYD
gHKsGygozUwDsAo0KjxBPuEfjkjXlGeZxLo/6HsJqsglR7HYGm0qGUHh5a6dMhcnIEvmZadYQjew
90ImrHE3pylWXEX238Z5PhU+z+fEpPclsCOqm7FJgAAO4iOqA+gE/KcmlhsNN5iWbqOi9BaxVme4
7ALyBZgZ0qLlvuKS3N0fP7CEkn/a6Qe4CJf3v4u7a8Sesnq8V5epIUzfh7sinPkdHSv22ANyUgeW
endA+vzD4qhdLSne27q9uO8B248X9Fsv72Q0wUPcc5/VdzPyHUuTXzhkFxt5bZ2igSmJvsTZFR58
kFbQ/UjbVZyIRWXJ1764S2Hl79SS4CkZeomT0RUqpgRrvnCwZ8inf4jE1SBLee6T3yxokKUdNS/c
48bk+uQFl2KzEeUhoJV8Juq4NIokvZsVe7+jsT0Wp0OWXllUwpP/ixN+WpmxnB6w+5H0tvOvZ41+
0Z93qGsGrmOnESP4Y1acVT7yOjH7ZIUkOVO2HRT+Ue7RrquE09oN3gtVnI6C4QqW/YkDhVfUzaHg
hMQT+H4KN/+LzwiS5EKPFL6OLGXP5SRGhXByl2zaaIqQOxlOEV3cnfHGLPlKlPFa3wWNHpfJILVy
1lBD6/vpftdDqcyVgWUCWSqk+Qy04K7pX0OGnlIiIKDpWhclmMTZ76O3ixriLHoV1EfCfXD4xUQ6
Whu/612WFZ7lISJ8QrofiE/f65t9FA2SenAEbu+O+3gNp88ktm2YFia6pSN5L3uX22S+y3vO15rW
YObnorQc+Wp6TkVFBzGewvxAIHWpHqAm8tT6wbk+nTuerdKggF9XBswDNncu2D35M3MaNwLK/E1j
WWOmjFc0WlSYeq6/0ZCKc/9iC1GLMU3kNJiIgUccb/ZsGIFtQ2HzetjK3aHwKOpPM+8x5SynOtYW
XLeqMFnL8Q4CLp8+GFKIUEXzuNdrxQlSIq4XQRWxZ68cEEY6hBJJn16FGVz6lytVgPgvXHRXqtNg
IijnA5l5jZ1KFTNtFW9Vk8ctf+ISdQAufoC9gQPHIW7eZUz5C6rsRVine1vXLyOumXURmUPAPogW
wpWLfkJ3wwDulsZYGt5m93+zl8huat3LSaUuCLcjjgq7dYP3B6kp/Dq41aiHThU5NQK9dqPvma+B
aOKOf2annFCRKhlSzphSXHrM6Rr7VRBnXIb/nhOII6Z8e8f3c9anA78GDoq11UwsbzlvDVhBIXzL
NrmzVs61m4JQLH2eav02xxCN1C9JQrIvFI5O8UG8R40NVnrppsd3l3a7mftCB911q5b/2mgsjjCi
bEHDW6zGyUxSDgcRQafMnH5n+meWJAVHQ1xdEfRPgP2xMu0RRgq9hAc4Fk/eb3pM9mBQk1Dl2BTB
lGJxi4P3NuzAL/lNM8Ow2D6KaSWTJr7/M62ixrDV0Ev7gduAKCVk0iAoDrKy1S63KlRhzAJM0iVe
8GbncqZ8UtTEf+CJ6vW2te+zfkOFoGC9K3TxSohieuaV7PgnZBv9iPR2gZIVQwNcUcZ5fI4x/ojk
ZmrJfMmEupW1vrlIKotGsy9MKC0idZyHZce6SHS2QD0g6+u2JEgXWZttyKIYr23meyBUwYD2ivK0
D3dv6sm4ZwJPaEYumAmUe5insp4UwCgaj3hKYfxocrP9XbPcmJAaPM9fLe8PdE0JHdSzr+ZK+h/2
p/yTCYZsV99/mVM20PsIRM8CqfK0W/4S4hkgwkBkNIeio3zrg4+ZEXkY0Hzs5oIKDmXBrD8oHpCW
N9nt+S0G5nOZ8jX205jSLKO8vkbxfGEXDRPQ44RRSfTwzYBVSRzBUeyxGQ7wLlLElEAPwjgkzFTj
rh7n+c8ChGmwmqX6BpM3ioBDAlWL8BARvOCviQo5TPvoY2kX5Yc6pDILv83GtIBmFKPhcXg4E8Sa
ASjE1KwMxl1pnMhc+r7EAaWjC75vxv1go5nTICCrOdPUgROOYbmp1B+ZXXirnuGlQ/E+WhyJWCJR
ujtI7BZDzZzGzscDxGtdoX9hsB2j8TkVp42qWUmw4rxwcS06BeuLVL9R4Y0ADbNbywVFe1DYUq2K
K5e7XPjkZx6hgUs5oangQF7jzGb0ycv5yjZmKeg3jRJOJ005J1x0s4pUV2exPw7x5GgJKeF1U3ZN
rEvnFMtBYW2pkxOjhRPsI9KD4aUYr6fe79YlrhWrWZwbz4VAtc+/udVyHFgOX+lQETIbgso6lH6w
sHfMFBOSZRrPx0NEyX45XT9s+TmUsw9zcUnaHK1h8EntLKsDJlNNrObmhmYGir9MeRvKLM0CcyvM
ZpRW8jpsH+a+EbAq0sn89Ku0fmc4XhazTzBwUdXL5zZqDn18twDlyz8ZWYk9z4cD0IIV8CeTPdi5
i9oPp31kR5t42EnXPXCdKBzxG1MJhW6+EtTV7U9+9Y8hSfOCAObiwbCbzwDLLLCQ/C2zg+liNv+n
ROJ5egxrUM/NT4uRPj2xi1AhnTsRa+Yc4Km8Z3RCTGh1O0h3aZ6WnPIwAnuAaLTmNVQuCuuO4Md1
FcsU3/X9HpW4L6zxvVh1UQ6JUm1AaA7WNive4Fzc2Ils6STlbCbbdxMDAWWkq6tQRzX2q8vRzq+2
j7Jz3ngqRjdtrS46Im8ojETpLk9rkblCslxF90JRmd+mrzcTNZu7alUg3HP4oT46TrYN7cdHZM5D
aFO22t5N85pp2p8g2Yyhih3bmdfe+RlW+lyAxzzhA9BV9EBYU8l06VDrN67WSamP7SH8qwqjjaLk
v1L4s06h75I9UXmnFKMLHGuk8WbEIHOVP/jBqRPnu0vG631dIzNT3toaKj2/9iHjzQn5hVtztc99
hqFzENTWALqwxBI9jthor/xYagB5kGXEy7ugNu/oiqzNEEW2A1lwByV/GkfnJQQhrcS93G9Aja51
D9d7P1Chx0NA2SGxKz0WBeczIfDjpdKCQYiP1fB0DcIZTsS1MSYVugOBTVFXfo7j7652ybRBg2J4
1Rs+VU7cKw3xdc8Rz1AabUmEP/KzZkvPvm33zIZVreHaZZq8icOQ/a79Os94myC8INietBKiwuXf
/2bcgfYOCYKR0LhwgNYM8UFynj4BHnwYycWbwxa3doVtbQKOB4TYDL5FWft+z6Ifwwsb0Ot0cw2H
dSAzw/aH8FJnGVYcoUaGOvhCAbNlJQ80MZ6HVsLcMM8rG9bTIQCTwwRMMZjFvo4odKFXeH6+5kJq
t9kInSqLnntyehAylvmU/z6gQ+bQ3MyBoeb3EHfaLyYlYu7D+5LCaGm9N7yHJ6QM9ZaNF8UApoap
pYpIl9QYsiZuC03FLIw7izzjY3oWJt4/TvumLQJDDGuokjYfQc9SYvO5A7GPR1Zil8DDmAIB145t
hQTUf31DOyVDYwh0UJ4a9pE90kFnpvIC9bTmwGp7UPEtj9FkujlFcQ9DrdyYw9Ry6/+4ukq71mzq
9Otr3yMUH9It/33smKONrCry0zdxE/Iio3hSok/QJzvZsawe+m1SfckReWP5WGCoA6SEPUi4UmDb
YuGeUE3qzyba+yYpGDDFA6zCeN9f0Y4WgQ9UWOF7YPEpbKB9/+JW+9+9OpME2g1EJ+lbKVDQIpJC
IoPdm8iQ/W6U6TYY9gFiqRW49iaUbMUVoYYVEPirIzxJMI8qjfmDTjKNNRY1s3vTNfuqNdqHZDGG
pWmcTeUZafJJfLNdEJ0k8N154JtliTimLLyltGcQtIK4AsAG7WCYh+JL00BGgxbAavZZeN7kGYDz
KzGz21vbN+rAvBKsrrq7c+ZiH7PTGzl/c+xPpCPRtrJuDbrbPWi7UdIjN2l7TMu9bLQtqIuuGhwG
KSZKWCAcIN4J4SrsscRGctgFsm4pe7UKS03Ml2WH1tHojZNJTQtpRfufKltQaBhrcBSX3x8lx9+o
K+uXrRcSuI9iRlNnxwf1sLnlF/DVMfMRwKx75IUW10wO1dCp84f4jAvExV+Xn3Wi6uSMiomceN8i
hH6/vYxQVQMmkVBZlbh8bGRq+Pv3Ez01TzmbPyQqDG52257OK462ZLfp+fbnNNqrImmbzGRF6pAc
NVxIYyUfw9j93921fkVtP3+sQzYRbJGQQqGZjPzfWeOeBpflxeAVwPRQ9QsMnSL8Y003nVLG8J+O
qyxcoOtpaSuCnHXDFpO7cbL3hNBXNoKLn5Bfi0rM5Yw9QdV53TSBQHNyza7XmeEM+pqLEU7J1sXL
rBJ7fl3jHYnr8HKDiLoO7cp3GHNswHZoF7k0x4wM0xdAF9KR0exdWhkxNvrNzSoy9//1aZG0MUdB
nV4PtMOvDGTHmaV2Z/jB27TcDypBn2eFntZ2TJEN5QSWMNSNFxQo81UONbuZtRY/4mJsFVICiPOx
II3jMixRpz7eOUcOB2nyi2PvyktQgEnOul0UqRBj5uFArL+bhYkcZD8xQfNI7wsrwxa3rkCeo8u/
cNocz7BhuWjNAMIqsXWqK7fuO0ygEWwEPLl/yYk+bPIXCJj9GgDWCH4IuRGTXVGQBtzVlXTHxVqT
X7Gll8A6h/QRXbBsiG76+9LwcP8uqRSLoEAPU+D3yjnrknfiirvzlP+HZCRK1EcS6VBLx9bgMiri
G8QHERH2vaICU0bAxgchiz8xh99LF8fIe5TgfFEIu1iPw0CVNVcN8mUHrX6GOn5CZrfgn7ICe44Q
CIzOovQKt7xueSpmakalYG3Z+4CvAzLCOBp92vsXfvwU+BRpnW8BtcH21AahIw0+OM67o2ouyDJk
k55dDx2j0tzEfoiva/Ixwh7FLFQciGKpG1i+FN4aRaonWLZGfLJh93+ADuSQDEZSpcCbsC5XK6tm
PL/VAmjvcWWWM+iZpx31AYBIsvxkvqMn19NVKJxMFENQqTSMDKkKp513cj30N+rw8Q7+nucs4RLa
8gG2vqQphFwA+sf/Q7Ydif519tCTyZ58LEHmtqnSN8Qvin4SJexenbbg7IZHxN2pWbYf7WdTXC/U
l1R62cxR09RQ6gk3HaG9+C39kJAmDRZSZIGekeaLlDGGHovVVM/7YF+OkqF7QPOKmmAM3myvEYnL
iRRMxxAICpUL/tAxhaMBoWFi84tpxEy6jcVdQtzH8C7tHouXWDaDQhnM94ctlEpxcJOGmxsNZE2U
3AxWC/C9wP8Hl54AxbSGtIZtzW+IxbwStiJ36oHLuzDgoPVMQyYc7V37v9unqSoy6gw5o+SlC+wO
b7WOrgLhbsw7xZGqTZs/Edzz80zUBiZnkHbmO9hZS37BLzUa/8d6tOKPxx9QiNSqvSf/cNWT0h/l
LSv6JMEG7W9NCpC1M2gCJ+CBT9WzlFiMQjIZS0uXbbXOw78KZGgqoqGq/66QGvWN+gVKTK5uOR8t
jynG/JfPjtALhSJfvCLV5I7Gp0XtfkKYsYn+XVNQ+nP/WuQ5Osy0ZNgW5wCRBKwDHtY5KA6+FYm/
1QCyM7SL6Q2mxZJOzwgR6C6vi40wPqH+SwO/spysy2rrBlPWwzfNaCTJmhp6mLy2CDF3N8w5aW9B
TcxjGj5aClXtWKB3DFZHyHx56Dl0YFVoi8IevtTTod13ZvdAOy/jsj8L2giDDU/HlJpjony4RZjX
nQwMtv8aSPswfgO0o31Jb94PFPaEILmJKDaROawHwMxcu3B+HO2I4tCxSCw4F+WK/KJcksgJikPn
ycy2fFAapKxu556l8iwjWRBSZS8KcMX4iJAfpYCcjHh5tlM7wttMenUbicH9P0LrrQIRX2Mk/7kV
XamaF737kP0LazCpurCPLlhIsfPowIbIFsJQ0vW549YruL99l61pnidEAtf351XYWvlIX89t+dYU
Hh55U0VCcggEtDY30X8nRKkz4cW0DRGpQNUUnjWF9iEL/leZXYtLVOCK/5AAxgmSRtV/cFlrrvsy
imtxrwAc/OgO8bvXNz2zOS3RjyGiSA9Zs2cEqBR9MwJ3zyrUNB1tenRmPicQYuWjDuaibTbHO1gq
kDqNeHHOjLSym4QlJCb5CZpwd5Yr61IcuFs2R2p7bc9zhvPrwbTuwMgO3surl6CwmKClbyeK1P63
GtPhH/uchuuv2Xn2H3QYoq9nCI0HcwnHNmqO5Ww02jJu1+Kd6fIhOPBpcdQjdkwLrft4D/ukz7zl
i/X3kScDgTTK+8ig0nzESexF9/4z5RrL+zL3Lp7oUo6CaXa1svxH0/jW7qrbwtp0MV0xNb4HdK/p
uoXFmoYio40dxDj9KYK7/4JIMKvDoRuF9SxSRzlZjPGvDqAqEhAQmYNqe7C/smqWuSlr1aNuvFmT
agzSMjY9qiXy95bQnM8NDkMlW7ZjWKNPRecN2k1Q1JDb3Lu0Acp5LUF7IZhJ80JGDMw5zHbAHIpq
wQxOLOhuu+TwsqctCcvI9Q8vLvXf6Ag+hzjogHit/CJBdByVQ+IMaBFn1qmsQypkDqdGsKez4RbA
8rIDs1mD9FBZufr5zBAH9rgfbBiDUOOunt6xbOX41bxtqcZD+SjcfQlv9/eJ3n5TedwElYX4Fk+A
4k6e1ZGZuKxi4YWy+NUpGvZNcN90dZa+kcJn7kOrwDnqQdAkmQ9Ti0L1v0c601pGEeIFDjkUUIJk
Zp+b1QVWUZPGvs29Q+uta5FfpjqkgSgCUCBJLTHvw4HmVzZ1El2MVNvAYqKjLh/u5wob+5OIMnxh
9O5wyjOl6+1oRFu3z4Pd7kogB8D6B0s/V4LGOBUBqkij9qOYxUc93p8k/RKMXssYjZsp1FudtS66
vjPyPDkYDXXQAFiT8mG80nUjz0weSNfpqq7ae0TH1SUugMHfUvUYciqe7JBPcrw4YfX1Q1xPKmyd
Jw3BA3VMSLbq3zusU54KVuiq3QmIHhdQlWUlvJXim24MAiutIzywN1Oxcx7d5SnuMp4Xb0PA9JvT
xWFlwMSgD0X5hvRmlM5t5aefJqUw/VyE8/OWkdd+TFngqIZTjDkd9RT0rhn3z971fOyB7Vxz1dfx
UAq1Oi0b/u4zGhC0bh0MXP3qnCk6yJqoYTQUh1+l/KrNNw2+5nKCHpC7TAVY/Xn3LNKhr+34z5z8
v09Q1ovVNvoSdyAacsS5Ug23hNcXJtecx+kVTbGsYBCkONzHc5jI/iaGvXrna3DINUKzsgEbeyaB
w3dZXJqHhDnjNrnAxc0Csq+OH30+AviCEbUlg6lRwbUvIOdAJUmOXxlU+6BlzaTavLz+vyvioyVM
GDRRC237ucPq2OcOws4mONScUTJoCbO3oBmsNb/g0ayY5V9E3HUWBl3GuxVgXe3s0a/W3NO5XIv8
huZ6s0dnOrl9XTkjwg07jqoPn6egVH5EuyqHS8Rdms8AkSVyfOvE0/LfPQqapNW4Pc8evEyI0isy
N4TwVWc7dHuAI6LsK7quQWUeCcrxd4VIC6A71kjxEpGW0Nwd8YPIjRJT4a8FJ18fb50qbJRiTe83
PSTmgXdcr8C+giyBhY7BWyGRw4kXaKcIQ5jEZEG5EkbCBGEahnYUUFb0Lvnm6v2dlvTyrRDiRFrX
yGbfJJA6ExniQWUJXC7f4Uz+UjjZhlzowunJDSZmxOaxlrA2Opzol6I9I9r7nT2GfP02sFCAx0Xi
1lu9tTe6ImySTz1WjK5FCZnNr77BK6TyTV68TfgNPVJ3/EAsqtudgQl1znLHHulbVPPHGRxNGJ/J
tmJfjBsP5TH7ldfMFgs5PGFCWZlF4uNkDcGL7ec15fM+FjMuYEYIqsqI7/BKD2qgfomGYfI9Tvmk
HjkUClln3t1wDqLcPmCyyhPyCfcFrLpq6tw+7OXt7dl61MR4lhoGgsCdIwWMjwCNE6GfpUT81VIb
U6zGormv/n9Y75CbchUZO2CgX2Lqm8M45GxEx7KKU3D5AaDm56jzKNU/lvwvZ3LWRgr5l6HwXtNC
JrMlTaf2D1hLiMxcaMEzxOnYy8GlKlGQNEaurR/h3Y4Wb4bkctT/Ey71MTX+6ZJx5LBRS/G3EEGx
U60Xs3FGGr3ZWlxcn51bEFC/PhjZCI0WcGw1eX0FDCq7+Gzm1Xfyr4MIE720BM7Dw0mkPcXdSdvL
+iI8rvMaMCdbZNwcR6lrJfUYQ8w9++QjbBw7l6sX5Z65mMppEnFrkD1phq/ApOgMC1FkwN1eSe8y
KOGa6Y+Z9jaKWo6+X54gr8kEVMHMEf8W1RJI3vCJ6EN0LjbPlux1mEaJ6bWGbvd8nrzK+4ndd1d/
vZWenJFzya7myVNhntItG7NDHx7QHfn6WvRPKxtPnGH3HXdLYA2gRIOKwAV4O64M5NSpLa4sXVaO
QgHk1qnitKmpMyhkm8nmCI9Y7thZzAqVqbUBtqjENsPApfZ8So2lsY58kk2mKzJ+X80ehF4NbmS7
h/HfPJf8oO/kufepZYyczvAKb2OCXd6w0mkkB722WVoOk4h6Tbn36xkwqDy4yPiRH4/QymkGSABD
PSHI57OpStG+HeHsMkCz+oG8V/1FbEerSfCQpCPz3XgkXjSSKjuHC28CNhxVQS3LB+fimfqbs1NO
Z6TTo/2r9F/pPKDdQXc98BZP/5fmJ3tEmFsMM6kPHz2r7eLvhSnzhCPFKbHfzqiFmMd65cpl9jKy
XHe3LDpHmKmgFoOtYJhQJeoD0k/YNAd8fXwV+TOV2wOXfGTS9sJw4hUI+T/jJRgckSXDclysw3JN
p1Uqadjurwq6zKksxyRtQB6s9Lripb080XLHI8AnawUPbxngrPoGN+XK069YRd07xYWmGcMstjpd
BkDwR2Iu5qMfVRuFzFP7jf+hjieEzzwnNDSd2QIskVYX3p38UgCJnECuk6BOmEhNrrctk6pjRytt
p+EEHosxo/r/NLvz60Zue6vXAv5XEsP/tlamrGmaPi/5RSsa7/+m2RYHY6ynOPV0XvzVMsxlcZCe
DyYAEU/ESznt6IR9Dtqnz2hvB0qZLwOjrmJdqmU01Zkgf/pfb879kmimSNxAGF06kWpH9WSpnlwq
ctS1nlyYFeEXhhSfM156QHBCUANIAEHm9j7piCG7llIEK4C7EdeEPUMVDBRr+2aVuHckZFjgYI/c
SCFNJ9Ejyhbfm/QM9tmMvIZuYgFX7tdBQZGSja2SSDURYXbdAwCLGt1PN+/Xt4z75/ni6D/pReyj
Y3opl7xlMuCJDOiYXLBoSexnJFSzTHUW6FTRslJyrOWP7JFhknHypr32xkI+20w0lndPMqYSUNBm
ft4dGf/iwMXdurCSFTs/WW2rKQ1ryXPQcm4U4VFWa+ItGJcZrD4qs/z/lU2/NosuemyqJQ3QQYnQ
KUK2PsQhKASRFYwkS0KwKRL4J8gbpldksiIeXmZn/7i8P+zEluakAeDE0i6qS940bSwj6yMtTdIM
5TFi1G7Jkeh1xmORdGj+Q9Ivbr4/21FJzRlTiA/tstKLG2CJVD8gpQewuqbQWkC1jLTGlLC4yKOX
YQ6rTLk0p4o0g4UQP46pxPwZcBYYCY0ZyXv/lRmr6TEWK+EnST1GtifKXKDpkdTAtOFyPEsD3sgm
ML6BIImVRycwCDuEQ8Z34RJbxMGiFB+7VbEHIonhUNuTVuruf2PMmqxOduYfoTUbN6AR2MYP1+XU
tcffuIl3w82dS9UQau4lUBO5naJ5azijhtA/bNDdobi3YQEl98szmZlzVB30/EZC6wrcflHe9jlo
Avm+5UYZwBP1M/5L9EhPkWlqx814LNKSxsG721wYJMV/twXmBoGAkwEZ0XNuxLvf6dOHjoqJplhJ
Ew9ZCp7xjMyU5eAfkVAw2+IvRroajKzXIYu5095Imgmixe+ne4lT2vricLTiu0AIym6lK+8x+GPJ
SoagW3u57qWqWcIT5T/DiyXLNOd/jQBEw4FBWsv10wYbjmlRQCueDn1B6mxQhWqGCRrIH4dWC99O
DamN6snmWUhkWW6bMEl5MV/8PtFymtVqqGbyYTeUQ5noWC1KlKMB2fn4LSmjq/dmn4uddm7TSAH0
SsXolAb43tYVC8eY8qKQAEHM7U6ZTtEwVfy+WceNzBs5nPYUOw2NLTZy1hsg8Cqax8YOLn0us2Q/
e5lpKfj68d3MXXuFZjfiJXIWonq7UBOkHCgqK3TBUzrWZ0mex4s6oyFrzSCX9czlZgMWdKUmeADM
w/MDMZHiD9d+CaXk7kahjwhzc/hvVIaLLP75v6Sn4YGCXojvfVk7aK5y3kT1CuDYj8Z+6FbelVYy
xBy8bP7YHG0Mu3XMiatuxksYm/1HnV4RpipDezPKhTMpPA3hJq2SAqLQJodnbDnSn5YcEitA6exf
lz6VzeAQ1w5m7XUJpS4hVZY10eLhkziT2kBzeVD91rLwXZsKT8aGCSuY/olw5cb7ogqxxgu2TJRv
GSa63B36jd7iBh0lSlekEil/Wu4a3x4jf9i4yyzraklIxoLHWWWH/n7QRalXfzRavytfUJTGZIna
RWehYMMyI/o+IqQnPFDo6+WXl1d5lvThq1Wo5d72Nxr7RSO3xpTmD6Vy42orhaypLOxUwBujlKmC
Zt1V0in2aWSa3YnDPDQDFxStfPFjbG5Y1RYfmLRTuyzWWofb9tH0efYbKl4wTQ818dYHFjf2KI4q
jOWNxzMirw2LYpPyPazE1Eyd3oSf1X/SRyEqvDxCGRqrfpD+1eaiTvVauzUsk7npEYGD2RRThgC/
GiQNmUCGJSG70Me9c+BFBb5VGqpoTlOOjVpGD/JbUe/h2AslByMB4CUmcT57TWrVkp8Z9/idBQQ0
BLOczQp/Q9TEqLVZ9OxzE3no6Uu0BKaWETOGERhm9NNCC6D8n+1PFDmNQMAgylk7GEH6FrNCFRWM
/mr8nDAPwjVXq5yoA/yfk0L4+4uUZkJzt7pfmOv1Deh7bNLspFt8kkAccKQQlDWvYSq46r2ndgc+
uGGKWIv5vyoUCV24AqKbys2qQyXIWwbtBJ0irPlEJbCWsFBPVxp4gxcYUDvTvi3dn2jqIOR6B4jY
aDgUcf4gYeAHuU1u1U07taCVwf8BELue+aEQ+XViUlWOrOwy5K9UuoZi/OlTZFxXcH6ZDlhjPIz4
qg0UnzB0U4WwyW2a1UEdl4iVpG5Wz7c9V2PSfUsdO7yVx6SVzqySDl6qrNTY2sI/F3kd6HFRtqNF
0mkbwyA2TFA9AEdea9HBKixc3qKenTVuXDR9VndGv3J7QJqbS/wCeHUuOLhBg+e8WrfSbZPuw/+V
SpwXYmV8+rASbTOLV/3SXtbJNUjqrRumFOpHhrFY245+YtRFfiw7QMwijZHajqqfSRXMKI8F7rV2
ElnmKQUGzUxX7cybEWlVX+wBxTUMk91h8bEA/8wH9mjHXiiYyh2xK0TmLHI7I5QCzyK7lujZyfXJ
NOA5OL/Xp9uvVhdQfSAQgK8InYeoIdHvFk62cR8N8OyVKDUDR4lCSo3H1p4hBL4ZsBvCON0JDIwb
/OlnCnKNlElFEP47daUG5rV1meP7ZxCJBe7sCdqn2F+CNu2nL3USr9kHqTW+mcGIYXSq24cJfpUh
ZRRXiD2p6atvIpAr3XRDZym1MqeiG6FgD4PW+FlwPS/PmDtEt4XIVikyfeuiUbMZlYQaAMEK9fTG
ZoDPXi0gQObw1DSQIx4RzzgUMnDYP/ypE3ZWi3vWrvUIcJl7GlFUwMfi32wNB49Q4TfEwTx5PNaZ
xk2mE8yirgwBLlKN+fbHLfC0TE+B5f4+MGaGRCk/eKnyg7F/PGzYOPAdKM1w+8ODTeo4GFu4ssQw
bwhUFaTmFpJVBVSTsUqsjmh0fTKOfsd4n83B3cPk3vlNv441zQeXyUSXT0xr/ki6lWAFoQaz03F4
XeGUrodpgZxvgz4NTP0A2/HnNFTpsspmHlfv1ZJw5pFB3rpOaZ00V41f0CEgjcMd2oD/3Y7Ktv/5
8cpYvYPl9rafnBjmI2fpxACj9LLUcrL6HWkfRqzNon+/wk4r+5DDyaTYunn6/lXyhZr7mzBZXng4
H+JGek7bW3eT7+XWTMtgnLsN639jZnEJJOvphJTQ1qKituj1G5j4Wv3YD1d2CuX+gffF84WZXJeh
m5eCU5sSgPeeryE7kS48t2X7suI692DrQMuR8BajrQfaqFA9giFo/llA7N427UMf44ZZ12/cmSPj
HM2B9f7jqSJ6E6hDDcLE5c7tKOzF2YRI+NF5gMvWVnEZvITIXJq+CTpaL+N+UcRXr4bi2MBc/xOf
xGoven1P5AU3osOuDtcPhTCjtvaVUGMOqgZLEKRUYimLBwemCci2QNqR4gflkP4WWaVG3suOaE/Q
j0TsY3ZZNdiY2Esc9dWz1b1q5p8aQSDkdDU7yEPi6e0rrQiiBnGGWdIaq1pjP4UvhlAOJckPYg6T
2hi7IPgW0b7KuixSPpxAu4JjDfJLK3rIdWhy9+4dUaPb7cDhZnPXy4QSTokdiLnYxhzIXElE2q6s
b3j9+jypMWMw918z/AnD/Hetu7QdeBCb92gm9/m0kFIptP33oNF9TqprugwLrkav00g5Yutt0EX9
psx/VQWhxa17D0IU6+J5mZUOBAgzo/XjmmxnNsfXNEDLoI9/i8qTPfKmzh+Fk6pdSJn8NyjRFy6v
UIjuq/ohtClURkMPjITIuqApF29BCVAe9zTewJnBv/tFvvpcKfqqlcum/KRXpprMFaEGUxrWl7BO
bugMmcjcqLTl98a4pJGW+vCp47Slb8EpVr2iuoZwbOdWTzyIMFv5CwBIydmH/Zp18wM3XoxprIkw
IwAp9AUBtfWeJcRLYazjvDpGVUhC3TCJOh1VB+crRLkTfX4snl3yAHqT4NeTOihsMT74BsygWySN
c8jUiOlWfzUJRcv2FgJJ3JdPEVnDPEGV83guuMZtQQK8O/KrWmHEqRn6hMuYZYisJhcngie3d3FK
yiuc10kJmGrvbbdyhPyXsZj+cKuO7sNUTn6q0SAks9hhYDeGQn9xJUUqit2v7CMVmSb7wAvCvnCt
YwDWk5J0EH2iC4pWqVwY4EDE3iOpfY4yqrXYuhuqZwyPWB3l4u4gekF1F2J6Jd0q5sK6nUF+OJLq
FdceN8C66S8O5Cwpqt7Q7c68i8oPfByQ3c3LJM+dlJE4V5bZmx+LYsGTYoL1YXLEPSwU2ydO0HUj
m51rqsWfWcLky336dyVV7YyGdsb2Wtg87SCERR/ertOi9I4j/fJy9Y5pCMJt8V+zdlazRAhCkC1e
XtvH0A3NrwrYasTs68dbOQw2Q0FK6O2+ZNywfPxsVgC3htteJRgDDBfs+faT1R2f4dm265XxV8Bj
HOGTLaIruUGxPyWS1n2yIA316z4xILGJxtaux4PndjGzOJSrjrU5jZXniuxTUQ/lKveqXCEe8x1o
RE88OwwPvUIvS+ZGEuzEMqf6dmoShF9yTjWBkWXG6Er/ryql89BKNJIqvXK5HyIMx7z+uScmIPek
kwwma4lkQtY+4uCJowg0Q0j1pMp4mdWgpb4ou/xuqXO47ABvMReX4JX5Zhbn3lev2vHzY+9pPcNY
KVKRr/B7ptmbzXMiBOQuumthPcS0Jd99cIid5cRCJE9PBU4HUFDiyv/z2fFTlgbVhlUxAfm2xj7W
jW6ENwqah38dKyc7m+xxVke6/rvupATdsq/mPSHd2sLXw8dpS8uMJkBlZV91ZhYoWu3JmSSIQdYj
/ZkBrEY9PjGv39KMUJZrwBpWO+83Qn6F1HQbpIUAtEhOQL/FbPBY0wLSknOqoBl5P4tGZXMIMkwd
x0b86qFmvBVqJ5/5eFjU47C1rRbTI6D8LqWk6LRl+MVRSBoc5dGVjDBskufmP8hmYSVDDdHJNDHG
arXi30+TXVpaD41NQHi+OwwvQG9i/u5z18fu1k/XOsJW/bXmU01PKgQR7dk9+yo8J/WNcHcM5O6p
oknMXdlljhS+Ia37PkqFRMVgKnUCHswDBh1DydsifFa5gXvpC7itflcG6i5s+ZzMpjS78FzPEWVg
D4utfwUR8NvArhW0
`protect end_protected
