`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TuTIgzswyfO1qFkkny/5zxOyAlx484Mbnf+ezNXCBatf/rY7MmjRpBC9C//G6svZHgv7O3ksv8b7
ws3dvePPZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nbe3BKnfOTiCQ32lYnjYz+CHLh5rGEsPGuwZaWw7GgleEIs7VKH/Rmvul8jT++TJ9xXQ2DLKYpx5
qeazr+WkkwjQu39PHiRPOBpMkGkDADClyAiH/zRFz6sd4lEYu7Q5sTuOo/Up4JU8Dt+UrwwVdK4Q
X1ZQAbIHpFi0LEpxYS0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YFdHTGDSQh/v4Vg+WZmCdlA9Ir5DRTjyT2fS/to+4G8fz7XxplMWuaxLaqGho4+uKXj5QZatE41V
9kZcIFml117itXp4ZBByxaQ8lPDp+FqrFFUFZtxY+uhnuxGdgZsoirnu4IXcC5mq/iIn8V4mK+2B
sxlMdcqZCHBRJno6hsZfuu4GUUn9jHjzxLUjDpsZsEMxQyTouuKRkrQpTEMhEdoDwN6BAgdsmPaS
f0DwQDYtlOBXJjQItd0yDs5vEwNyW56n1jzzBJ0UVmk778KVUdHVGyVrxBrVs1l+TIq4aoCSJPWe
uDXKmB2u/jdNlEDQ5LDy0hfrEPGNR9N+X5AWBQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JCM38LfvuAakigUxdj6+eDxvvzGJu/R4HrsQuL7CyEj3U/n8Z6IHIkTOlbNqV5QEhtz8dEjF429G
A1qxL5Schwh0Dcd5aOjzrUOLc8Lg2Xt+mknzqi3GE0sxz1XBu0avjtDuOgAszdl4lzGyzntncUqT
smHo+8GnPGh2xVQn6uI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tMd7bEBVIZ2I+7kShBYOfQWu3r5kSFQzZkhKAMMrVUYKW2uGnyEXwIq1mdyZxqQPOYHXh13edCTr
7EmAUb3vHwMaW5inul8Up0+K0iARlSdJ2mIi0Ep4pq8ftpjTyeYtCw+X8tbigCoAw+nK86wKlmK0
mhS/0GNdhXqyHhPLQcxd9y21fDA9QGdvcRMPq1wWBSJW5YgEWXZS7q7owRIwOzYJCP9a+7q9KQJM
5rdrefm4VmBCWzJukdwhYLZ+Mqq2UeNvDY1hOyjmrMOsKYkG0MOufeT7d3pRKp2qhLUzPRRMlmkA
BkeBX8vI5wJemhwP0oSx0UF2l5KRoGMatsJfig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6240)
`protect data_block
u7an3AF13MqRlrXan/6lB1tM4AasUjS2t3HiOgi73PkvLmEt19WhJFmlyKnpKy/KSErJcNP3QH4b
beHCn81BHmDFrPHU5AZ4OfV7wiejKSNi9XEO0Ojgbut0Xi6F6v6iTUlyRdTEdW6tIOZyxQSeKs19
/RnDoaYmfLWRMdIATGnbcp9ARI/YVwKOR66xd0hh/utyZY9T57lBKMtdKZ2nGT2uQ4Hv6j6jqdMo
9GNdn1iikd6+/8x8JL8sP/76ra8H+R026EFdyhZFclR1FhdfSSUJxlhO8L4rKB9IbxvWCtoA4sXO
lq9LdQhEaHxnYSJlTainSTsZZ5v4crPQ1h4viKVnH1DX0E++ZVFrTteHHWokA6Jf4KkTlLhKhHue
1NdOE9B2yDQZOSqly7Y+FS3Si2vdWqG6CY7dzdq2lbYUfFhokB6Qp9UwxfDMEM8MgbuhOJ+9qtYt
gpGalomzwVPh5O8XOuxmNYYDhZw3bmVs1iaRrC0w2xR/Rnl2obDzTW3At7C1M45NFbtL7RgtI1AJ
khfQV29K3DjSOHVRCf2yiG3tUJ/g8JObDlt7Ghy9cRJkrW3AZqaBPReyBe0Ojv6A3D1y8g0iBrQ9
ayr6Fw18RyhRMiImcb+BiF07rhOH9nRGAB3QipRPp4w/6BxSwW1puc99YsRxbovqHetw14OnC4rz
URppXGLDUknqGWwg/4QVv6CvvCnDSthCicUnrRiFDmvOMtxUxr/zKcoI1Wb2rsg7b19nsUa15QCh
cv+XFs8uaM6107j6KrEuIVYGrGivTRV7s4z9KACw+jxI+Z5aKqPaJlAKw5ETx1DD7x7MNSUMzldl
oT6zWdYVZYDcPL8UX+JxAhebRDvkc74oBhv35j4PBZ3gAnMJzPHXgjWahb6VomSfvqar4TXmQf3n
P4nyrhPWmQPOMoHlg/snT2EGlfNlsnOLy6Q1WpJbGzwW4uvr+KhNwzMBVCQQpv07kv/EEfushf0Q
Sn39JwzMyGfZUx2exNzXDK6g4AGhwWKUbiP5H04zqIoK1gFQrBhx0MNk3D64xG7bswefltvfXi/f
RVtkIeAsXOD5NyMGZHO6ZHI4GVnATYZCkDhItxG2LW5rfS8D07nuJuAZo6Wrz3nCW3TniNwy88MA
J8vPbzkphtGDKxc+YSSxH5ggw6TQm2vRpQn3LswxCgELNtcQ0ZnPeFEU+ercRJeBOQXJOUNPyBE5
azPrAzqFFBmd6VBVPT2xKCjOZb2/nyo1Y/1ePRn8DA7L24ZrfG4mWaELlXiEBchVW3N/ssCyDmQj
nGG91LZCz0DyMCXF95Si6LGmYlUrVAh0iUmrsJiyVYFyhECkYyQ1yvfXsYSRLFeePqobNY74gCXT
N8U9U6omGw20islsvkZxW/tqNpkhR1jwexpnAfBFX9yBGhzxaK0eN5rvuhKwEsoDpIjE7TkzORN/
ybZc6toMdYWgbteGp64JyPZC2hlr2LmlDwKEavxt/a6EznXaI/e+8/nm6QKNf8/NzHdCIO4k6vu2
iy8B++u05tkiJAMh7ISkQfu0iE9TTYmmV9sjM/OZR9rJG3hwQgbpil60fs/jDKHzuVi0w0Mn72Gd
K/ZuiRyYX0glHS83ouQCfRvgEH9W09+Qnk237RdpUBLsiPUPO8cn82kFysvZiT8h0/6MVpoUqez/
ysNaHhxBQXyKqcCgf9CjLYvyNHaL7dI6jrnKKtvuWUh40psX7bbOTyLhsL4wMbi/2Vblyc6illY6
b+kD1SWGB0xI/NJ8HEiRU/yUd5DEyzErJcbkWfZ1LMjBKwfwvZFS/kQqYUriZnyPblAH/y9w4XDq
TGhOlCMreQBLHlR5jGJkEOrMlyxCbktA/EkcKETL4x8g09eRl6PuzPWHZU1IbCpR7uCO0KFi7VFp
MJkHsfVYgj+4PsTK/iUx1Ogh0D8Tl0CLvyik/2n6xugjDbikqHZ1F5YcB1hcnmvYcvNyJ6R2Ku8q
gfaETFXXIVsJ6wqWq9UKCSu0wr2biaUsoRnW5RXjFzUcvahYiyosAHn4lIK1ofU+CLHHT9Yxk1JF
yD7z0dPgG/Bgy3e0mUQrgjkvvXdb0gqoiu/8WjjHlTSVsmj6XLV/wliGR9fJHFCwbTHoDgAMvl0/
y10Xeyo4HOUWonqmm1yDANqdiECbbde6okbCzNaRNXp7FIbbCo1ZgNgJvRYU5J/lMmv+BdXtJSNB
KkYB7nIr1uxrGvAaLPMa3vPQMZ2TvT8a1xn2gNr9QTQK19X7mllKBesTPU9Oby6FnIFEffaZH1t3
cVDUghLMHWZsmpRMo+EtNCyC6E2fKUjsqyy9lR/5nieMO9MVyoCPntQLAyLtwlOZ0+Y9xhh609Hb
d9fRaMJ0P44PYEau+jp7+/VGLI/2WKXXkfbftWsjlKbAiiUNdEPrq5p/Csc4XyvbL94lc40X+6TV
Ue/5/IGDLA+X7oRnnIWXB9JI+mxHQLOEYNLo4ob/G4zFB0l4DNxzyu4w3chgqI6WY2/62AJJ77Jb
fu2w9mgPJWQ7JH7KshIaic2UL7zf8zeR0sWJngZ2TrohlektHz5CMp9FhbjEw0oeW/+0J+/7y+LS
hxX+eU3XR1WrhoRvCaMNRZlkh8JoGe5VlRHTz9PIWgm+N5Jg4kaH+v2JIC5U1RNf9PWnu+znnOtF
X9oEBLu+1Qj3jzjqhD0Dxj9Ey391VHidkgW0NwxP6mvodvfB5bQAtaouijr7AVJ8i/3VHYZ35fmC
PWLGotRA08NX63/vaEascTdBMsQAFKWV30DGWQAu4ZZ/KWF0QwYXdtlugexPUWCaP+FR0YLJxALW
iL5AcJ+g1SKKOf9dl/9XnRxQ/BY+WZEDtgcCQ6jfMY7r27yFaTad431GFYCboAEJk9Mc7/Zaoqyn
5HKoyVDgqcAmFLmRom1CxqkWU7AmuxUielFUnDw9vSF3RnhUYRNNm/c1RLC/+VJSMUSb/Q9QnTCS
uRH/vudgnDOw/ZGas9w1wzKZ/CIalh1QxkJj5wbVi5cYnmbbt7N42cqiPQzsQ9/5Wqm+KrXH3gOC
vjn0Agn+uWHS7A4xBmgq5xtIbAOkmRfChu+ObycB0zzD3u1vwvTPREt9gAlL1Vygkv6Hd6kaG+CX
zJOG0Y31bzfPu2mI/ywR8HxGWX/o/x8YvW5yyfEH0+UJQhmOOXofFIQHoH0FvJpkkdooJ1/IS5n9
QyJm4HnU2FNvx+a+EtyKCbXJAQF5V/HKsV5Laqf1PK3JQpYYpBHxgoS96pKTNZzw47XOT4Mkuug+
eomXcW8potGA6mT8evvDiMFixFA9bqAhfDIQp3Z336AiLr8mD177zTlG3TNdI19ERzNYqPR80XDz
VxMqk6PMo8lDT/9bSn4jVa/gM+/FchL44DVkWTkE3fDlp8R/iwoxmLre+spQPWiyjlogky7Kb+DX
yzZqCH+y5E5vQG/E9AX8TSEkqJQAAUh4rnx0L3IMSCrmJEcc38PSdAKbB32n3kznDNlX/1XmuqxS
pNQw8mBX/GT14C7m+8o+ynaSj9oV4/dAJufpCa+rFvmf6wKNym4k0E5C0Co6BpDPmI3jCFFi0pWf
1hoedGnTltjAHALIbWVqWQlNuPUrgAmF7U++7pu83wzdMx+mIUgPEdAEdDGxsDTnIgJpuL/RFdWS
dLpzsMbbkjUkR80xXy4/Vjpak/H1a7RFbWriYvIv9s2iEeEiQZ3soNlEpdg6TXoF9716vJ3qIZ3l
b0Mp2+E1ZUApzyGkgOt/CszrbBD/jPRhGOnYxmj7z87Eq/1rPoA35eqKBDftEEw27Pjjpmtsiu8I
3X8uWlVC5InueROrV3B85RynwTf9cCEJzNkb022tmwh+ouXrSEF8uTnnV35j6fUDj47JUnCItU+d
LXG+udnf056ojov3Jmj7z7YJveYo6nwlTG0+/7Q2UYkWNa652RLUMlwRn/lm0gRplwCxlKrqk9eJ
THwMBmbWPsfyXPMoQ9lZAKT9UPR1og+BY2a4c/rzm21bZz8gDUae8VBa2pyKK/7eDE6iV1oW/FNe
rKDpUIkCy4tzk7R71yJxaxhzlF8yJJGqkRRlTmiIhK0Z37RcuQcJUVNOkvWM0V/zPXQk6MpitAPy
fcy1f9R89ey4jMtyyEajW+E+d6GCt78nhOMXwCOot+Z8VFI5VIdBGA8dLKptk8g1BWxbFRMKbEDW
sMoJqkVOs/gy6wZLEuM7nuVUzLnCIav9AjBYMs3PsHBDhYnVKWFb5/vPKq4rRA6iD3Of8cK+7lb+
Pk03rYQhU+rivNrBUzbA9PeLcX4rz5bfKOwqP+EYjn3vV4pj4eo+eNH9JN4L5MUEJt3X7IzjX1qr
Dwd/iEO5qzymS6cQW9WtDXfRp7C521cnLN5SrLqRgOepk9PbbBC+izjSHbQvFC91GdnvYYRLvdm5
NLpB4ivtyreGwQFKTZnzNiATBaaQO6YoJpFlPyMwqHlY+SwLXZSQrCCR5+9CgpGDmZYom72RCvYU
yyHctsNPcXrmfJpwTWTBBayWAbSnNC75c77LyDJ4eEmVv2lvLuqwCImw2R0pPl1sjoRMFogcsJQT
pEm7Azoat9UZWDI5ymSEec66n9pAzifWkCBrpGLZpH1qYTo0LNqLK4c0iDnEHLurxIjWX8aOBi8T
wSRkoH1jT35+6iwH3xH9op6X8aATbGsv7uSJWIA3UT3KE7Otmuwm7K7SjKr8TfYv2oq32RRJAqJL
D3mxYNsPvn8puwtkTRNAZS/kQ7vUUeVwGiDuvo/3tDkaGnpJlKgwZoGs36EzhO+KXttivZUoyyei
8YrVPRHZsGDdS/MQNKMMkenoyM73ETdcsBEKzwckYt82LEXCzcwqH9oD4CogvjZL9cnc1OoIqRuf
adHF8JMfNiaMwqhaWbaNw3IVeBekHd/SmE496QXEgABBtpq0F6P5pHedlBbirMPP1+CB3KfhhDxG
i1TmOWj5bw/4j/A/2QxU+83Cjsthw1eP8YrO4gZrUusuZ/8wxO/NK3UQ5kYs2hjeFZyuwXNtcCCC
St8FWyWLHB5ambTyzGFsvViaP6kIJcOa7MDEP8siWVYHZ2nfqdyIkmTzwTw4wEJ+unTcfzEdeKIa
kyEKIl8HHkmZGAnU4K2zz4i7TnNEWqsK40ID2OZkyFeg+KENoOXTjMVfGib6y2QOseAcRh6duzj4
Pjz+ckGAjZUIwG/dNGGTwQCKTbwFMBb2y5R5JrlfgVbupk/YSrfZybeWzzMstclpirxGm+cRYQnV
XGrP5I3CDZWyrk9ynrVCGNbSm22MebJ2iOeOWKtjbGMf4DO4Ck7tVWoQg3khA2du+qqYrKFvQmTN
fj1/U9w65+ONVeg5q2TerDxmrMiawqwMAEqctlkJQpiv8T7KaVbAKEoQe1me7eqfcmDIcCZtldiV
GL4GIi3kqTrUCqw4F7YRs83FFc5rly/CbK+0fEfh/3yqkWPOdvOKdJwKvBcJeUHr/ehWEr72roZh
hTjm00BSRrvotGlRXJKgNsvCpBBGtDj4dKLVcF3bUEAGrOLFeY6EHrwg5qMwCwQa+CMsi6vIm/KW
HG7QRVRZs2cW6Zk+6OQXBexqnNeVBghD1ix6Mgzn91yLvx9FWj5RcctsejYa4MRnMyurLUSW6bvQ
MzqW7iFD0wQiLZkPgvLWwukXGrhYP9TI88QTTBgiUTF2eOUn1VYZSQ76CXMJ2UTdjxqMVx+wWKQh
Gr4szFDxD4PUIHD44PGVsQx2+pPz0cwuEqliGz+WXlr92wWoO2k2zEqfbdWChYpHMnCyfaB8yXxH
FrRQB+6u32uHcFnEUe25RaWEjsm8y2d3QgPj3tB95fwYmEe/N1IPp5cLSlPQq4UOVUEbGI2OJYqz
2dIzye+t0cUD3vGSU7Ln3HHcqJQnORJwkUJW43PrNxCpzUFnpDn4naA9M2nhlfyw9OqjrvZWztro
bES19NEmPrbcx8O4BZzcegV1C2qKtEW6baVLpxF5kGK+pVRfT4b5H7I3+SITcT3H9mMnDuxVbTjL
PdJz2lmtcJRIf5Ju1CqoDWJM1tfTNxFmKMgr+Do9t8MWvKZ5U4eZwd0Jyo7+2YX6XuYKYIXBpzIJ
78S7MWK9FR0a6JToU5Hvzdh1TMoIfzWiDcEyM7QY1fgTdL4UfyVcyt2MPfHvzYHCrqpsxbA7XfCT
4KfmJgtT5XdG/Y8xBAoT2WmVIiTjExNSPXDtZ4j19cg4xaCNTVEX5DPBija6O+8tbS4rfVtLyTdj
xwvdbnmR1OiRW6g3mSSH+xOLoy2eyUi08s12x8VX2e5hYIu1eN1K/DExxXw0bJ4h6n/E9gwiiUC1
71ykqM31xMHq4Qkp4qTplvfi3VUHTsa5ATjE78iQUdA2j+rN7i8v35BP2+847Fd7B+I8zs6fAVMB
XIV82Hju32SJLd9sbzaC7cV+qNGnZmkMTpRwTIPjm08cebJae/EsS9ywuySnItZKofRq2PgI65Ej
OBPeMhSivL5GzR3zdp1/G4IyYdvoiM6poooFAsq3yiWgcR4MtTEoow5siaqE9fjJHFOuC2C9bwq4
3lxKaCEA27YIHUW/sE8bCRkhdwWsWWgEJgZHwvUWe1AbQlGnJ/9Dctb4LjZmY/kgrYcxzM1FSyPy
iLGMgmqIDe59aifqhRKN1kUoldEObbcCzKB7s8QYhtvDfT/HgD9o4hjDwKfw9Vb/Yir6pt/xGPC6
12s9nEOKUZg9YTAqmn8pCDEwbXmQDTesATq9986pEYLSWbnFv4Xg1jH4DCr95khAU+I2wpLtlJe3
F0zYWJ93nFLdTWFRAhpE2GZzJmTHRHguRTaFqH1pXywG1u+v+7R6Cz9OIueHIOVZgtJcagb1jKES
FLLgLx0fRuViV2fv7QtcHiQxk9sfQFnJql+3aA6FkSXwYZ9LsH0D55i3t4srAT1jXp8DRitePghU
PXNrQuCdUcyjcreUf842g0XRNA52QFxl2j072T+DtK1CTVNkwvVjfdfXeBkz4xFaBs7LsxWr4MyV
4OjXht7xX7FxOFD59FGs7ueclXbK5FL6rGcVa6Qsb9JL5BzFacMZliJ643K86pUUw/I5RGesySdX
kkGia+zinpCZrzO1ZEe3CzfAYEJW55jPX+9XEXvu6U8d/FYN7JIzH8LR+NOT/dQjPzYpfb0Mo/WU
rTesXqNseC/2nhoehrSOio2ABu8VjV4FaDuo4hQccwepllmhS5o40jisx0ncdaUpPpeSrdyEDW7y
6I2rCRPu37KCW+DFDze0iqP/yciI7OrtQ4mqRtMf5+r18nsN0qq9f2AeDNsv+k4HGIyfhtSZ2i1a
aQVmVurs6w29CAP/N1GVyTleUhODHK2cZE8XjptmcutK2n+w1t+spXetKjgfuhYoFuyyfyhUbPD3
w8VJhtH3tF5f/TRbla1+YTW6afqezIDUMtyJavUupl7bf4NOwoxkoSl9BHQ2t8dKRgjeY9D2p/X3
T+HNM6S1K9YzuwCUjfdwrjUVnhwQ60Ir/yFRkt/uPRWSYTOGvOKlRWj/20v2UXvDWhyKDeTzEz2W
Ae7CITGiBihUCsfAdb0X0fE8fWMYf4oUbDT6Hw9GMEYlygh4PtmBEITVhYE4RHToyrFVjs7nESB5
KwRFclfWoiYxKumzYmveDEpOkR7mrvg3AQS7ZuUalg6Zfj6APNNchlwohcjcGLFwdJzV6cWgS3qV
iDFv+6awbROZDVfq1LUzo5NlXa6Fk3T0fXSWe9BPKDtZWSPTEblo6HZ1l0GHPUK+KLnEnLOKPskk
Zow1KFoPfbPHs4hZ2Ix/x2W0KgqIA6yzcupTCk+yldMwEgTk4ebskjlaaFv8tXd/k3xZKAM3JfNT
mFNj86JWJ9N470WofmjSc0uEKrXi3cSETZKdVWhuO12i0/8r0vQoy47NMjctHg98A/1Y++EXcgF/
dE5tltf9rx5Xb9LS9RpvIvPpzjJUJRakTU/HP+p6y1ndwYhtHOm2q7rVp52IpLUdAgD45VV1jkcg
Pj8r2ubjFtu6RW8hBsbNF8xvtum7e3elrAHj18i2+1/2k2GJNZ8fvrj/x91VWHsfcQPsa/BaCK0T
GNSxWl6I3Es7XXo2HUGu3RYMFqQpmOq+JcfiDJmZc6fnx20NpqBnptgXZMLpbvPpi/WZGOaiW8Ww
A3bB/ntSoQQV1faVq7g7VFxC5yP1vRJTKrZClO9HvfiaiDIjua62nuUxQa8cw9lcYZBGF+4Q2cET
9Qo4TNh/Vhcpplc161Bz+0ug382Qj1MqYHFbzMnJJO6lTmlj1SGLK5PPnF49YtlNDMpSVvxTcNOE
jiADntshDGEBVJPqh5mn23mAOPKKXeu+vobm
`protect end_protected
