`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p9mk9oDYGr8pmZkWXbY2TLDcNbG5E8gje77Jb79LHblLzT6z9srp4YogxjZP3AdpB91kWPxyMOW6
yZ8yldjKJQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mVXEkppMj6g1IXjCy7VbBKs+xRMg53vy4CptQMu5kxBNHV1PdY2Z6vTMCczc46movp6tA+re7V/F
HsTTtWCV8ZPfOv3mcdhM4UeGfFJKyzETnvTW+7FBhhQEC7rVDuHV/zQIpFu2woT92yIODVDJv0OJ
d7TknpWbiizNGWwk/hI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kaEPvPGfpEJgQQGZTZXbF/2CvE4Ypzvh7RT2RT4lopARsSjuV2b5tLmuzYSb85Q5AFDGlfRWDwtx
F2YZzMpA5KuWPN8p6nQWyhLNm/SzroKHii7qBz7lYa3mPULaNNzH3dQ4LQE55pFWYPOfv3yGdzz+
x0MEF1ydRO95dewin0KqN+iIoWFhfzxKJvwhtWiiI/X05UUfC8+LXpcJqGLxKw605Jlb+NeKbbhq
fYieug+3ebVwrZawhJ1LjKOdIJ8rUBrE5RUDvZKfy1WLh7meweDSbRCQB5rPDK3OcggQilKZ2mNq
8WI66wOyhQxGZBLF65BiKY2T7DqYxJCp5hGwRQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CVvJhNJw6EHSDIQ731Kbkfkwh9Wl9VKmiOV38T/SVAU+kI3c+cxqP00ao5AoKfnBVtld7H9d2J6J
kXhNjYdDnAvSRM/7oTsMkgQ3b7EgkwQVLR7bm4uQPlxcIXIdQ0tZoHzgZNTJUL7DL73vJLbed2E/
KzI+61P+AYGjXhbYkqY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ga5Bitt3CebGZAmuyISY0yRlSG9x1Tj+suj5BLHTSTSYidEbK8uW4qCTr6BxF0yV4Xp11LL0s44p
pTF4j1DpdFDEchCdBhPTnweZZpfsgl1tF2onzxM6huOLdb8WUzx98iaDFlYXkwOae5tqfbg/QqYr
LyzTmB6gN+UHIqqd0Nvja/wQ+C8qsyVXUotU7XSAyQnl09HX5VboIooc80WNwl7i2epmVdrXOo1U
vnq8TH8TcTYxW0QC7SWveJRCbce/nT+MzP+z7RYjxYN8q+AXvkoPoJzcA3kTVwwvXpW3tNSYC/EL
DULswVBWDYJoUSH86zvW8e9kh4GPJv6rviHyhg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32656)
`protect data_block
GFUOlaXsp9nvniuf9Yj+35P3XFkM33Rly/Cql6L+SVOFmDHwBnnl311fReTRdQswrOQzkIK9mLV3
Y+dA2qHWprdNKpYEA/FKxgvP9cBaoJrnWYNV9lVLg0aeJ5CMyiLrZ8uLViaNWnQcGAEK1EVOh8UL
zIePotyeAlUUm4fx4kAukivMG1+ioQAfnSS7NCTp9WoreSpneaw0J2BtIBwDvzO90Km6jK4nCxmL
y6xUpkGHEkXeJVC9VJ4GfBtb3XU5LUPMW6BWuNVnTDodSW85M1IVYLcvA47nJsdjT74DatyIgYUs
9zipUpHjbhfo1guYIveV6AOOwzclevEJzodFZNIs6MDOl7Ue1k63UM6tOBgRCSAVpdTtX43KSdyi
W8gSSE/xRO2zd6CEtdTMUECMgz+FM0B8rdhfvw1+PFgul8ga9w47Mlr58ZFW6w3gnvpHAXW1yzwo
ZWlth4GrpB65EaNMZGfnnMeFy00Qa+ShgUUX0ogN1bQoXO+NyAmZbFFniUxaCvsyhRILviiQPiUM
z9joSRDSoKam7aQ9M99HubxmB/uQcJHmoCEmfkeyXp699SJwCFc5BlI4cLWYSTmfbDOmGPqYAsGf
Y11t8WlliSLcAjqgX9O7Az7cJvYB0B6F/fjcIl0Z4Qy8/c+9y9NSpts14y+eecL3o7CsTFGYCxts
mcfvGzAD4jaRf3eE7U62zUK1740KMj8i1V+dUZ+H9pdT2BOhyQOWt30MzHy/bt1Hm74dX5t/TkQK
OyB6pSWgm/eVnEz+sARa2+v04N2rJC5tA0HXAyR4AohGrMuxgbzhVutpRXQ0+dT7+puOzOnglslc
6GSUcdugLQRCDdC8vaeLrPZdyI6FFtxWl0V5XkM9sAVNDWc7rwo5goLkzYqMwdGfXwnmlDOD/qhg
xQ59aZRzFo1TUwUktuFrnMqJpiYjES00iA8Cs4o928AIbanp39AgHKzL5g5CWLiDax+O0A0avJtm
GDB1kQnIbMHXOKmoIxZZ/RkehaDc6r3UtRYqREaJId46EcNdYFHXUAnJATvu0utFCOcMPs2Bivo3
fTJrFGJboYO987BWLtP4TOQzrzqLQ3cghfIWGZuAAONScAf/4CqwqrC1PxzEPfNxgWLnoCvO1cAm
4v8mkhe6yEC54/HDXzbJIRAVexllKZnjw5FYIgnyzgkGpZv3pTQ8cP+BNMpwL+pre52bX7ZfHYFz
Z/v3axxsmtz2XzyNPpHKB8n+yFlaYXt7yLwQLkdOs6xxFSL5bFf9VIlUullom31Lib5XsWh5bd5m
VJuUKcG2wLmgcrlVtA0qACulzxVbgznOq3wKISC3nGZy7q4Y1CqKEVUuXvVdJQM4bdlAqUzKOnvF
Z2llXnGXMHdNpJnBPYNzd/vdunDO21Zm4aghBDU1ZotyfIKNtiWvyyctK4cxUcJ6BipqhxtmjZAz
+pOV1SBbqnBMr4WdvNmon242BUAMsiBhu/otZNFoydHK38NqIlAbXYS9d10/D2x/Cn9XnXEKLK4N
hNtEEPDnCOg10GHtVARfC3toVhbWL3fK7jos7yBSsQxtGVzYZqBXvf8bd93J0eWP8eyHYpYeB24Z
JUzjNn5s1C7uBNKYcw3OOGUI6iHLC95nJuaSljThX+O4j+HlwRUdpOCNgX2pws9WVa23bVvFFd/F
NUwHsacvXufCrBQnFvn9082Y/2nCLZ/wST1gE7blYRsHouXCsHD+Ca+QksQcOl3XQ7PQRYeSM1do
TjMAou110MAB3/b2SyIOb9Ue9/qDK4CCUZ7VCxxlfXKlT/ubgVHNJbG9rV+TyHntRFdZjt5IXYqi
XzP7iq936Uc+LXXvZbOj2Tw4SK9gU895jH4b3BOwIyhXqrQpQjrAVTJuTuDZb7Z8mHDIhVtN/p+k
5RvZ9iFnh689QcqtGxMD9EHcAv+jkvE4fs3aChn9D8Qstg5dhXT5++NoKYNpEdiPYNYJXKPo2kU/
1NkgyB1Alp+6af9pSiQF/cCpOF0YrAWGZoY+GRBdAU8IR31+r6Yv7Fe6gPHA9rTvhhUdOG4WWRiM
U9nnPUfh4H37StBYotcgmCPEGaX+t+w8QZCsyi1gHKm5mt/AT3LWqhEamXTl/RAn2YitGOIi0bEK
s3RrCofyxJJQ9yDD2mzb+GEmhfq6NpjokNr32lDB9S6aErABkdqPY6KDGvgAaimH3e9lkuXHW7/5
mdTDegHSn2eTA52aCNBl99m0Dj/5CNdH7yntyvZ7vDSvoq8uM3ouzvc1KZWwjAm+oWbpmh5bZ7Jr
l9laaq7ij1rnk6BoAQJbRQ5hwwBlwi+GQr+yLtejWMG12aP5b1SdtGCFCqiGP5QxfD1irT5HqJst
WMl4UWOeti1okuC8PDkPI9mwHRsIByul8KOhAn9Bn9HiG47sr7b/9A8oY9js/SS37agXjo3Fzjig
b/R9i5J4Y38Uku4mwYUqjl/s/hNfUjOPnD4VwVFE4kEPoPTqM16rdESFfy6HCl6YiCNVo2sTQzUm
wAX3yrUrLsDU357DXZ3n6q4s7BQX472RIkkuyLHyPlj5JoWt19KCqhuSxY+SKLAJ3gzQ7Gc+3xNY
+UtvZxy/l9r35kvBExK2ZmMZTYkQIJDkB91/dRfp+HtjmH45UZo0Gv7Psi5JC5iXq5QHde6rNJvv
9Cl3E3gKlTZI346mD/dyJL44mJZ1WMLFAtCHDLRTHgY82n8vLRYvp9iLSa4XgWpnUCp+sphjdy5T
OtjC23CERotVZflihiI8rJvJMfwlEM4z/fUqy+7Ii90jKsJJEr1GjQbbA0/EzLkFQrjRxuE348ma
jqvx2vA7zKZYI1cJjrmaHEYjmy+0TdxMldLeaH15WM7sJ2Uz5om8ItqtmzMbWYt03QMPeCvWUmXv
rxFzNpTCRtDC1hpMOtkX3EX3UsEXhggiit9pycCRvnQ4HbDSQ/4ugE4GObty5kZrpYAbyo9MEhYy
L+mU2G6p92qHx9560fpesWTDTiFwrPksBy2i9KJp35q0Z2m3e4MxnV1L822Sb9o29PlIBESXPtTi
73PqX7GI9pUbJJGT4IDGg5pgkvdzJQwhnYcg4UyARnU1xiYdCaBHeSK+HPnzzor/0FNUVcshRV1Y
fmM23qJlOfaNE4XKZTby7CLYkYYEDjBzZY3tscXRr8pSwI6zW4Pk9WMr90F0z40fS9bhzSEE6Om0
hG0Q+FBEJdf0Gl5y6fXOw1F6OGyBfvfGcAm8+cVY6gjCoDXLoCo3i64sHT8jRgNbfXCclqP+Mj/g
2UOnDMOhEPdHlu4VNxtHiu/zQvYBOzJobM7Z5fIjnYB1TQ1vsNMgcFQbRvMqYkIXA3WZ/4mBMf7H
lfwRg5WlBgaWZOpDI1gLY8NlJxDtzwCQXAyBXos2x3QryjqD9N4FboB2Qz3MjPO/YlSUhtonp2CF
uaa3Sja2XFk0qjZM7MEwzBbqt7cDnJiBQMukWgRxnxOKo4oA0WXNu3nFP2d+uko8bpiuvmJUesLC
bjiwqELal6KrawqFPKLLIKipReChhx4cs2tM+4+cqHeIw8CYzqRlM8sj1Tc0n+TjtdHorDlkVZM0
1MVMOUrjO/HP2kOD/XKZ1OJajoLoWens7tG89ojmqQW2KtOIXS7h58vYTP/iU9wltq9Skc2xlq3L
Byi1P3j50rjnU6/zUHJwiGNvzzFkg7nYkju55rd+JTKkBu5myRg+T8VOTtu9i3K7+PYmfuQBfqYU
7pGjQ9+rn98G+o3IEsgPv3z/lXf+S8npKA4NXWdAZwAHhSyaHZL4mNlJsxa0qCVvLhRlxlhH3QPu
IOvTv8LlcjyGsoKziHALm53faD4Xd0YBcXvn4cHuQ1uw8jq9nvyxc4u5PyhK3+i31+rUb+XbM/Sv
ewUi78bhNKcEFbFPt6FHYjp3G2kpcSm6HsfLDcn5mBoC+8p4d7BUMuGgJZZ/gmX/0/eOGmYGYjOx
7NNRik3UfdR/UA7ZN7ehnHi+9ld0iHUDziUhU39iEmpdF4Va0u0JW8F+M0bydAPS5+EEECuGpyjo
2JKNqXXAVkyxUXh52aeN1kAyFYTPV/Kz/ZBY3zkCBZBpTgyfYXjFZYq8iB9+drVZYwQrAaZTe8ty
RqGi+5YHC6eqmXJxhyGf/I74xSRm+FQrje20QjAsE8NJq+72xoKs8zi5X05lUJ1nMPjWNqeB9MrE
2yL6BsR2P5DbhvYudxssOVPZINBUXvsxX+KRrH+kbr9gYq5+4yE25fPKqfZ/GzquTCC17UQ7ZaC6
wKy8Go/pUZDy9EtybH67LigexrJHrDrgkgXcc0c3t8/jJ3xCvEhZrgMQra21f0J8VtK9iD8+aKra
FU5ImN4Usi+W5y8hlzuO+oq0TS8JOT3QpYZCzTGGlGJ1PR2tjkBEjegrdqH17q6TP6+zCBuhVegB
7QdKLx6m+jeup/gyBD+r570fsEX9MyHyIJulVpdz2Ltfwz6V63t/mUM9IR5OcljACsqkdqs1OLxZ
4hNBHsg/TtSeUtRoyBg0ZckTKTC7urRkGzygJV92J4T86ejueXXmy8SRCQVPm2FtIorgiUZPYNto
onmMJGOPOlIXjoqGZz6qpu/M1iGybBxUYASxVBAPbogxGq+qC4ITbkudC2wICFBW77qOYyF7G6d2
dKjvMRJU8v2HuNWKAYrtrFLJPpzCVd6yffSOv3ZzXBDQXj5briW9/vQEAAwoGgvrUb1X56ZFBLFn
K5LO099HTTUVbdgC8l8c5eZGVdZpDHUNMGi6EJYRVTqQ1SVvk1eJa8M2LGesV/xMLhliwQU+2Toz
Rz7ARCL/sja5+LTLXFA8u5BWPxZelVHE70bIfj88Ng8i6t8sQZsC9Vgjmp/VjX+lWlILYPnTiNjv
gxAld512KtZqgUHzExDG+u5cvDFJyUIUFx1CyavAzuX3rm9zU5d+5lUAVeNi7DythVQGGmZMy9Uy
RLOXO0Ka58TAoN2WufFs/ZXUkrDTUh86XchCzvLMV7tpum5G3kPclfgYTNqtPt+WriS887hX/9pJ
oz4ZErpyeNA59ysZEsszE3Gesn2w9UyxXQeVbFgp7+YV6vVBymfGdjoATMUJlPfF7ydF9HZ00fJV
f+u0DcjVh57osxTbpkFH4mpoUSn/WSPHD+XGJxmpzupdVlwfqwFKemc6XyIwczMTF6jln7/giGkz
0YRGftw/OCEfWmvtnZQ8OIhG/XUpKyokAnPa0blQoNgY2ppcoSIE6ie1JmMGAy/QEN7NN3LghGs1
zwIdDKjzJjqL6eDc/+imDlYfSn5aHqLxAVLR6HNzKExTUaK30BqZtJjRUe36hTSmmBfh4CFd5Af6
EmO9Loy+myB7ksmZIg2v4JaWD0xoJNiroFAt9i7N4PPvI3g8q0iYNWHUmmAy2lQ49FOzsTjmXl6w
RSGxChASJUr8vaUrWVabkzxdctrmIrRe057N47PLFt6GvPwHbsV5FGo9uWI1XnsFjxKTCkfDuZtp
s9RsCGQ7NywBa2/JYvO/4bN4Td/Us0xf7ihaZaCtMbFRjWS7Wt+6IjLk5DoDfed+5HaV2A8ax5jX
/WJgon3QWaCJ9aglMObF793Qx2q0pxKQ4Kl492tkrh+Lv1c20Eg72gbNNb5ciPVqcbePSco9+IEw
MVCp89rCg1ec/vdhOurSrUH7FsbOdxphOcBPyXIR+D/73D9BtZM5w3ooZlAANdI6P37vbSRQs5c1
B4a3mCA47D4setXN5h7br2XUs0nlaqu9wyDR3ZqAfwHP0kewJxTlhvtgorm7JmCxDbanI/ccDA5o
0XP28j+zURJy0g15L6Nkn1FqrMuvVlS6xqA1HDtuIxR0x2IbueGIhRaYyEZj/F5N2rL31XoesIpr
nE49CHIVX+EBwoOVoStdAyUMWxjy+cy1/PsBTAhWfeDfh4OPoRYKzsh8gZIVtiH3yU9QMLd2ujIe
PddS1dAKC75RCQYCr5tEKbcDby8afrzrzZcB12qmbhsmMFTKspQb/LHAtE21qigRl2PZF9zBa5bp
427bK9Lgi5dcq0fbwZJVYrpVX2/XNkE0U5VzG7u4xxOOozLPrYXBChOY6xgqhFyrCTB3mxnghqgo
cYw91pJ1o8lF5t2eKZl37TYLVxObYnV1sbMlG+ghQYEY+b2/gtsftczvyeI/qVdJwSVox9GpHmsH
Go6M9zkod3xPTASLx3giE/yiJls7JqEQH5PFEcDvGB+YcsxrP/VIAe2qoDQSGpqwgfJaodL0Pp52
GuUf7BkUEburuFwWSV5URnWD0DVPMwHGUeuB5YgbUsRrOrYyPVlE2EHyMqIwtUV3gQNCj9xfNIcS
fPd/VwAmHZg7i7Y19lWzWI7nqLTNzlW3QrGj6WKT6a7OMFDTb4mjGt0LNeoK0GI5M0pus1aLe5+z
Njx21lflLewsuQ+T93vxaHIjXwYD7vWRIkAUHlk6+eYDn0E3IDDIicDs+0Sv3G4OSc/4FT3JJnSu
n8JNBgGd/TDg4mClXg8Tz5ZtUWi+ievggz3kN0/JEQkflKY0PTZz1cd9XZOGkgLHyKKW5n7q65Tu
aLKSIPpYNtLOAGfrJ6FyHTOI7jy/lYdmZUW4Y54S4WpOVEXSOZXNd7l/dZlfc2VhVRh0fofRmiRK
m6j1bN/T0U0QWe1U3ARkYNUKeuHSCw5XecNlhe3KxcsGXgA5ptL40PsGLpHMWGV8xbbCb9ccfqx4
VZ73Dqq5usYtLEUKCSprRgvzfsCWk4HPUijC2BYMOTGX4AgP+DUAFTvSB8hs/qiuAtlRO/BJSNkT
0WxMFB2E8DLk8cZMvx5bXJ5zzuoQBPv9Pdv5bvkX3NqcSyQpLjRkkdYFXdDRg6wg45vRhhmblTTB
XYecDVVOOU6HHYQyS83x71ytKTdBKiNgn4ght1t9Vr9N559XnGXxxwhARabbkGoTidKHKrD30Y6l
64xsRV7KArCmff8SaHGo4oxhpFxnluPZy7EnBCaiLJsCpmMvIRjsUtPHDsh8v7iOgKB7AHrxZif0
hRCogLUru9+NaeZigDbxg+yRhfFoB0h0xi9ukc7wMvdHUBFDkf9oU8OGMsd1daPn2HXLCZ1IuQJa
SawiJc3XRPCaj0OF0AydmC8pI/eqW0ROPpDURY074TtqYUtF+GPFqofNur92/1K2BMhwzUIQ766Q
zM3QKBiyPFlLrtuXArrHlaZJDQ1GCM83Bchy8tVAZE6lsVQHvMa6h/9tUIlU9g4ZMhWsk2EGmmTJ
O3GhAUOqWArirRHw71JAj22mckaYZObVuk9L6/wWKwHDtHIhiAd1SXFwTeK4NCq2fxtWnhl1oiVG
ty0YeDcnDro4zmK0nhIq8LWGGixtb4thV53+hsZBdBiHEx6iKc8/5djk0tFoQGFLvAq1IBo55QNS
VkDYfZHt+h2hWKcvgOFzZmNvIbZF8/pLky1Yho624pak2W6Zg9lbWVyqrfhxqAxQ3kyhuHr/+XbL
ONng/eLXF4De5VigdOcLKxiwrREvC5SiQLZe+4pxkFJMItqjUVdi3z6YhyZ3RwFHC3qvPhwk1qw+
w4NMtBUwC774HUuXRfft97peLjV4clkNFEqhZloC0BpBiKLqtG/qd3/nfTvxbwit0rB6R1AC30Jg
ewu1+CJXvoTTecvDJw9YBhs5HSxUti/gsTeU6XRS3ZB0AKF8NTYL88Z2ot9O7Uwkzg8sTXU4bYAj
iDr3JcmlvTIHgWyxGApizQG7OPX5ZlcwH1yihATZ84ieNXJKvbGFcGuxSc3iH0DuqLJlK+EvJ1r5
9T+Nd3JuVSl89jb0y66+XRUKhsDT8nAuoK9RnbYa6gQeyUYt7MTBlvcrLUOaFsxmMAgtyH8pTDth
BfIYwHunDqFrgmWsfqEwfHvNr42qvwVhJFqZVr3BBl7CjTHy2bLFgvNMlJ8vqsVVlqqKJhqPYM0o
+qZ4hyMfV7cIhZOPAQzYl3HR46yVqOpYUmJAEXjDU4VdvBrhHNLZ2bhqK/K3jcFkTfl1KkAkwbpR
R6qbf2Y8T1smB3BqwS8NocdAUPHGePsHcdzfTLWRfnGzjMD++/hBi5k8ug6Yg7vLqfNeunCTU72c
LVsune+VlwI8vQGSBoHeiwqAn+gaKdgAndHGIO8oZJTEaSoXVomTP15rDcfmbJ26llTpWNL8cjVm
sEChKwgE5PyZe9fiUhbK0KIX+QWAlS2ChAgiXyo2jGvDAnNcwc9B/uZfuTQjE/wseDNPsuvukbuX
TFWqyO8debMRjJpjFQcXwa680nTw73SHfFxLtk716fNUaGSJ4Gkq4wNtoHp6bU3IJC377ws+OCd+
qQ4oji9ekJKmzqs5tN07MMIOtizFj2+NRk4CnYEfCeLW+kmqV5sWPaICKnhJt/5D9Gf2SNCJ/fK3
LjP5urLBkIgkolTsjOYRMSjoLxSInDmKiZ2ZFPD4ejONDIOiQOdhhZr/9PBHBY7IOMEHpRbhZ8ZD
+sSEUYKhWaGkXaI93odHHD6jHar5Qe7OVZf/CCYP8ykWGccYgkeJrxtrcMuYL+RqZlLZuuCB6Ljf
cjTzL9l7j52yalOB0QaMkYymzd5u+hIXUJXtbfm39lEi7n4CQQclHrd0WuefYmwTep7R7Xs2SkJO
Atrt8AEuduP4qDfIMa1O5u/pokQxDyCl92c0+EBBB7Fw1pXrEnad0rdh1SkRxn3miXoEZXWgONyL
PpfrJYHaEkNWS1T7w8xA36trCdRTsFSq/rA/iRAWk1vITQAyx9xQiV71ZTbAg8ntw8d7wzfBkPbF
rRMdBumHLc2WHAdcPEqePArGnzoGu47DoniekD0/WzZv9/NKM5HkTbsaZYPUc84suhWVVJ3zpSfV
JS4rjQIiQGQcSEQbVstNoBHuNfiPPK8cMbX/NXiu+AKJV3bu9R7P9dmG7ir8GVnvmqvfjNg8lGhE
HYV2V+UZlapgqWj/CLa01p1AWKZXSAVQuACWjn6xFULdUXJ8F7/ZwjjVKCp5N5UbJnjEZADGH1mZ
Fy7KRGJKUtisC2i4PF+fCdZ9hA9mC+IXr/VrDKGqHgB6nr9/D/NlFDuKppdKfrmq35PCfiIkuxIl
CgiZhOO8IhxAxur7VEILq+MWXYBnZ58B3dBBaHwPFGLRDjPkY+LQA9Rtm6T2o+hkLoXowt3BLX4G
QV05tGmWlWQ8G33ltzwnSkjht+lvHo4bO9hE7Hha/1F8/70O+Mxt2TG8tpjo83S428Zc0pFJwaB9
et6zH7JpmYAFWMA9jy7dkGzCV6BB5QcK3RzEYL9kB8Ec1jWKoqhrwqF8OYfg43YYOxRzRF37dUbC
/5kD6DZeHzwZyrW7288awpo7dUdBv1ecYPkfcmq6Z4PIx7M60mFVEoMtrygbA8zasM8qyaA4Kxvs
7CgALcC1/Y0yEvyBTHhnZ0J4lZBJHa88dDEtep2G/eFuaxeM2KBzRJQqBe+k10BrEWihCzMW/prM
BAaa13grzc/v3R38zREzZ9q1Ezt1WxxrCpqDpd4B7gPTuLhowCl89wo0basrggcdk7cL67ShQcfp
1dRe/fzisiPr+PVlYq6+wMZpO00RsIuDYHMbpZlNL8i5ugpEKlbcWMrZkFAiMYfIEoSUBLLtb5jj
Kg/RL96pyaXyTwDtn0ZUYQ+tn8QW8RVyLm9EVgKVSxEANY4LXTNuFvnR4ppEEEURyvimVq1ynnBn
nAJ8FRLi7aQyOVYsUqbbF62ppxp11XQVNnCNi0iNzN0ZM+nBGwupJI40W6klrQOYMPaQu4GRXNXx
nI/tdr24UVOCBVTUcL3CK3HYWAJW0IMn8uXnnFeni1cYntZelEHd/tL0PcvOfdd4F8Q1dmtr1NXg
d6gYsW4itF3D4bU4CFqVYZTTLER6UhwUH2XuVnG/b/ezEgu5aim+QKjXnWTNTDz8FsPH3rhXLDlq
CWQJxea5j7CN7sutc18JeplTvKnjAFXr1N7qEubtpHydsPBSLifBDE1WSX+w+hITwWGm7SbghkW3
YYPvb/VdI49G2BKyz7HpH1jQpwv8ZaQbhR9Etaang+elIjqBdywb9PYzz5ya/UX8J+rogpq35YdR
DuQCdBafd/ITzev5gZBhfjAtiMEwSSwPvZAW8xt5Hcw1E3S0Tec1mfm5DSFzTDI5Je4G19yZEHai
16uNjvrN+A0Dvz2xIBOPUFwR8Lhjka4KlGECeYXll8CZVXyFsrSQu2fTwc1EtVzuil5cKeryNDvD
DDtzroo215xVpPSxC78Mgdk+u2iYEA/N7wQCiNxRLpQdb0ib7D0hiQKRkfmpOdgOroscm5nbZqWG
RjshSMLcbPZbSzU9hoo9WCTr3EaqJ4wXuJhmdjxCDet7F0kYlNeH+di3HYmNEU2TYA74/CtcXBIw
sYrF+kAFdV9HcV+O1Mo0/JJJeBoZYlNbOxSoBnBj3wekPeixjCwt5XYH7JouqT5hR2opLW1T3/lU
X0duslGOHqo592zKYQG4QLq/13N+4PjH12zrrcAZZmPvQw1Kfp81w2esG4rI5LFxssk7Zh+I8K/H
XrKKPy4uBu971xpLmRoa7Fl0VmWappV0yLFdwbsyThhsifc+JYoJDRDfHODOXNqiW6MHTNG96nTe
D4wBdJJQztmLxI8w5QejTwApT/Hiz+1+kCcymnqLN+7g0vE0ip1JY4T6OCkYvuTsimYwxwsP7Jxk
frPIh8sJr69nrOIx8yjmmkTTpflptT+Huakp8Y9ESI57sCNS3zwqHt3caP8h0/gi8ov90tJAkfaE
nZkL/J+CBrG2qegt5ub9gOnh2idXbPBbSRSqQFDY2E62ZsceQzIJWF7wP8DtZVLRAx4yffuZWeT/
lqfUM9EZg+vnxF1hxJUIKtVrvUwrKQ0oOgWPVwST0t6LlA13m+jmyRXFwqbQJNQXhpEzootLGNDG
23loWlsMy2g0Al2imdrQM4Vc2TLPOPwHiaGMA2a4VJlTiA2KuJ63qfh/FR17VOrRLpl1urwlAoWG
CoYltSN0ozWhZE6bb/9lI7uliXFrZObBJzlDd5f3FP++kivfn/GjPFW34Z+KLPD515gnQMZTqWBe
zem7y/lSgI0imG4c/sJjZoCkcrrMtq+RxwA7tZJLJSITpS67SvL7pN5caPs0x1t/b0FkeDEFq10c
EgQC1rBW9Oy0LCLFIurbQ8YOmyUxSdT7iBGS7F4uf52i/BS8AdNJoGOsCWSoYFite1NSl3+ZEjd9
vGNKoLWBLfzPyt3O0c1eBfEJhhT7Db4j4Xmr/hPJlej2mFqy9j5ZcQ/TQHYXmMN+Y3lBDmWgGBNh
sCjKRfXjTF6WaU2smy3SbrXsmEeftdOY0fey2kbZ2KTx6JNYXeB5SOQVXlya2BFqhg/gfCxzmBvk
enudwKRE+dRjF9GSb31xPymydVh/+93sXe6wNMxPZlcweQWxt2cRWvtFqqGd522T9Qq1M9RWdTgB
p8ozV5KjEl/J9DFBYod9zSyCOlAhHVAi+1XW8bzI97EqHSKIgI2DBc9uFKez4NL335fKNKafa5E9
BZ+yzlH9/tBe07UfX78xsmN8YkZ8eFP6eFY54x0pAA51egMW+8Qe0vkjoBSN/L6CvhiT+7xm14pB
PjGPqGrMd81PNpJXeAgPZ2U9ukP1Ea2PYg+X/8x32512S7tqBVyHUD9kFmHT0jC7gPi6X2+6uGbk
9vzJLuy7kdqJkmGfHQ70VOzOpeZec7Ytn+JfLJJ3J+e30+julJUpfQunXXYPaQMVxYPq94RCtIcd
HjimGr2f+h7Objl07fQ+RY9Dp6wL/A5u8uY9nnASyiNs0Z9xA/4VZU/g3b62hqwq7lxbHmvyyVNM
TY8rINJ4MQC2rGG0Aj2zSmn0CAivZguyPwn45L+kkk7FO7uLoDP20mlEcvC7LED0k15+COV4rDzj
FGFkM4gvkSWQcBgysEIp+lPL5sIk9eWkC51C97O4N/3cHyzyBgUu+5U5hqQsXJIN5dPpouUAwV+k
nSfHnrtqXl/XWYySTCcA1xnqsCKdMrpVyzaEZIumlZjHpWmmkFlg7nj6lY8ShrwiVMLEsHOawODO
YlvXUO/xHtKlHia+X0n1ZAw/1CzAS3+gNyCeWyDzgKhr06+nsFxqmOi1ioOdSh5Cj9w2EuyyCTgs
8q0XASW/wTbRVBWtpNtV0w0AgCWM2Czufys+uI5T9Fm88pX156Mplr7EUUPpjDYFRvEBo+uHUjHW
lYnk84KcmMQaieMcXr72gzeBIg4HLdrfG6iGZhM2fy8Fj6r2oapsWat1y0yW9mi6NUeBA+Gh/JOp
on+ZDmHgdfTW75wYLjyT5IPsyJNbyqoHk3O+x4iIrSwFOFjgr8+Umgw95kAOhsL3Kgmo+1M47lTu
Do75wvyTtNPUlKxPqPRDtCtL+HiNipZfdXlbKwsndHV4t67uB+35AV5hSON0Ezc8wP42v1R8f5sW
Da+QM70ukqd2GT9pNBLxp3mnpvbtGswuV7uhWJXfL3L6CpIe7cttNMScPRLf3q77PK6HPWYCDEL7
z509NgQr0ojk9kw9A44m6EKPpm42Ecf3KipMbFB4PNHsXCIM4YtClzSE1b4dlJZD+rJvjVnR7ahj
k1IrSU6IOBlcUvOtK6JnCqVtcCAQdNcb7kW2C3Xe17dkfgXug2R7CSAdCwqzFrPnfTYIS8uJrobY
S9ur/YTsqTdeQGNRLWdfB+vZvPgp/Qzmi2rOcWwxqg378559E4M/lGti446Yttn823g2s4lJDMQa
FMPZX8eJ4RPwweUWY8ljA3ZfYVeeOgRc8JkBWjuuZwd9i9QZlJWbQQROkSh8ZyAk9qgwnGFpHB8j
VpgViKNIVqIF1PowCE2dNKWDuAR9nhyIVR6mFWSGMZHbt5eEXugCVplwTvcHTIkbe0BOgqUuZjmF
fqdVdH3gdOYCqZnqigmkvAY28/+CUPKlhBGzjSNLYOsretXbR5LnQ6o9qVNf95MYBHWLYg9Ko8Sr
44YODC/apcouJOiXqkHA/6gc0DOs1YeNomcvHdE9/v4zVMAwQ8BULQL+2KFaLjkVG8/eTtTyooqc
mX67uU+Uu6V8vcGT25AgSAyCdud/rSU6PdEs7QOSaDcSZQaX42nzP9O6a2FHmTFaTv6dCSCoZsVi
dxIYiHxWuV3vlyMYrCo/t16yazDd/klWmyDSuDrhhO5oUNEc8VRl0G8PYNyy+eNgkqv2BaZM98Ou
Edokq0O+5rzI7DhVT+dxHLgJLwwarVgWP3O4mg8ayyPNbCLBbrto3E1kYExfd2LA+cQ6hh4pjFH3
VuUPbMc3toUAM7jU1t9b/KqyQZ680pI8s9PdHuQJwJFld/RCFSsORLmf8qJ7KL7an/dS7U94WgFr
KhCo1pgViOeZMCyuTtclpK+b8HWrLT1VsJXpz+gFCBmkTD9gxVvmpchso1uc7R39IYPXX7inJzx4
Y4N4t7uCQ5kBmCPRGQAhAfcRblxqWlAyJwhUtxB/eqXox0R1/JthofmouAjKR/Vt6WYKzGQWGkf1
DxlFy6Id43Ay3pboD/k5jfsFeVLqV2LNuW2IE7Z8QQIsQN/5MIwbSgAa12sMdilD3wHvqNZJixDZ
+6YvqkSUUTw6OVPOVBkQPqtAD5f/leGfX4zFMFg/qnyjMXvBbmYsL1515jyvrGjQWwLQNAF2Voep
xNHkvFADx/eJE+DfhJGKjJK4/hd7V2vO28jTmq4z2JIjmcp/lS41dDhoweuJUJuERDIXH3Fh6mSU
F3kjAlhR+/yOjTmpGucVzWUVjTXsh3iDaWau+u1cMKUvHaBCagpq+d2cHSCoB4Y292XnP+NSXxZj
fxoXbC+lzEqHK5nNN6E3Yu/8XTP6sbZ6qbcvCWCgudXFoFukAH3jLjGkR0n+zkRS2D9o330ba2TS
s+OLTd+o9E4rsWeB0rbTLacbHbQd86jDuBDpCCcQe077eymRWO5LIRKWsuaXtY010+TdgF9ENFRj
LiUBSVjTjvC3J06RVPcfYTvzuftvo7Fwfc8PaRlyy7iYXlACAirB91tJsroGMc9+rP40IMiOcht2
6WiGRbKSw6NQoCFr3HP8pz7vkK/X5aYtu3orkpxj7rT+OSHGkuYaltfCnZZX+gx68p5kaepEOv+2
/tbP7+hEPQjXCfPhHWgC93w1ppVZTLWVsC9Xaa+cFS+Zn1QLANL5YymjvgtR8PUDzvnIifecM+N4
6O5KT9wIW+S/C/zSEB/3262DsaZaUKlxVr0HrkLLfa9Ytrh4FMbhbRrTUbt3UYCnOeXe3h+AwoeR
rwkIbjPRQ4GRZaxFlXHeaRJSaaICEPoCmmamGWYUlVXhKk4Snc/28seJeAHAPWUDcbSNP11tGM6x
USg4tWC1yne1Jd29OJkqIMBLUlpa0vClcG1jFjksPal6JgKK8TuDmUfWHA2pnlhunS4VFkPd4643
WOPS82eIasxIQ8g9wPio3Q/kzMSzUqh7BXHpttqX97nzy2c2F2WErxsX/Ip0mRBB/bizwr996qm6
HIk3VS5XcgeF3gi9DqMaKz4TpideGvxdxe0h+iguZMnKnBvVgSoG8hTQ9W5GbflkZ9GkiPx5//Uq
13XPzEj4K8WuY/IsfvAallxUyWiJprMF3vHzIXWaIfV+0WtG1qVFfmeAYzxitmVaWaIWbIiID9im
qag8BWGzRJcyrNQHI69mCJJlnhtBnTkKKWDrN1ccTTaKu9rx7xen0pcxHMLR8pAxMprSiW+22NrJ
TvWgPGBYr9UwXf1NB8s/DJ435ZooS0SwicjybVPNI0cpQ7OL3Gj6A1Zp3UTGs9eXwvrtPmeXEIeS
9ggjkIu6x693HsP0WShhz7UsMnIo7Buz5q6QcR1RLXGTCYWKXta3pS8cBDXYPKuFEzFObzva93gs
j6J1vKnNzWiV8iGG5eyo4UGcYrP7eed6QAHX7Yw+6ttYqRJt+0TLDHRpuC60p3O5ePo/ekGuDVyG
hItMSZuaPU9pLiBY6zS3jt4moYHoNb1pKQHk4S3feTaD3v+bi8wMQvVk/ONKscr3z/zS0VtIjsOR
d6Dhcf2arPJSXdWBk5O3Se7ulG0l66S/jt8+Nl1g2w5L1ZAxsd0wvKcNO1pexCUM14/xZHF11t/U
4i/KYDyTmD2KWxmXTFhdni/HwC8qYDMw+WssfjpEdXP+cJczMDuHkQoiwJF8R3SdU2hV8wU5jM5c
/ixvgOcxqZDMjpn5bhmRACXQpe9GAq8kceIh62n2pjpvSUIxXq0tlH9bORqarNOIGFXOp3uG1c+9
GGkbQWgHZDpqkM16RYR0nH14I7uXc7m175Zi0XLdAy61Gwg/SzugMl6aozcsyNy16QAnNT51wVtj
V64QN1sCkpAOer3qSM167kgCULqGrhHCKD4b0U0ckc0h4m4lhYXsOjF2k0jCRfwctE+LlWkxAZpN
7lTPU48/1642DRlnbOh5+c+mAi6K8T7Zd4faltUtPGvCeU5vEgwNi4i2CkTpKiYm3X9vY9V1SsDE
JNPEouQNPaACWx3LvV3I+tn0zJMoIDvYRlaNzlXJIkzQmHicMFDtdxe198R38B/mVYpaaCz1gKAy
yAl0Hmn23xjyIXbcqZ/BcBo4CuMsGm3XlfTkNoaqowlZFBnzZTVao7dFcgK6Z0V8a8gQTNTGrsPy
gotaWzCShbQToI5DZc7CAQpl2moxOv52dgf8LPyO/ivfdfPRCy8AfBORXOBAKTMDNXNMoAPn/LAy
LjOEiqj1Kk4gRbond4byJajW0Lh4RoglpDvQ1bBAdXpfOUOqF0U6oNV3E27xMsW2pFESh6N6oyw8
XWpSz3yHHRnWXnHhnLAw798dBZCK+vB1rG1DCuu0X94Sbjv0Nj933c++H8dmEdwFmNTWf10ApEW5
cPEBnM1Rcg2aS/2YLKsOY8R38Omt5T8Ff+OEPmTOhh9F5Xw07Ysx6V6G7amjKhV14JsAD3wwaOiS
gnHbv9es35KdH3YirE84/dEajcs46rvt/ZqJUgZWn6veoK8ioD8+Qz3l7yZM3OnJlYPJv3OcsMaz
B6QW8sPKvjuxauc8CTEsLoZjrYbfEGFv+OhFDYtmKr75reds3+I8GyMHiG7KM7rjUsT6OOecq71C
K6bR2K6AZNoFjuBfBXWVSZWXJbobGQtpomRz4/9iELHPqL0VyuAMfsNr0QMyYBJ1SxrQa8GqLdE+
Eripbq4ZbY1FO4ItwMs6zLwRg41hlXaCe9/7E6Qw7aT1WdzaH5FBwS/Qts4Yvno6igvgISNo5nzm
LUGKotCuVwDuqyxS0c7zlN2JPG7lR9Bsg+XB83R2aDEhQym6GABLdOzNYDtwvcyVdMJ1Ko8KzhKF
50oB+PJhUz75BauAD0aahAAoYZd3DdNTIRsBFAp/F8Hn9r2vNAPRNar8lEMGTYhdeuSvAQTLetaA
79REFot1c/ikwoQScl8QANUfR5SK+8H8Qqd+Sp9TxgwQweX78hdL3YBFomG+j8nEAkFE/2XXbGJD
BcbNCshiN0yEsE5Ebfax3lbdn6jB4eGfdsSfpW9SP25covyEvaWMb/nKOO3OKABsZyl90hEdgG+Q
0A1blQm6E9n1kpripgX87Ynvf75ND1t3kNrelCgDLj2ihFHw5BxWKaL5pR0uT5uhE1q5FvCN22Fi
lD3wcA0Bm8NDBrAPNTncu9xikv1HT3adoRAeJkYf9HjXzUrsV4mwqw/g22eFw10ZBh3gW/oBh9Y1
Avlt6+d74318pvXIMebYnrDIsGDXQ7PBtXqTz9jFBGDuocfQlEgJwCP6CYc8DYSjEW5PwQ3b7KCO
CSmKKmw6SsTakTjVHL2CV303/vwMPsiZ99FjIXzYM1zvSuHYMt5pmWftQjP0BvAg87Q6SFVwSGc6
hbUnctnYILcifEt044Zd6lm8v+Y/gg9tdtOzv/fFa/O3Rll7kDQ9BroHCj6Qln21I8+S4Rsx0oGv
jhV4HjtQGrDoq0cf/KxWjnh9blXcW7rAUXiJ/MahVq7VGWakfj6oDgAvT4J22sZ6mXXkGCeStk0w
isNQQ93P38201NuCZk3ha7Awe4Zu2keBm+K43Io+x9+yject7G0IwMQKO40KDiyjmixpSODYambf
L5uGKIOxzLW8MH12M//wnThw5nzFy7vNfIiCzyqbFjML2y28z5ShVC2ZkUqjxtjTW2JFymd6ix+U
Va2Dz6F4my/7xjQAr/bE6IUQn44nA++owGd95AH3XYwfGCaRSBi+Mm2v+alhLXTi+o7sF3YxO9vU
JQbBFmdekFsgNQAfvinvs/u2tLCTzcy9GHPiySu9ngvb1yzCsCOPS10M8phaKCuAFYE3UsOCrp4w
CHGrIxd58cRUgXrkDZ79cDIb6W2J5a25uQsaYmH+IFCbKWgi1szvYNroAZiey17hqsT7s8pd+4yF
e57B9oIzu62Xbw673lj0YikDwAsrjhSQwpOyx5S7yC3BZVliJv2l7RtE2dMwqN206gBDAB3Qb+m9
VWmue4jW91LWPBW+hB1IcXM1GvxWUcdLVgTbuBevfyfaj8fe63hM4SG0xbuRTPomQ0WaMDNkdoHA
IEvZbth6K8tf9PCgWEB1d+JkvMCdDxXJj2F2rEswkaI7/QLslLQs9EJVhDV33aOiiqeJ2nn64w30
YvLv3n1GDSjOpqmVQLn2btZkxJfVvX5abhwmyHRYjtoaMYNUd0g4AH52ywLS+0sDheK773yIb0Kk
Wkj9BknZ4A/eAR2Kon6K55eAilHKFeBDfilrzizG9uKgTM4BV6k0Su/DRj5cCI8NwewtNQB1SgJY
7xIE116oqTA9hgoEHAaJ+UAARLyKY53GS2sk+kiPJqMb1d3AmmU0qQiozXG0hjso4jgkXqgEf29V
puVbvz/vbCqqfb/nRUIvSCkhAjxYWMNJcPp1VZujY9tl6EJk2nxGDlwh4TsiFr4ErUT1j/y566ls
uKB7g/xsr00+fG8B7+Pt1+MEdnbfzDTOJtohH25ZSsF/XwiWf6O7AbGUUAJmGx2Ltr8mb4o3QUwU
WljsBT5d2NFT0dFd3A9BkWRzGPY6XsOv33tM5RRB2s9dviFq+obgEO9qs+Fuv9l4U9cvKcZ/16pX
5XuWANKDD25MHpGpGtObgh5WWAC61AS9RXuXLCAiLKHx3X2iE3JXDHrfL1ACK3Lf/8ZCnqnF0ShL
85Mg3qeuE1iIMWpYjTfqnF40zdFF4N7e22ybIXVZ8RIfif80NwDCFAvPA6xngtSnkDoanP4A/0G8
xn47CzPecoiHSC5HHIb8Dy82vGn2yQfsOQe6xYf/sAxsRPWt8sz7BKIGCv3ysrrQPm4uFDQuyCBH
oTi+l4y/IXslruqkRvOcPkCUzpBHH0wy8N0wSxVKRaF6qGohzt4W4hewFdjgsmn0xf8k4VK97/23
e9KQBfVK4UbQGbQBwP2LUzVclV6F/HNG8BWcBp6nlh1iBwMa/5oGVU4CocEVgl9/HKWgQczdgrnz
8KWSHQLq6U4JEpl183tHYg2LGu58jzzzw5fgVVKCj5wi9RkMjdy/o5b/95sHwG4z0Ww6TfrR2LOH
HTLDI0IQ/xwDSf+l+7Mb9v8uzDFaRYwzppostwuwRFVWQa7HA7fUGX4maIdXj+rmv2ijX3vCPvPr
Uq4sYBuj+s0Tw1CbbV3fLIJ61yw4527eoXX0Syr7EnBvpqRYpbkjtji+04XI+cQ9VFFYAI2nySmE
TrmeOe8VffrIXjX6kBB7d9JnLmX0gbaPPFoqpEX9PYdEzJnG8ncfjzioFtXbzerHUucjz78ibwbt
ROeosKcJO9hYovz6Z+8xKuXA0onCeVrx7UrJa6SOQFLgp4BqD8O94XDxC0t+u6sQZWmQiVLKc5Fb
YEElTOgzGgXgw807v0rslrfblJvQ7CJR6HyLceCca/6s2IEYy0dssJR5kmP19C/GQoCypxFt0wuG
QDMM0dPZci9TfMfmtGdFzoGu+A3z/6LGdfIDjE/Af+2UcF3CBCGzukn9OWyL9SZrXWHTlFE0ReX9
RDwWR6tI3iimaiEPdvwm8eY5XeR4E19u4JfVc8rYTj3cZHHA2Sa+Y5y4lnAOYmgcnyjPOGaldEFX
u++qfX9NC4k/gu52wXSweS8QxkEapUZUMlelOgxt3fedTjka5PkU56glnBHPq74YCpmVHCKslE9t
9WP9mFgJ3ZN7TkiVNRzVT/hCBH++QO/Kw/JToNvZAhcsyTYcuxBJmkO/Vkw1XVG3NiVMf+v0d5zI
CulzFnpfzRwM8xwhGnh43MK/NV2tusY5eYXkr8vAnang6tl/skwwW4wdcjYPWQps39etOnb+GL3l
M52Ha/6aFEw50tbX1Op022TnAuKm18SJSHMmDF7MJceoHKPSd4kuqkzUo7ss97FNUyZA383u5bHh
kTczjd7RZDDDdaz53q4GGHOe6jpz1HArxaSTxtEqbdYbjvHrT+6LiUi3Czr4h9mckHeOHdgyYkXG
j48yqF48ZKchEoISZclVbDZ8YPFUBry5ndhmV+ydRywGXi41sVbtj8V0lerV5XA38I98i0Rf9DFG
AB/PtN7GQ+h/iyFW3TA+eNV4X8Vl9L20321mg1vEYVUJCkORpLWfzrX4q3wJYst9w/GLepI4LJxz
nH6+TPe9MJGRm/izNpygvauFghAUrCLhmdekq2BJE4cCXB7BySfr5OvSw9M7NrMaBpgXZFZrZycA
1s/rA1WdF/g4C9bihiv3k4tFU3eMaIbPaSgMg58UGeWf23qXcVPWFY98jJcalPyLRh434lnzDSr+
pQfRAKulS5Fdcb5vZwV0Sje4VKuwaTF0aHvPxhX0D/Yxi4AIWJgCU01HparQ2002ahMbQWJ2sGxs
/jOJHSWzj25EKK7Oa3WtMRAstGyWsPq51BJoMNMa46JR+8OAsaUCwgCAO/6RqGvwchB/UlSEvw8Q
rwrpOMvMI3HiSc5OM3h5vIn/ERNVMgnteuuO/ORoA7/Dlw0JQpECMhEJNyn/nqXrEHXtfEN1CrLw
rqpEQE8dU4mKQSU9TBSDx0bSsiZg3+zrGuaiRZCaphsaTWcEUUiw5QyGXVpPrnYZ2mMwp2M/u6Zf
5JByqUg7Vn9M15rvmNQ+H0T5/gSV+Fp0z7jRdBG+jVsHEvzy2s4utee9LMNaKNLSzgfVuJ/eXc7j
ADa2u5XeLYrsrxmn0V1Nx/RDHVgwD62r3689PSlcEaOy8zIO5FHpFciP0uED1ZHhoMQ2jHuwS0bR
G81n50Q/xJhE9oVWWh1VVqvlaXC4SQ08kMjRHu2gc7PxkTGkf1YExHs2pR+NpMZ5vrSHwNEYY/Ke
/ahcMCCa/Atotp0Rty/fCrnrcyiJEZy19gOyRt79NVtP4Cw/m3cRmxiWsUZuaVKsfj1BUUkPgQ6j
56LN9u8ImmOUG8kh0DT8tuOvdLaP3QRtEKZ06AuV/A2zARXpWfP1GmhSkua755cAJX1F2hZn2ZnO
DKv8w0Q7unNxWgGHvw/mGXWvujIIE6sDVEnzWDvgCeg3jtW6XCVyBjCkNLrGQgkHqF1Tw3Q4U2I4
R+fvcFYnMnm34qg7RSKkW6WEB6bk/I6/mf1YqIdxoHAUce0BjdcBMAGSbFp0CZAjMlkoX64Wpbzx
KXAfYZR53bzj0xfiScwlggnUwiEqkKuIYmqqCC2asr4ySmUu+Auew1tzlDHTImLts+v3HqFBKayg
W7NBHR8ypaCkBRfL78vX0RMW2PwTxQOIV5izOFSFpTfWx2NsUQRkRi2MkP4LcxjlcoPQz8YxS8Bb
BHFs5ZBw6zO1rTKchQfQ4G3l6CU9fGRy+PeZlQIlYsR9JTnDUgweaYuB8XY5sbc81F9trDxOiiWR
G5ip+aK9MBh8Ieh+jmmJKuvjUVpsNDO5+i6aB/4++iPW+yuX+Ws9buucz2zYw1EE9zJJeFhYhIbu
aLw0yB4DN4FkyR9lR+MqW/lNsMJFvqzIl1KnNfQhiUX6T+v+lOexNUoH65bQ1BDxdzDtr4IzZg4S
m9Ua51cjweFn3U+7alkR3v7RNAXNGoZYjvoxMGVRER0GQ3nitKprcLKZ3hkG3/2UuMIyOsJQwNID
6j+Q0CWApTqFtRA2zueCFmq7dW5gJCmHyCGqitZCcSdH9KyKugJrkzNi5sNja3os6KUCErlX/W3A
Pzj/6qxbOEnuTCXY5NJqp4tjxZL++zfQ5PCQWUUP6yLS5JBo77SU6HTVCvVb3+oUY9xLeVv+JKD/
ENIgYUq0bbYbHEiqVWM655i4P8agto5Rd39Wc12q5Kg1qx41EJLzBqGmKn4vwOOu5dNporK3gHoa
j2Lcj/e2Yra0Vk5h+dUIyikDfWLUMYcFLROM4zGj02N+fTa+RlGAXcaJAWb+oVanSqnGCo+JTljW
03w+4CA/va5FlBdkfLKkti8lCZD/sIHsWk1vjnJvVIpsxSxl6sNoaPT5e2LldOddgUnIWOCPPQG8
YEcxMxIasK+y6jYVc/burKncR0wq91Tzc0lwiZE7nr4cRZQwEG8But/AEkELayQdVAdlDgpIe4Yz
SP1EzMD7q/O2yaLzsw0KJ8PwYcuF8jw4USH8vLTS3lNR3QL/wQS0yW0kb75CbZhWEqhUC/MlRjMF
/pOVlDYsxgD8Jj6z/GxvRzS2ov1sWZmhs2s4XRuGe1Dprk4qZ0WlpOdTdO20xcIgFvdcmSUtvyVr
urdaV9tt84QYCB28ZVdNwJGDF4mPWAn1NB8hwCqwSFizHucsn7QDScppH+6xF/7LsD6gRmU6DAcH
Yri8CbWSEabKBN3mlhZ8uv1xE7SBIsdQzFd/mpU2jUzOYUwB4IhHsglOa6Krh0rJxpyhXjwhWz3I
dzu4ehsXN2Vw5g5YqBsRda8eucQZDOCzkc19W+1lc63T0b8m0NxcvB3F0kVWnxjbl+vrleUtDG9/
dbSYrk5vyMBPOywynPlAmIizsr4JzziZ1k1jRZKIJZBWXAg5eq/aH+kdGdDOmG2i47xZMivxPxWB
NZCpsqIqy+H6e+FRu1j8Kbu3unpuskd6H1s3IXHF9iZmRyZ3P94sX1m7Cwu7Idkp8czTbWj4NJsF
UuSLSGTCfLSDJj+O5mdlRYwgfDirFu74KFoO1xZBxMhynJSg9dSKCatLrfd+NIHmyzNWeSP071uA
V3zujN+EEj3mGyOvkerUMPd6JeQzhBS+EudJTVPU8AQWnpxAXQo1x2QEaNwBmvB+K4oIbZ5LYxbX
lhkaDayLf7Il+9ay/lAUqaJoYk0dvkQLA+eFf0fP1cYoC5UWnZ1khE5ouEYn5uon1oNWGEqKWf+X
eDD1NUOSnksU8taWSxjwbuN1vXU/xxTYAoUhnuP2vbswcCQLYpYC/8lsZy/yEd43r1+cbRbt617m
WAmauE1I7gCQyEEe4tbp0py+q1Q1eJQ90N9n7lZxyCn9D7Nj7k6WdOBcgX69Tb9m1fmEWQM2Rcg1
L4BiSMmMF+BWjyZTaSNY5vEgquZQ48z69fnuf7aMHGZjZuONsinSIbzI7D9NvfgNR2VM35O+Rhpr
1C5GkTVABZa+BcPyrYIF237nvoPq0sEQlCukfL0pzEDmnV99EFQ+JOOpLcVmmchjkAc6nnxYic4X
LW6PeY1MaNS+3OwA+xKHcOqDe6670XbDPJPha330K3ZjARShUtFJrWhi+7QL5l2JCJcSJAC5BXFG
JW95hWYELLJQ6tydScMxAzpALLn1egNAcdvEIf9PMeE0iZRlB9IhuirHbjkdWdSDRcMSagBf+QRd
OVZrnl7AYW8VM2/GEch3ND7Ygk9arJGmp2eRyy9hpG0NLc71WDEjF071pp3NdzVysQsuGhYgkJTm
eXMHZ1wNlLR7fyb6gSlbBNbGvtOBYeJzS1kfWkNNZKSMGJbbVdE8XZP1dNtdHku6NsitSXFWAUoQ
Tj8XzV1EEIESqMnaBXTK+69bn13Sr7XhhNcKeDcWZwjrjRmUsJ0RRfyyrdjscPrA5HcSaqCjpHIy
mVvcHSFuDaoUYz6AIhQ0JGlcD9EclO2Q5Gnx+UZ+Ss8qUDdvf9o475V9YDJtVWCK+05hshGWsYaz
ZY7r0yu1gDs+KS9HSl0VQJaeCxQwvUW18AhzXTxCMKrmGWe5xhGJw1y/qxPT6xgUx29g9EpGR0T6
5+HpfiC2bWilJSDNA6ZC7MaBXfPSQYs9yGIp1khJYR2Y6AniYqw8gjYCV3WeME5IKcVf14tJbnUr
dUYI+9INlz6Cjpc6EeZYyOUF4V8fBGLJsnhTTi+/kMm5bquuzSPagOps664X5ibI8e0hhG9ioO9A
/8NKInC72LhHJwJR3uzefSDLOl7Dg9AcB7HYjWFfEMHjRfJ8hXe5L/Ro71gMeXcod73/xDx6XBXQ
pVG7p00WQnkKvfuXIDz5fDdfo1lmnSD3OfPDcqJ9Zx7CvBhomRLS0DsqtyA27fHFbjz/nze+JnaF
oWNFUNZtZrckOFdyOSIo5c8RGK6lBt0NRfFCgMsweXhObAeAdVDTYnEmyrf5p2Izr/Gxcagm0dOZ
IKMa07W5NKIEur9wamaIAEubgZNASLIvo+p5SuMcEAmodkerty9jUZuGhKbiWIYjS80BmS27QS9z
jrHqOHIF5aPgjj/luBao86GQRxcBnF7CWwZPKdA0MDjbgHIuWyLS3tnvNkbW663wkm9ie/lBg+X9
l0Pbtp6Zxtg/U8CFcMc8hqI2y6hV3ou9qHaemym5Z9RwLGKU6qETFCq2hEYrQRt7Ftbef0MxQZQt
ukwt7+VGn3OhTBDBTxmdcc+XvaF84OUdWee40ZwreOW0Ld/05RDeql6blwq9P4RNFnBjn8lT/ihv
9uHU07wJA+h2rC5IgTmrlr7n5/Ow5p8kt0iYdzEJvNZ7oS7JLpTwXzbjK2kdNzPMRL3+kWtLiOqT
t/YtvJw36523wR8KgHj1zSsAzxMl4VIxt01drDtxjy1ScZ0c6VfpTGopo9dx+sRWzLPToXjFeHkI
/lw6qLgud+FKeTJfH17IcQVtEzgVDGeqmYdUtVfpVwgPOZRriP2/cKCQgXNutWehzQg+XS6p9Spf
WDD/vBZDgurQ1UDsfQ/2EKRCfELM4sZpjD6ilMShWamJDDLUScnWI/IDeYFHWPwH0bpHoaubO3hJ
ckB6YRIP3OkmkF0jTjppfYTUrFKr+s6GL0NPSwmgdj9jemVGUfvEZaAdi0W1eCmRPV8F1sFpnbU4
FSxpMxp3asf34T1GbGMhitEWvjNN6MaWE6FQfB3+FaRkP/k+ywgVGbeOLSR8ba5xyYdTXixkGWED
5GZFzPIl4J5QTaDV9EMtU+3SUbF63zYQG5l4Fpf5MSIG6K4iHXfsJCSAIOIVSZgNxZAyBmfCgzGO
2acchpmqdt+9FsNvF/gRjVOtRQI6mhAI8k9wCUtIAXP2MP499EpMPI2+QXiOA5CEqfCGYbM71ldW
UxXEHC2SI6A9dYtvQHLDjStg2JdLtmRzSknGl+v6nV3sOdkkRAnlgHdUmAUXfeSkI0c4Qjlo0LhY
+KU83nt/TRFXkTaUCIqEgfgbRFD8MANqTnBW9yl244J9V0C1on2BRGpvQ3kg9D8GtoufR7bhECBY
jEi/HuwJsLWKgnRMGjAixRJR/DgKCE1NwDRm17XCUQqT98JP33qzXIhjrNZBh+fcUEOIiZ48Cww6
YS+Kp34xBcHNtD6YEKV0hJG7qlCknixO/dACI9yjFSnuIqAin1MFYkHKchSvFjBLet6pYtj2f87C
agYl0BBjoVomGKgKtjmDTzEQ4phwa+htxr+kKQT0SZe7fgmaT9RVU1ZPoZjpXdclzO71DtznnX3u
cWopsJ6afm5xaagsXpKfmVc2MStMsh4rrqZG5j2rsfW6cuYya4ChkEShHy1dNi4VDXH8PAyoidmk
cZVqgMri3mr4aL1X5M9ZkjuBfJr3GCZnfFRN8W8f0EftUieoz/VR+V5F6iRRseE8dHqqL1v8Lek1
ckPkabbXORP5H09uLiTBSn/Ac6RyUfIO3dFUiyK1VeHpM/OXC04VkqbCIUR1MVa3U8TrKYJ5tDe4
4mF3Olr30WBu0nAIUDPOZrGGo610ZgpiOmSe3GShE7X4acBUGeU3eS7sThxkA3f1hPMlGON5tZMp
vG8wABxQzcGw6PdMjunGAryAIE1tkTuGUtkz8NvUtl+PAsj9YPBIGLv9XU48ARQOcQo2cNEOrAMv
dVcPlH0zpUfo4mEt7avjgNA79sDftqkAkK7N1OWAVBC+a39XE5XglMjENczYAcl+O/QZwm80UaJV
SPCtVl8c3ZITIZNryGMuL0Lpn1RjQFrPzpi2e/bxJj33+mbuISwC7cmFAFeTolG7NuNADL87WZDw
s6dMC5pX6z4Tlo160tAPIfNO0o+ls0Hzjx1JiKIr43ScveY2lENC2+NirR4QgEcJ35XgGNGjLpYb
pdrpoXKQ7TONLu/Zinaz5UF4cKynrqc36Zzo+BwNLc6adUoHeOoARkfzafeBQtCE+/ncSaVpKbQh
3VZrekcupyS1FldF/7Jb0SB+VX6Tg6jYNo4XscHIq2qrWpJHUkj2jqYrpe9wJQLquW/+Fz0hCM37
vILmJaDwLyqOYrICoheox+/GKBMNykuUgGusK00JRZ7tdDzGdRvDNSJKk5Mi9vpzJugwABQby3Xz
BtvrWLUpJsfwukKIIRUxVxeVkJG7FRQEr8Vt03lLb9CjhxpFRk+ps5cid6URx2avtxRcd3/ky7E6
oUfIgC0NiISniNVNsxdQhBliDDSbAGKc+GR9ck4CJgDj59JyBpIY94hpKPWzXGgIChYWC/hjuFz8
eG4DVomHZ9P6Tz4cpwEt82HG8MvMEOFVj/uPG6bZPu1lfS9WMIMXhnb9OiZvvhyio3VRQaqHnN2U
9zedV1WQ7rwSceXs4441UB8liIqEmYwFTWs3IFwaPXRhMVZh7e7TouElacq0rv6PnbE90j+jMaLF
rvsVwbjp0TJ4sL3X1JokZvn637AEfj++ybOBnHQFo37ig4tzel+psE+aRSf8FmB+nPrVXxbVqTpr
9w+YSfsvrdOGX0egG6556bdBFEspMXjlO/RUQL8UjAJpcWZ2cVWjtr04INiBLrgQORSZbMSjsQ8w
nU/s4xu5deXzVQ8OAQANT5mL6Gmuq2Wm11BUeLRmCzMguBnLl0Ok6VIgvROuYIjrcyk838GCSl3b
mr0+D19LskstHRgcdzfbBn4PcdVFQvnQ3CM3gbOByzpDZdSC8wtn6XTL38jafVFheF7ghahxEkZT
uE0kJD/312YYpaYpGcqUxUjwazU5pN5kK8vj/HzUcgLs1i8fhiRD156Bq1BPVlYAUkSM8ANosc7S
TglZ9fXuh2l0KeXNPrdFeifM5BJMLgPZ+1MdvPe9LHYdt8ryH5DMw5nieKwQdsyKSClD6VoXwDet
uCFceCNhbD/YtpelyXCRh5e7I+WVSJM0YnIRd5FJTaWi5U2SMHTcd1Rad2PiOaBRzUj93MdH/Bt0
183CT6rg+SNdx3rFLsRUYBrFnjkLj7gxIxV9uoRQe0ptM84WAg8HK6ar9eZ5tkXdIZYzKno6ndlk
4zzs7HcXsZt0m0DCXFMyhehk1zA9MUTKFTlmK+fzf0JCHnmjjNQkcMDBWebUcuGhhtpmpUxdvID/
a0mzznaZQDpdx1fPpfMOGxlNOs0YC1rXqp7GvRnmBVtCoO7GaHH1ZoO1PfgHlBGj8UgXFGavVQGY
BE1rVnFSUa7lABa2EBeEhyDU/wgk+B6m2AUxhN9O9gl39E+qeaDCKSTx6SpbNGCx81I7M6E3IniT
/Re8SWc+GTAjKxmugRnZsNIh5GgKy1OiFJ6YYyib7FldhOfaqUPIa2kds0WwnnzuoPm66NOAWDbN
wXtl3J9sALO2FrfrDmQhCs4P9u/DTdGcu3NX1bQkRryglppX5cs59Nm5mGmdR88ihpGo3v1F4sAO
Ap41lXSe3CWSkKydGqLBUFsF//egpZ/dLIcknq3Q1rQJiNgUiptd999CAC+YK72pMqqQ12xVz1Gg
C3OmsDOSW3VdCPsSnXg2lgrfsJb8wKMccPioMptiqUkUyZFQcK+gsww69M1W2FcI7LQUs2/6A8f9
hJBaTFOW5Yxo7IddJ28QJaJ6k4oF5diUXjRgONJWBiC6j9Bm/6oD+7Qq+3G5FDcL55fDdPj8Wzu4
un60Jmb15baFUxy0Z9rhlQ6mnwIp2IWy5O9LAFdW82sMVhrJ54I+9MRa/l4Vw5br8GsRxI60hGLX
sFxeCq4Ko4q9ZZPB4tDE9vnJWe9jr4BDg1SWshsjJULNzANMlwKI0EfUhS8J4W195jcWVuJNgHV7
d6D0q20jRmxp2FwXhsu6CgLfxZNQco6+YuXgowQFVcUOkGM9SHb/8f3eKEQkV5F7KbM0ehiN3BN4
T/PuDSdqYpXWErlNf7wQSdJrC2k8X4gXmwSVqjmw2ggx/PF3NVJUl3H3xTXYghOabSQREgph5Jy5
LFvmCfBdkOd7U6/Um9Z8UfspPNIkW7Sh2lnF2Jhw3okoQ0LVBjxeUVHApAlQSm48QyN1Yrhs0xw7
RDYWUN5ZA07uYxBrJuPibNxfCBa+czfQeBDG1DGtPHm7wxXmY9M/5SVeSprVl3dqsQrr2gCphI1n
+LHhJexN1PIm53Gd4ULcGAxubGL/S+mfDnyj1bV5LP5/FweaghKpvJYaeco/Du/ToRbDn7EsQf0S
2hlvV+Iv2RnBEDtCsfBLczQRxQLPTxP3yeqrHHUIfTCLr4IkEvE5mkALVjw0P737dM6iFKCHQMvc
1a8JLOyP7oFzWHYXmyDDGpqs1R17FOTMYyrMwQu/EcIGDy01/zH1ewF3vGFBFsErorcjOzPHMyPA
4bz3B/3bS2oFj4B4XPHdJFgJ8Vh3yiWuv3bZQq/Fm6e44vlr8YWALVzSu4tXj1Qhx26elmqoE+Kj
ZFr/8DL6iDVUXxIn0ujJJdRE3Yh1VXlBRiWq08cuYxm4OpbLevE3qcTFfU5bTadh0VNSDqcF4VQj
NcpMu2y3wKdM6wDvtQ8YEnkQVtHeb0pxYZz61a3xPg1mZB/ux9XmT7LPaqA4EVfYYOSZxt93/Uo+
5NX1N64yiyEmNk0tp9KAdCJs7QeqQ8WwzgSglqT2skZdlxwkB3w6Vtq4NtmvZen3ulSHLJ3aUEZs
9UEQjukIv/vzBKNhtwpjw1f1eMZdpD/0WgJNwESEBjOcIQ30bNrWZ2qcDqIuPTGjf3grZ/mA4VHl
T0buC+P4PKEB3lxzh96dXPFPfRtpCgKDn0aO4l66hZINDqZg0aPLtJ9JW1KJmJiqIJla72rrOtAr
UfI95nKMNrU4GUlIpbJT4Ru5dNushZ8wQFfHNnOWzX6ptPD0kwwhzq5Ho7k7h9idLMCPPibb3KDY
7X1sZYqUuctuSiy5a2ByBXJ68GdPqqA9EO+coGF6GTMQ6VOgsfWHTWYOs2BQy8Bf8xR6f/6CWGGj
OesMGNDuUoUlRIwZjjWSVVSX803yPauWAYWuYNPPFXUKxu7+uSm+GJlOAbyVp9RNwlkm9NRr0YTD
MrkTZRgajj0hnYgyEIVSgjbBAGbx6/EklJRXxJ8Iz7m5Zgfc3rQvmF8xJgmFu0I3/nx4IDtgtq9d
iJWYbD0CpTYaSEy/YNMwa2gQC9NJsOLmHlXnunR/QSnQOfw7nn2JpcUF5vRa2Sjo9m+nYnZxepO+
zmn3WpNKjVA54x4duOaVvG2xKWIQMh7wEPMpOtbGEhlcIcTBeFz7Az8UzSPuY+hL35Vw7CXCx0bW
VA6xFJ40KGMvgMFOmaPXmztXHbkIUfkdzTwBmeHq70J5BQpU7rjWiqKFitAzUXX1pB+Z91j1yvEk
YkgjsP/4kjPknl3W+eczONV6dtJE4pGxifOV2ZqrAr2r9Zn+PVVs1NogynOZBF46sjXs2CmqDs6+
QtuZ2c6JDZPNq8ZGtss4TTdK/L4n8VckGehee9bgBD6oqOyFZ1+wNthiA924cA2WJ5JBTrBqr+1O
BFUXq0EIKEATAYPhMw5W+QJaLlxT3ZchOHFygqHp+yTH6EbralrHfQCcknda0p3mugku3TiRFbPC
3LTioRaQaEZY3i9CuxRVJ8ppcPt5zr3ek79BaMfg87VnBSsPEcK/uWifDyuZImt0xTob23swyxkf
Yx22/p0dot+TqGV91dPdFhreSao9aGRDYn6F8AJKRHUrSNLC5cX5Fyqn8fcqB2aIj+F9iCsv2Jo0
u1xwek+0GaNcxV/ZppMJhHGCWlh8w856VaQzqUfRkN9bqicnfSo1zCwbNEPXQnPN6deaNL+dJLFk
mwqOemNfVYeQLRgL13PcXfUjf8GMzEGVaRtgJcLHRDPjftDxflmZ4JTcUdGG/RRllz6n+7APyNAt
c/LluWO4CnNKv194pv3twb6QXuTnsLoD1lG7q0gGXfOP6mHYF+W994JiSblhfvQ8MRbIWTVwcKVn
kO0yKQfObTs7OSPjKNGgMBwUYaTwiszTkPxkpOYOtMHXTIOIDp3XtfGHX1mgide8OciGBnsNWshG
fvYqw0GD/sH7gKO1IMeYoPD+xzkREDUMG3caOSrVe+Wf7NUb57QQ+yPxO2vinFEmbI+snnNX70su
UYG5wy49DgaDjPmHwKZ7l9PKVwYUFpUWeFVG1GDXOx0brNFiWlxJMgqpn/wIoEUQZqls2j0NgOcH
u388Oz+JBlQbEuuvOUmdS0wGVbqVpNetMCOvSIcIh4S0QJ+d/M0OnjWTUCBHLBKV8i1AYjAVz+GZ
pV7rY3sFyW13lpEKat9K2HIcLz5pkuiE6VOsqQyy4LVgP6CiNRgdXi+FHRz0D1gs1mPbsBt4n8yP
yelt3oal2+gfTV+kshaf9Nf953ErX0z0HFVGY7Vr62odvMDUBaG1rFPDYnrSjHDX1kxgFa37m1Vz
cgL05AiOwt332bBY/FC+Ym8NKs/QwTXBqAlRP+lpTwA8qYmfSkeYXHA/4FeZTb+LGlG46NXcv+8X
VXg8EMerb92hTWYfI69dHPonmzEYLXPile2dN43VKMiyH5B4wCnTrdZNsJ8OOv9D4qrJkIT8ulS8
GtpB/1LYrS6aZta0oZg4PDI/9C9gtCnafLBYs8tpDU6j2YMMfyW19PfEV1GPs6RX9UTjRuzuOs22
wVwfK80SJLRDqHGSfuHlrv7+yPHA4KTqNMapytLjPsaTWWsrh6m33KmnL6MXtSFejOc/kudIz8IQ
SfN7LJSM5W2sGTZrR9mxc4dDFPd7QJg0VEqzzZgpvBYQZ3B/GIhROsTTsyp3mINJbJIAnPA1nUST
Zs3upQKkFSLKk959ccdoLxDaKXIpIORm0RbzrRAb2Pgs+022uQaSgQQqrPgf6rZ6vinzjqeEcS3h
+43y3mciwPf4W9CBTG/30MFzwMMVP65mSk/GtWPJV/Tv+xc83VoV/A0Qvy4OUVG0SaDPFifk3ksO
LnFSM6UbxobQJK+V2E8Dz0qGmMHueS+fkCmvuFZFhy159n2mgo69eo9odM3pFr3MlMAxJGELvsLN
6oyuBQYBEMTtTe8yQ7Q/Gv2rVS0FBcUlVqwaiq4VUlWJCc3N7U+9/C1iwgml93JpbtQc20Vgg7Dy
cmw29fP5fRqhHNvPtF+e6SPAEugQ8fUYumFJn5zjMWjY8DEU+YoKWsFhKEj8TghFm2GeMztynpke
/cUY/HxoX/T6FoXmZvb3Af0ZlP6m3p4oagFHREOYdyElGfOEukBxkHhDRuXhGtp0ssjtJ69a2zYP
gA8NpF8AtJVdZuu57o1Xt5P3331mVTP4gMILgitlL+/mLiQo6LolaoqK/oUcbpcXMOxK2Diif+lF
YpH/z6vvLMtf5QV7VRFcz6tEt3LwZ+bXQ6AiH1mT+3O4zFo+1Zu0hWGkos4EM8uU0Gf0XlMBLoou
Iac0bsWVBYopmfbpLYcBNdkSoCsCZ7ToMCZ1sWYP3spgSJPCg24whYgu3rLfWT8RKE8I+62H1hvZ
BmY18HKGxrOcqycQTxX1x2O7FP3ZYy5XuZXLZLxUzkIbxqmRSf56NsA6pwB15ss8xBn7avNK4omp
s7cRqyT7Ik7mM8Q7taFJs7gys3STCqMhvTx8CJB0eMbS1cmbmdvM+kEv/y0yhvwcyK/iIoZ0dqBO
sKYHNTyOUHf6xlbDMsClUShhJ9tqZhEZHTu8eI7uHgcLp+NEdrPxr34W+ERn13MFpRWTPWue5Tif
/Os0Jsv09u/K666JAmSj+83WDgfIt1SkgXpUKIZ7G0VxM9Y8W9OFfI4cayj14MJWmrY6EQbKb0Gu
p6TPaypchGSuJu/D8Dfsg60WrmlAnNBkcUdlIp0yvzJksofFS+Y39fdfLXckh4GHENfqbn8LCcHy
8XnwuaHUtGXBxdgutXXLn0X8vvacxvXiY40QgONU+W2R/HPbVhGijN3OVC+9bb/Om+AQYNb0Ybsi
gYHRkmu607e+JQFjN972t7a7IXqYVGkbR4m4HENdKy6YMV7Gr6bjYEGnn4lk5c2eSRmH8Caf/7AH
TKZrrny5MQwqn9Bk8CtOk7iGDh8/Q2qXpPK9+wZJMVh/9QMhc8O2Z8l/AfJGwDyA2LfBf4QPhvw6
e6UqAqyJNnIGX/0t1PT1fdw2laYrSxgUsFElOpvZRqjmx2vXvHC0R7DO/BfJnUQ4I1fWHoAT3uG9
h2f9hsKyegovRteavYDZTVdqOQoFAGUKJ5JIdAneduFf4uEbR6pJaraMo5Z1Ws59YlUVaZbVMRqI
KvF+TXkTXJ7El/DeLcBE/o7Ai67lR3+YK2KoNSDRZZmwf0X/3UzO7FIPExuQop5Hxmk3mQCM2oHb
6dFgiQjGxCvkeSN1V2fB4R/bz8BkezfNKBgL0lEM/PnkhdHefAfs8cgZs1ZNUDk0R2laLUqX2EdY
ZJjstGWCg461biBhT/mBxXxa4iPJIX+qkhEIAEM9Uj3g6/BNbYdYZjUN2zxX6CwyaRqV6K2/wqiF
8DA+ZdH526WdsbPwhAY5bessQoFtZUJ3AcsBkGqdgVi5aJB8EBTTuHc5sZ50fAH+uXE77VHrx2Gc
5dnsNfTLwd6SL3XYdeSyh936Qhxxwty79/tNCX/o80CrkXM3B3vHMZ/UUXT1OXxk+o2uJd9Xo+JA
GOWoVJyOXRhlexl3UZUmG5tvj5BoKxz7bcrdZ50Vws4llU1OGDVpF3u6c6viGhqlmQg2SMGmJsOE
jV2D70s7wf4NzuUEIXCfCTkRTBI51I419ckc+mNVB9udf8co2sXzZnWHUYXk4Dsuj/fKGpO8m9SW
o8TetB1vGzX0QhZcE4PZPFcgSwZ7Cp4dhBOs4NR1E58v8awbBQEWo6rYeU1lDAXiXn63lfhjPv1x
KakrqnDTB30O0tVwR8tnTFrRrbpnoNGZGzGQcHd3IQfL4vsJ9uJAULaUBraA6DDRNK6JvPdKvAzs
Aspvk1uMqpKiZKQNrKfA3mJ/v260StH3qu6c3RH6fTpSBBK7lPYnL0HMDa4krD+YORbLbfVoL2Ni
qzmLaV+chAJz5UY7xcPqaUsl0iC2pRIT8esBH7IKlB3E3AOBubaBILQYHJfD2oVnlqPQHiTuQCzR
Dt2kxqR0AEjuIf3cBCubEG2oE9bdilaPieizBUeoOhpWgdRYShugnn92YJdaJYTZNKT4PuhYNoUC
BqWzMzf3tsHoTMVYOg5gEz+ijh99CSjkDFkVuAVjxPqmbUVsQJ6VBx21M5sfbUG5tqGS+nr2VKjp
wF0dv9ONvCGHWhyDE3gqM5cHn1SeclhVe2dIBjDoL1OHDzV8xZJSKzDDNfRt2uiZIjRyc6myp8Wb
GRkJoGFsqGMNSC+fhHBXAD/xtzUdYl+Tw12doHVyju3VwufBlk9eNnkUgpZpMslcLV83cQC1vU3n
ngw1npoi9ZHCFSeopN+7CLmcvLVvAyb9xg/DcO3DS9P7FABsDHDrgflwZDGeIlVfsjACfiEKExwW
RZb2FcG4mlQ0xOjj8A3Yj9tvqbkHV3vNhy4V8W79Uqd4Kf1xrD8CtPk//jxvLY2bQGVbh/EdlTV/
1bd9PvhVGxQ6T2q/Dwva8i2sfW9dJyoJOEioI3OZQWAc9Axr9LZbyMO0Zraeai/1l5p8/BT8ffrG
zU1cWpfCUR9Ka1O5DqB5L6IDwt+kfWe9FqyalD3v+jMeK4V3uXPKY34I+QFhQ0XgzVJaFmilLGfn
RN3JXgfgGMeRWbgeqFFKF0duBLdeI+QhJaOUY0mIbRG2A/C+roT56vG0oWAvEjWp1tpmpzeowAbf
MX9UOkA3ppgyTSHExaMRqtSPW9boY5mhEtL6J2rlZZ6g6uqJG/vi0bWBudJWqgEMSw/s+gl6TwSm
zw2eafu2W0dCeQPAGjIo6ugs4UJHZ+1HUE0uq2Frw8T+NJul4zBFdhxiTcuUzKgysHHnMsVth5HR
3ieQKVZL4rA0obtY28Ivp+ndgDRHEah4PXDf1S3Wy3vi7xqMFCJrLJzGy2VKXyoMd2U900s5jr6m
YEWwz4C6877610Y0ZhPFw35UC61JUI1gg9SasUGJC8KCnV5pnHMrBPaaY4VCjTrs2ZkQ9gortswI
xopyqG/NQ2kSDPvmnniGcvi3p5W67O+HsHB9B0a630Xwt/0NMNifJAdITDJ/3NctS3FcyB8WJVds
PvldVBqgUq6oayKvGtcbeDOFwoRQYBlKB4iVIQDawquENIcJXetL9k0iw96IovXVsVeUTz9Rzldz
D267XNKZm2fq4nNnBwropr2FDvnYFUPssgOYXJ4uxjgV9IWvP8d/ILYhaoIjMCMxKnRMYXGx23Jc
/5JOd4WKnDSuwaU60o5OJhdsjN15YiCqPwM5ARHCddFPzcuyed0a3qH8UJ93765+SoYAGnNuO9LQ
H42ZLImeTZbWgwamXcYa3ELeOWJdyP57wmhlfuFSei5nds1vktleXQM85InB3eH/gHwJpnHA16y1
eMsx+NANuFrCRZ9JzmlapiTUr4l+XfycC83K3UQKSZr1YvGngSgpSsBu6tMwl8s+ZhMqrrlfGJ/N
c3FiG9ANlrJIuU4pisHZs2UgjdORiwVL4IPWkfOQSk+09tN1WHToc6BSwUEdP7+cDCI/kXvv6oCm
4vuPPKScEFv0cFvwg/C62PxvGipEnC6nkPpaW6lsMWoXjar9OHXeIgGGVOtyvuOLLjPlbWIDK8n+
pqZnWTRwUig10EC3CPSYtRk+6srwGhhHe4P2hgBLdb91KVweayoCF/rYT7ra0KiXQIqsz8LGlWzx
O5xuI5/aaO6cNy0NURJDayX2Agd0aVB8NMMjqrGI3594Rhj+LoQZ5F4lb5ugQDgqDsK4pT6f36b4
cxeKCe2exvQ04F80ivNHuO5ywPIn+n26mRbOrIs6blx7Bcr1XsnYfSJnzeWaBpmm3spDuorEF4jk
Uj9bUKMZGm/2pWDLZNwQTcqo2CcqgP4ZJDvYkZuEQl0ubefintDn7YTUwra3/6lFHv9CJ0ZLJdvK
VXMQ9PnsbqcbQMKQQsANXpR1hmn2/rcX+OK5mG1v7oeg2JXgSGOTi+WNPz8Iw7Zl/sq4yJoyKgMe
FEvPsQwLeCDoEbTLK7LmUUZjbw+ycISUNU/0Er9rEFA9Ax3635xgddBu4gKR3aeaaOLJpIVa7X+J
zyJtJLWlW54XMpeMnuKrg0IaEKMeR8N0nCeC+DVOO1QeZjycyevjg/SLNP0bauqwacULCc5ccGUD
fLQYcL3fKeppkijfeo5nR3jkU1ab+1exr07Oljs4QnO8kaE6Fk+/5HKDi39yGXY7xyi4IqKkB/FR
fT9Vv+ZPi4HvqdaqQI+AsorFskkff60DGFWxAULsuiVX+rIHqQQZggwT21jus8gCbHYpZpw+Pg/y
Az95NYjgjOlf4N/TfoMw3j3Gvsa6HflUPYDPjek7Pyaf/cRWKEd5Pr5hZIKlMzl5NHUx3sR0ga5x
MyvSnVZGkZfEgC0A8IamHgc3UNup6N6XRk1g2BLYndonKg6oTrALIZ/2fAw1NND8JVYWx6h+HxFN
uD8DlZJEwfKAm2tmWVb3iGj2fNg6OSRHWOjKzCN6Dlk/l7v+n3gEGpkxWWUcHY9PX8HyulNpwJbU
M7+9DK+n4iOM4atss6sdh76ehEkJaM1/4VszkvIRLFWiFefkwUaeHzqBLSP+pewNKm5baAd5Rigv
I37H/tIKvv0BwtnCK5+/GrcP/NGk02r7msbtINSsP16Ig/Ey4dH8Ydhtpab9cQ0YNt1QAiEOQIhq
B7y8ZCc6TUwWYsqRHKa3QgcO79Mz5qcsmMaO5Mco8NBnkNQ4j+pBnrHHsUStaQNC65OncP8rsTFX
+lNuUfSi0nIk54ONAXse3sq3j4xS2dOK7/1w0fBLglNlVDGzU+AIAiAQxPP2ftwr5won6Nn2HeZN
ZLnA6eKVWZGz3GYpRd/wyI5SSZ/+PJh9NK1nBr4O6oua951K0ruaa4ufOkzEbKiEY7vUXwbGLAvk
abRXlIxt4S90miymWfORxegVYSqFqSiXGbGKzNLvYvNdQO0k4o4LgD2T6H5+figPwidihXHFJRCk
UPAUOD3xrMgNTHR/y/eugZG8/lLzKhWNpUkHA+O0O8x0MTLak4kAesYvnZVqA955KoilOROgcGIn
I2tUEQ3xmoF92r2sLyYlSlMwWVHLBj33Ps/Np7ngI2ebgI4+JbAnlPHRm5LB0WH53XyDNgLaNjUf
qBd2FKO856qKqz7uZbmSocWthsJyePdP9tcb2Ps2vDwJgIC2qZ7eGyD4kUCZOIi4QCmPyiXMEcxm
Eqav2r4+pdb6e2J4ZaoQ2Xzeh9akIxxl906YoLwPum+Sblx5vsMqktGPnLeNDnVm7BP2ZB44IYd5
SxWtWXHTuspwrdX2JlITZ9QKIazykfLVh3HjnwmYROh0rxv0qXnNZuX4fEK/wdnEz/uyd8a0WmGO
OZeEmZ/nYGWMIFlpBVAQWANuOyQkktBO1DkKZEZTVFaFaPZXqipdaG2lDCsTauvWBAiU4jMaD03+
VFgUvwgtvCNYuxRyJcShO4MA8kTkNQi/J8Xnuj+eQlAQ/VeUTAJ+5m0gC+xU6k2aAoZ8J/OlBwiK
wT/FkuLADHLRQTYip0flCVrlB/urySFdaArRAGKFZPNFQCWmuMLWu2oP3ERAcxFnl+cQNFjzNza3
lwv7F7v11D1qgdSPwl91A8VnB9piVWZm93UCGdqvx9R9IYOXJ6y94NUZq+byTQOD0dZNCj+ir/Ps
vfNE2y83Y4IN59HSY54aC8Lj5K/MRXJYwvUgmWdbpu0FY9RSPhvD9TF1zkfn99+3E5rm34qhP4Xc
tYzg6VRAPyxaWKOavHj92IuhLxFC7axapIjS2oRfMqp4TG8YIuAJffRH9A38Yrmc5B5C1gRBXMP3
KQMwvTIiviF53mi+UwQPf7jSvzxtsFXxEgEWDoVdVZUUjq2CRMNpjf7uN5qyS86eaSxEErBwPphb
M3jh59q9t4hBIg92EC0GO/NLQbdAPQhrpXxrwMXLPPCd6x+kkAN/a6WxUgLc3Vi4E6jjvoVoFa1H
3UZxy75d87JDQlq1eJrZjpxao2H6FpuHrc0HjkG2cbqtIRHGNRAeBNIqKU8UfGOgGnmp0QKle1Gp
+wQuHBYDDMecuC7O+u8OjnBTWPqouq8cC4TkfpklpEzxYFGGRf2k9aEU6LUEEbu+lZNKx1TnSeDP
UtEeoMkupnZsImkdKDFNDvZdGSPCqjyVOfQjWcNu4W5G+Lhk9Dy0taI/bNCSl6MBAt9aGMizR5Jg
nLV5r1f6yK45uNgHuIJxHJ6EdCkHlxJHbndgMycBaWcBeQMyLvkPqqSsjYWyn03qd2u7dtI36JUO
Dw3jZpHW4XXoYL+HmxQsYMROFk8M2eM9wTo7cwVE2AFZZReC4QDLiuS5daEdspE4Ofh+NNw8ulMq
mi8ZVptmQ7Sk2TcE0qlRLI3miqeR5V3VaHXkwa39uErBQxo6LZuPbS9DJCF3tSaWgOCLOkznSRmM
TjDsLsmEb81+YcTaAp33leQ4RKQuYOlThNdabG4sq4YsutJil24QhQft24zKBwciyE6Smk0kAS8i
akCcRHbSagVg2fixaeRgaXUtjd5yBafnbuwwo94zW9AarMPTFnw6pLNEfhlWXibriMeKPgwuoaCC
JQryXsIhi1pG/ohrDOI+uCDEeZGcF5sBfE0ogPYmc+PZeJHZs2Mmeq6FFzGCWUluyW3DYedY/IgH
0SRGDj3vncD0UcrD6hdJ3UPqHt4edeu/n/JczYUfKYWqN/dKMkLtiupbWsAMfVqEGhkGdxb3EFfw
RoisfhlcPB0a+nYoYPdNl3EThL0QRpzaWm1Sk+iv0aPMGgX7CAoKtB7PWK88SF8KD6emrh3m4PTt
y5pCDjdvr0ceq6LcRPQqS93qLV78JwU/IP3R57rPHz3l0q7s+KrPial4XAabtj0jJsMx/iJAPD3G
EzFw5sLt85Wfz6Iij/wWmCD4W21QvLPv/UKumpe3yOjH7cF6AWNbXnXsDxLsQWPb+CYLR1m0diEn
K7lQRloL2wBxne0DdGYTY2jrRskXUWGvTkkTnq0OmIDamr2fXWqQ4fgs0trZBWEgIIxwe+sJHs/6
31aIwQTf/1Gcb0hzVfbkADWNDVQisn9BzAgk5l9A5W4mXoL5kMWOqwrk3FgPFai3xKmWA8wqi9xD
EWaUhmAvzuH+iB17inrxW4tmdMiSEC7j/MkiqN0tklwpd2wcmD6QzjUZhZB5f/W1oQdxbL1YswyJ
rjsxtdYKQhQ6XQAsMtAcF/vRqlyBnVgT9nZnNjf+mlZnEz5X23k5df4oTq8vwI9Vn3Fn9JjZxOU5
U/R/bRSN/9KMp8A+qGbwkGkBADU4lK0FmEb3pPTLlc2YzCncGJUY5N+RJbgpXzI4SSrPilWehQA0
+vO6Xu/no3tH9pVwn0ms7/vmQB3FizmlcpbyDyRkUP+aCuq8qFTc1EHGN5y6e0c7nMC3uMU/tkV3
KeUBJvCKSBqGH74i0SruFhvGtNObYK0bNqZsjrdfP2JnUUMVgVbWWbviml1ESTw1vR2RXOq11zY2
8aFBut2cI/MjG1eBKuI/joEbNdd+v6yBWJ5EbVJszArzRfaG7aQatnvCRuhws8zVICochza7trcc
upF1GnbDDBSZGHiMIeak7uKkVNdWXFLqRsRZc0BKBYyLn7SuW1GcTJaYXm6WyOpIRbDaqIOPibhO
zN82IebEK1FeGTrnKODf+o1Rpyx19Jdre+q5SRZiimyFJW6BhlpmxJKKUtPYCija7CWWJp8UeZDZ
mbfwDVUm5W8OvRCUjYMTyTRaCXKSZtg3iyEClbBBLbuT7abgaN2ZqXiTx1G26vO42l3qdHmXPE0I
mOKOIHm0sSAUQuEaF4ilwwbQumHOUlbxXxbQrdZBVyo/QhiwEB9/WlCrpDU1XeT2oenh53+8pfx+
XE1XCrwJS9uc6hs7Svx+SR7lcveY3luVqun0VEEHc96K5MNUpWtqb1SJ2bdSuz/VK4c8szgTBBvv
e1rbW/vJYRv1eX/JAgp0DmUdF0HlpFAHBvDcmRbWG/EH7nw2EbKmYrtwcRABHKKJfu5Adxc1SoVu
RHDDeX2BXUFvwhQavw87XPmxnbonN4JS9uu36tPUX3HMDmS9FiF4+/vPifNpOMrF83M4aceuSiD9
2MeVpqO0rPr/TRaQEhugICfJpI5K4uFfhhheiE0HxqVdZoTsDnZAz2USwRaX/zxRS2n+BHmywe7W
Biu6OtNV71MniyRrzeM5xyLJDOODQRf7xSX40okDfuTVgXCeP8kiDSZuYG2xuv+Ok0t3N5+293NC
+gWEoFvO9pIN2R2oP+uvxBZRGA1MUlRy2jLXKNkjRnsfewW+DwUN/Mgcnfua13ylDO8mYUUxFrgE
rukjmMaYKNzgGdC2KgTMeBUWCwNkRS5qQzeG96anMp/vpb5PgYnvBEmJp0xcdzwT7T0aJZE9JK4f
cTzB/wb/2f1Hyvt5RaQpPutcerC+yrbtcOKhPvaXkhr2uqt/L9vs+8NDSqvM+zTpT5E16x5m1U6p
U2l/HTCP3/r57oyJ0CKPUWwdN8WuAFWAQaOLdveqjFAQL67nfn5OWfxgAB7u000EdsX6VSSErglH
Bx3uE9PbeKnDqBtkAgdhDRVnKbXLGtELyRjqY1wBcAjQU4vSrItPOVySabH5W2k67z5nckGLsh+V
onik+UjuDf/AaY1TwiaiRxqCZVhk+HQDlvKJNYhzsooeM4kMEyWy8QcHid8YERYAb+ds5GgTjJfE
ZldmerEgQN9dKYCMFhKvAN3q2EpqHHFqoGkoHT0+k075jF2G8yCKy5nDKFvhwnCbcgDG01Rkne0d
tHfH4iE3DWj0ec2d+0n6P5RE54YKi1b2TpqXvlA3sLm+sq7yimjajzHH3NwsCnJk1nE4PM8v7JhU
rumVlxs7gT/7ueiCgExITcJUFOl0vfsybo0rikjS18kEMzcvKJyfr3Dmrztz9xHNjVsXNP0Q151M
NAJ52mRQl/lLBJHz4GcFdub7bM7AlCgfs3/V+keRqR7X+NcZYBSrYRQQkzMOcKMYpUK9yVP1iaZK
/DdyVVnhIEraI3gm89qTXjMMyzirxZTUL41nAZh1mjOKIcJm17gYSdDnKMeY8e7SFvFbi82sSoUd
tejbVSGgJY5Xi/m/rfW3OORThdtqnk500DzIpAXGpHL76/2VoUDQJZd+lRT9uNvJ0q3IRgbvsydK
HnbbR0hoeya2HBThdJvmmS7Izl88I0Jfe/BvA9ho+n7ekzx0dC6tBPB3aPF7o9h60ONeJR7s6jPE
yjUcZyrpkqbcRPOqXl3/6JuFFA2QY6Jr4Rm3aT8zcJHnnW4Kc2O1tA4ph8QQ2V2b2NiPobF/y7L9
yPcN9c53Awou1LASbU9bybG7/vieNSRUzLain1BO12jgknDjGfz/iRChHzE0+b1Y9Tqjk8AeYDTL
hn+3z4ozvfS28UW1oh8iPENmNuJ3auPVwyd7iVuk+Lst5jPYEDTRBOcEye7kBEUybjYguX0+PEMt
e3sbDcaM8JNQBJTuvebM8zr8oXlPNuH4qOY4F4cN9poj9RTt7NYsN5FBbo2d+R6IwfPkBG4NPY8z
Ksoc0ThhERynlR03PdXmW/Z5eEcnHdfeSSAFC1OXtqRm+DHcZcDFVfudVPnX08iH6kIld5L/Kt0l
34gLMgh23ch8XGkEwuWs6m4IMe+fvhYHk03CUuhVZDy/UibHjjI8Xgb38by4qK3YiV1dUIF86I55
yhdKdYeO4pFsEsv+ZOr3IBcr35/D80E3SGghZheBxy1PUyLonnI91CrNOuMHwcnGVeOFwr56FxRE
6fnYB9+7IrH0byfFs/g6Jh0/XObamX3oXnGy1EStagl+dLw0nkcFPPQ+wqOfuUzZ7y0u+ryi7/Mv
GpvFu23AcXpTm4CboDDNC0CJ/cx1s98ico2YK1YFKO1vX8yNGHR9fhdCCZrh9Pn6zgnbdMgRHUoj
qVzg+DAZD+jSWUsSOSPrMYWFoZ5WJu0WIQCrDaO+dEkw+W4EQBTYGm44szr7drSfXUyXbDuv/W1i
47qJ8TwH9YWOs8Nk7UPtljwO97Oae95mjBWGzLn4SVwSrBEnxxwWuZLDLxLbCmbWVEPy174KNZHp
R8S/mHSyc7PvWDjOjYetXi4b8GjdI0FJdP0Su8KepkPtMfR3K8NAGyDVBMWZZDqWJJ9IAqq8mof3
cK9NW60p28ljapPGHcTWDiWjjLFAKa+baUBlBjqMFi6CjrXLbmNdkFT3vi/2gzfKdspSNGMOuG/k
Uawu732u9g/kZMH4SKsAyyqUTvEDdXnOZ0mEDM9Tanov/5pr6y/nS1dErkSg3P4mcGNveFjAiI8D
wDjuNI3chGR8TXEJSL8Ei84HWRUw2TdZslB+bypmZUOhBhGRwr6BoWlmOgBuvYK1fzB+3fa9S6cK
4BA/RrL8dKOjbyJpj+8hnbq3fCPasv76mdEX5T4lvg7qTEC7LeJtklMF4Qenb8VrITIKNgMKpEJd
RdaB3YPqaapOC2yoCi5c2H7BPmwie4Spkdd8Hm6u2kkbvEgxkAQd0WjjwCizTUNCxl39a9KN0AP/
KSIj2RRZrAQiflHCzeDtcn8CZSfSetr+CoCE+viheBImLOMhfYKEaxtQ5vMHfhtWQsb1r0ma7Lal
pVfqkn4NCfEqjxWPfcPWXr0k3tKpMu4MjVyNARdzsbyDslfwqLrbUvcjoK7pFV8RES9+gZvbKUb3
UGzAMalwNH+QoHyTjZ1y0IPNH3/JonvSr+vC1OiTsa0TYZvxi5sEGGyANKOiLUCwP5tVByrQtLMg
PJBYaAlCmegS5ncUxaNwEFTeZO9YtB4kdPZyAcHyivMGS7j5JpiNiH0BwlNhPg+dN66T8UjiggBE
vEAnfpEhHiNmVjLe18lre7I3Ru1qMEhJjjeHN6BNP4fpHUJhn+F0EEyEb9zM2BiEltzTJdajIVko
xLkFSQeBa4gF6OzquOCQfbhiFxo4fFvvIpBHXk0yg5aRw+cbZb6Qk7crr5YgNJ5D5D1VLtprnFtL
Qr0ZJ6KtbQlZWbYXOFtDUeu46WdTSCASMvnkJyyNMbUlJxePqtzAZOU+QZ9kDe1JhT3LtpZsPB0r
AZA6gvYlvf92JZARYVat0TfvnewSnk60zpr7kMQco18Y2yGrhmUFmvPsFtI7ZwDiQ2boTKYB34T+
SqVupvX5EO5MTDvJHJ0tneSLB1yYTbjNDfKTSaBpqGkRGrZfBywKGjn9H7m+BJlHqBqDRrBGs+2P
5ltocpVG6JSCjbLxORw0q4/j3xZaAS70gq7HUzgAqdzHLx/LtWn93xaZyOWChQO3+GUXiObWC7kB
q1Qws7842QIbOrAl5w6NE9iHhNf1pQl6iSHSonsxAA5i780Zpeo8G8SUZtDNsbfmV5H8QaeYd4bD
eyVlixmdN1cZ2e7XNdgw9m0OLmJgg/lyPN5PWVVc41ASGb/57DZNHdBh4iqOPmupx6PDtd9z5lii
6SDTLXUY47QCHsebnsuE8UixphBK6M9jmF2IE9lqI9LBxBccQPXWXuGNEv5hYGxUmmMpNZP4ikmt
3U+a4eWiagMCrwwpJtbvw6ueWhT6X3prkQQMyhf/F4+Ug9az5WkiuavEDEMxHWHCQjnol/puuRsB
e+ghlOfVgmoMedcLqB0diPA+Y9XyqbeVfwDBb2Ewpd8kv+vTXzXqwEu+jngpiRvvXfaFfDR59PyB
PXKlsqLJ1yo1CuEqHsSA/XSLKhH+sksPYp/Q+typpKfmHSKksZXvHkX2elAr5VhtSLPOzF1us/f0
e/kJhSnhK3ijgU4byuGgsRaO0GahHq1iqj4VeAuwE4W+9I3ICRC1Fr68dRcwBX3WWyfG/VoQ4reB
+53JuWDrN22m5GOh9z3iQ21jc/oIJ/rLBxT8EnMXrEVa78/W3kGQrq8Z3riEdZtLFqHOLlW34964
ruGwj8qzWxSvmT9G87wfOnDM8vsSSYo/R6UHg9Y8o6GpkWisxxcXexi6dSq7DY1pD2v9slVbqCWl
FC+BuKaoHcFjA8gEdpYIudnQUIYFyJrsfkPh+rACguBzvnL/ORQ7UXP3ryAAWpVNzH+kaXdazCDz
ry7xFyBHMYwPB5XShZAzvJzt4+K9wgb8rrpv3B5un5zVHi833E0zH696zNsAzaCabMDQCVq7LdWD
Zksl85thw9drK1j0yT6eIfCCiEeeN6+mdvsYPcr41uPPTOQkmpnDgeKFKmlkQNQ1c6pnxVMhOxdE
dJDGqNL5J7aHSrHsqUCQfJdG6/sz15m4AaOSNSWgf3HxbY81FG4ymPFrhFtnXnu70z49pWa3vG7c
+Y9JM4pfz/Va+cYxA+OYpinLh2jpGzNcsgJmMtfegfJJRmH634Z7Bh7WU8ACTxAIWkzjp7BK5w96
hWNdTZ+uhie5Z8E7l8ukFI2YyBjpv43Rbe2vxVZrl8wI/bpfW6szMSztwspxewzoSmkEBbursz4O
2qknI5SiONYDfUdMQdHKPlslq8lA8mySsshmb9H0jh/NQZVGr+pfdEqnbup6IFZ2O+XiouifrXOi
jkRgq2zhdm5IfyhgXu+4vEXfW5o8OFZjzJ8Os6B7XFYFzrvBb+ozYvp9nv//dKQykHEv2XHbciXh
+EzIs6YzqJ3KQXD2tfrxfKDTEfixz6cX7qQ1I/4thokmKZZQDib41iEiDmOW3vKNKovmVRsyLOW+
ktfJbFxsiyig8Cymqbnq4miUmxjzosso33+cr6cDP1ELmhDDiZOJPV4WUcxgpCCCZaGInHUcoYlm
bvFU1Sk1jBOeFl/u4KaXh8DiivWAH/bHQNJaVuumBrom0k31Nc7kv/hxOq5mXwnbY+QqDq6KkCo8
bLdjb6rBbT1oK144x2r9NFRvl58OB3QBT0GWj1AIYMgn8o7WqxeH1ADEWvVIGxsu2RiNCU4Q1Hys
Z6fnuwo7pGX/J2gv0azltitQWT6+BfeAwanmWQcYE/jSdtB8Ju1S3ZEGKiC4wFvZNEgPDHUqBCSp
Yrgygi3OahV2z6NeRMsZChb4H0rp3a/LKybIqn4a/7/cSuHeH7pgx90wCEY163PNWof8oyofaE2v
q0MZNUvDWs8rmtTkp8e6OaRGp3UVQXzWW+fS8Ni55LgX4xaSw8XU0LHYcL/U5TP6p+AEsw==
`protect end_protected
