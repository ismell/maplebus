`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YdPUHEbVpmrRFMy5BbUuH2UCjaSpbPEMVsts+v5dT1IndQ5NejbBs0G8vAg4suXtRslPbLBR7cIf
wqWT5hRIYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BcP4tuSTd3xtaikzwM+ec/FgaFt0i4J29OX8jvVFWjBcPIZrDC9wYh4ywYH46KhanKWRt99og192
DEd26hPC5iQTxlRFqSniYNrlye1zXu0tDWJQ7FNEnwZcG9ZoN/CNSctpQr/SGBHKUggY+qEfb2TT
Dwp33BGM34l85OZ5J7M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dJU6T+Y9BjYjcKJ9W2rDB82E+BAYCn6cDj7JjtePsn9pkOKZj+9Q18BV5+xQPYWEDQwzxvihpow4
dtVC1JTbxFDXdOBMWpZmVgHFYHmpq/JghxAOE2rqE+n4wln4Unuce3LdpDU2qFgI4z/fjBghIaxh
txdVZZtj5LAJfkttjRmUJqU193mSFL9jiUQzXixjv8adwB3Dyqda+zWTSfN3AuPISk71PtG4fTW+
8pg9lU/u89sVuNGjVCQGgtDug0P6oCsOBcxY59Powb6ZMX0bTwoPTTy6JNnOKH52viMTSsK7zOlM
y7CissMXOQHwhNc7ecaNVb72gCyjd9TFs7cTOQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qfqMjN0toCr5CJMTnUHTxN04rwXKsRTHawjKpNMbNTALGpFlWbMTPvxwHPNFZA7exGvSSX1F4C22
L4ggInD+HWrpf49QAIUpPdWr08kIH+t2+aTpHfVCBRgpcBkHDlUiFgURf/EUOsSRBT6YGf4DlVTX
RwllEAS4P1Yy2dxot/U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VLwYmT+2XPUWzKZMa8XZG1WNv2NMkuaJvFq2LAqmIlsQucdlMAQ0tsJAUN96C+sE6vq+1xxe5HvW
CWWPoaxlbLnwT2tmfZ8gASgLYJpZ5qAxVhY8nShFxseKx84EyoU/XXuPuymaDWvaSx1APXAEI8ZK
HtQjejDxM8I/vfCE2qJziAalNXv+F2OwzlKnVnbAG40VYUzh2Di4GEpTr2udiono6DIN/CCNPeWz
1szJRQ/LV0TBuH2TZe6cLTB2W3a0QqCTuEe2nm5ZjxHNGt20LjT9SWY/zkvCDF1MPKHCVRv0IMIO
VRroCAZv4P4sLmgfKaNPQjizswst6c7iTfLQOg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9552)
`protect data_block
Y4eZMYcDaeakDqp+0Ti4pwUSws4racnxd3P75//oW2M93tqCAxx9sVtHGgpcx7HBJZYdL6ueP7CL
+LfWQFxXvmUGqxfuou/oxriKJFael6GaVoAClJLRRtHUQjoJd8pXqpuRnvXU9dgrD3C8NsLFLGXx
JFccdaa5PXMkzv3T/DbH2nzhz4QL4PTh0JkBrHLTRh1bsTg0wNucAO+81OE48daZu7mt21qXJxzN
ErnuRjime/t50zXz5Clx4svX9ETzQttYRFaY5eLgryEUfZDxWw0lL4MJ73xHvHsIwi/N6AESZ9Kn
pos8HvcvKPpeCF1uijAajXZ/NA8g1DHrufKstygb9DgsANmhQZ6Vr2fN8CnOa1sQsHyUdkgBYRVl
H1SAcKthruTUCHcm2uX5Z6+LSOE9DfKbzODIa1Z6KoAAXKH9vOlUAVhQ756Xp+R/H593bP9OPRUP
LcXRuVBJVaZShBDsb7sEIa250d5Lzs74FHlBSq+2aSS6T6SkgV9cNtTU8hypUkYEm/+IRZRS8xOW
9WWOzf/g9x+PnJVl1WkNAoxH6JYlM153TcGgfh9fc3n4as3Gp24Hur3886hofG+RgT4JqJJf2wAT
wR4Yv6exY4kP9BJwyDBg7PU2Ulc3tLWFGik2dtQSBghW0QrNZMCPAarHiBq/gHJrxGEi9agrrO8W
b7WwZbFfwmRfqa2qhMAkhvDeU4kX2dVzPMhyxcrhgeV6e4Wng0AX9sr8o55H2t6gPkIVMfCOcCSG
gSQvtzWLGGM6CvxUIsmcB0/crJ8NH+rkI1wpGgpySz0a1maKpqbn/9LmeK1IzRqn46c657dla5LV
4bCQdgmHDvl8XtXRtrNWz2BdaBRnjW9Xzmwk5eF6NXFKICC6H6924TVZMgI/oS2WyB8PfgNrWf3f
v4fUR0SEHisznuWcHmIrwD+GBDFMJ/PPcwPyGE1NgUqVoYmoKclORvWrSsSCh3tG8/rIEfHDS+Gj
dRvyDDqFCbynR3IXADjiMWBe6K9MJj48UbKYaexiMFfSWwLg+eLWkV5tltPCctrwyEWCeYHGHh8k
uA2nDS13hqiu25DlGH5YJItSWN1uiKqV/7x3aWxkWB8mia7429gkvffhUebR/cSyF8BnZCpq9ilN
eS0vnYKWpM39msUKmm8TOQ3Do8jvBjMJ/eqbuiZcQOlTJlV8XJ6YlBCAXKAsTx+2vBKdMjQFcz7G
54yqunu71FUK7eYQ1AOKoMTtMgEfrqAIW0iOV4reEMmPfbbZCnxR4doLMURbEw35pFRiA4PsMMK9
HSJqntAUgQNQvOh0cH0TYeWRkFTs79HyjuheFVMJW0eggQwIh6f9MlrTJL6qDrb6ZgSeWCTV03Z5
/5M22l7R/SaRT8l1K+Hh8wwQWUjqxNnkE2YY2r7DBjUJsSVrdSfx78WykBiLT3esR5+KGpS0mgLn
gvwIHJpMk/Bm+42oUMmOE3QxQcRJhm/mEovj1et7m1nqkYxJeuu4q1aOmYbehry7KOkkUnZCfWiZ
b/vYpc1C9bMQOppl61uHFFzKm4qy5QBUgmnX9FQV5wPdBTIWeomMTaYIXehCNk+ZxcWp2COEcpaM
sJ0EmN4kLjt/QqLsN3nsjRkrtAf1KewZYc8XqZVrn+dCiS3H44x1VNCN/BpxhsI7giLudYRIwcFx
t+9aLgSRNVNyd9O6jJEHyGP2CoBIwSEdV8OfnVpjjZPoLeF21sofFM7B4aLC4glSNeKdcIE3MfAS
Lhhe8dzSp9gKa1TtJsAOVUcNOyrLZPG+9d5C+FTTSft5/BPDnqNw3UjN4xXuXhdBRWij7d/0kPkQ
h1TeUUhXHDpJCvACrWu0XspmZboCIXPb639k1EiDnZk7wZwVdOiYmNwaTiNDEyAKwqnwtKiwtkkP
OkcIdu0A6sxWDfNSTNFJt/yI0pQtZtixvBtyX5JmmFYJj49BIPYiHgK7pjDIY7RPHbecGoKt2/DL
pXgW+O5Dbs+ihnGMvFYa/ySlywCE4+e0MNuE2L4wLlaUQHhoHOWwU3ataEg5oqbTYfD0SaU8MS1l
exCl+YPorvWLM09tG9zFTW9pJA/LKlQgal/u79OX5vQbfBhYWaJmTdlItWBeDDXNo1N4PZH9KX+Y
yQfWvND+1m537cNokVQ5DaLjTKYhGoRzfx9HoYHKxaBvUoQvTTeUOZJxXGBNUlHcDPb2ZykdXFpw
4AYYi4qADyV/QMs5wAaII5oQzTD2D2agj+vH+ZEzFFvUzgvvMBvOOkDA104xMvzYzIuGv5RXXZLf
7x71CZPCPCNEvFGSdmyjWfmSFBdnebZxMMBOENciWG2ioNopYA53yLx3WVkd2QXzKvdBCRXBq/6X
G8lADkKjAqJ9f1aMvoiAgLBF8lufctJvusdcO70uWULlxLy6i9TN4mo9CSdL2P+2AO4sZVuzLkhf
RD99GrJFO+TxGVEz+zfWxgjj8/itn4oWnLEoe5/C1E0G+dsBrrps5Gsams2/Rf49b1TieuxFgmXl
nFEYE1DDje51VyBVKBCqCBGauxd0eUw6U4FgC7G0jPKd+jrwdLSnAZxGiCampGyQA4IU2BAkJk60
8Np8JM7sEOUgJSrY/ItEkFmw/H5D+sxza8jgRTSi9HImA7pS9XOAA6STTdxyfWHxM3hpYIzXt/5o
9QhHXnp90XTgnU4Ee5X+TEY5lRNF9kLWhrE0F1A6w3eUqe5WVlId6KatWnqpMVu8jGXserp6kLsr
rb9iGOaSFBJ4Rm10PW06ic9sgzuyXBRqnhbnfwTOQ/u03SZo4F9W/gBJvij094EUbaE/ca1yIsFi
dSB4qNWLkiNdLqPsex6Xd+vBsosbLdeK3XFYvetSTVIGA8NkNwhFyr2zS6Pb/R7hc1MHrNHTQ2kW
CK8uOr2QhIG1NCz8tUav2a+VxyEsLedxZJvczDE/Hq5mvenSTALUNMtJvTIUjAy1aY21Sq/YqCgX
Tz9z0CqXcDMIC2aIvF0Icup0Kmn+IsovudAPuM2sNhCxf4YUQYVcCW5PzOjKOlnS72vNVnFiK6/B
sKYeuPwUpVYK1BNraxD1Xks0jJj1F8UwNgNebhCaLAw5o6/WN4zP8ic6VXC1q/OlFyfelAbpulYQ
e91mgg4xwPy3nKmRn3xxEoxsfVkmJ/c+4uhUoFKKYQ8840fjsOGHeFM0LJ9y9BZF2qYmhSltY/8A
jHb8Q3xrxX8aXOSrPwoQ0umK0Mlgs69RuZ0krPneOIm9Kp1X23ri7qJrs09PEBxiG281mhBbH0V/
M/8GF41kCjsNbdkNxenskuQy0rGOL8bx1o1mjjZ1WdzJZDod20hNSmG15qWfjAaVyfLiqBanRy2Z
cfRkErP3xmM3Y84puEtsj9juh86YddGZXZ0w7tWq0DoFT7JmUCfbtBEei2kyJ/5C7LAFW92C+E+S
3lFRLxLSET+/j4rGZ88JC2UuXZehuRNe1Fo+AvfMx1oAz33G0DHhHVVZvQ9p7xodgLzCNpi1C9Pz
N2tq7rxLc5fRIerG2XQ09zbqSszGj1hhQaj17zhFx2b2HpO100FAw/eGj2ph1hJjgH85HV2DNRK/
eGujTXP016cGdjrjluUYRtcDY7FfK/KoMDjDP5jltva/AvjLQUZrREOBWYHfBLfq9aWEwis9AnxX
GZ3GQpWNpCtVIdziFcQ8QNE+GfGL0URef1J/bZ7R2xZgJcyyeXjNY+zaNH/Oy+Wt1enCq5eOSZQq
2Hev4LGb/AE6RJQZCIJM4MS4qs9wyQZardXGI9zP8yT1p7w6BfQqDmTJYTTVrwZT1+hoezMqWuS5
CRfZJMrVRl0vO6zitLheydeyFCewX9L12JHjBcYBKsye3YUi8KlJ81AR0kQiUuqoHUtZSHugMYR6
hk5u9ZPJmq0R5uj7RaRNCIj0CrlXGJXlD35A8jBlSFTLEuxeS5GQfz42wD/PP6sX1Wg++P8ZK2Uz
B+UJrAeDt2AQxhPLTiNSUMJzOPxtn8nr2VDq26cvdf5cuZiv8F3TTy2HyyBmo0ktuJ/3GCig5vc+
dwBqxqKWQbPY1GhTLfepdHDaCS8RzmJQ+1QOQrQugAMLMaxBdmW6ZBqLtzhOYxy6Zm5O/nBjN/tX
tzz6dN/+kgj2xGrQe+xufHvgyiZA+32pTHGL/FBFds1Ty4xw2H7vJFPTs9Fown0RZuryz9H3dbgS
2vHf0AKIzww5qEBjGhU17zaMrtI32kKbjqVmLT61idc3lZ6W3yt7tgejCyLlUgETm3SJL/J0Fjn9
IpHyrwYVF/7cjSVxjh66tup8DWa9HyvRXidt84fPxzjxvYB/9CgGLZIDK6ozoY386/HmPsjENUHR
ND3qoU9JqAcwokmVIM/JVuCA2NREFVYOGS7R3onfjhSgcGrcHXzuXSDoued6a4H8mvY2NNMWSamo
6W3yCtvGH6ELRCYUTeuDapVLC9eGZPyh5uZPYo5ci8RDvCN7PW8Llg4c2Y/LNR4geyjx8T+Dhebm
wf6IXxjhkCwxEReWOiH8gwSN7NCt1B0K79yUkM83Y/M5BfC+KCLX4UhaUD/oA0cKNbZ6M8fIp635
O+X5S0jgbaevyRZmKpbsrvDJ7PHyxejE4d9ygYTPkhFSRYpK15+Vd/knx9zEmakAf5tElb+s71ST
hfqbTsf8zh4eITLLPdD4kIuF9RezVSjhkkipDZ12Lp8PG7ampOLXkZxLZheoxl3ujXV6gD+D/4/G
+oiLSJlNKVGZxAysqCdIF9g27s6BXk/Epc18R3wZU5SyFZZ7n6KydinRU2Om8n7pL2pBgF94ub3R
aY9ydxz32NlUSpy2y8Jv7/rAsjAV59W9xBoWP7BfVkD0RJJxXQDdywD0ypVhHawrR+6lliOOTcVV
kSs0eBB5xhvZ0vl3s1h814OcCA2/ncU56gPvqAyK07i8GjXJTaf2h5cHhBGprH1ngviW8RNOoDlo
yoU9dttHyJknpOWoxJMh0/fBLyCR9yRtg8bFIWMohJ6TXzKhgi+9DWP+bQ+OGeyraBMQh+z0HOD7
riirFY2UaGMt7GZM1+LbUlFPvsGMWcq/iEuLMijLRmdCDgftxYOOyY2Bx84U45QT69h1uOcDky5Y
ZCnIVbjnvHkEsgQk9h71lQquiFjnmf3axWFH+FZvgEYwPHsobbi00qobaU+GHHM8QEzAbUPSLVDr
FpFKjgRz0YKwvx2MnWP63/tA7doHAXrH/E8GU3FTicnpKoVNCnIImlOhUDAiC5St+yxnakLT2T/l
nmNQLO28YST9oqn0JyvDtZ8MHI4TT5XXQaVARc5sO700BOtwbup8lCp8yj0j49Gk4TMap5VNJjcZ
b/naAU54uda4SLCLob/UnC0F4nbiRyY06vhYp0fxwOoXsxh45ZxYKFkO2cljV0FrQ2T6vcK1n34j
h5CfqU/HLH3T9O6MjVjV2v0vmOlNaFfkpBbjazUCqruwCBlOTEG3FuFBwMCmKdYWmdV4Wke91UoT
yMiQ7c2a9/4xaTJ8xPgWqgKs9EerKB/Hfmw0Uf9lnnqIa9j4XbuEu4ljMGPvS1feHxnZ3USwmFu1
sLOuS2zAA7eLDmd5sCt38zRCg2fa3EH2/drqp3dsNivdNn1bci2IVOacpcAJJ7NzPyDVDwvzXlxp
1nlS/GTLvgNtbePV49jTHucYGbCjP1TPfL+9Z5DRGr8HevOKUFZ/KxbNALkjZMC7ZNFwtL8RBeKd
zT3+KllqCoud+KV48J1ED11BdhoW4I6P70DRtF/6ZMEVJlXxrWsINrTSdcC0ZWw+/f9NnZvdjMO/
CipqJSm9DC7np8nRBHfhuu8KlPhigw1kKqb2SVZkKVeItMQG4zdSgrlH13jdTfo0H3L10wFjqI8l
yRKaSdO6aip33NX0jWrv6dzdW6Mh+T5cvKQ4tfNxnKzZMbKcmW8PoAwvD9zWaDYLPsiWEpwYHgo5
EVY4NBV5Vtth29m/nsyF5fcozIHnblLAsm2gTdcO/hQYzO1CDJmFeBj1c7kzAtBQiXZPpTO/RBGn
tdAiwywdum6IYWivnIupd5mYfqR0LBPSyhcwRDtx0gv2ACJUTBPnwZpK9Q1iPwPtVMiq9gjHVeg/
VG1bCK+EXUrwu0neiBWj9jQbQcI7POGdTVpnMphmAzKnGke/+2cwElD/zs2h8382+jpG3silMN+1
itPwYb36U7irCeRyHM6aWkhKOtXeRNUOQRDj/aT2089E9XDyqilUwCPVRHubp3iNNqV34teiaRzU
MFOs1tqUx2SYU0dNM462w4xNvEiFvnashvozGdQStcPcV0TgTwACeecGMSLa+OfGI3eUjZ3/p7Ub
OJXg8rI+OBGYO4MvheVBcXQeEV38rzbaCMrETG2ztAsmr7ygsY2KTh4+p+Zfa433FDrZRII/9jvE
vSzX/5Idbjl+wDiony48MhVt1PrxnT9T234eMcRmWMJdT8S41KJ2AeW4hJLuNCFFWCCrOYDr7uf/
BaQEekGoWMP2Wv7PpD2rF2jGF9JzDxKMusOihTbQYWv3+cHFBb7UqyERNNt5woONnx9nmQCdDkJc
LtVoaMCTeE0iqhvphARkqmLy4nERQ/uJFOB7Cq6qAZXg9KvzeFD1wwc2b4dViXZY4GyfwFKnkwYE
4OFxbBEKoawSW0tk2OB0uQ8NqsRY+5xqFG0QaRfp7LC76kJW+SZHp15Q6hmuQW24QmeFs5efN9YB
v7zvgB+TGOd7YcNuxJwwAuRxPTWMKEFFqVfPOuKe8UD3YGbsK3+xq53BCN/fOM5tQ6ShJlMh6ThZ
IDtuD01gtdLCoVUlOFsl/o/WrXHlgnoc8LAYx/Hm0r9ShLnv0p2B7ReTm54YV5oHblRO8gM82I/z
yI3tFWj3eu5kqQeCGggDQ9g02LyzErRso/YjKYckoX+46CEgT/DxYew9iDUxajeECPdcE9GSsxzt
w5PGAOgwyha5e1BFxMQwvYziKVGX1N8RciiJaUzRrLK9z3sO+lKzZNIWlv0fWy2CgdjvbqeqXwmf
fxG4FR4aACHi/beq3TfH7dpWnItT3yDbXT8mdjBrIcg6kfQZqb3ZLG9vCDpeHMruP0eJMP/WSpaQ
c4W+0Y+nU6OTIF/eDTesi2si9iDLvMQHBCvvw+JfMBPRU4OZDV490AtpmVcbUCXbY9mKhoASOB1y
/qlfu6gwJXn1UTZS5Jng8vcrhZy0j+EOLUJg4+Qs79Ebwuo5W6N7oxzmMJ3I9DS6Hbu21bUN46sH
BcdXaa3WrjP2F5QT/i92UKE0lSP3POAHZIVReM5tmGPtoW/trmC7qSLuTmcX5SRJ3Fm7sT6eFKLH
ffo+TeYrAwYytYFsFrvS8GWad8yNgDwD9WB0DMHFue65bxlQJMDBbU0DA0jx7gtIGoeNQt2U4Ek1
tgAX9PNzHq7DLFgIiunCeOe1fWVJLfuiRNAvocHOVCQrwQQ7mwsJARnRIeIMCjQyUr9m9kleCBli
XWsMJlvBlmoxeRQkP9yGdrM154Zl91J4fQEdkSGe7sOoyBB5Qvk7aG3bH6CQVnWwiXcsCYtYeF/R
qf/SnArAe6rl1LtboNPcCy7UT0vvY/f67J37YGGWUa+2zTmRYsz1vLV+dm+bn44M7K6zigtqqEkO
86k1sRsLs/LbNkr224KA88Tcgr8gu1Ws5Ysc1bYiO3/E4lzvgtzgHRU78dJyVt2b+VFlH2JBShR2
ViLVe5ZDEq9WDwAqtm9eF9R882tlHRMvk5LKjRixyj9adPeknyYzAhOIszlKR9TlFaLG+Ey6eltY
9hkmyrZyEzl2R7pYHzyO9EpqzK/nhEZKPYVnboRfxsBp+V6kfiHnATh6LQkoV9H2HuFX2P1egNY2
UOH5hr06zRloMUyrjt4dDBjmNqW7eopMt+I34PxMDEKK70OlX0oWFw4p/M9LVem/ZDJ9SPKE9/Cz
qsJygPP2kHQYhymf2vuPoDpbl0d05SGQnhir1CZx9uQxKrVOTx/nfpKfkjVkb7YRMWN7zyPJZ/M6
SqYteUKdY610FVL/Nu3SbVUbgn4F13nQFzF5xCEBSPZL4Z/oExLHb7i/L1grMi028J8syqJ35kPT
CwvdoG382QaH5vc/SO+tp+gh1IXJXlUnchu3h4vVkI4m/pAVqK7lOburL8DxDUxOmoLz7oI63x3E
I0bVlAKeLsZlMnSUYjVqUqSMQsd9js6QNUeM+nnbWX9/3PvoPd3T3uGu+E/vKRIhlmojklTzVIx/
0tQEHkPk2vIafRsDafuyYlx8MG3yK5Vid0yFrtH8j0P9aoOmTSGhUC0/l/yns9W5c/RdMreLTiqG
ENpLNU8UKwdyBRssKeVvoGxSR0bdxwZDCNvL3XmoUiMmySEkyKJZPxkob0nsMilSAZzmx49nCH4M
eN6regEcCFonMJPNiDhd+LQ/FiRLzYDEVG9cpOZxbv0/UGKi6eE+8Ct60eNX4Vy6WlydgyK6aGGa
Qh9TjL768GbXRNqwrhV+ra7DvILJUChSguGDDuliKLrJKDVJDnJcpFR9i6fbubClUjJH66kENm76
7HL6Z8WdTaaFmzBPvBiHVtomsJ/dOc4y2Tl1rZYn9ogE7zwy0yIQ6fF907Z+XaejZ8UP+X7ZhMUQ
00J4y2Ya7ghlWKdHsxyTkbN/Id/TN/y1ulQd/Q8PkdC0yTnJpVcmKwdoxtQpsk9FlZj23FpJhaWC
GNadMowpL4W1xQI58ltK5oVsq9RrTea9Tist6CSBigsXbN78reSu/fhVNPAYMIpxKNi6BeVKU/dY
Zx39IpZOM8pbEt5yaTx/ti3jZpbIWs4RCz+tQOV23t63M0Wb5quX6Xulvgsm6+fvn77befR1SneV
OeMqBoV0drOf9D5kDBteesNVdMaKxPLZMeYo9PPbqTI8AysZb02tQ6E8gPsPIG2gRdImYLk72GXs
XJ4pE8HHTTHxaA8BDvhGMh83IKZMbof/j/+eMxDUGWjLfJ51BjxQNVBrJ/lrcoz36E7pZoZZNVPL
zoIfYlxlPoEt9ffUsnzFJUyKt2gg5Q/a0pMi257d35XkFoKr5iMENn8JzJ5jpC8Rn2MuNhpr9dco
OFBwOh0vhEH0BHq6RMwPaIikdvOegto1NR5idUMr4I0xxtyb0OlyjsbcSwMW1xu0BKRbcxOqDjVO
zKx+zGqDXdcnxg3VQbRTXSLKENs7dZzjrsLxbQcDI6nt29IDIO+o1PClDuxDtvgJYV5pZFeSXqqu
qB4E+alrJ6XNo/QpcBuXUhC9D/ZKN6810AtQrieawEd3SbqcefhKbvrXGFbFWF7Xwc0Kn7ke39Ev
l2pm70n2dUwaR4LNr4wGmH9nvXF/e9HoUo+jIFbN/v2H7cZF1DodoHCWFYYsZePfc/5dEKxnxkry
EHhX2Rs7yJFxUE2eU3i1MeTxz25klN8hP1QOMfd8LtvpE8hAK8ikq3VPuMqXbiDBYuGNp7vENrOy
UeCmmQPteQ3hd+BUXWOQ9AvT5wUQd9fUZij9n81RoBKqLVrsTfc/CKxOjKo7M2obLfXmInE517lW
00qLTyjFmOCu8oEKyXUtY+5ymburehXFV42IqIVV+aUe0uyegyIlCJO48UDBu/P5ENsjLQPWPdM+
f/h/5Jsp4Srfy7zORfv7B/rQjjkkuanRAD0LVYVgz36LmlvUkoq+sEgUoq3a6HkMoWnftqrPKnbe
7I5YeAz7S39uZJObTM+qjAPHp6UfXWwvyprGtwnI8UrrjMX5X7w+4Q/IUDpQKD9jm6vpaTol5XKB
T6sXOzSWJr2M8uT1bzrUl5oNAxatVEhTuyJIwxtadUu08u8jRuPCC4Ffa31+nmQ/+sRMCmHDeT7f
c8zag7d5P1ut+zbt0xWgBi48YKubIDPLYCloAHbnOJ5AmXQJYsNM0TYXVTteZtV9Fldj9tL1gzaR
NiXrBobFUBZnxsEYBZnmTdugPMwez6Eq/QJpdcM3rDNk3N/h0DjPjIekS+ePjUESVClitakhjoGC
kgGcIZrYs9yAKGqwofuaaLSlMZntxvXQqXw1CDEqlxE18mYJcYvgQwmrJVMT0mjiYckp1Jjw2uST
fPO5hzX/JJv5hJgiIVl2QSUpyj6pZE6Goodj/v/jrKoFP4tj+4yvM3njOye3Lv2wLJCY2JotfDXt
zKeinkcFDudC5N6tmrKwMdaZ3Mz/3Yf9mRIVrZTMXGNv9ACtL/QyiUvjZpoQYb6TbaaLoqiv1Ask
M9RT2FVIFn98RwjTvUEsgzxt8NLXIGMSoU0SByEFJoa2YObpBT/7gqgdii6p/NGbUn7DmzjZGFm6
jU0P2KKB9d97CoBVCMvrDgccibPLtTO5NEmapO5kZtojl/hSiu676fA1rZvJFqKgKCPIVPI2GIli
cCCr0XKkpkOHcnn388vertcxk2yEKzqF19FEDU26rF+uDIhcuIcy/V8NYeABVvGKPH5k9xwsgRmy
ugrHSbb4qtRSREt1VwFaFUHaV2w2qcuM83V2s1wOI1RbFo+blh0bsl/0WqBSyIwx+dQz/7NnKwpB
4yJA2YZfbbJr2jfH25eMTr+X5agjZwsg5TZ7IYcClWdPGiOIlivvWCkb0XCF1Dhh49+ndBFyFeHy
k6MI6M0rR44ucmuUELqzd6dEHIuDDNQFDxmqJSjTMX3nmLfL0ovGN02+pbEjCqUcDcSTKSfVhyH6
VKI372YUclsWNNnL0K4++RcPxT+a6uCM0F6Mkm6Wd7/JYX0UVLhy/y4e134CCTixXqIEVfWqvq6i
GhEIGixG9FioOkPwwVAFVMD2Z7NzhN6JMmCOHrBWQXZG5MvCEDwClCQH7rf7SPpS+4bPGmju4jkw
gLKWmNlENUXQ1DPLF89mM0CgYsqkGyMQrI5CBEt2eW9+jQMTAnKOqCuef1MUoj3IXo6mr+mXqYDT
WGF52dYYfLwSlgT8OQ4EAgfJROCU68QtBbNN/RJ4yItjE11q7n3YxWQg9F4D/IjPENLwB6rsyhqN
hhY5l4OfPIAsjX6ZtwmSSJ7zWVqFbceZnpY3KD2uxG9Lz6YX6gpmafW4Z8Kjl3usspFJxWdWWV7G
danB6xdhBPUKwIo+FUMzsUuOtqnkqjgqwCCaDi+8bZoSPdxKjPmyp7eh0fmJWizaRd43elKQFCL1
U05wopvUCJtSbH7ybmV40ImoHTjkGgeQMQGvi8Em73HxqVXja2LXl/tznuglxRNaguH9afoMH7ve
QgXcNmAdYAVGVRdKlwF9Gc/jjWEGUui5EW12ZkjdGFENe24GCUTXd0fmPlUrHd8Es3/PIapUahM7
YDyNBFgiStx4Y9WmgnJOEw+g2/2fRdXwHRBhAvs+XfGoDxm9h/fwtEDOrDzgJVvjAYiWVeu02x+w
usoe//57CFQcukN1/wuU3MfBgKLQVpu4hsio8pinpuoYPgwKt/YcGSvG6CtClUL/3JnYBLYaKFfl
10AU/4Rwgg+kHKsDaNFOoopA7ta3u3+hhwBJWICm0oRqPPM6nfnisOeBFghVRqI715XM+tMHh95J
IMFQc8dr3TqJwfDeJfJsBTUu/UhvKoefia/VaTmxbRRdpXS/Sh8JUDUEFQSdzt7L5/1jUfiEg1Zv
NW6wQFNz4jocqRciJZ0oBBY0IYt1Dx6UrHJvTgYQYJ6EaAfrhnzv4xbXRt8br4fvVGcF8pZRlXWX
iJvdVIvQITJPSWNNpGwr9Qkcgw9lPsXBwxuvJlw9btJN+K9yfxop/kIshbgtAE5Vr5zm3QmTS0Wk
MVug8/C2mGUTTv5ybnFCzkElA+GKdG4ZiCvN6aGLW3+fi83Y7rAoT8CSH2luJzWQCYspWjBlIlct
nor+W8OWPh/jKf9Z69VCRnIYAITshux9/CWxmGB1i8slJlOtAwMXWYjbqH4TRdwwekAGIJN7mW2I
MxenJ8NduLu3+X3rX4aZjvoeN6BBLJIEmNE5R0y21xGPZMbhYylNpAA+Qtlad3T0QmQw9O289FS+
l8cbjBCbz2rjwE9SMlTv/1/BIhTkF4LDCl2Jfc3jtvwNu2iCasN4ELT9q8/QQVlg3LkLCvDMEW/G
eDQwnEsvwxkNLNX6Xk7P3cUTj60FcNlkmcfQanbrJsSJVMLoN0u9+FIt1ZIvCFWMBRQRpOyVBD76
1oCAZYv/jDGREHCkDVwIN31+QN00VY8MtOYp4RdsEoT0SBvNCBe2/+a+pRxXbskkpj6Wh+uoIKI5
0UzH9kqTeOp/Dv3hLK5AbFOflEEJI+VxqgVyeB8ulgM28z68bZ5v/vl3TmWJlRn0dIMLcX57iST/
R3BnKMMpx+U7Aw00nXv8G7ZEziSNIMw3G6RkTUJCMqPXoeT69/5ftPKPzlKNFzzFeiJiAjEW38kk
Qug5w1K5BNoTAPDqxGtB2341Nj076ufdJDm7MnQ8vOaEZFIcOdspggFJNOQok6CLdxy8ZCL9xIWh
DG/xoNMsyh8VcDte9YckRJTEmxaszQKC/jSwnJJw4XLV+XgRgXPvocgBrHhP2u4lPsrlJrV20vtx
U4JqC4Gh2A4RkBgSL6aStgCwCq5WQsD4fgSPXUviDF3yrYmT+mzpkecmHgrL76Nr6dabt88qGJ7a
htTairZu2uexcsMo+3sPDZhbHPV6X0zu+RMYTt4Y4p5zQzsVXBVOYlLU376xaEm3aXs23+axZE15
wpVR2/Vbp8WHw5ltPeeO2wKeWSjCGacky1x2Ipx/fS5wKXOEb6r2EPHdLBpcIqo4VPLNl2puon3M
54zDA54fgLDSaX+mN9T/CnXU+mAnTF0s166JVTFovr/3
`protect end_protected
