`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gjxNsCDFkC9M22hEUCIn5A9J4SEpzi7/2EIXwqj7B+rMuUupqgwNCW2JZsw95TSkCmsvLqSSQqyC
V87S77f4yQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f58/zXzeGXQ9vWzEHQdRdZdgO2jFCxslr/TxtXLsWxLbFxaAPBn++8h9AyzMXT8Mu/6Df7oE/y5R
fjgH1CxiWFJBRknc4BuDASF2DL1eVs0jO+2jqalmUUvVjErb/hTrrwz1jS0/xDWx67Sl+45QIkCE
+WQ5BRjnn3TzJ2M+u4Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ONwt1LxmBGjLQoP7iZpm4qToBvuznMYjhxFhBPzDRIc5dljyvKcQW/FppXFNGTRWtxyygCmP7uFL
gvL0H0wFgnek632oiArDuIRWY54vtDWURSqSEmHTs+iba7UWIL0/e20KP0NkFQHvXuwgujhJas4p
PDvfsIuUnovWEBkq0Iogm6eijGLiefQi2sAuA3wydFUYFOcWVOf7Eq1Q++/xwsYKdBoIXg3j2KjQ
CLJZftds5vS7unNvevXB5d+DQHah36zsY/Tex6DdAPGbuGs0fqz5O+GOjsfNWHqfJRp8kxeW2tN8
6GWgwb1Q6B0u5O9OI2EPG1g2uK/CbAT00PzLAA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uihvvqZxSdyREC5QfeKbV0P/ZCuPIotzXGusCr7keBCpbki0WrNXA8dTkxjR8GXOg7P1l9mnd6qG
w9uFqHdw2JEI2gWj8F0Pf1zBtemX+Fc6XhkGgw6o2PlXSvQPdAsTtGImc8KrYBWs82A9HCpPEqvO
dPtgPtNn5LGcSwR3RF4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UfIJpkd5lyq0gGuDqfkQw4tLJn0aw0PuV2RpnTTZ2XKRQEmSmnQWrM2cynDysKoI6wwiYVceW3BW
vrKbVYlzUF3fmGGVnRjxXRC7bpce5vTv0wvFNq7Xo+8i93Y5TJokZxoU9bQ/YT5dxRcGHfo59bDz
U11uKxaH1ro8q6BPzXWZyrglFLqTbd0B8Bn2CysOhksoNhPQX6xTIq4PcFiOgIoDU+dQabA6D1Vd
NfXQC5iRKfIewvxWxLJwhfCYTNyB5f37TKIrnKuKCYK/FZVkVbJ83hkPOiwk9GupjYbbe9uG3ooK
5LzlbVaoL8mqHc+viP9lxurOGK+B8fPwv1D/EQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 448000)
`protect data_block
e0PrdpaQjt+ktc9HCrOczRE38kqN2vQYeAzwlr8cWJZSNlAMmT4oUXnEO/F1leUdSCdsDBECTK0d
kuKeRHCTWgXwi8f6xjwDXAEvsgPHTDYhQSZg1Pd4GKUMrfD8P/dbNUGFknMJ96z6QnLKG3MUxS3B
Vl/3TK19OHmlcMhzlVAMlV/QAE8TU26gXfWLJVffIu0Ua9XDnQc444g1bS5EeXP9zeFgUrNtLSfk
25Em4bA5t/qP5Oql596W30DkrtLHVL6zB+QOplX/zrOPz4Z4x3OQ53LP9DredTf0Mf6Kh+lsPRNb
POYsArI3Rf542zb5EsGQ1o/bHxvyE7D6fe3dtQqcn9DUeLjQlDnXNcPa01+VvoYPAVfp16dxIo8b
BWsHV8ZI4Te1uF+VgvNWgc+5Lx7JLZAb3fXfF9HH8RB9M8DWKqPT2nNE2GsICLnuSaz8Ytxp3iN3
emqOIEaJtIF31au4UcsikH/nDsDJmT8Q7yqmpms0uAflhbuC8kM0Uv4/pxEEpQXmukcFLJboI+m8
dJv0vNaGOchU3RYFwqdsyeCo/ZbXos0lrEKXtU31x7uEt3Q8P5WAEDCmDLYXvETj8fDROq8uTRrU
DFjODJ0uxzRbdSzCzxNG4ZRpckJ32VVRKqJyI6hZNwP/LG52lDHsl5Iwg1oXlVRBdmODCnt75G3n
wPTAKXHQPTHTKd022Jl0+iAnHvweQmCguULvVMfrklGJ+CyJXNcK3JAHBt/2GJwQwTk2b/XWnOzw
efCXuVMccyY7LIcxYjwuZCWBli9Er7UrFbZA/+DuLJ3j7b57xrtZKFgwqYngvaErbBxLM0Jv4kFR
U6XE0jQOIWWeS8SD9vyx7c/RPT3n/st0N/zez4uHF7iTr5qs8uvlWtWb3BoAcplRQ/e1Leaeo/MT
T9iwuEEo53GWKLoLmFwvS0+t00weyz7KxVia0H0CTjsBJYaqWV0KBE0y3Y2HXjVFSWdCw69TFs4q
/34vLy6Pd92yWjSreP7vOGIYU02LmNujVYZgvxzdAUqTE3odrP6yDIVItA+56gKaXVyFctCo81GJ
v+2dsjj2VnZNT3NXNvuUhYBbNl1gzk2WYwoKhnRl3Hf0KlZYTi4UiCklatpqUTmG3hyhBjL8EDW1
OujZQNt2hCMNwwLxKLmEVg5zl+FImcOB9f34gLXTD1maaepK6J8JmvaJwYWw+6eEscGHGDjV/yh/
chDJh7aR3cWSajHStlJ/VwaDEeVacp9HXD5I17wxP3m2/Rts2o3TgQDmssCt/WYElEbgOudrxiPv
xvXYmNof1GJFD1zpxHwwNCbUBD1etsvR9z/RKw46W2pUh0Gw2GvmH34XY0Kh6ah4VY0Jpx2wcjIB
DsJyFa2d+8fQ6SENY0AuJv40NltjXuAeSluLSlzt3luwnTBN47VV971+EywuvaJDAVHLQ5iAv0ZA
gbhtXp1abQdNbc89W+vCdl0Gm7HETpWl8c/OL0BxnbPNI8N9VglX6ppF5Lnp1m15iPx8PR8UCBht
VO7+B5UGI8XScL/AXncSjYNBSJQbnFiVfxL07l1mD9EOtSpFTmRyUC9Q/RFtjkU7ErG1shPgAX3B
evEbNWjOkkvDDdbyRAqk60RraMnfG6UVPtxgl5/mfROHWAhl8l/3brl031TUF08A47Sv9WGlvMl7
K1mFyx9H3w7Ae4ksahksSK8dDj3U0sLJmpnmEP9dCQ7xS582xmwq3jCQGBBbWfF+4PpFO0Qv9idt
APmobhDZxmQfKWeY9y+eSCnmjaHIrBY5vwmrjkz0QANLgVlBQaF/8c91tuv3HV6wJN1p+IidzqJV
Amuj2OjcaGr/dMyqidM/duKwfqap9jHSJZqaIxL0esEEfI7ksLhokK1zgBcqHJl78KJxg5hHxRKH
D4e0dFMYtPjunFOtlmbFEmjTgZdhC1z18zHYrM/FZjyM0+SLfoI8FCrp5rWFiI+qE+jxz5hWJCPH
hiF6KMsdizAeUP2LS0qdQlQMMm8m5q8OOvm7MKjT4HXSJsXGTYY7Ve6yISHCllrELx4gSRp2fdmu
MQv6yAlhliwqVb8Y0HRjqii12AnBCylxoVHLufvDuh/bkT4zeGei5NJb/oP11luPFkNoUWC1URLP
4WxQkvETpoBPbQumFm09bbf9EQiVDADeYwka34iumlXYePU4LjgeRLQXAPZ7EovwQnajVxHUPp8h
v3O7Hsqd0msC1XABz86T+2B7OxAk2IpkZ/qkpYPq12R9kRXBANkV6UoOHLYIr/38jUzUjGLz32px
/YikkF9c6I51CwTSBMmhYifon2Nw2/DMwFUeTWg6ABxcRcoUGXhdxVrhR4M+Ltck6J75vslnW3nG
Rd+H+9Zaeh62fzzH5TxpmH8RmTGcgknV5GgcI1SqfThBbDAxS6xYCSEgaOjourFUTU2d1jBKqJPC
oA5huqrQOeLIyDoUkFfJ2U2RiiP8Tq0ruCONJ9kgcsLWXhGyIx6OfGwBGSp2dSxkhgyWf+l7jyYn
HxRPkNpSlAx8SJ8wVS1XW50DBa/p07Tw1jTV7blJU9aYsUsXHqPYJqCvx9w35EcSvJ+3klgZN4m5
0NLk1AGAzA9UxjOA0Ohpb5G4qVAvDxjenl+3M3pgAEzUhv5LvYEmOX89wjb7twCCul0R6O6WdnvO
ufVFBou0NCUfA5CSrvU52uvKdyWclMOVRTrCecXUyXMsQtS84kcqNjeE9XVnGmfns2KMr+3knZ2T
O4BNTAFehpgZYAmh6Xomt/SCAgGkDmAZA3dCXxU2gUfhSMXV1sFO8CKYDx+aeEEAXtjZsdBKpqps
BSNB5QrSZrFlLuBa4vE66/sBr12PV6aHW3cyumVrXfTpfYyulLZPjNgWzlkjTCcN2utr9Yv3XcDP
yy7JCvDGqEJk1bEOhY3/J8catYViLmkyGrB3C7Y3xDrF/w2jSAF/IuiLwOrkrlvgjcKDiE6GFbCw
uIVFbqTU9w+TGMGX0cffn+G0TUO2ie1qrsAP6n58eKT2MONbs9keTHsdz12726GY/DRF4YO7ypGb
UKPBhh80ap4eKPyCbYSMatZNUb3pXI3NGGy3QEV4+SFZxSUs5PA/o6RFWJNRWiF5qG4Vhy3G8zsh
xjDHieQ7aV19k6c6rF2k67P6ME5CGVcghIDISzTh4JVtobDR/LoitNN7TW0zkAkmj1YjdmgFuc/e
dykPH8BjXf+/XBSOI6zrKmLpoLLMV/4rirwPY2wmVkOe14BnqrO/8FQH4jsNXeI+bTVAqKKIaqDh
Dd3T2gR0s2VVhO4gQkWlFYOQA7hVcJRtxASj6S5dl1S+pWoMfilzgQ6xBz8PWsgA+Tu1X3Cv6YQT
MjB/pvTyYKBMXH1TJM9ZKFUreRPMv9DC97fRsV9jgXKudr6EqUhTh/vxoFwGOVS3o3q6B0GuT2zh
Zu7WM8YdhEHYCoeT3PUh3ygGj2y2x5++9Hrtg/CElYUJ+ZA49DF+/+Irrlb5+5mOM7OouAsJZaeD
h2GEDYXjKlvtM9NIm+lc2ClgfVk42FZJD4xPAapBSjdIMHPYN0iy1CBbmTPuYFIvYVTlOLrQnz9K
FeOcGVo8QEURVJhjlj8qTaXfzwETLS1SGAFmr++gmhTWG5Z3kVJNgxIKy+nQT3Kayl8K2s8M+wMf
vlZdFKYEAypbtUkn76dOo4we00B8AMCTvXCIr9DiBoWUv7312en22wbdp4oRjHx4i+RIchURqhRJ
7GfOaAa+tmvhd+b2ZxfjO9MCDHoY9xzq7B1JR+dOph4jP+H6Ly1gV0DN2eRDVHUG11xWfQw3Nzso
SAfKJGopEqxvGZSYyoH0hZxJrBG7LxqiR5T+rHTJzivNxD2oIpIK5yZ4GIydl6x6kqXl90SOuyQ2
GThAXxD3pz/2b9/932RHnB/EO7IOg4HWCFmeUQ+ZH8xG6Qtx1izukqCDGk7emzJ44zuHz3MYYQnD
R1HBZKfIeARAU5VdzShBqWfY+FiVZrysDG/F4iiJVt3RT4UY8f3RkyQewCahR5smqi8vXZit/BD7
17D2Jt0sWNz+/wqskLDcqbljfK5Fv/AHcD+BgBvNiNqK16+8vjhfsaQuKjCoQNqyeX9P+5OfFgwM
XK50XnF/cRh+UjJq2QN6xztK8z4Yi7GRPB0bci/Ds5zBSJNWRwzXdqzY1BlCJdYkI8hIeIY1fB54
ZwTVfaCAk5n1fxL773+BB1lHsR0bZNldsNF6iM8jcrhtdn2fQgCfcegO6Ttk7Jqhj4LesO06rU9v
f5KQkPIztGLFq8zsJDkC6ORSAfp1aKf3Al6ajUVOsDQzEH7PGUqk/oDXDVFZLGUpG0hEwrssXdr9
PH90ZcQOJfzdbI+RAZouoKBdtDQJGmt2sErZBaKYIGCpsiB0JGpiVm9A8VU67fukQESbDBhXRMn/
MqLS2TKkdCthnjoFToxn6C16X8bAiTR3ZBlvkdbGGS50WV/4BMaAgD99CcRhJrXCiNOMr9T+4Zcd
BmwAQOa7HdQvmWkP8NSEmD4EDJalTqhVIOsvZLumTwuJ8/TFODfQ6CCphFQ6W7QoUrrUkrgGOzvL
3UXHpXdh1akJv76DOYC4i1SoA9xsvi6m9sDXzNoXClPZMgrkX4W1VID9XuHNCY28NnzOOYyVx0p7
n60blduD54OxicoPAgZodx+L24CZ0vlIlhNCEnAk4zCgeFCsqusrLBc6qI04mPhKIve4iN088qe+
MpQh/9mOoqN9qrP+m1pspO1IxMJLg+cMjQ/7xIYhJLZ1kW/SOAS7tL2nXiYFUvhIvInWye9++Tp2
GcyDmuN8epcBFgYULCIClGANVLMmxEYqr5VJxRcchsB5/ABGyMe6v+T+4YG/4pVm6+h9C6ttBVcp
TxJa04c27Hq/xvMGp1tqLUaWD4qSoyaoMQ4bXNpBRZNUiWUUbq6PmMSJ1DudUOt899/asWCGr/4M
1aDeF69YJzaOLmyoTAOR8GFlN9xXR7aSS9py+Zi8HTWKuanJUDWAVRpXwYgXTxdH4Ub8DYNvKMCA
yrf0oLqJk27Fce6AdoXJC+96+2mdX42NhQX3LLNZlpdX/EgU4Cd6vUPdL6fVDwq/Q32a4++5TlT+
UBpw0GsvqXJsU0+SPfpJLFMvr02lkRLfWGZvfQInaYs6PY4ltDW5Zjz+h1Rqvsifdu2OLL/8Gxal
5URak0G82/cmyxEEvmKQUobp72+Vu88Dj1qYSQpbxCOS63XfIkjuk/uJM+p/OKIM9EoxcWc6KnRG
kGDFXI4fz5urpBMSEVtLSdLMCyXVaZ2+8N+VErc2F3jcdtrN9hxIN0sVh3amKGJWWDCIvW3he0lw
zMdZFm7mRVgWqvCu99+z6ClMH4B0SjIDu4gPws6fkCy5ZNRagxXZn+ottM6eXQGWhfy1JaYyCOOQ
YvZESsezZAF0pMts7LkAJVuXDkM6gdm4R2sjvBzTXOGv15uv29e08Si8+KwZDFFd/pakzKITZWHo
8uZeAFfVkt47OBKBbRFuQjAcBbGZiOspQid/4ZRaLSmZ7BVuT205DSSoZTV/ur0FXUsxOXGNosuf
NXbfatk0c4nKp5WW3tVkTVjqnaqNRGGQzAdvVJKiKe+gpz0KUy7U6LcOoAv4aV7EO2hzF9wOpSo+
ZnwL6aAxthIr2YBLZTP/3ZOuecypVenXkceGnhLgqzfrM+E57lhqvZ/KCdoCaUwy0gqdVjinTUDW
2eA7fuRjph1s+oDz53PnGMai0c7QYff9feox1yERzRDSqc84b9NfKqFRKgZNHrbCOlNe72SMFgQ/
b0FD2Eem4Is5cgYe9kMchH52SCbVdb2RCeqEpGzFQVOjnrrrjhob1VxlHHXqMwUJ1q/3G+um+cBV
h2GdRRjpw70H6vIoDDUJR+ndx80HBdrEnf5OJtI51bB+cZgt36gvcKxcwiojnrjX5uicTTYCVz8b
UfYP3kDemeOywYnB3xxbGccU0PwXh4S/z3swVA6d7zFhQIkcs0ggv9oHs387pv4ckrrAjvXgfsJX
nScrYlBKoXosjrUkEqImNeFa61DwzG8L0upnf4iq559nQvH947ZnfXbg3skZ6/Yj2gt/5CXOXCBY
HY1QrN2yKizkuHPSEXFbYKBhQY/09J1rTdTFMDRMiaSRSjPcWlwVjIWizRe26K39yS/P7lv/OwTt
MJl/VBRLnPfPsGUvV58fb1mZKgtpWzUIGTOhnqFHbhWSGJ7EWfBbrAfNZyC64tqgUrw5Wm3wPObH
j9ZYti/7nQd9HXk0LJAX3B164PpBDQujWlGudEAfJlDn3RVA0vq3csRkK4fhRv3Ss+YC3GDg/Gno
WwYNmTp64i5PoFZuPkNTIw7JtYVuzI7dC5A7ZnQdB5KquLRnRuDRlfKSBhPZJrwFMa1Js5oUM/9f
m6Lj3RV68/Rj8QklwF9FxrQs4hL/zP2ktgyTNmzHV95sx3ZOeDjKwGeICBVsNbWP/DT5H7vfrFQW
OoOxiB06MmujFE27t+wpaF1i6g9vHm2L614Ba1IUn9kZ4XW2gUChYltcLd6iYCw56LVPTvUnenBf
fJkTO56CYA72G08WFt8uuyCxjsBxlIiKsQvHmEs32HsW8KCeRxk0XgcmeaxLZ/Mm3/F+qu2uwCv8
vlWbCHnxn8bBkbvolirxGBs083Uee3gfU0ZF5SI1KgiM2vytIIT+bsxfHSZunrqJiSZlz5o0kVEF
8QBkryfDQNCCbCNWWE/DkjvMrRfGnc9T4ca4AJ2rVIeqkjkObTN+NhhcVvNalKPkW7zy3GnA55Fy
ZvRaLjTqXLks1+lYMyNuL0bvgF8u8mPRdUcP0vUrSehZOzgIXh01d9TXnXEaAmnaP0cFNE54n8rl
6wehmtvkoBKrSrN7imApVu5qwTSnuHwCH6xbN7S+ViuTRecuzfIUJfNM1QIXTYlF7s0l2A/oOJR4
EqUpLf3w6+awyPbgh6PQd/I1eIb/VvdABrpyWXoDmoz2Z8aU7EE0A5vw0BPlvjL0oQPo+uDvCetZ
ByOOX2hxhMkr0+TjSNShIHbUCQ5dMDhxh8oXItKgc9qy0ZEPvuT3D7BT8ESs8/e419qHs6s5qM9A
G1nuYV2sTQbFuCpnc1Xb8/DBua8vfkQkFvfv3sFJEGwk71doyaWCSlDxr1zz7q9/NFGiGrHiGoFi
jrMleYQ/WzRnImjXUeL46lkl82Y/fm6TMFwuTmzT2ZQQ20JaxLUmU8eL+gEMjlhtZHZeHuOI7e8l
0qpKyGE9+Ml1ImrmKkBX7CDyGcBVfzU0HK1aW6RLuzw5CzoUrsL8pybx0w+Ipkb13zp+XvINGdNv
lheuJxeUtmZfJQvPh6CSfh83HllGwdlh7im9U0TGiWavHk2F0KFOgAIhxqWT0M22YxnPFG2JIHyV
ASviWRal6BKga76LanUYiAOnVcRzomGr3dT+y0ryf6+NxEsujSAELJL1tg1n6SfR7GI6ZuAPTZg9
57BOEdcLRqqPqoOdtMEpohMm+q0MbJ1gIM037VqyFvIf0CLKyNH1wD03xY3t41G7eyR4gHrf8bj6
+ZdAU0kM+eTPFTACHeHhNXjAEUzuSroZw6RqxwWL4SKl1z9UnlMOnMvYOMZKZCQ0ig1OM45JWFHt
RhU14gfw8l0IVjmBLdFECwA3wwDVTGy1JWGYkZs0UPyQ9YynN/mldFA4XO1SSzW018xDNXbOG8vk
DMy0U1mESlpEiU9qtK/M1N+Jvpm7+P3mG2n7o9HemJmCXzI9Q7Jq9bcEAIxMkmgjPGvF2BNodXXL
LTFJcCaWbZ8sPsBN+sO3AVwulQHYErq7e3fdMyThaFJEG8BAhmzkLJHYqvlVhZUmvfKPllD7hcHm
GAcQ8A8wpSuHBf6LAK15geNVIXSmZ3H7n+G5XU9CIWL7BO2F3L97iVo1a7AZOJTM+sa7tsmWcpoP
mB9J+Axk+QANt/2kVkum4AIgnYdITdSOuwOMy+pG9IPwPb/yHfgZbuHbOplIbac2cOy1EUsjj7pm
RsroFfBZUcg88cuHcn4oV+FmR3InXw1Z5sBMldBorFxdK8wrAgGHAiUlNJd8hP+S1G9rtdPM5E3/
rjWEW2fyOpu/UFoRqOJ9vTAuljXFRvbTEIBYNjoHgGXXO+9a+C/PktUI8ZeuOaf52aqCTq5rI1XC
3Q7gh90PpSALgm8SniJURxpabwkTbfF5Cd3VBhRlQzSi631QK4tac5ACleuqlmhwlDmr6kXrKD2T
H0ilMLEiIkRrYjIiCY6fFTqVtpsx6JCm+NauH/biFE9+cLtIh8AmFHMVEeFsMmxSFrLSeVBGKBIM
Jxm+FGEReJl7AsTwblY2D1niJ0KN9NkrXiWSmyPCYCHumxltqS5QOi9wJSc2pnc1aEpA3g2beMfG
/lVSDcSiusH61tiO4gEZokaUNP8RgT5RzFTL6fUGVPaNTxvYf7Aq+lKQIeLgu8xv6Dr48gjpJwWo
SwvlKNVUS8rX4CB7FbPzgLO3yAPjcJiPXw+TfoUqTyIh6TRs70ShooTwPhUjndRJbjFnVojnt2fE
ERhgrdsxGeQXhZsJNl245R8375W4BPe7ihF89pTkgmXQdDgiSs7knkpRz3l4jdUxOh+yew0VZ5FY
bpw8PfkJ/NlMLE6mWlU6GPkhH6rwQ0uZpeAIPWRMzrs7+pBTI3BN7ch76/b+SYMLoNEZOWk0f6Hy
Qo62nRmwhdTlxwv0+mgtBQVnY4W72JoTTt75xKfuVnZo8V0pC/5Bg4MbA/fSorVt97Zsy5TFfZyK
h1W0vwVwpimP622o2Z3/rjaRWvRj6sbiS3QBfalgK+ldxBIvn0vMgG+VUNDlRBHmC2ppknrM+qoA
p3IkSzdGaO8FOnTnSDh6g9dPihRcUvm1ZugFJ2+GPWQt+7x2f1Qjc3jDi+y1if0Wg6GbP5PeXUDp
jwzHqsU9z9POWhF/K9PxO7mB0iwLdtuStANN6NRLSTcLUgUcWvdtzXMSxLYs9cvv4kjTMa6BgzPV
m647WmuTKTwjeEMsRHp6lDMAwgQexl7HAUT2CSBr9tNWMQfpuUx9HoxXVgTWMLNzfxa6ZIpEibKx
qtmqpLP4LiyPXB/dqnHZ8yFCfrLiewBj7I/YC0KlebIWcyIJF3kJOCcM2zpytb4+4S5v2GrZHkZ9
3pWT9pTGUiEJUhdTj/h9VE07UBdHBoF6LHl4gqzs0nMFL4ukRKKruWyaT3+YyiEPqNwT0SfXuy5l
iH7/W8tJjB74qlAImO7ZAYsPG7KyF1L2ba7R9WyJ8Vm2YKtJqOH+D3PwzPOrGP14DNcm5h8l7xNR
bJVayLMOz7W0HY9S8wFP3JhHQLIu434tlb8kHNVWz4KPWkikOUNRQY7yOp/bm6YLJLAfjq60f5Jc
o3pzzWvctr64mjST51J8B7rEwUnwPsn4mGB6HMghNL6/Jfaylg5j4zYhB912z36HP7giTvbXiGu7
jjYFSpI/4yJhz2CPRo9KHlFZ6GLockN8z5Udn7kk0pr7AadqkyebcAXmUSh8H/N3phG99o3qI7VM
D+fT4NzUqpQ7yz/OIYTtMFNYUxyPIS1jYm+xV7hJis6C0CYWngq0dUhs4k7olOYXY3ywAuTPJvQ9
kCYEhGf6cmQCsp4INBJAbawLva8IMjSC9nSvKADyQarKhtcj4MOA2SUrSWFEbWYrhosj0RLUcpcw
8WikkXi25MgW5JDd4HPQ8lRG7P59ZwReb22J/3K2kKi1gn03n2ZsH37bRHIZS4EWwlFjqKlmunmz
e1VPqSTAmOfl7jCV+H5RY7rkyv0nzAy8nK/al5xZfOmE/oXQGpMXYPRxD4QhEYizn3agM8ENlK08
FYe9rvB3PWdzrzIsZzj+W398cm3vzO5BOCqxe/xWS42WDvAKjaMSEb1huHncTH0qBuwgh0nDsqYH
Uylvo/NqfLdbTxLhiQywcw/QOAW87s+eAROqKbdeR2x+D3IEUr+z85hCrKHme2iakeNGhYPvJ3lq
FJvgmWVQiurPLOP9ScJ/2w5RHUKzHoExgaP8wWHgdSKgmk/as6utn3sEFZS8lhfqpg8u+oBWX7DC
hdmoULJLI6fQx18cyg77cZS0xjnccJUkz/VL8PTCOk5GYjohmSs6i8yHt1MZ72cTHxtVW3zYaJ7Y
9le6VgAHPGLlQE8bsRZweo9gi/e4dBNmvsejznoKdu+L0hLtQYkLDQ05FXYxhc9bamJAtP+aQ1NN
wDdZVnB2HMjrZeNUrPPYDsm7nbMmboyS8ZlBxGEBOySZHsBZM+fBfWM0JGbH1Qp/IGy9Q+UrOqLC
stTMCSSEjebFCJ8BAeu62XYlllya9WB+cHje3JH35sZO6rkAaImEXf1SZacEX5ETAAivh1x/QfTS
9fAV6qjaBsxr4YjO5/+gzIhDlEf2WDOnJSsakDGDo5BJbx1Rc+JWPptMWqM7bQeqgdahkRC5ZU3i
2W7KODPysl6mWDrEKicsARw8nC02gqZAHxa4iLg0prST395H2U18Ym1I5RliTwyv6sUNHXnjfM4P
aQfOtWbkfwco4ZShKDPMhv6IDWwJGn8AzURBxsrrT/5NG/8EYj5DOpjaCnETga8/g5fR6xzYdjgj
YG2RRoxUGb5Y1qJWu+CqjbaMH6w/lYucdqn3EefLpv06kNJNl7KYXPU2r7t06ZQ8C9ZqMarqYAy3
+8Vx3B4m+Q3ITOvuOaYOjPZ1ohoozeQ6tVqhuQdwhapzASwDEHxKlTQXGijl58BF8xvtQEdXSk7f
JjOYgtk/gdVGlxjK2uYbfBm1MN+GETiGSdxkMSxUnVPnVMo4EBnK6izjdNlFk+aWsN5RPZgFBYYH
lXcM9Md3HNDik/5buJcLqsoa/vSob2+I35lDx/ogKkedQz8Md/od1Fqlv04/O1J6PHujE8sAyID1
9E3y+Xg/ubLWG8wOWXFhyLOlWJKmHSl8i6LOMWtjcxAv2omXr9kJHc/wleVpixtrS2roMhYdopVq
eNvcZC/QqMScj0K3IXEgRb0tThKSbST7fJyyW5dVDsVOVumU8ApkrQxi3cMjxs5Ywih8oI7BlxnS
6QEYYUfQoxjVkGUehmgIvsYiLEKIeXLGuVbF+Vg0vsJZhHPpSbrtR3AbWM6Qkm9Ts0H1+IeuWjiO
AJcu6sV89cLVhoGWZrRi+FTl6yOsz0qKlqYgVi93vf1472yM28WPqkiqjMqbgHGOOZBpCxfqcvf+
jhA1QiIqRXXoT8AaEKQeQXbBtTmRRnHfRF9M/xMkOLpgVR74AAKDVFOjy0U1J16dqSaoCGHSHQLQ
+wj47WRAQHgSXEcmfNad8yu1YngJxXVKgxOx99ipVZEqETCsprTxnF3CRoqo9QQIK/zcAipUlu2f
kQbXP1dqYgCsQz+CSnt7Buj0eew/tEDzO2xJBFsc24PiKTv19+w/mVUDPaNzDqFG98VteC0jNPkG
oWXHVUPJVvOyFzsdpyrco2SLjR3jmnMpsXdaoPLBOyv1GY8mriUa2ZpQwl4L6KetyfbMLC9i6Gen
Kzjy6NnPIHYuVsH7tiMf0TekPPxEdwXA5rYpnPy+CGfQbcc8ckjRo5SyqwogIT323uBSmOeGSxKt
hqGzIyiN7yMlOEds1UU5Tttm7Hdtx+X/crHpPS9OCyd/0bbWBdkrt0SqpYkMvm938eEt2Vc6kXEr
ceUPppjQexpyiRjHWVe+GOdvDEbp0syArbjHE733fWh/penwnNKQUB3y+enw4/NxvJQIrFC65D2g
QUQGNizNdPJTmdflPwEbHu804DJ/3O6ayokCgioUySkySznObBJx9j+uk+ppgDZHcfFpHGV2AAb/
Or1XhzJ4b0lijOR2zMvksGcbVHAxHgMdKM5zKtk7Vnx68BUa14e6ztKuzZuzSH+ea2AYqxqpJrY0
tuD0xx3zUuswTvGL5zCI1Is3WTqkyM3PNolKTFH3T32K//xKFZ/R5ZMHOxqT7ZEM0nHHvzV81/iN
xnQBZyBgXpu2CdNyvvKmFi6/lCA5giKmWQHB+S4nBlJWaqAcAvL1TMK5sG3gGZBv9qfeswqcaQVS
F73FOzMLqV047HpexaqVFz902U0sMCTs6RFeMaJTqajAdX3Rvf+86gfMw5GOw3t+59K6+dd/GSNY
nXX3HjE/EQZQ2LoZ3zz2wlWUN8ZsmuGuuV5W8XGzd1JyRjFMyEIKiM860RJ5TBdhshy3sMIxuPBM
375vy4CaKNxMmTajuCUrmyNV0jJ1fwdZYQe2FAEPMw4rvrIhvLRmIRVrlfsS1gyj0YO8Py/4qUDa
MhrCP6a257QEly6Y0VXh/iXitLl7Fs6aVM6D32PpRkszgGRUoeAw7nhv+hKxEu5uRoQOH39nZbkk
lEnAn33N+OrepYacqXLHma/qe1d5/PFuU8On0BXFicaZ5loPHXUD/J7SAs64Dh0OpmrB48iR15E1
o9JD3AQhLqeC+ns1pZMN7QWKXGD/ty26P74bn1D0R2bhOqEwrpmBUIut+MFdL1j+cfjElj/Cpj9H
/MXsQbnDEbGr4ZG13C3ILKpPGEeZqHiktk8tfHeeNw+FALgj/PLrYXd/tYF85X/d5UhTsveI0oSA
e8BdGpc8Xnc4y1fVgzI7c+y5RBUqLnUIGTmEVMZUsIQqf8KocpCVa9U+SsRkoX1cVkGUTUv3YF2g
wEOn0oDiqw6qg0JISmstrAMtd2eV1UnlS4ADHJbM52JlUi1RhKeph4r9xJ+87FOrTIBMGceIhQ8M
oag2LxOh8w5fV2d/iCxvaf3/BHZBWejyWj1CQX8pb0tpSTRFbUhm3vmBi8aLNTJvIzS23/Mzda5a
AxvbND28WstEdlnQ5eLSTRMz0QzcqB+HYrp4TE7Tr38hT14JC/oyRg70Ngnw9IWbBs1X6r/jzsbf
pQL+Yr8UuqaS8W5F8WKRAYq5KMvxgfFamgDLiTAlJ8izJdnsNwv9bqBlRPq3NR7Iatvtvwmedl6B
SAzTr33XY2rp6bME8lPXzleavm7XIMIk0Mf2Cr0lF3ppaUjTzwLne9zKOAAK4NyzHLQf9xUy82xq
b4/fRl1fZ0tx/Jh3PaoRTXg5RzIHMsFYny2xcYaSLZLkmiar9Ix8WhKC5Q1qcWscVDM1yE3ypXjH
EygAxsVntAdvBBxMJ2fz8N3eolwpijovC0bTZsHxzTdcud2V/1iyWTFvO4CeZg07XVH1TqbbJ2LQ
+tTpSK7UYiQaQu/cYK9SpixghfGBL069S0y47Uki2WJAN8Q4hcjbOO5zFsP4pEuorngKRDhdFW4k
L8Z1nvGU4ZLxRp2/6fndjbB3LUvaDipmZym8U5V+M+JyjuXD9UWdiQmEnX4HS3u1d1SmEVtMGbOf
UMvQstHA6md1r3pUWA6dR/j3f/+d/r+TOwMzfSocPaKEPLOpUeq1VaNgEwLLKfqcZPrBcJKpMLBq
HEwUdmiMbXUHPZ9Q36R/s5xDbvFMX9FoDUMKKnkAgaAMgTq5bwLiY/dcq4whTFo4CgEOe6fq7EZr
DTjEsyhnVWTx4HTCDM8Cp6jJjOFUm65n/aLbqmxaMVqWLOqV8jbQmXSKb32CnDVItdJnD+vBZ8gd
svZVQX8Ss2C4ZDlh2qtoWD7Jq1201JSh2bZWwh4LFVa2Ax9tWA29nzKQzooW6xFT3TGM4WFnRJBX
px3F7JNKDCSMo1y4+iJ75I8ThIWO/DTJW6GI2OXSa3Y5Zj2r88dXJssN3VV0uwgHtpxr2vch/2d3
gK9puLhclb+JcSBgYUix/uzzZoSz9tj1QQxnYtD3YJI+ju6r4wCT8jG/w7YOTxPr14KbN1Jl6Awb
VRkwCUbBuHE6ey9ORyFoPbgSHhTGK0w2ekfSbp8PkBX+kRrQOuXp1IN24GPFsZDG/6olfqw1wGK+
cO8Z2bMVfaD6yekKav2rCh9MOFXJXCA/Vf8z5H3A5nrpGthqBZjnvt6/4lBktCt81ZHERQjGBbS9
g/ODv0dlSLyH01cXf4GYBii5XEwY0F5oDCc5OaQw6hyoc+ibRbojv8mjx7X8hO9erHmOWva661EF
gqvWbDfao/b8cVuUUwtq6ySUevY4Cg6xpPuAJrZCrxSs1TUA5nrAL6wFKYuHBCShlwi9i4kRWTjq
XxH8l+2pKwFjBgKa282W/HzJDgn9tWRyTwuCRWaM/9R1dHMM8S08L7zuZVlejkKk4mJbPtXxYOD/
+rQdI7YC5CQ7BG8h5kx7GPiXKj3SaY1dKHzjszCUAa6quOSg+Z8Q2naFJ/LHDj9+3WiA9Eo78hO1
DCmpskc1Bfobd6HCX/rdbJNYS+o3jRfeN4OU/n7uS6qrQhzR0yzXdqn+eUk5z+ysMOqbR5Ab4S5i
c7kNOH/Wk/ybgQDbM4SPTNf2a9bs5NDsESnKZMc5VH8LcBuay2aLHvc6sbhFMYIqrtx1L7w7ixx3
t7/47iXC8OMYdFkYxlG8NhGGsU4KARQbzL3kdh4fBrJwDV/T1GNXfmekpgBLz2mPi1fbj70NO+U2
JfH1JWNwKbxAWyd+7jrRnDJhHAwknmAdzaXDN7BdaoaFdzDVqNdlKxIncUx9BLCdD9JUun7DWXY2
wgRCkfZ2P+vjMvoOZ+GmUt7IOmWcrrm8oHx7zEeGi/8GsBKmOhGJMqtXN8xYoOglfEXbDa4jww1j
PmgJLYh5kXk47vzMVzuwyVu5/nKtlr/GqPWIXuzLB8PxImIG55UA7mxqY6Hbgb5YqiOIkkMx88pg
8+DN7OBWFxJqLyQZ1dI7IHrtqFRbuOD835inpdtwYMmkRCCzD8a55ZLxF62Wxx/I8T+c7yoKHWyf
p/3fMN7VLAtGOYmyP9PKHS/xjPRH9nc84Dhe4zDHWLwHyICUL8Ep+Djr8cz9ube1n4evnNrpuA3P
pqKbdn3A8/DOUAHs3XXFUyJAn103tVWEeqU9ZQjJWH9JgMvsmamJ4rUwa8MIRFSe930o282fMaGk
SrUKsy2ZrEOFxu62/KMQwbtolwxrWkgvYlI0ZJfo8mTBHumB93L5tBH1ebaPI5Ue7TF+T8PdJ2TV
+n8Psm/LqbNVL02HCMxi7cv6DCqU/PWUgUyLCgR/z+gfJrF2eti0zj4IKyDEirnP/oJMkRwLWI+8
+jWXjmnLNyl4QhGUaMbXWocdIq+RplAUUKtoSDSvMIru3rdQUR/64orY7K8BnY0diyTu3QM62MWk
aSc6C6we2jT4qZ5zpYyJQNNRSwpJdpaS0qJ/lFhsw2s68Txtz/PQCRzuQO10l7vnoxv/qhoR051K
f+llo9AAa0dBviK1xDnKiN8xO0F03+4hvfHSQtvLxjzW3FgW/XO99UfbeXcPo6KppHkiUy1IVMf6
MO1hRokcwnvIp8sl3Wk/RpSS9tDjJcLJdOo8d72woZlSK9Ol2AXQTnU4UtHk3I2VU32iIBWqOpm/
XCw0GzffBtmKXXGRmOi2x+JPXrHvj4NOVDue/Q944bXb7AEln7PyVqpA6zR7sn6vDz+KicSwrLZN
kaUbvXmzlBefHKWlJqEFLWaNFSS9+fPhIjvqFXks3w2g1ydjzLCVi9tCQaoO6vgAnXvkSiOnCM4w
4ops8Rk+ybhvTwqv/YPbd/RMpbcm+5VHMsyO+t8PfAd0s1GvcKpX4graG0OuFvrzmkfwQnjbpQlc
+8CfNlShyTHBjB3K8bX5xKnv6pg78lK7EbmOYwpjRFId5/FSVZoEGw0wvs0bJ7hkGMTSGvHuKehw
iewoc44jPvX6HmOLFpwiuf5YoYG6l8ckm71nt+A6dKg+iI8Km8KsLDK0zMvsOoGAVJRakjVW6YW3
Whc+xeIGxPZwrkdvBDGNlfZsmrXfPIJIt1aB36eHDNWaI8GDNkNUl+DUaSG48Qjehe7rXCBi6LTT
DTlRCtaH1CytB5g67WoqC8u3hDEGmd/ja3kUYE9OEE5ugbR626MhD4UQlysg6diOvIMmonmB6l3O
ger/KoU4yz4J+UxoouYqq1rz0ymSIvmBJEPesCc8ZyIjfKEyruAmHUQlASFsRkWEptOo10qn4VM7
sAGNu/+7WhAcXhG43NRCvAHVBEiCJFrBPqCMTU7/b6fglTyPjOs3qfVdOCP3SGQNAuOf3Y2AyS/K
e7DqwsaXifoeQHLwnTjasxrO4u/j48BkCzp2Vk2k2YGR6LFTqB1LwpWFKteLk4aq4w/6rRXjq4cG
x/m8ATmElb6C0glUsw1akRU/o27DOjSzGEQRLMddW6HRmXXmoa6ha1iU5o6SiiQ1YGFZh91VUjET
XosF0zaUz6O8qrTmkxehNnzNGdlazFRUSuQsCRMCbXDA+bQ8+a+1AS8zPbBCbZbe0AQTlwHFtO42
DRr0lmAlqRz9OjSAhrV+wlyLjLN3NvqGQIC6R4zQr225kL3/qmXwvuXMulj2RIPpRdwQJ2dQyMjM
AfmOaxUuGl2ZIH0XPpGKUCh/O9paM0/pzTxYNfvkxPKKiqpAHqtTGjGgpqYEoCOktIccC9ZNYRQ2
d0VM69fE4ddpb+Hf3G893p4TkFiM1Ve8LIg81Y6XO7sglyaqpY5r4B7VC3V1tpRj41yIK9Vpnc91
u9QNE4TDJRs3rzh6kv8PeX+fciE/eY+c+KPcOx1noy/lf0WCoG6iFhQkJ8FfDIObBRJfIt9bau3R
lTXDuDD67CTOIAKj3A4q+Z+DdEPDAFoC3KtD/Mo7jsP6kExkwwhPYyGOzOx7lFtv6WliHijH30CU
HtWb9LuDuVtSPyzXpadbdWF096YdHcy7ekw9vq+ZtlB23vyyEzD+yJGNIZBa3myXWx4nBeOEaYOa
BcTMTVNLTLok6fKDpXkSiWkh7Ga3Bzk5pJKX1oqyrcFLiUeuVvzwMUTfVgl8ZUCzmh9kW+BLTyRD
HZDcIepEMZrWzO43IyI6ApnzcswomAn2aZZ+qen6JTcxHxc+sZNVxfT/b8t62wGsF+FlLSP7zQfP
TbLRtazBA+7rOGfD3GPSPzFZwaJVXLEavFXhq3/acDhz5sVapt8noy6jmoYumtfoBSjCdJ82RpV+
w+62f3HJZOQQS85HuCM05XTI5Sj1K4dWCeS6+UUJ0as5Kcp8spm7POrInj6iLAJwCNge4ACrD4lK
Ex2S9Yc2GZl5Q5j0SQYbefdU7zgXEjKr4udKFMvUaQAKJt+y9usIvVSLo4MCmZkO5t7Krn7RQMTC
S6ivX8tkzeLloLTK6bk6kAADLIMOGiEhCuTj25lnPNLL11tWxgpiBNRAavHao/gGUIyI1X4QfbUp
e8ZtddiiW++vbXJc6flwUWCvg794DDP6wMT6Kg+gDbjL4UDuDbEycPFkODPPxmh9eAdBIw76t84K
6xJzMSWDmNMRc5D6E6agnXJ2dRgsbWfrfMJrMlg46jthgw7nppwup+3hgjW6fNF0A7kwxwA4ItUh
lHbi/3ZXwUyrEbdNFgZtZhE1julOL4BDb5EdI4ThfqW0YeyKHP6HjRX5bLKwbGDEV+L93RUW4oyk
/TobSCznIyk4oPAOUGuoaZj88r7CoJO9DYdWyR2N+pmScIhrMlK6bkzZBBHbfzY3zK3kMo2VQMH6
zT7IbSh+EOvUAmL/pcW1tUQU3cG1bXR/gZ3y112ISeEDHyaYTAOuLnqFXcBlOY9JBVKcZiOWfqvI
Fz3Mtq46YHqPuXAoKuvX2k9Sl5HBnYevzfTNd2wcFZ7F9zbvXxD5fpXPcedl2o8Me3bwTkA3q+SH
Z1TgSGdc1sd+C4MGS5FGXiyzuQ5CBgkBY6XY7N9h/UM4U+K2EKiktDLgOrQsUM+mcDenWChDeNMF
IJiqkDig8ZyFYRJqWIXPmm5wNEzBsyHaOB+3sSPeAjVY3vsqvd5YsuYJKfu1aWhIE+cCMwt2RZtQ
n4ThaxltLRM/yYxLL7dUFUQh6DROvFhnhCOLvwBjlsCPNBwlBMEGfzI6q2f4HJ/bakA4rnajUt9s
f1kf4cgvrHkoocl6wIx3ZX6BKMrmaFItrWle595pcF3sn/yxi2tNKcSxBmQGmQ0ojcu+A08Ocav3
HezhPGeD00s1XN6og59PNtybm3AtHovlaKpRrGuDG5I73c/P1MWRmy/LsS5fpQN/jdEUpUfvV8VY
ZSkr2r79DAcRS0yr28kMlWJb5TMuobKA3hFtg4uBZChomXrZsIKTqyqk/s5dx3ZRmfffqJ+6b70K
sy6lzlVC5Apdy0+6m/+VG7//GgqiAXhfeC20yKdEGPRoGXL/GZXtaa/BAfYdSdtPnxSzD045T2F4
CLbPfDypojA5EB/0HMz0mLfwbnlmPCiJQQznNpUnm7gnfQzf/vXeIkeIctS3Py9mDub73ptkEhf2
M6Qx1ZBVBlEkJXNQJIWT6SJuDObwuw00aBqBc6Zfzxw9D1tF0WPLd9ZviBXKuk2OCVKT8GhK7PVf
PO1zkviSTo6bfZW/Nh/smijwg59IiNMSaRfgFRhREkdbM89wtF+mYWCn68YA241+TfdU9FAANap3
GeQCds8Sek5WZcW+pj0PsUNyW6jsUu1ID52z0Qi3VIpWtT3QfwHGYeq4WlEZ9BKT41aWX4d4tIcj
U9nCaBktRUVvA2jOAwZAgt8lnQlwmO+NCdzpdbQpLXK4WZzsUo0mLW4uwmVXXbj1f7Q6viI8wWIp
DlNLUwbBAl5AbA+R6kiwCcduppfTeL3pXAZimnEljMZ3naMQb21DkyYWXwhN8uan1OGjTdo96Wrd
yHuDCVKmJ31Z62xnpN35Xvyuup7Mc9hKs1VSwt+9fvnu+Ios0McEwqfdO8ugVA/d7NjEuyF5TwIM
F1vZOg7YMLvQPqz1FHVsrv8DFI06qQqCW8+US4nkYSehYvFukREK2C25it0TILGok0EvndZLFhFc
1oSoEmEedeRwBOqnpkcdlNW2SnXc/xwzyUhEJ+ZDUiUEt/Nn7n/k8CiolvKfy1iVyZW6hO78PhYD
WJDNfFtrDHLz8aII+o8cHCifyBlR4GzlIKLDm7GkCASLB61qcFvjgqyyg5DXn3fqKtC3Wrr3KKtF
i8arH79y5izt2QJu0rAg4CBvzi9/TNjN04elUheKFQGm64vH0BwIiNke/62hUFejYHMHKIxwjK44
zPW3Qq0XXFWySNY1Re8Px806Dhr+ZO8pPkDoxczIYVrInoUsVmEE7Rb4GCVcqvoKAoXV7KUDEZZ9
MJ426B49CYobMm4m/azYaj7XAfF7q5Od38olvZQL8KKr+04nxUy5gmEb+xJybtrKbceOctyylCrz
0CN8Rnl4NhE04ahVcaXCGZ9jiusWbtFWn5DGXQt0d7zHZrxbRMp+s6qpAhql9YFkw3sQSZUTw8v7
Wdi0z4nVWbqsBAEzV1yqNkBce4OEIhUivbSJG7DLJObDknE+B7wQn+0hpVId2kn8nUMzlfHqrlet
/K48f8anekxbUmv0yxcynIbS53kQY7SKe6o82MyCvGjlXAo0qW20lN6iSLx46fDcEFwz1/2XPs3N
bxw8bUwxlkzuJZYd0km2ZKbcGDXNhILj10CrM5P9WSF1Oa/fyFOE7+ICGhrkufkENPmJg1BBVQzU
Dpxo92hR1HgZXHZ5kTZU1DKykyuZdaj25vBjb95n5ZXZ5cUIGM3rgUlOWgnzuyBJiIWglpQvSDJA
BrHmnHO9pevMHUJxOSwkYXbobzFoOSrSvzW/colIkuINxe2gwYYNN3b4oQYG/SDyTSpErmMfdyNZ
nz+cXiZXpuhGbwu8YQUVxv35lUc6QXAZbPz121VTxo9lfCiAZkpcCDdje51c1mNWE0Fs3a1XO5Hm
aD0FAJjFHM5P764IyJv1WIAsNyU9ww4dJ9GKEcdiuEefUGODQQOLDaYYQWb3eIOYCOZVLQKjVC6+
o7pagDkJkqwjLYx0qPTc7eR8SHPi4eUi281JRa6scYN8tH5WU0yFPYdf2YC71gyheYHokfKj0EBi
9k7p4TSGCJc5tLpMex+s4yPOAeeldXvor2rOVRUm/dXySHUZK3fHvKd7p5rIjYMahxK38Npd0Hzd
0ot1qkpFbKBlufv6oMR/BTXSU1pEpR0ftnzwmYYYNBNbOF/LzzN1bNmRx/jVlwA9JQ1a5kVAcoEV
Mvgzx0eULrrckXIa3LpCs5BeDNmyg5tAQwUUNN1Ngyhb+Q0qYLKyVKd5QjHbJ78jirGtP6edLGr9
9B3f4M58SGufEamLeg3/KSnlo0Gy74d/3fH98ETf9snJ9sGCC9jQdn5KMQ/38M1+3xwPCfjeGefg
Z/Ybm/i0VS7deCXu1nOZWUUHEzo2l5w+tKiBjue3xCcSuVizntpgmOBbTT5HBaghqaTvioLOyZno
dfJkEupIuYN8LsJqthNN0DiXf3XwtQ0mh5q8WVVA3LRNadWAUdVZfh6NraKBL3Mbv9Foz5KrYLxC
/Cd1oRds8hxQb2AJPCbaEtbMtRtYa8dzZtOYK9OR4LyL7sKl9TYrhef4Qa5X0tzwLPjprc2mefWT
iavByZHHIMan1EvCjS0b3vrQXRIn3wCx2P5HlrFdiyA8njYINXXybnUXi1rRguM0FgZ9+/EbqMlS
ccA4dL0UToBF+yRdj2QhlnZwtFrHEdXCsVnMUxR0++GVaoSt/hO3SpFAsxXtBEvOVJ7raQqKTTnY
Qiq2g95t3nsxZKJITyFi6gODPYZk5AhxNCnY+SkjcWKJ0XFxL2w/2ACsHPSp7NU3TFxhOe+Z2BZG
ajgT95W4oAjW/MVZCqrWS00tinmS+yI3F8oIodDNkvX0LYr4jxqlMVPBUGMy2FY7ClHRxahPDqUx
OKev/3qhBZDiPw/kc4YNEZoWsA7gz9q/6HwsPQmG5D/6bMvGXc0ZYJzx84QJ9FJDanr968zJI7fo
7fbPu0ZwbI7fJUpPAvXJEHuR1xJGnabl90lyMSHm4ZzIFJr4r3W3k+3qo9Kyvg0XQ0U+B2lj+f5H
DaGnyvh7SLjTaQ6oWEEXxGvGDDhHHfRGxaCiJboSt7lX502YHkDbXq4bRaCJRgz35kg0g+KibjgI
OhKsMfFxT3mVuWk8XzUTPZrRmAlycN+DV02lAU1M/tL5hJUAh8nSNlo2pZcnbFLIytzTuzrIORTS
h5qZvb4CLA12JKH7LRC/V0wCnStpl4F4AYeEWaAri4ZQaPNJ7hTLo16jFT/6JZPHaU+JB5vKEi5X
TdhQRkKC67h6Ijs0d/9RJV/VD7O+/616u6sHRpP5RPwcKKWDxotAYwmIWOp09Z8XwuK78LVyaydO
Uwk2rz4cR1qVr53l4tkBo2gy9XUK2/7ohrhn8+4fELSrm4kbx3WWRqxFRM3NxMrj2cNYbky+gIdS
pWk+FdIi9RqGGi/9D+t/zHv11o+/eq/HKZB+oEYTiE7vOsIERUmZQkFz3k2lVE5sEXiZIYB33F2f
9WTpBb8o2luatGgN8JRScymTWKSrtLCkcyWRiigF9I+7KPrJ+aCroNAMZ507qwaIGHK4NJnvTe7w
7PXxoDMgP6OYYWBwg5qBqgKKt6nY93ynQkRb/8qSAEVgo5SRA+yaOttNrQAle2m+n/Hl7SATFPEj
l9fsPXM0fVej67UNHQIdwh2xBbGa6G4z+5J/g1QSdkwkDSchOXlI5q/kr/rPZSW5dNt+tqExJTUk
4t/Hx7p+uQAoZcr1XVH1NZcXLiItxsNNEdUo2JqlAcR6RxyGahFeUSAYPPFn18Crff/nqALl1uK2
IiAigRmEMR1z5+DXR8CzEja6vk3NYMTc6yG/UWj4VSwmTXe22Pd0Sj814kAJNTh1LR7SqaXHqVg3
ONN9zF87hZ5gJ+ckaHR0dfNDaknx+KFYws2OSFkschNm/5IB6EepvhB8bvSzufcP+zws7dDXlxSH
iGqUgX/+2oQRLkE6w32FW454QOgEOBOKdvuCOk62Z0hLXesQHgAuJsq/3SOxWDYm15U8sPsNwcli
V0Dma4cxSi5yO2kk6Y+DzJXhoQbZekkpcAz7L4JgTI++uCcEeoDfaFYXJFgVaced8Q4S3h8bn36Q
IyQT7mFOH3NmudD23LJX2DricK140OPOhOy9JvwYfayGiFNNDhjtsTtGGWscgmyP1AR8iZ5aqEJg
IeuoGUqlLtudI88gbhO3UHZNqd3IXbYQPFd4HZWvI8pQeU4eYM+rLXZ3hlWoI+P3lJDGKPB2BzlN
BH9/m0cRiyCJ8ZH6nVJeBjZe5RH334ssd6u7yDKpi/M8n6a93W9/sz1fRhozOyLjbiZvGCX2z58A
1akI3Cvj/0ThBTJxXbeqwY/gI9l659FfCpgJGAxquHbN9pzYuQJIXNRHXSmqnli8g4alCJ2Zhnyc
W8xdvZvCiJOqIEBbPvsKdGJo8Dym19CSufGDZW/EPOprDnghI1D6V1+DlWszWpjFNQvd81+hEGd7
Gz5s9TS80r0U9GLEHBMH33hVm42OvpYYZs/wZaDPzGOH7Z91s6juccxGPt0w0hgHYAjNHvtgjix+
2Rtx3ql6z4tez5+OqcQ3ebUuTVLQT1ExSWfHnQhJVDlT6qlFrUoqCxg+veWMuLSYQIp/FCobfkcM
eyWytAsYWzhFkXbR6+/UX8VRAru3IWjyXQppg5m7QbZWc6ndva9fPF4eJLgRObCAc5d1lX/hHGUy
K/6HEyby+ypoaeQs4Esr+h6rM1SXNLYufFEA+yvRb4BVms6vNcRMudesmVj+ohhH7ZGnbtfdaQia
LsuwClDKkDLIB+o2MgRZ/ZTtVTyiTdUfJuPMVVaUfWyh38jvFXciL6ICJTrZXAHyLbhIuzcvOqCc
QXOQe3O6XKHTzqm4FFcbwVqsvpPHhN5XBu5cEaCGiDIKAGddMadmz15lW4rnQO5kv78rZXjixQut
RfL/ed/aay6jumBwbsaPa+g3Qi4tldmxjYQxBD/x36ofB5Oo36fKA8xJHx+Nvj4Vx+BU1GMMFQDl
0WG/oVuhPApWCfxlqnm8mnhMxpY2D6470kRYWQNRx+Bg2lZqXsgvJLsTZYvvZtRgGBTla21gBMHn
TzDTzNK6VDzb9bDEvLkUMGFEQ5Zk5dLhM+6chQppIOYvYofwlDw4zXdYZuNgsVl9I82RJ8CMqjUV
MJ+48l2V+76Y7KNqqRnMEowE3BrqpPHNqAPROw6G5mLcW/nAPFnZ55XpXQ0T8Txs3uyLBB0in8xC
yIvJP+MLTdyB+pVGvNI2Dj4v/8rCxRzNIpFNw29q2zqe/p2dUHAsuEmtNWlOWkIVE9OWdTArBG+g
jtRpn0Tg22OU+omoh5iKgBueHfQX9Mvfu896qczNxpDoNbmLYwx63+hIkVv2uF2obe2sunKApI0D
zhYjmmcevBnkEiyZ/h8rQirt9S8SWHxIZLirWxc2sSOq4qL5Cz/uSppTqCLIBRrkuH7d4+TWMBw6
/GgkOtbZmiN7kJqJqJHMZl8yyeVYqxCQuKFDs2B4j9rUy+bxNjh0bCepY4H8zD93MCxVNLZZdF64
M6KlQD9IMc11fpAQm6tQtxXxMZsp87/yfy9jKk52C6sSPK2mX+rfo1ykYy2Lfdu/BJbr0fQSnBdu
+J1rG1+C6sXGfWVLMAtNBbvl2AwNCECcK+rTfFbGpqX/Plu8t8nFSE12zaBw1iYikd3JZyZrt8rA
E+D3GMhh2ZhqJXCB7VwwulKQWOQg5cPlnwn4tj0CZv4HFJd+hEbNYpJyrecOqa1XxyeBIHLdpWBJ
Z3pz7mR2t30wGVRoiIi7KDib1l+7s5HPW4Jwmoz6Ha6XZaktnNOelaMKeRbI0cu0CaIHvO4R7xx2
zQ9CAFTbGQCnTQBHpFxOVQpNRSJnmB8wyfG/uzwI6zoWTHdc/m/+WsghtOCsyYz+rVPBYx4Lf5RH
Bf71FHkZPjhG43K25VPjtwYBGlAoYKzcT7a75NEi9yNrqU8u84LKhnW0y4Z941Sa/GpvlNE05MU8
958XbqQXFNs5WjLIO+IeUbTsutNTgQ6Myn0KCx3hi05yXqEjbqctd3QVhGY4Kc+iMwTmlLEcZKyQ
S0KOe9d2oUaU6YYEtJqChjlLv425PrzR80B12Jg2sxDjgEKNW0QkwawQesSP8L3Vjiy6rk+d+4ZA
+AGUVMYZ1Y8AnQUh8lebmk2CShpVI1H8nkeCFKbjTf8uivKrq0aTfQcjURzctw3BETGPYWBHm69P
i0KuUaLJJn4VD2Du0NPGKyNtBILOj5zllydY1xsKPS3pM+ATQnOOKYFKxhQFPhSjg3UuCXI+rdtB
K0PSNLokYgBUqIYhnHiJew3SLnQD6bisHemQIcwyN/IiUg0eaEd30Nc54QRtIQc2Nxid91+qGAkM
EG4gZPZoPrhRRwZCZtwtSGikIV0rcjyrepD69I0XpirfiPnopcaRrMn0y0x1nYUoUp237/9inOtC
rJFgVCTVHBypqnIQQ2IUwPGzwqi2RPe68fAxvKV0dV3fJO33NTn9Q5RCpNnZI+jruSSsr48C6nM5
91gx9YzJuFmr2uh16+aipqcMJVZS6gxJZwRtLs2SibWMXNdQhc+lGQaSwkshzP0POt99GcIUMiPF
gTmstx+qzYeqkJuYItgHGHXKePQd9HfSPvps++WQXDUKrDrzabTKJRvJ5Mk9PSPph1KLtYEgG4xC
ASJ6N+u6pIarAH4/l0odNKZUc6FfdUfyes5dZZlja1pTsQSIixAg221r5/ma2SHP97Wx84cfuEG0
zGK660/SI03/C2VGdGZfi7XBJWdKZ2CQ91VVkPzg5uQcaj0sixJxlxkwH4If5lZ6sHyOVRFD9fZ7
r+hFpCKNhWvaPLxgJVBtX0lra39nDcLQcQVZCM5yvTEXZDJWJOr59PFVumeiI8d6qHocUdkC9+GA
WQfkdtusoeYrZ3RNF8bdx6hnw5PTKXkibvHPP3mVYB867LIOXso0OxfRajaDcDJn2hOqf6NKiFIm
kx+elnMGjxgETGNtLKxmBEVohP7mx4KYPjIPAT2U4TNoOLNsYo6D2WxmRIuciTp6rkHR/nVk5zfP
ZT4JRfwOyxa37zywRRgP6SUF8oeT9A6bAFwSDc+H4TXObXaRCtM4JcYsc9CxK7msurW0YFXjjEED
urVP9odzvnn92FiIttKfOdhZYW7X1FqhSn9IYzmDl+aO9zZOyZwOH3mxfWnITlOJazE/qI+HSC2S
JzJrdqbYThnbDLconY2mCNHbvGcM6DhKVeko5oZPa01QDIwUj0uYoXKrXdBv6dX6ovWRe5BcLrS/
itHORXv0GXmbMeoCB1jxq2xJIAqk4WPB7W/cMXWPxDLAw3TNV9aL+3rsO5pIJ4G+bNS8if0OMqXS
DikzTPPaAr9jIL2LxFHyQd75UpKPzTfZZHN74DZ98wTD4Blg1AkY77losomr04CLoe/f3Tfe2eQ/
YA1EawfCAdMSVE4t6cmFQZrGkuTHhIrwyHB7LreRWN7r7ybDTvSpAKxkDbvSjPpXkmum2DMsTH9Y
0UIOnu/UHIdLB3xlgpQnkmVsHAoNCYxORLXCR5B8wcT/M2V5gLnxag8KSh59TzvCLuZneZWV7p4S
YsmGHiUZskNF5xksAOiFooPKhVdpdKkC8IoNiFWe3DifTFqaj5x/F1+Ah1O3KDL3H8BuyqHgNnUz
lO+fGOtQZLekExVPG14uvFmC07kDzWTZAv7rLN2SSPBwMBeJguhW7FeTGFEgL9a175zvKR8o0YGG
Mshp9GKOf/xJuxkLzG8C5TCgor1Vvkz9RQbVtF/htT4a7sJ2Y9nYjwL5aRlnVxwoWkFIRCsZgLmE
NH/KUMV+OHkvS5Gc4NuOg3d+V3onjylGW7E5/J72M6ck7Y1MoCFE/FBsk09uCDhYup2A1o8ez1bt
Tx6dZpJ0tUxRODm7E7M5ECNO5SXfHHr5q++iQIEFs9lJRTrba1nb+Yejim2zCEbN7EDW8LYlfZm/
TRyDPXlyhj3NDFJWastk9WG2EkeK2TCFt5o+2SCzsNei+i2tfZJCv0+fwS9idTvOlxrLVEIIxSfD
1GhUNCvZZaK5Qrc/8BM1iJaU+1v9wCeshyWcpomTeLrvM5OjKGnGaAZ6uub/2BMHM5Ub6xA1hX9C
8WUkisMgAPEiw2dr3JMKmX1H4tLuNBCxdWYfAeEl4n4U/MqT7M7Zhogqii6AZ36CNGU7hOPAjzuy
lZvvmrLrO0nuN7EKol8FuYF+zhm/J9CjfWY75F9gq/tyaySqLMHI1tN/0561LL6HFu6YSBo9C093
GhEn5BGu8Y8lFHpRmygF4eZHCIRjNqpmWgWvgvNPOBfwAPckynI12qLSohQdXMkQih2elmJIWooP
XVd40CEut4jQdVgAVtigSOxad/jY1sc1T7sqIW6jlWAJkoda4azfRS1jZbVOt5wTjtQKv99n4WoU
05Rtqzi1FxJL4NOUkV3NHb4lRd+0jiie+Ve3gq5K9v5M6TGMc0lVXa6UA2qUQuDh6Z6jKtj4LWrq
ZRIrLeFge8tQhVKVo9bWhbQmWOp81pE/0B9mwlU07HYw6Qyt/3Y3U20xNReKNdoOpqcIPtk2WM3J
a0lx0Zw2OHk4xyPMGqZHkGvSlTCoctd7ouriW/DVOgKRmV/8wukrXAZYtBGvA/ZOXLyqwzntezk0
dtDqQlNeM0EKg72BII6rmq/D9F7UeW/X6JFx5/z9Rb4JkTCbp/ep8LHxH1/GM9yqvA/ARJT3e4wA
U6uO9AFRI4UcDUWJqqWq7EKfNE/eE6lvar/SHJMfvtYgKgy8UWxtrAING9yMGnlvxctj/fBcOwmM
fMpoIfwxft/hvMznj7P6acQQlYYBaNBpT4b8stB5IbKbGYeBsG3QAJZcYuR1e7u6e75DbjMWBBlS
8fw31yUEKD8VvOjefIX3n0XjGNZ3H+DpuJrNalzaVueeIpoAtG1N/EKsltfYlBjTg+3/A8j6sTjC
7C/ZP9k8OvzaDSw783UpKJJ5ZEOLMjTdeLC8sOZqW8jV6yFACsrrxN3QRYA6+lS4eoPcsY/VDYjg
2pxv56pVEgIRmFHfIO5pnVLL4G9yz9oAMq63WLr991ORPCCST22CUe/ooPRbY1FkMIt/WDLq3RSF
ErgEhHALYhriy557ODPEOX8VvC5kyIZnwQHvj+jfuv/Fd5PYrAraNNBR1wZaTRgfvFa1K4QqwUCd
Yn6J58DvDp+OeUuz7BOYRNa08KJlnJ77uS82TG5LWO8Ph6EBxLULOLNDRl1UH7fdwoyuJBwrWX4D
5dKaDAp9lfdJCXxniifY8qWMO0HVNy8PPxIjAgzVLKLDp1vgMh/YdDPVDl52vkxJQT78Jlt2Fet5
gGMEWqbvUB33A/w+QOKSZZRs1/6z8FaYwc3UFQXj09HDYWaXirYdChkdGtcVhHb7BHCwgAg48yQg
iaz03DZtAhj5KaWE34P82uceU92oYA3ZQNPtIOkXaz2tXYTRsTEEnsrKGwtJAVzN4CrctlrS9zwT
N/4MgsbqAkzXoEfP3lB0f9R4roYvxtXD8L2D8XKhuA9i+2LKM+kd4fbtAZgzlrN/tLF7QrD07IzV
IcxThsNTm6LBoXJkTCPFAiG/PnbwLmS3xLSvBAntvBhyjJ2ToobYfWsvkfFzhffy0qIiiFPHF0/1
W8wNDBt7FKqMWmc9R8LMb4FzIDDYVLuA40+ixwlV47owGAQ4OWsjACTvyl5SzpPTvqKD9WyJRKba
GpuK9IPjc44t6wh1bReFQypOyguqG8L7TehsvR6bF5CjEGFPMEecwzbbdKOnl0gDnQZ49Dtbcr8K
4V3LoHbCZCgMlgeXzrcCewWHxXMLv4qYSAdPdOrOZ/lv+uCsJXMXGIOvczA2hVpfgu2l70q6oNQc
6iEPiPGuojZ7xr324jUH7FF0kEFH8WZQLCOemfabU+xLZL5w1NXxZYUIPe5pP2oDwAxuGPK1VeMA
TwcQv0u4bZfQhv/G6oxOwJflmntAU9cS7XHHz61tYgbVn7YK1v4ojikpdVToV+vLSMuKiEODD3XO
w9fjo4T83b9uepOhm7pN9o9NroQDoJR8woXV4PJKTUsRXtCmHCKYrSzGZhSgvWoaUICzWBW3iwka
bqRT32kZToqwH55IuRUI/zO+AW5aOwRtB84Y/qviUDUQdtdg+tj/xefAQpqyShrUOHUYxrHcOP6h
vjTszorvYkWnrZiBRRQjXwJy1IrLWDh5fSSYLcGiM4jVNqL+VjAqHXLRk3nqHtD2kyg6RBCEmLxu
0ckkFhHX1Zo3ih3Tl8x5qdwvFQsd53YHweoRh4NmouxY25RWCs77IRgF/OSJZhGxfv6crOoLkAzo
lwgkvTlmhOHsQb03VBPUwxtMQkL2Wi3mP2KGwWXvC8w1HV/kw2dL6hUFmfoAe4Lv8Yy3MraIQRAR
mRIpN7RDb/QgvUxiygscVL019+cMQ2Kt0ZxTdcqKx7IaUKiQTFO4VD9mNbBq+lSNvZQ1huTthEb7
JZKvGo4op9utxKQ+s81mXArQwvJzLqPm3LqrJfDxGVjX+wRXoU2yudpns7+LbfqfsxufxjWsXb0x
eaQUinP9V5cNLgByueY4HVkmKzq5fxnyWt5vJm6EIGuNw8X1F03oo5SzVymFHlziDqQh3iMt3EKZ
kR5bSngcsAD60bOS/kM1R+lEkdeg1Kw4JwRtIpSBID2LdBJ2hHUTn9jyOgghDQe/j3UbdxEAAq++
O5SUDtRjI2SzyeS39jrth9JV8w9RZd4ROuSwptvWXyjT809KiimN+TD/llbrBtpNnR++zFyWkt5Q
PgjblPr1DAhA0hEo0MXv14JUdKekPwTxX61SNk7zzt0fJmTJZTWtnZzMZERjhYiSPaIsiP8saNjS
qb0eQWdQHxYoGQE2R5jhKybPFSr7cH+3tGeC+dEfWg+fCBUmU7ae/gAHx5TrVIR9/oZOQ2fIdksV
lTBsi/yLu3V5fCgX3AJagm5VOyC2oscfT7QduXkivvXAWjZiXBKiIo4ZnbZSKsI7v9WIcfxFzFkr
KhNvD28UY+EBUPcoLA/PU2soGAb4LfwuUj8G9uRZUtUdovIbJvoHtzxUiNV6dxMnuy2YpEhAXNwH
tV236CRzhX096In8vGGrwweBblVJErS19Vux6am+uuA5JJBkODMIbHQOQR2HFXcclzauNUhhVvuy
gcI+4MjruSOCZdiNfF0TuriL9Nr+h6Zgnz/G5PrC9HhEpdTIanZSaJX7zoYzzFC5IPHyl5hjfHGM
VXrCJDnRzzK3U3Jt73wnHxVC3yk1eqjS/qG7yjVg4dNZXjmvb1RA0o4pMUNIC/ecE6EaS64D99BN
VaVieCuJ3WbkLhhg8h5cy+9loYmtjq7vD3ctUopsvbyHGOuUqKQjs/+PuJYZtTMPdcABBB25wEak
P+M270Eoq8NWTbtm/V3EzuLeElY0PZ6cr/B5EqNqfbJy0EahSbGN+RpLJdZv/eNH/22J2qZzoNgo
gC2tfIGkJ7sF+e1rOrXQUqu82Fy9IF8HcwrI9Z+wrPYYM49cdUAW74LvGzWkcfhprtWuGX+Q1TJu
PE55izWOwteVN4UbrRewts0EX81mEFR5xx+xH9+b8JZdn30Sbda+474j8BSei27t4eVUO+7JaFKx
AtomgAlDTUOr/wsSfini1NS3ACC6uY93scguMwoF4x/HdkGmoIxnFlC6OrzSS+PkLBj6hxeQG7Fy
vP+g6tmngoAJfdGW4KU8aFCITkq7kIjmb5lBVJyzZ/D+RRGle2wFm8n6Gw6CPz4XlsCOIBeF8fWj
/i5IICV7rXLspePelj9M21ENiah7Vl/A9X4gRP6AyCVc78U8OjbWur0OEZrCTsqyIEBOkBy2ESvk
wY6B+cDbgWpKwkTyvARfKXjHqpZ1/C5JlpKaO6+c0lDnUo+8rfKpaDQLQKLKfCvbQ+1XFwxFNBIW
Jz+4Q9vFMSvwRJlxJk3GS2eV1AdxtyyPf3V5QkGV0XWZL8pWxyyQ6PTEMSEBg8aPAPSSIwSyh6nF
ZY83iCpLXQqm5DEkVOBh5khZfWUMOjzOF+IoxZI/lDEYBark6aeeuMktPMDjB0D/2D6jkn4OKMx9
G0OSlMsc+EBwK9vpVjmtYozyZAJhf+zCjmXCC84QJALDWaFAa8mK+173E1M29ymg1QCW3R+iz6/J
QA5P6SoEHJujcMqmutvP4l20cXbrU9mqZaY5pvW/hwqil9S36qQszyczCIhtwVRIgeJ5mt4qvF+g
wt6fy0uLAgdFIUujgQsYdEVXDYYiHNVY6SVFFWGspeRlznNL+DzUrkXYkSxf3WuW3qBma+0ZdtwX
aN8Kv8V7ddnilmSoXD3J4RwBjmcqPpGKFTKuhBnwe48GY8QuxcemnizDWMYwltocZErVeaHwepsX
zVPlfF7DbQx+DJyElx6pa/0weXinZJTUJTTNe56Prjf1uZFnIyz/frfePkU4x6KbVpigZTYc336y
k8VvoFbNQyYxL4c4cTP+jLh0LouiZvjD5FuyE7HI2ktvGKxdEaNG6uT/AWcQOIipKXQ1EyMhqtov
/nwOlXpKG/02QSis0KQNatY+pUI3D7NFQ/DCrQ4wieZAqXrq873C68wEQhDMmt3RdDT8jgIQbKWw
j2CjZvbwgl1rKNfhR6FmAM3jqayTfP6Zx51g/Zub8j12wgfW563CT4vGknxUYCzFT9SH4U7uFUIT
ARCjk621C2ot7n3gxVoKFFEKj7jgaKiBgpLgSU9J0LBM14TpDa5I97tECp43V/tL6f8HgMLLGyxK
ZxEupct98REz+iqb0yR1MCa5tnpUcLCdAicnIcEeZEnUgj/18DzoPQF5ZP0A1MLDFdb09tssDnm/
/oQ2QO8JxscM7aFofYEfiIbPdcnxZcg3GZ79CcglG3mF9C+4J/e4wPjrUBzHuist2JltMaWG6e9Z
wJZi/Lf1P5CJSd8S1GxVl1o+aXDauwfSmzw8Nk+aIweRte1HW15cMMJY8jjirA7wDcMqOgEU+XaN
tNOGCn7i3tLnthiPK+XDOTqcr4k2Yh/OQKbH4oTpVT0kzeE+BVdCi+ddb09GNPHYc0ImGegO+LU9
fdLOgAt+cBSTLs96znc0hs2fuXvugy4sy7bQG4M6HcLyGKW6J6X5hAIllYkouyWDOXJLiLBHwsi8
WZWqbL6/sbgFLqKm99AJg13mG/IVJTgLxRPxpSMRL4VuxB7bmPH2+LLf3YWVN0FNhRgj5pGQyU7j
yxHGCVggVEupb8dEyBWJx1VeXehaJAeVv4IqTYZF9nSS0rSuQG0eVV3GhYrk8QAAKIl9kJuRacgW
TD9akKTP5/rBQ53AdYX/MOOWB3KaA/7+p6+GXWiLssGpwpoRAYTuw3Gz1h48Y1xnW1V1bloc2SU7
sxVCVU3DMzQBCGlQViJ3xnbzjxNCDqDMTOtw3jY1fnH2o5oaBXrH5mylivgQfRmarg0n6gdaPNqw
j0thEpIuuCnfM3sNQxXdQdEyYlr+kLdAApwBDr9qXDoSQXBSD4EJU1zYU3eGXLTX0MoioLOlScwb
jnIfiMlrWBJuRaaPCzkhop7Gm6YOpbcd3BJLF9wmGPicFWpNYkqG7gnauF0iO2vy4mqABXCjubsd
+EpEBiZ6OKwX3HDmHKhGwuItMqwoKKOyxI2RsbrkSAk7EDEfruigMsx/cjbxIxqVOEbO39WIOHPg
umFi7w4UztYG+xLCKlqy9wdm3yaC8VXmaRQ3iTzYBHce9fjMFSTSJeKxuY9IpS7RnTXvDxCg8V03
HKAjhOvZDg9DtVggwcs819ANTQXsNwtEPhcXy+Ws3piIHrxxboKjBp6agUcZmzyhlSi71tSXQNhD
E4iwbtRnmZ/pm7QRkqNZewHW12DcqpMzDptpFpXaKRIrcUNzfYI6gto5ujmNcLajhLie9poTS3Op
WfvGUUD+rcf+sg9AHSLJGr9XuYuEoK5U5l69S1SZU4Cghw2mlYXRFOap3GUftUPCMHBVZrZK5hBe
Rb1pZEXDXjwTmsinWdINaX/tuKIUV2V2ESE9Ra77Cu5XOeRYyVAes72ALTG3NiCEH5TdAJDzPrKT
FcE4zGi7gSxjKtrw/U8txjYzQcNjKVYZ5bvd1U5KPkKts9X37Z/+yzlE6D8ZMnm385EqPc8Dv5Ie
dTUyv1DrD/OKrYc+Ul9CkioTvA2x53tyQCy9CIO5K2ratGU2O6bmpnUL06hxZIo891zaScgZrmy7
3pQG+8HSzk8AEtI8fQoaD7Xlu2VB+oTXYnpIX3YPdfrYAUVFWS1nczNkulcTokDyjV1d15FZ5ejK
7cGu6FW3AAdBQwDHEWmjq+cESCv0GWsJ4pUl6AAYpHHKgHd8tCkX1xEUbb2FaAjeG0rYBXVz5vC7
pQZZ6lcduMX7jWnxJ5ZdAmHSqh/GxRE/13ZMqxgzRVNMfPvoc6bBr/BYClHGMUkJNwY4OgFLQ2DT
5Vmt5uenMyolCjXJhBMN+MBVzC2vPlTZ67yCD2Tws0RbzF1mkiqwSuQPg/ApAE2lu+rqIleZyHti
sbFBDJPuCcIQgSs135kNKx0ZCFVmZk7zLM7IPUP30sq6r1AShnpnS7LavAkTxQBS8RHfFKe5eI8H
xJCDShgCi2qOUZBPUbIS7xBJlA/vdKDyAPAAMT06vsI3lIXc5/KB934IbbNJixOmzGbvslB5rdEw
AvPgsTjkko2ZAmwhoTuoylgg9cjpEuGwI3JwMZJgaiD3kiudJP+/kYa6c1s0iJ3yrzNTha/Wrs0P
fyPxRoYvNkCXk38c6VF/EHwWMN9WxAM8GHstrSBKKae9auKoBtZG6qWaA3xcjdpxLyDLzVZ+srvv
WQMp0b+MBgveX5hw3ariawM4/j3XHZjz6aCLUCZA2HglrFDlyRSAXmUtoIsGGEHNk6NppSlmWv6R
y10tzrXz/Xvq6eYEIBM0WzcWjNit8xMdGxOKam5k6AeuopVsoSf7jWBbJYdNPBGLW9nf8iUnecSg
m6mM9YJ7Qkum3JWryxBYEFhIvSi+yG4SOCmkuMQqyNWq80+RHJRNOPU2PzAubLqXhZyangL5Fjjb
nWBggk+3dZAqndi8AgngRND1UCCMRFwa5YeEjD/vJlx8J8mTUIvLs7ta3PvqiiWcABoklpMWaWty
WxTZn8tmVEWIsx36hZwRZwPpXgodL2qMKDeHD7cxEGGmKfyfhX+pWUmFebUG6sOHNklaXVKkj+zD
G8g736oU7FTCKHyOOXQuiDwxxC2wF+6bbh4JaatU5sbNVjiVjbn5R5kQrxdd7m3ja1uR0ZKR72lx
u70kEZIJ+ITvoP4JQFGQUHR2L1MH+xy84F9wj4OkAQAlJd13K5S+SwOkCjErHcmQ27KlDySpKBYT
mhnMVR5BMQNE7nRlNIwJqIm8CRiDOXvzRBRH8UD4sp7NFOD5Ax0E97+JIfiDmU5yZZIzsOaWSA2U
wQZWsl4yqPf3kWe0YoKNwuRXYyrX8yGeABC+22k/lG8ujvJ5IKKI4ErcEkdb7xwBEyer4Ai0osfI
g3fNj6lUmaX07e1M7bwZpSDxKKxMd/CwJZAUd25tLanakCTzFJ9ipZC9e3s4Y9tYfmK857Uaizs5
bJHOwUyGETIIjXKh+PxoE7l/VCo9koPrrcyCB2dRgtEnHR03gwfH1H4D0x4PH6WiCT7eBnzgnbpn
SFtCxAtd/8vxEx3neo9HBLfsIeGr3pYv8JVi8woEYwUGMzAsd2sAQzgRoxJU/WwdedFl42criTQA
bSeeOd1VLDm3Hr6fCEA4zWQfsqk+GrOrKu5O2bYDFQUv71AMQ7ruAbDIZ65rob8acSe1sDuwHlZv
6sWWV35niw6UDCIxFEmCknxfhHsNYtRmsSiOG67iFrZnDLKgzOVdyURmvr2upij3nLJmmcgdYIGh
hvM0Aupwtj6gv4dGBM5DcBXItfxSnb7pIipT8ZuG1q1bGdsPuUY7+DA9lMm81PyABIzdbCrCV2R5
cl7x2XLdw7IYwIgUfobfE1PMnyKOGBjkTJR6fRMFBie7P70fSZKnEINuOisYRq6SHl8IsZaMu6CX
Ae1FLLVpZeoz03TNP0A73cdh6m/5rvuAtojIMeyZCRFjzI9QViv59dTFXPfRaHQ5EjD+UIX60jY5
1kybTqKD3fJqwlOSzTyPGDr4fqBhKeXmphB9affxh1tMoP34oeW805UZaPRQ4noNEa0CkQ3sCxK/
lnjCI7Hoj/zdb1DQmHuej8xA3ap3p1U6gBdn3jqBaGBTat/HyKBX4yXDY3m6Vzcpp0QYGgVgbvVW
ixwGEnoi/GUWpNa1zvpHuHcIDiegSqEm1leMzeaqIU/QCG5T39mOPtJB9Z333+k2M0ZzYIVrGu+h
IIE08+0G1W3jIA7+QgCtekTdho/By1dDcxhIFpqvhrtNn2Kg7Kjilr7m6QsronK8U9mcWaPzX7Fk
JqMmEGCAMvFT+s5oLcbJOQWPj6qXKrPx2CCj6msSnSl2Sp1vNA/r0KpBLDPxBHQU9SpYusRy5fFu
lCoIY+Ic+FPOfPAQb0y+bHj7J7M1woR20IgZi9BBPyYPLlTtdI4OZ8P/a0XqJphG3Cf8Ju/LyMM4
Vm6scX3aHasxPZrslBgqRXqJ0sfF//uptzqYdQ4jEBBPUmFYHQ0RMeQcYQM6aASxCyZVUzhnqdQO
Mk175cw9biAdArwVyn6GRlG3buiQDU5Fqflu/g+SxlfLMQ9vYws1oq5iDM3CNKiqzUz9AEifUb/0
ncekTvbWnx0vw0m5Epzfk9mLXfCI/gNH5aOB4q6FC2m0YUMYOtFCnuW+xeZ1XFTH4ZElfNTwPGVS
R0OZui4JAlzb5T7UpySUGYun4X+1X3Vggb81qH8LT6Kggd4amhhInEo8da1qgrg3bGlCfZW+NqMw
xuEAqndQpic2RdfZh1bdym7hGzYNGpez9yxTaOBoj5u/v6Xf5qXZ/XxehdKWonRnz4XulCm/noEn
rp5vTjT9tmZa+8mpCuAG3r4p71xEtPRMMiJg+hwXqkbNtwMoEgJ8W+QN9CzyI8QsmupZSv+t6RTP
CyPmwqYV0oA9kJbKE+C22m6krmVrsSPLNJWXOafmW9/kb/hdccBaUnJ4fmdQLzQI5LdfZmvpL9B8
GdfCtIv1R678AOHPAo3owOwxYRWxRSkrUvMWsSGGLD0ZjHiJ7i128hHpjeeAYtMjQVqmsIS4suR1
Fv/hS0J+D2+sLTdh+glq/UOp7AigtwtByCC1DiTSsxtuWzH4BXUoGrfG4rOGVzyorF5LL0VhfZLb
etmZfmAXobVLq9hND4bo2bDR7NsxQNGLpqV4Wz1cd0xfvSLFDgiCkNbPZ5UZx2HsORwf/Nt7XrIX
Qsg7wjPm+gb2zb3v3yl/hLABoKCM06m9mKpgxQrqHtkbUoy+D449uyFLyYGaDaKe1y5Tn+MCJxH7
wGzZdI8zp1LKZHS6b2qw9Tllb8GvI8oOAYT7Q/CNADrL8OxwJn1Ax3ZEnK5gppQJ1R0YO3e2/5If
J+Ntst38z9nTQbdGEJB/X2Lg48qKKRg52c/5yKdU/gq9pMqpLZnZN9y/wK5YGTx5lTSO8NfBE6xg
fNgarfr37BVimrHoqXLB3zrFPyihq5G+cEnnJgNYvLbuqPr1uOKUjDO2UDuuym1EifdX/Accqm8B
3WuDqclL1gkc+X1lCZqmbT/ETTrcOpOaA2egoF2XLutb3z3G6AKWpXaghaBnLFq6lVRMfzj3JN7v
xSaZJJiuijCoKNBPxRCxIvs9LkaWBRT9Z4SflZU2hgenioxZQwq6jwPd4YurWYPrq0Yo/iDNhTBi
MxfFx2LIDLiLqf8hNUAh+66LYfR1ffwHJcREbmv/veZsOSJ37A24tdL5Vj0qdjvm4SGsK2JPmvzH
L/w109Ef7An7DdKe8YD6PFsa2p08ULC+VDMAUsNbdiWrs9wgsxSb5PUSQZ75M6rd9bBSUP5wwszB
Ph4PJDJlN7aoZCdZZwpBmM8Ski9hudIT0wR8uSeKedt6TPgnWwCBFrHxLX6dxI9npL7IkIdP1Srz
J4jU3QWwJtbsCb/cIKCmOnzJvIV9MW333AzIcE72q1b6D6tJPmux5gnDuCs3rPiSpFFulTjgGA/h
M9ef89OsUeXPflYmuR8K86Bz8vp2Ti1rKhthyBT8uEHezphVVKF62Rn+x13eC6p0nLtiS0hZsPAu
rZlOGL2Qy+Q74rFfS+BAktriuVxjxivl520BRJJTb4bSbf49B7gwZ5dFTMUTERKwUvzJkNfedC5C
pbT14o6IcMs/EOuGKZGnkG4sNfutsa18os8TgX/xSzqWsmfPjqOuLaRCAfoODSCiZckkJDf7Gs/h
OfIUoq9kKvgewNjfJOA7uQIKir57tpD7s/3YCFYbqt/MYVRjB86ScmsRcCZi01FOBK5qVu7Iyjpl
F5TBuaW2Hw5qIofDqyAv5qPVOd9QhoxLJK3MujZqxcJirrxUxsFc09sBtFzRt+IsbwRfJPnKoqDI
xKMaN/n+gnKvqnU1u03y9EoqY8f6WLxU3SbxrFPIDiJURjlUKTGBkXx08nAiXd3oRwUC8fMbFIj9
hoY38YrkVtwgQICQC/zg5y3RbhxsjZM0bMrwsv2RCEIqixVYX/HxNUKt1/cOFsR9YWNNXngs4CwK
MafqA6LOJxWwwL2IA1rnPKKHCNRRiw3dk9rMBRbaNdDBZdojSqQGwVc+fGCV5CUlOmRlUSTc7pwc
vZPBzpXndVuCRHPtzkdkbMIf1haNfD6v+cE6tnNPNWDT3l6QJerOMCoaMCXroduWsZut2oYI0B13
C2yClXO9M2U2cPPIvdavE4dvR+WRqn6Eblx5vLahTItvcNaKBgFQ0AlZHuXY55EYAIT8Ld6Bgqoh
FSC7fSBLEM9OOsK16A71hcmYP/5xMe9/39Y+Zovu+mMqFzFTebJox+5jXmLSvNh7kvIHpkPKZM5p
lmOHC0JjSr/dtvv1e13YAiTJoc6cZt1IC8dtfwQILdN0QwGdFEFcCx2R868mNoiRf9eQewdwWzRG
o3cfi4vD/dj2lmDFTuhvTmB/nCxKROn45Lmek3IWXdvGVo7lQDJtJpT1ayZoRYsIBDcKA+qD0wF5
gax4Or+d2xZqrk0ifML8o7xCJ/8KbPHN36UoBby9o6MFjusjRy2iZZxKTb4EJEnfEvN+Rqg7+NUW
aY/oItqhKHaA6zqrMeb4gw6ZEFVVy9iHggNbgfILEZgutechFMfOYu9hEx1yB43lKY896OD6XFUn
Qt7Jb99jfEyQz+pTUvbF/Knjef3Y29Nw+UiVUqEyjcEXWRAoiQQQ438E0AWuQq9iVPe/23Z0LY2L
ygmL8P/8ycA+lPUrjtrT6kY0oq1/iex30+Sffq0nIAZKjD6Ta87VWlkB/ysj+JZ06ot9S4w9LgRn
3ijzdWABuGqsAFKR/BTWaBNtkm8uhYKtkukRp6ZisQg39EsXrramVZtHM216tz2d+EWZAGaTQBRW
/TaIVawXcZAVLPr8W9plfh8EywJyaqKwuN7LmNbkJTwKqt0LbgzedWW5/2sGEHiyB5QD+aPHou67
PIBnXu2BC75MKU98c40qCHoI24wcQhht7nh0xHUwZT5UTRA7CBISIfW20exZz96ON8mhuTmSPU3b
sBpVHhm5E7jHn5xZgxEHoPMYBam3x2aGD5luMnH4m77g+aGFPrMnU+UpZ30wFAqwkGaKWX+r79Or
+1xf0mGDQ9T7Fy10q6jLLKrst1pmpxDHQxfMc1xcWS9MNSrvRkh7LM1vnYg+RXY4+9/LRTNueotf
kdMzrIC76DqM1HPEBRebNh9pmH+hRpAhjOSfnd1foNrWtz7Oauq4IM1IYduuIFr61tf8cP+mRXB0
fKHNNHvofLZ7bEJoxAFK2H7bvl5/uR1a1PEpEMCqBd0Vl72iIeBAPixGjsIjRjzaBSfZEFY+atUL
J0EBPI6AYfTdVijtIFNGrC6g7NvNR5QCqqskSCQmUsaSBhdjadEFCSo7aXvS4TwI3BFoNr9N6lf5
vpvb/dIrjj0FmQt7HJFC1wsK6ypb/HmIcI6NNLo1HulIQZe0FRNTUI0uxpO25zQP37rBCAtcSjnl
dLhcT2xgSuXzUAKEdW6qCK69hTn4fD84gyYufov4KaAg2pz5yKd6ytJ+3RPA7iw4hb433QGugBXb
AEBM54B6nOAtafLRpo6XCJAzmpIGttjnht/wxiEn96jA3GIkqYIZToqYAcbca5juzT9yCfh/l97h
r+G6XvsKCI3FzfVdMgp4Q84aadEzo2dWj8NI2GEY+bnmLvscIpUGLYtBqQdC+jXiDnr37YwJgPdB
vUrowgVJQT2U7tKXBQPHGSD7vpsmoBRwNETMYjyj/dD7M7fWY5tYgeUlMEfGLNT2qLg9kMbk/LT1
h9wgr5IWdp1S5SwC0CaR+E2i0o8ppyt18c9dDmjp5wD6YRSJW5/VxpCEfGByTFplWqpg/Y8QbgpT
iS2Ym3LmS/JZZNDDju0yJxHHlidn+t99x+lrAdw24zQqZi8v/49rf18Sd9nF/dXSAQwUoGDSOHe6
CjFJthjtCx8uuk+L8mmrkn0JyK4bH4WM2kp3SwWrjTTybuT2D1GdXp3yG1w5n4/uBXjdVxkbygU+
dyoNEwxy8ogcRFXY+3nAlxWFu7YqGGFMd0xOmT1/ihcNArvSIu4dHj+OFVadHIpK+9RdrR0bv12E
k6fq7roEJR5O1ksG83A4lih8uuBUcckuctXVy4dfPm5Ozit17sFocz8jMU0LXZne68Va3FAdXeMb
iN4I8+ymPChPmfsHx9TW/3KU/ky2+fwfGJtOh9ByQJteFR2SSBx00nWE/Sd2Z0ZLJI0aiG2ZH3e3
YlkfC9Qoa/CIeSv9w+ROnbMUrRT4ndVUGfPHLX+WD3X8NcGnsKXKQhH5Gn4W0G4oxI2q4nf752hj
hqkoh+g7jksFvUXM95DBoa9c9fCHHMfjxegV3t9vQjOZbuNcHchdQB+XfWbTerxmc5T5+EVJ8jYS
CtRxPajk1ztv74METroKtdohO5dD96PVdo7scSB0DNYVTx81DJs5jJl5SrMoLv6F8OGrXtv4HGrv
TURNPk3T4+nhEOXvGW61lmh0/yIZT2DdfoQ1FE4j3KsfRYqGyIx/nUqAIhdJhR7PQD4VK/JZdlNS
JCkU9nE7kZMHVFEzarfr7a27jVXNODRxWTvyxaAdGVncySwegZuH7jKhsxvi8PUSLgmjr8gtWxSH
hDudQueLO0sOhWvQb+4GaMblzayUpJfYS18deXcv268J28nK3nrLKe4fhD/i5xxeadS6Azgo4Rzc
/RfZYoEciiAgLygicLTPX7dzFId4kqo5jZx9ZZO60kv1DtPn8Ayy7jW5upJW0kz6hVTv60li6c8S
k7Yy+QefdsEKcZhfyskJGxOqUvZnbPYvzpsHwrJZioaPCW0rEBUlfbOOBKGaemePDkEq7bLzlCmL
LB1JNDW7RizmcmyTi0z7qgAej+NwUaGDO0OIzyYtLg7OkO09xzzo+EIefN/BdBFuuEa3ZPMjL8x9
X/32KrB6SaR7xnfBqq8SRuk12z9H2jZhj54c6x/iW63jFz7+/rDh6ePta89ujc6REPiWoHJDPWI4
0A9j5DMDU1Bks5RIC6KihzlKu9RNdaNf24Ra1Tb9O2/iFzcemYEFg4r1m8FKgCgIdReVvgd521s9
dCFye43mW16sFCxDkZjXIpE77eaFBTZXLx2fV7nCqEzKv2D8STbU/tZnXMt9dJf2lnGogYqG0DdC
kuyv9a2F3iurE2USJEL4IlU3OKrRXUlxDe8KBDmaZrpx+8H7c4Ks1FhwEf38AoPYPWY0W2sgl9nN
ggKHG7H8CqcvZZpfDHdpBs/w3RRqe9di3Xw8/K+oduBpCY+cL2sp0Sbj+ojqSnBX75QYodMJOVHk
7TpDhkw/rf0NZpmTkDk8eiw0mWdhl47fBncH4wVxbOCAC/pIl2i5aDS+xT0kd/w2QblE72DPS3jM
S8nqACDE4VJBOlbF+Fk320bAJsy2zyxVHmnXjpW8iK1D9Urpk4S6jB8c66/0DpYHvawnrQpXxl0K
ZxqiXtMDhd7O6l0ucQVwi+D5IWuVeAtFcjettIgsWQ9OhozqXPO7v3NjGTO+RAJy3F/S8VWS7zU6
0BDjQlSQ+BZrMldVjETI7WCAzLUJ/2NMPiODqPnZIDpVwLzztt11n9mdaxGcGRSl55s1zK2I9Bmw
IFJxZJQ8tB/2T7a2BOkuMqPujohTYrIW9uHtqQiidWjjkkinm/msJwNSBHtfJ8T3dARKWW5xBELt
BODlV9GVfeUmXeom35cUfR/e6Dz/tL2j6lkq7hMR1CfoywTY2XjSzklaSflAVViifSP9uAssqlP+
mmsd7GUQqJaiD0mvx4Uz1loTokV+G+7MiVsQtRMXgO0jMAULgUhZuAfy3W6ikCR9cwS89pOT2C84
iI2Jr72IYgA190Z+GRImzmmmDCT2wN5QVS6xGQTrCbDOgz/G/KfhS1eyYTlk5mkC/owYOplP+kqC
RHpRaU7K9uFJEP+9RzAL4fuNMiNp0jRFgWY9dK4/JmuqwJkBPfCtZknmMHjQqHj2QDQNjPKwBQfh
0h34S3oOO8ug+Tn1mqsGAp7A20tKxRLgqF/Sl+1GZrIFkFkvZCEeD8cBxDhS0OFI98WctmFl+7U1
P3+RzcQACiQnnMnv3k28vI7xwX0Z1rFL/oX6MoViGmfFHGtCtL/Vx0juJOcGdz5gAUHn1hbb6/jY
SwXKCrknWidI3WYheuf4gVgxmlf4YukFCI2DWccIYzEPujiLUMDchIF1fTQtJO9PGwSUQAl2ILMb
iDCfifCsMLnocpT4Qh1CGkJOmBUxjTw4PCmhrqAuVpBqFcW0bVO9ga9/X7QaIkAO0lgfek21DTC6
iX0yCrp8cbmXANXZB1xb/Lz5jqtFvNRATN7JWjZWUxOh6MCBNHwn1zS2XI4hOhf4PQ++ygz9PI2H
MGrrht/XFCRTJSS10I7rBphIYnsapBwgwy5j1js7AKXLMqjwMYaoKRlcpx4YphO7wr6pQ9xYaDUD
L8SRdfdKzyLFWibC+u0qkVHbFZNn8Dg9EKqJdYy6lZJKFql4nDmUCqS+4Lj++DWyA8XOjMEVA5nG
Tp/zD6hBabsb/dqZA0LV6LznEc4ysZZrLBmBnTEBlPlZgP3zS3P9u1qf9VnquSj10m7wXbpjjshy
7aBaOY6fC95UEMsydo2f5lK73BMF4j7ZiJpA4EGqQHJDCZMOUa6R3G99GjEnX3F9KVboAsgAMq2Z
Y9e73aqeWCcYkqa7S1NYQQ1DQ4kWsBcvQ0IZ3ZMnMCgMSZ59yC9a5fV3r0yQsl/MJuwjbTeoSvrS
VRsiV+jg3EwQ2p4nn06ZAyG2x3T7ctbNrUGsLPaENDPJ1lIn1ZRNnUoJgScr5GW0i7CwvanCEgk1
tA2LTwK+YOrbROetgsd+zXkzQ7vO58Yk4vTDvA+PCnx5RR/iMzOqOAqc5Md0rQ02UJn37hMNl85Q
R2Ax6ZqNp9qTQWfnEjeXP4WpXYnqPJaSSdMdSr2gWuy+vTqeHjLJylacTSa6WAuR0Sx+EGkXS32V
Q4Ck02TXkFUN9KRZCLM5BGKKzNc/fDeZ24I2CnvQ/ysf6/tSRzKPr4bmZwTciPSmdSTyFI7DnDDG
5/6v6cfgoIxCBpHHcaxyChEuhpj2403xyCOJ89tZeAjdymhCLPBboKFTNgLzpPqR9Kzor25rTW2K
Pm9sZ8Gs8GltpWT5QVKujk/DPuN55zul0aUTOg9NhQna6qhwlg1oLqDC1vhDh9IWFHC33BMvQYD7
n3awjDtc6O6Rfr6r833WKZBAELhwRscsk1FJimFlw6POcBizKjMXx6aDLMer2S8NeP2ezHHbb0kB
zQXBkgZqsE6bPKNHMgcDqjEmK//QLyJ3FdJHrnvw1+/d7D8FbIyK4vi/WixF9RyTa8fHGfII3Y5P
oYin41oRYUytV4V2qdvKBiR3HYNsKppOE8qopZBHLtQJYuwCk4Gh7JS8UU4nNBRKORhaE1I3HNHG
22yu4Q8x4RIG3bjkRH8pq7IjKj182clGTH41Y6rjFKYdAOk0AnZbt6bIN5Z5POGlP+Nk54BOR+K+
xaxQ11leBsbRRiXlofuCIKvCbCUIHClrXe2raQwyv542eRe0prifvJG4tR7nZomCVaLSyF7Vq7T+
APeRuo3FjWa6U5Lh2WXP2Ta+4G8PgmHP9O208PNYd8t+ECq3ylYPz2anApfoWwvNP99xBqX3xFxw
+aCT7JSKBJMup7Hoy8zue9uNc/n+g9sNGo8yL1hEovFqS44/35NgsJZebAdvw0c51uma7nJ7hlyW
1VJ0ehK7oi0u6MIIcFJfSklDZHwHcJlxC/hXKiQxgEZYfimU7e/1o1WsBUptkCuoDcSU35HZ5aDP
7AD7kM0mdW9rmIH03qsBHcLiBdbUBao2fC8QQ6eTzZ1DqHV3yLYmRouWIQYuZjB+ctDepGIrPzqk
16KoSfZAKDvH1jIUUT4GC1o9DNAHN8UU4J1YdSVcHuhJe8aHW7Jeq8QGue4KW+JFrgM35tAZs+24
DYLVhsoEGSdwR+bfsIZEP0jUbtAEkZwGqU9c8lT+vXCxli3sREFlsEczrv5NASaoYlShmRyRScpy
k5khtkFQ+XG23H8+AImMHj9sp4c5vAUJVbKTYCkXQu2r/PH+MNI355rLVzNw1iMbqjHyLPmq+dTy
hg8N51CSDQm5WBSZ7Fke9IpLTOVjSVf9sPuaPVgBeGwtwbLuVd9fHu0e1wLRGEPzk8sI30f5S0Y/
tX3Z4GHpvl85UU+tEDpUfpHm88QZ/QdOiKeg0vPDGiM6hmk7syTj0k9jl+JJzywo5uswIdLLwtwl
43vA1xymUT9v4tyspU7sMZb7zuv42EuMW6bCkgN/YrAN/XVniuddIrCwqGgJuLUeR0JLB7zgvGkK
wfzLVrqO0hDS68s3QAuiZamcNVVjWc6MkveY+wwLkxqrKuSlkX3Po/4oSWTXTnW4XiRh+AcdCmIZ
WkePanqYI/5WoE8Lv3gPOCKKDiAvlXrVILsOTYJzdOKvna9WjGAtVKvGekBbn3UThfd/OThRm2lW
wu0f2rfFubUXOGQCeIUcpkOPJOEM1rtMetLP/FIh5kjljQhdVgcSgFRJNsaOhtx2P/S8/FVMTOSh
o3vC1/LWxYEdqfkhr2kDzPvy6uKvKFtCD39bcm2ZquwPLHpVCZ6iivr370wgOFzXSHwAhpt97dyQ
8fHDF+CDbOc4GpTLvAG1Sw7psc6BYHSyPc+OlSTHkdsQQMwzYyEXwX2GNV6zLmOMgpCpHHAoLWpn
W2cgYnPZhZXjll1hKc0zjNzyssVZty2i9GX7FFGPYNVO64tggJ1hErtXZQEycMiOmvOvlDqT5/eh
xkIEAD9qADAIYJnPYoSYM9Qhp0TzbYwPGEEOEWbByyj3Sn8Qsirb3VPWSBXWnrnTa/bjDRRqNL8Q
Z0qaKeRWCTFt3tFmJq32DZpJzQaGztF4RsYCaObNC8r64aF0kEQeqQDeaUxabUWF078CVv1aA3IH
YlcHC0P0MkzHXy8vuow6oNrTWpeB2i3woZHNzt+VZjgEgFerB2XCSoGkTiD753856O6rTm75tPM8
RWFQL9z8WjH5Kj2hGdvVbbPCKUGl1lLyBpudkA9MZlzLXJmBGAzcqSXWfX/U6lESKJ7axBRIv8Q0
bonAQB2iu6f9Dyh1kl/XmlILs3P8DgT53qW5H3hvRJ5lagk9hBDKkM5VG5TFUGZNISX0/LN+6Ztd
LhnbIz2S9MHdeJsngO/QkvpsaNvGbnPOVSaWMyFXx5ipGO2fCACEhrBBpH1pIttKpmoSnoqUBj59
JjMwWE5bg83mHyBd7VTpbEKIVc2PQ0yth/+K4bu6ou/qA1SdoaZmfR77Z/2W2dTtq/2N/krCZLuS
KQwpeU5Z6pNKofb+oqhUxT+E5jQE+ifk427F54XTv+apHRngJClWO9TMU5VaZhG7x3zniyKrTYSu
4iis0mTma2CeWnGMFK+q8Fhlk6mAVoMUULEvfozdOeV6cgvgZKaQwqeNxKLWYYS/CBEiz3aJTyKe
dFDtw2l5BFva5P46wKGiX8zz+33oSE4CHCo5y4IrhzsLr7zwrKCQtE1xzZaHovGWRnxKHMHPZowj
8OqvZ0i8uNut6VD0UWE/M5l3WN73L+nC/PUBH7kfbxIG0ckNFJ4OKYPko3wbkwBZvZE00/0rmAEr
GoSjmHUkQHVg+AHMzamE1YS3lGcvVLVub/yYjCEidU07DKVCzHKtvFQCKx42ZPBZpsSkemnWcBYn
vmcG4gnZqLfHsPp8r3RqjERrY4dKQQCTxnEJtaIYEO7ZDG7kOcmrAAtQWM+F17FLRK1TFvVnWAMt
qBegIit8rV3RlmYJVEbDm4KmTxnkHzlCiQVsN4fKcRTuzXCJ73OyWSRgbXIwlz9rhWR9Wps2hRZW
TCh+2ttGApQvEtjFM8aIzwb3zU0usn5HZmvNBwCZ2cEOqij270ge9hQg3x3Dj5Sgho1kUz0rhTTV
VkcJTGb5aMAVdw6dFz1wFxV+iSoILH3O+xQjVxikcQsqfoUOEbgVGx2z7jPmEPJFlv9yBvjn0hTp
D5Q4tFB5F2w4Rw6abCyIJokp2Isikz+0fE+jBAkOaXR1O/ODffbCmlqC4NOFV/6TwXPTDbJdHkY1
VHRPwLgT0I4GZWbQsDrStD/84P1gVbG/A1NQc8CTedGxELi6G+h1WRNNF8IQTJu58OVXNNbNgOlQ
Xzsr5MqchYnAfVOyXDfRmTK0UvFabgVZXyntxz6BfxJJG0h2c41QafnhZYAXPV1ZJWm+ns6wfRlV
yo0UhLLP9AMjiLwdfZ8RSYbY5nTfQ3xlu9gVPQ6cXScjBlkL5AxG+cIOOzZ2xsB8nmoHf8MrNCTK
YBv6N6aOek40v1iNj9ZG6PoTB25ImbjPdVJE1zEwOBS0I2JI+FHxxlNLAseO9BOz7qUifpsR7wk6
zf94an9EUZfcOkNDRvxltDhHhMR+LkHcYGy5Um4bcXEYuto8JMtKeHpIdVZUtW5qEKkNTb4Ey4l8
Cu9Yz4s8fOQn8zuZ6Lmco2Qnsi9Z+0hWT7zlzy7u8C/B4jaRyDppcBfW0tvwaiCE1pjVD6mcPWcL
RhYSpN3LqchEad3gYMcs0hrPT4DLsrb73mV9at5P2jO0qkcazncCbQynfOsHi/OaC9PGjHiMEdQh
ixDNu9ieQMZv7fxX9dz7r8PfatT/kZ9oGXKD7ZEZD2UG3/XpSfa16hS3L7vfLoTm5qpdClK5canO
+QbTwkN+1Nal2AWQwhIesdumNpEPsuKMcJE42NSLTiGs3rBPtfioL9c7f3n2ybNq2DgaoY8IhZaU
4WMA+5rbpJhOHP0KS9mj+ipnu66wa3oFTY0SG2EmQdc3sMKEKmcgOAGxCSCgV7p9bOp0NFDHDpSL
4Zdf+KJbgYTd8RlCUwbmhgkCx7LZwkelqYSt0BNVpnY4t1kyJk3X9Nhd3CiPQh1Ghrylg6bOyfIl
im+4Ak8IiMqTCYuxIyXEZ66ZHhIVp69j9BtWgrzoIxr1SBZPrkUI/+Rg4p/IQew8hrhjk22+zcLZ
/GH+K7T8KQfopSfCA1kqgnsm1ABkxVorIPQvDOzCWds9r7PWEVvJhi6qe0vz99K5N4IOZgBMrMw7
7/FMcb1RJSKcOxWWoYXJ+eRixSirZ5wlqLr2Z5iFXejNdCSeUWggMYjpoM/wdFEQAp+ylhKT/hvq
/2oV2m6l2s9b+Xy5HEoP9PicYrdJAJClAlcFL9D4Gc8cpplyenBiqVzkb2nGorYKITQnt0nZjiOm
ImdBMB57p2dXKYOHrny5Ge/e+si1hWR9cpqo9jEJ6HCGTmQiFbmbUQ4CQfzXv/ZLPE9f3r3W5G+n
k7HgkfM9bvdsolccrX89/oprOA//pSl63dmswn8qEoaRzwMmQa71v3qzS9PNI7VGlWVxDo8Er6Ic
IalGUhR8iDxQTf/y7exa0OlogFkIEpkEpItYEYShKHvwwcA1yIeKbbt+XNstcHuR4NpvzWwu2e15
fPcWPKjAo24Dvp7IpY9bAJ/mtdQsONyT2U40Rhk53MpLsZt8kGjgQ1XH4kp2jXbCnJgeOQOsGG7f
PLwBoXsVH4dc4yUYoRKhq6iq9ZXot5cutXneqXzNlNNmOWUaaSgHQVIPX8wknAL6d57B9b5brHCg
lfAqQZSP1asycSd9CRaEnaAo8r3FMiUjTthwi0Nyar/4ve9xGVJtSIgaYJY4+iOKAKOI6/iNc+HH
cmk+AnzpDSth8punxLVTm+gChgx8JA8nSC3HvYBMMerL7TXdgI/sGzbCB52R06TYbeIrUlubpL4/
JyF93HGM+AOzSJzZahboD0Ts5yvXgmf7b60u9fSxL0fPYm5SVHtqOhrHoK+qs9fSeFECQWiVNnFJ
wF3oH1feNJ5sZZxADPeLY1SeHj7/CCRVD5B1V3rlAZs6Fjn1JCm/cZBpl5vndUXQNiOGBSpOAYaI
DGKq2lg3tL1rLeYbHV0WDqyJyaR1BnRdX4QQw1CkIzoFdCJqgTU8N8t4ZQhTsHgzmWldL3oqENlC
Dl7Q0oUtsfwudQGTaCrfaxlNppMetA4tXxvuI44jZaeNBhr75Ql9MrJe2Yitv2cUP96YUjn5hBhX
ACz/ecREejqHaWEbnwJMLW52/fsTa5xgckLK5PyQGUbuap36TyR2iMmD+i+Jo6H3XDeR8NsJbz34
KNjc8CqImgECIDWSeTd0KSDFysIpaBisK7Oa/8Nbz/AhccfPw+Msjh705XT4hGB5R9Es1BHX7mKd
DKl2dcxqhUjdCoPgUj1m44JjAlvU9CQwFTns7Q25HB0u38iunTecb3D32MbeUikD14MjK6Wvc2RT
bJrRAdKgGG2quJz1u44GMZAC2tUBKmLxhOZzSocBkB3XjBfFXUldR4HCjypMOrAoPMNgbTunXeEY
adx+9BgtJGQ/iW46cIshDqCwlwvhtsCnSxxjci0KY+/n9DqViRB+Zl5McSxR8sYp79GevtmddWKF
ixYFcidW0oUWgxLa73qi9LNcefZKqtlEWNKSpd2AT7qwjf6p9DstwH3C6CFImzr7CdF05L4Y+fl/
Azm9rdx4r0DKlQBTlWfxyrkkKxJKmEG4CpLhE4dlbJF9zgqtnTS9+AKC7L4pLr5L0pimmkd7VS2g
S7wVpik9gfHQ8sMCXLHW8l3MwSFJr7vqDY2+xTSsz6FtfN8wXGe2mbiD3cZOAD5bPcyo9FKNyR2/
w8Mt8k2DUljEiGPTTHIU1kyKaZ8e8rdDPtKJD0qK27kSSVcABTThH3nhzQUyKO/sE0WTqyv1cGCI
MhuA+tWoawb1oLR1F5R02upnzqewXxKSGswPYu+MAhVcXGcaLLEVjovUcFEjOb8gSan+0cbEgIM4
xp8QVKqBVQb2crB4+0LXNK1wbqn83h6AnmPil9qkL3PCdAa4pgzwQinV+Yf740sNes0hyuO/Ijbb
hYsxCf62duZGJyKb2blLZoJmTkv/VJgWjIidh2n3/jYf4/rzkehjYDc2yezGtqQkB668o/z6x8VO
Vp4w14GpOtjZMH5LQezXqCnZE1h5QWnpvKlpsFVvtmW7LDCDJppj8r1iaTdJE4/nqAMW2TZKsgKh
H+X/EEoMwMzmsZkwK381T0KFLPyWZrtRdKPwGdKlwzJAbRTpY3jfSBzZpSaFE0Oa2gaZ4ZB0EVjf
GuNmUiCmgdXjF49l6F/TqF9APZ9I8kMrpyH/OeJbKgIMDaq4Na42UAkXGzsKwAQqfAH044JL+KB8
L+HGc6eCv2TpDk2VT6w8Hh6O5QlxL5m/Y1Q8i5xAsRLcjuYOrTNxOglZfNqO6g4PdCBmE/1Z6jMe
9DSKe7aamnGVoLW7NsIDGY4JABJbIZe5NhjC/xOUnB1DVuw1FP1CrnjGiAiJOFo9uyHeRW6pzEJh
G7dj0ZJVfwfRIoWW8cJizgIBLfeojeUUdd0OMGz3hQpAJ9OEF2nlFos5Z4SkP92S5y9OiiKUo9Sd
KPFIUJ8y5JoiQOKtQLLo0U/4o/pMW2ue4RASoIbWD3D2wX/ER6/dBxnBju1BD2AQ1hxiGghTx8t5
3XnP1EUj7grewbKemlQ5/0NHlPpEOY9fq5ZJl0P7EQ6gb+huyd12igS15ET1IMplY52x/IbvmSud
MfdgFqQB8LTd4j2XvclNT2fK75jY+1EZGKaS7+xfZ4Mi2tb7Gk4IHjHVwcv44p45RpKysp9vZpZm
5f0I658/bsmR8pa+Ti6JJnH/Tz1YxGc++FSGJUlp/zhE6kZ0iIv0xNXHeRu0m9QhG8U5yPeFFLQv
cdDp0STYRZE9+OVOEtMUGhnOngvacxNP7z9k14frtl6S8xugX8Fyk6BWIAFsspVUi0KLwNXqER9v
MvHCigrAlKI51rU1e4gRqZnVAeNWMDokwM0pvq0B7XA/2bsf05N7F540GzUqFPELmySHNXl2JRNJ
kV/a+TEarZG1FJcs7d9rScHRI//tmipbtJf/P7eOBVf1QXwo+zJrgX1s+y/O94sPh+K7wTSQvsnZ
yqbvDJCaHvT+im7uSJiJ16i+477EzC/6r9hLqOQva2TcO4H5tOyiPT88ulOlJw+GgSyS/Mil1C6G
straFlEWTJ9reQoZLr3Ip8miC3gyJ0hSPIK7snqAdg/C+N2fv7SiNYKgdOaxodDSc4OTbJw9VpbH
E7KfgAd9duw4Dg4RUllP4UvGzjs4QfOMPZrsEimrw7cXKeevlV2/e72lm/3/fZ2ZNBnK69hmCnef
bRpb8/czqcpHrrhwfKLc7dGhd2BseiGk525jFUMn2Ef1jLdmbC6Q2YfSRQBDysjPhjdHtwbo2gFC
ECnwoYBZ0WjjtJwi9VMq3bUTc6MGbO3UzzRGeN1CBOBjHSD9spzyp0Dzk4KqE/XdF0inmx1msNU+
274+L2dGKIuFllVvLr5lwWzgTSrzVNN0Sn0yYwakJjbgPpTmQRp61viDgyWcnslNntaruGGZLKto
L3g2tW25ocFxzecCDGXU8MLljk72gcEj3uVT+3sVMddzLg5Dmtc3kOEhHUTCYQ3Cb52M/Z58+WPK
FIoh8404lYsI0gqyTFVCRNCsrfXl9JtJ2KatEilUvwHHQR1gD0qwLD8aNfHEe/kQHcZBwJE8mldP
AdsGMOGvpgFBv0WNjv7HLYifTptuXEvGkYztxSAB48g1vHc+NqEAMzLtXCKLOSKszyRii0k5FzoE
EAV0LW0VLUVzczOUOExm3kDf8O6ufv9toY6o+q24T9tSzHnYX4QSzpEwRjAhvCowPxgCgy6+pklI
UiRZtsOBZEb0o4LZ00DexWm+6m56hUzcuNUzXASZ00MFaQ/Q+TQRmhKbGDIvUZQr7pT0JI7XNHNM
gFyWOfhRFp+RlF7FtX9vDAV94mH4bCdMUVMw1IBRyCKE4beg9m68CX7MQ2TxCmscdlMFK5zPLLgu
va2udxdHjN7BCIFljNFdc5UVoKOz0kITmg1b5Lc62yxjJawc9Mn4vnjS2zVhjZEMeVqEjFDgNNs3
cHUINFcPfvzm/+NpO7Zw+qCl0hz3eBd7KyCFT2CIalP6vwOh9/2uNjz3B97u8Fvqa9CabvzzOwxW
pxIuVyyo/gRCzWzgDxA65ZewbWQceMdIYYe0pEP5N26rWFHW/mSli32oNwgSStjFJoeds/fBjiDW
vTXvg0HRgV63d7wAl2PyEQRDxN0Z5iydSh2wMbqU/KYxAawzADocMtOaIdZL1Z/hi3p+S6GQeFYB
pRdWmCYS1EQKo1AsC49ArP1JxEoBqN8KpTadLUosFxllhTtkfWrvd7RKZfIphHuGUZyTs1h8HQYF
cWlfqHOo/dx9SC2qQGbTLsLleBNJdbzJ30Ickh9sCZ38VmsIRthMP7GesqZF9dhoT7BEImuc/PVy
8HvZCUHOndeheHmVnBKYCgDdQPyhhIkUytabA/v/YI9+GfRymk03O+gOKJOJhncerwKRdwdRTgSE
XIldZalBdYrWuXPPRjsLqwC5eWS+VfsIVjR11jhYyFDh/1eavBMYIJkBfWstVM8d5wGrar3LG6bb
HUyfzn9mc9kLv64WjnqLbCaeIulfCubMtfBE4PoFvpCzmQQADJXg9iEiyou4HgsfOTrWPrvxMU5t
iWYeab2rQJ43K6S4N/lQoLwB24KYRpM5foiLsejAlzjseThWo2ueURDT7lJTakLyhxMIxyPtzy4B
/tABT/oAlpWBGE7LhZGHhi8oDfsC/1PGkn3FisvnFF0/NamDsG4ZFxb0Ktph9nOrgLHYp2Zt1Bzu
KG8XsvhOIwcJFLUDeXvKLIiyoAuhSMyMnkRHIdvRsDZAZYKMbFZ31XQ/Ps+mmTDFvO0pUFcxrx4p
grM/2dbl0L8tT/VaIAdXC4/sVuXXT6cr0Nkdjrt2GFY9oWu6oP/GrLjj3uhDxcgNTa6AE7m7m+bl
W38ELrV8bAeLCDTu+HGaO7SegK1Po8sO+7DM90x9r/UBomEGQUJgxeoqmii6vszKhfpPqjaCltsX
l5Aq5PhrzezD38My6O+qhj95JxS6HDyBOWbJlvkSW2XXVW9cPlAqVESVbmGtxtc+HTMkXya7UwMW
w0X4Kok76YhVo3Xi5c10DKnrrDAZhAmbAaaJH2y5t+e7nOVuhgfwi7YR4Be0GljaNe4zwiwZePAI
Qx47mt4UfHH4U6xcAsEyEXxsYTMD8C+QXT+QJ5H8hmK6bYZO7ufv7DrvNT6oEh5rF54H1LxxJ3Qq
TPwA8UjPvJKHhRFdtAOlQ2QXsivTn76dOGCsflusge99u0idvkkzhNlw133lGs/non8bYdZv+CX6
dxGcD16b/qL0JDQCAPDNHHa2DrJZXwit9EnZorEnU0IVtXCBHC17Z3F/Rgo6Gq/Ht1yFT8Sx3eLC
hZMBVi41w5YM+mQW1StVEvbDUR/ytwe9DIuLl6aeE1ZEXx/7PILBmdk1KAw8asBVnXwCfKZEnnCG
zTx/3e2GnqiWBPWBCjAQYrhYxk1dML+EXfN9HQOpxwtYhI9HIsyzjPr4CjYLNrCHmajA2TZhFZwN
5vhinwYINROyUHlz+TVOX/Pzd0o1hEDOoaTBO3ON+ua0q+K1SPm6UNRoFuYub5vVQYV/VxiMOPst
VGmWuyOsR06MHwvSLzQmtlh34tk8nFCQ7Jz6/u9AY9BOZPq7ECcc8cd4vpSYSNLW9BOnTWxd7w5u
TJNAL5s4SbDNsOvfBR8T0LNbMhYuw0YrxSh0oEBpkTmTxjk0dmDFJEkyCAO7lTOg0Fg3RH+ijIxw
CXR9exLETVLlLuMcE/uVI4+wg2Z8s0tw0S09SHEoru/Xm0Is5WswkEWxD0U4tbovFE2A7c5K5dnC
wmaDS2Fs3Ig0IgCwkO7slXuDRQ9v/ica4rbtpehnQ+sOb28pwZvK+Ue7fXwcoumfN8hqjqThXQ+1
2eEjq4LPSirKgcuphXZumfUa1z7sFO9q9NVMfyLOsE7HTf2YERgpa4Fl8zGvbzCHO/seq9QuZMtV
LEofMYft6OhYR1OgUvIv4dRBytDKjfVnCC0OU8ngBgdwUGYiyeLwezsogtFmNZ9q3VEkETz1XUDb
nNJe6MSOgN76b55H31gB8EvlZBxvcvmM0VNjvpwIj2OVzEmU4G/CHAhI8NTwxoeo710Xj1hA2vFA
Lyrvr84b6+/pOV63sBgOsJrt4/6zU90iorQc+lO3j8MLvkpRtHXZtH+j7b8LizYSpt10autEVl5+
lFwuQnbhDexEDaWGw6YpMnvN7/FqznSd9blIdbVWrZKbRPo8XSHH+dKRmsY2vZixN4HhIYawGZzd
kdGeBDCU9k3ux45D6vCoU+ZayzdBm6uKW1xzuzL+5YGS3YSeOt6OdriahzMJqJB7bjIWPNmXBVFl
4gCRTUMpQVs5hYBATpFef3orO5tYSjU6H113Vpc7lg5oKicjhK9NJGiJWdVzlyN1rngXuhHzrYe/
7Opb2YxQdo/Tb/WVCmNVpWjh8h/QC4fQizIg7x4nxdzImZdx7iEjiPts2N2cB3zVaLYCxczYK6gJ
IS+h22Ka7QgOsZONGLO+fJ1R+uM6am7MkrSHhOekWWs6EOI5gBy168LI+ATSZLHm4NdkIrXFKCjq
lU7G9bqcRA8P8QllMh6MZxuX4PyBtX52NSJiPhK5SGeM4tK3iaxHr/9F5OLEkgT5PalGPIo3U0rb
e1X8P4jDpFaZ6GbmQ9cDGwsiLc6sHDkdYOHt0vapXTjht2vwsMrMFEWnFPjxqZZA2rpdhcMLyyeq
Ehm+ICc9+DKTuEwrGfJR4wX8BIduSXikgv9LgFfuDPaM3HmiiPJjgrllx/oMfzY0wIuJlk7YICBO
cKDomQKH/XkdGudfss5DZObtvpjhUFiJj3kT0PzEPSAvgNjy7Axxfrz42uUFZCmR2SPDgItZoRSm
eysWst2D/HdgXXp4fRsleJTs55M3vXyev++iwJahHFOpQ6cd0foesrcsi3iX57sx6eJLftazSWBU
Ke++Eb7u5jdiA2/x75tS/JyOsrEK8C0ZMHasicR4mZYjR5yWEn2BO2ceznzq8HeK1mOrCjrSOIrS
c9F52tIFVLUXZoSIG022ZmxLMsqut06Vml7s5hjLk7x9Ksfnlmh9qDtKeZU7DatcTevQxKsd7SPh
3gP1fQReksRYH54yeIRjxa6VThzl/tt89x0oE6x+fKC1+B4Zi/KdFtu6ApPHoUcifJt8n3tXxj+L
r4EGCK5175BiLchZQP2za6Anit6kCBo6eKVRvUiLdg7plRO2WAEOkeMizcU7oRDQU6jQwSnkGbD+
+sC+3L1sW2+5TbJr2k5N3G5ncBCEBUlYK9qYt1M526nNOCOv1SSGIufkRhqiy68D9he0z/f9ryXj
gK1kX1LshezbLAac+olYeFMbVkLWo2zmI/Swsk41+YKZRKNAOtWmbJCAXNYxH+odRPU/UtqAlbVb
4pcHn1aCwZYDlNeYW0hgEUtyIYr/R3rR/x+LVdWvcye+t79W5NI2TPqjFvnTGGV4wvvUCK3LWVDq
3+m/TweNTowTe3T720zfW81HK+RGFtW8BHXsro65lpp+mVGUjFKGrIjT1oFECXxn01mrFtsqByU/
9/P5XxzSuUovnUNztZGzx36BfxOtssPavi57WvNiFS9wZ63teawC0gxsAyy2K/BTgd4ucDCZaQkM
IQVoKCA0zcn4kzaoJ8xTO5kSizLkuJycPPSM/9zLzAH4W9Cbba8aYPTA2z+fABwAMdrEZOHMDqAH
BNAGQ0DuCI5DaR803BJYrSPZuiNATsLHyOt/6ODExX3jM4HMZpQC1prxoxbbfbV7KCnh/Fe/KVyU
v4hrxtBkxD4jDUsyHbULlwTM6EtLgHmML1hXuoMS9ZzNr0FAy/5gJmgoVTkjOBbxpG5Mwnm+CO30
XUzkipJInD7PWZ/j1wFvD6aV42rvjr8oLNIdi6ViblsbOZxNw2hGcDthfHypitFEt63/v6qKQv5Q
hKENKAk4P9poAU5q8Gqu1SrsbUuK73+r9f5RA2UD6o8JN5FOKh1DLWOJ9U1xZz8SKsGjCIH3ox7i
Q7WFQUJ5wYnvz3kHap+wLf7TYYI0XmTt4lDFcQjESI4Qee769S0QxMA+5GgxnffOvLLPTdWi81Pn
8YS6ii+rEGmog8gVPhROHkrpxQq6KP+w0yLjvNKavyFs+Yw7X2j/svqBKPrLJMaRj4v2VQ/Xg2Lq
xkan0RDbQdjcf/9dfB0Rsf2fx2JfsAdaMT+fWxr85oNHKX0AuEcQCVMiq3Sz+O+uDtpxxoPy+zWm
VYUMLBg3zaU4fckzSgkGQni0piLiZIWk8njVwZUtBwQkK9RgOxPvYCMfSrDOCvJ+84WjHVhJrRZp
3yE5h4MAontkU+FHQ2eb/O4yqtSbf1S42o9ORLPNXW2IiCWka6srVJfXQFXKDqJrq+NH2punJSUB
AIO93wgUUMS6l4rj4OjKbEIFQcUlYFsjO6lbRX3UFlPIcL9cB5RaUUuwBmN4O7Cc28Ybx+evzj+W
Rp9CdovBazso9EkB7N7yg4YlzQqVnElS7ZtY0njteGC3FOIdNLVsPMC/LfBsBybbAh/res1w9sYA
l2Q1MqB7uHSkBB0VO6VvGrAHxWFviOasbTtl7rHjnNc+1LXw3iy/wG13iM2sxafgwTql0O8mM0BT
h+dODBbhNcNjFPGdSMjQlOIRcSymJKjbReD91/8XnoizEKxPgh0DyuL//Hlwo4o3lI4nxH66WZZn
16qnJ9ssl/q6kugvb9aR5F4FLAj3vGfHK4IUsmAe3QAwmDl4pd4531TUBGf3tcjT5RQZ1aQHFJH3
vzuCQj2mfNBxJQ0hwkTg4LiVkvM2YnH1oiGdLFI7XEW2eK1WOqNYYUzLuFgEexgp2qr73ANkLvsN
fi1BT59XhEMf1QCPKdvZh/NvOcp5vscf+CeCep6KebKa3HyfqXUPbum3HBWMJcJfgdXStatx/SRq
bzRCKJXac3MUgbyT61vVvzvmq5acr7QJiShuD8H+8BsOCEvm850bEEyTyzdjbFR/uhCbCaCma3Ms
7gyKai8J6H3sap6z2Vjc+UblADXeRYBITNvLqfQ+Jpv6POXyHvwGkW6qVnNiueKwCUjkFMo63PoR
mTcXtneUZQ0WpMyp9Cscudo51g6W4upi42MVEesI3a8+YAAPHtbnjoQopZyfcPqYbtK+hjVtKs9e
X8YFJ/xVE9IhL9MyUXJTCUSqeViv3Sdrbrg5oFZh3tNNhPfn1IJf7SSMNL7KC99G3qe82xWpTh2m
ngf1qDmqSUjNWf89a1JITevQk3r6/SElaHMrCWTSaYDcJyEdi3OC6BwOzlF/M4AdZo9VRVgqZ+1j
2ePt5fJ6p6+BSymBx1HzwdRDY41d0463kdIZ6GiVpz8nceP2qfMRrY7dAvEmJL2suXeMX2OkDceA
JSffloefz7pHJy5LNWNj7o7i8dVyHu3PwURLu9LXGs17f1PHXIWbFqxmw+QHcwp1pzc7GFl2D0J5
79JRqAXBFzzYbOlMm+O16/tQDen1KpoB3vamMYI1s8F5sksjzPxR/obMB98oZdaxneh2m2dJsmG5
an5yKdEDV17jTj1EOD3fbxF2NkV7+SXkMHctFqaoZsMOU3FeuSlRUxXaYReUtcvjCYVW4LBWLYCP
jmXmInuh+GvnojVoIE8SMsFzG91mocE8cbARxH5U1B59Qp8vPw9Lgscx4t8+2s4koI+jjtlRWB1m
R97ia3e+ECzBG849nfk5E8Sg+sU2abPpaDDjDixt2pJ3FEPt9+RDIjskIsKOYykE0vJua6PrKTDR
Aaxkrt8jFLvHkKWbu604+91LLzyA0kJIePlM/9tLGyvAOSPfnwTjqFb68MORCYuyN93AvI4KMrbV
WQGFuFGuR7zhf+tAqhNidvvFlMxNxlghMFCS2ACbQqYE09id6sDD4jpgXPg+ORNjonOxxud4d3ro
2qq/UCOZlqYOb1G0Xqj3qFBrUGPCEZRTpWZHt6T8SB1zMKqHeXjXimG6MU6TNRestJAhsBkA9RDy
Kg0DYBWmwuiLv0MLZU9XQl5Ig9nuYENDvKwFSTrftct6saoHs92tMMTdY9S003eJMmqxo4oMit9E
+RrB9rnpG/V7/QN0d8av/4wtoYMZRlzt28ilI+vqU6I3Xxm58MlubSnAY/kmxcs0ysojKQmZjtK8
AQex2IK61gqotzhL4odRFwSDEJRZ2QRj2idIh7ZOOAfqqwChsBcABpjPRKsRVRDdmy/shz/yn7OB
mAPEpEHsZvE/b6wD4cXKZeCmQ0LnSipAgSUAwBLFR+SgNCkRDB3XeiKN8eNJOWsy5zfatGpUJM2i
/TdNY5HwaQNVzXJA5W3336Kbjy/T2vUP3z9A3lZ+Ixa0ZXm9vRk5E0pzFfUlKd83Pb4/6e46X1Pg
irA21sokAsAcVcKPq6UaA56R3iv3QgXN1jSfAhO8I1Oc0vyiYHIWgDQNcAMnTgkqYCp30fgRaxC6
XgLKqq8v/8x9EkaOIvf/+A0xwZUI6UYDENuSvgbsBWLzZukb5lBA7xU7WVa9InoB0pO7Qgb2Va8a
mBK8cCOZOZ775547zSIFx3Gb3oF9/Cgve0uFNtNCWuxj9LSHbE1Sgn697nPda1fk7I5mbUjWoMWy
kYSstPf4c0iTgjzcH4q+mLIPLK1xlOR7I61i2i0o/RvHxkcXPx/HSrxu0MIZIHWbUr6+EhLAymkS
4wJ/GxroP82+RH6Jq62AStD5AUOdLcUpn9nz5t4AmVsL0rgdA82268+0OKW1iCPRerDvFEewfd3X
MMFfKm31+ucAc/H4+6apwiXCtJkftEfrB8iowQ93SOX+1ByXtbe8ttHuVndGlx1XDNBlJ/PpabKL
ePzbilQ3Aa9bkNPiyMAlbTxypKYrnvYNZvuYapec2xExYDP2Im3O1wyrhQDZ+7U7bNjfxkai0rUw
/wi4RiRuE+21QcWSuCo2Kx6USQPT7j54Kg8nA9QMmBoBSBv0H8r04oYQSXYUN+3tITVeJcDEViLM
7KCdt4bQZFBYAe0tDsvGG1x/JgoEAI0yCBWl2jZXO0WSXI5YCC5eZ83YFKk+0m3waQ0YuwjIcMd2
W3a2Wad3HTxSqhBspRHSunXFo9bJF/iGghLysBTZyJTj3/BZib0T7UC3bCedqmKvZIeWoX2/n3bJ
xCtg9cfmj7493PZVwzFN6rayoHIWYJhiVwGjKgCShrtb4HOOzRVcx0ZTjk6nPDwUCJuFevoYbogK
bb414tVEEzH0Xylwqhp3xHULmY5OeY++pylv6VnVsNkdQMWBYGCyU8ZyO2mTzcPqN7btK5w5YE9X
RBZmxsxiT0mGtqDWmdXXMC1kvFwGS7PUWvdzSpv+FhC1+gACw1TpimQZ1pKxBzQGbhTtH34GkOh1
xmxfA1npZPv9wgtRgvak8iYWQcWe0YoQqJPVqWmbXfcuztKvVL2hbfpF3w3qJvk18K8hfH7hzitX
fIS8Z+L3jahYH7VDS5SspdRJHSmJ8OthQo84cPuyKHsjrPm/ZUiKxwNXQfm1dsokXt0X6rws4o5G
rmn0mBWhsPi+SuMvsq0oyg9bQT0ZzPz2ipvfVi82etxGaM8B5h2HprjHRH9BbfUho8oqeddSiWK+
yM9J+S/lQ5cinG1k6p6RaphC5RU9TnmwBI6eu5ROKMxvSYPn8tbpCzuqxfZHkEgnki1z8rfWoIHb
AxQ4AQdd7wp5dxsat+I23YZkdfeEW7hVwwbqtev9S7bHMq9yEjKHi6aBjgzWC8jPG04R0uACYt31
THXh2LjCftXHqat/LjXtoxOf/M6fwnE/63Zb7TKiY6OXqqT3UFFgu9upKHw2+H2IjZMqAj4wsOz3
Ugoa5hcAuO8g31Y2GvD5Wm5Vw/OnXc511FKvPu3mS/KbBlIWE8jYRkWSo8Ku9dZdjeuV5u7zxIKp
vS5zZkFSY49XwtJDMs4MsVJLXf2+L9Gd7SP7JFDpc9enp5JKx6o00Hx5lxpqrWtEAu9fk/7OCCLa
oKI6oVYfvRXWiNDhjyv24qvXbh7Gc34PnU4As02ovREHEU5sOwAMlrjXZYQj79uBuHCdfjSsGW3N
X2h83blzGrTwfC4UR4dMeDRaxKg7KkznpfUAIt77/WuZnE1DXzjxoilAQ59X3G2TbubaG9hy94bs
A661aQEPYjIGvKENoqZxOw4ojR8Nl6UrUrOlv+aPNdvghesJNzUjvrbpBs0XpD6QQ64aRZGq/O4R
T0IvBK1/YK8OrLHJkAd+GDlOC3gTmZUCCLrOzT2U2wpQbNUhXVZAdRm/W+h3Ts73FmxUQ0cT7b8Y
QdzkPxMYQ1SrRRjvnr/gOvL+GOfwVu603JK3O1zrNmeUAdYzoVXlePspDp0K7kse2r1wiB2mnCWV
e83Idvhe99K8qILJFOUUtiChlUsZKaqUnR/Ogyh/o0YwEUfBK56fJf7uvp4yFxPSqotY72DtxIw7
axFKXI7iq1KZv1YS3AW65XJm1kmT22Y+y1ric6jcj1pK745CIhjJqEMbaZ9LCSTUOmeAed1FPTbf
M3l1t2LsxP+xTmDZw0ZhfOh8lPuptaxYk7GjBsceRMRBR0GmUJe/TnMbsFWGqvhxU7iB3LruCWo6
grvzMN922AhqvnDlJKHxEuHoVcIGsiNXkrkYQeGreG3qSeTfI0cWfCJq0W8c8Wyand3N00b0qKqT
sZYiSLaylOcxPTaEaJp3r/aPwBKKs/ILyHoVrwjCY/XAgTO0m2QDMEo/tQe48b8kYK4J77p1ZLqp
jXUFGqKZvf05Suy+pJFpsXrpWiot+hqcV/vJxfo7QaRKawmGh+T7dge4nfFp+JsJxr5Em4PVT7Md
2W4Q2KT92kOp/xRllPokqWtL4T1u1ttswfLB/hTB8KHvzpPTwCbCFsVZR0iG2fxy9v51hj0PUj88
sksSwq+bYpPAEfn7wfeiqXwWkt0pbrlE33hzdnEfZxTDLxUj3902lTJKE+6Lf3OMi/9S0c4z7/7R
WGHSLOBPsxRSbyiNCwEU7JV9k+4uk7xSjdJdmNZH/dUoq0SSzwUqnv5ZEP8EmyKF8S3RNYZPwDoz
BaksnTxtHPq+jKLF4EC5vDceLMlkaQ5GldxOR6JK8xFyOnHodaZlqK/mIxcGidEL8dkJGv4/DUWG
FTFCz1liWVqZvBOUCaNbfHw9BXJgmagMSDcWyS2p/f/jf7qVLFyLm9GBJ26E1jWZ4+py+ONG2sGO
vaObVm9MuBPQJI/Qy4O+0IvOwcH3HTLu4nGUIkMCP4RgOUCZeEG+eElI9rJlYA6/MbM65pi52FLJ
maIMnbcIslRNxC6GFe2KkTtx3dRcvjj+rmYeBvI7nUwUup0t5/+wgM3pMxulyofr6KCnwZppVcy+
DGsFimmZpd0ppXnwdEK8vaCNM1QtLsWg81sbnRPM4wk1h013u6nrQSX2i1+Hg27wvQ9MjMd598iy
T1HxI+vG8mlgVACcurixKq1C2JhsWIbdDtXGMRXf90olcjpkj4R5MzLGvQGVJr8MQi6hoYn1iD9V
kLxwqW5YHieyCB7wHDpzCeCubjhI5kbEAb/mktpUWPfGbLeLZm1/fhN/NKTQb0BMcf4JlY8phuCj
FitjMjwWdm+/Ew7T/3LKNNgeN3Rzgpu63xPv+FPiivwkjFIUDEX6Oc7ip1k78nXmq4l2czOez/Va
N3TXH+r2tBmAEy4c8UQDPumJwW7pZHkt1VxOSgi99SnqpPuAAYS8MXSKyb05xxFmy1E35xwGWvzi
hSFr6JG07HDXTY8naQ2B9Z5724s56cKDCorY314xZ3iOxfzdf+1Xpp/SSD5q8diTQ6B+T1PWZUA5
lgL13bvrg8d01BPO+Yz/5rqmhrZhoAb0YssduNKNMhJ7DIrrdQkkigsJjVKLk0prl6D8ts7SGK/z
1HZpp7bggEvtxkOSAH0/fnjlEkIuvrwfezMkAyhbkZJ5kgZT09L1rnugkEZDuiBG0MDmhy6ygahD
4tY6dMyfgU4kp0gHf2oumulxq079Tvq5aEpJG6aqmKQr5mkMgN3VJ+nkp6uJ5FZN7PZzN/gxga2m
VkVRCLZssUAj3A+LYtIIbilDiwP2jZyZ/dQOlb4Ig7voO5Wj3i5BdZ8uTXQJxKG3QqjAs8aqIZT8
EKm0lL3WZub5cjhmYJNJeZCuWQ9pZQ8OBU1uTeZcC0f39BIrNyPu40APHK0jgPp8+BoSSATZqKBz
3/8OeEIaR/mAl5arsua4N6VGq0ukrdl763GzVpbcgXSaGbXqAYCoLH66y9KOgTBdV4+zGugGsN+L
S0lwBEDJe3QFF9fAXOluIxvFB9ZorV7bUU1HJoD1kBojciuDp/M9sdwry1rkLZZSd+q/AkTSJyVo
8K2v9tcv143LLlCi90VoaDq/sKVrLqsBJ/cyAMMjlprbINNteSzcXeVylJWIAOQZu66rxvjxfNb/
cQ9FOlGy1kV6BP3j06uoW86prX0sewrRr5YienF6fPdh6ypQTT3L3Xod8/FPBmeLhT+FRXleM44q
n25oHN3ireoe898nq/IsMMOVags3qHd14Uf0JFv2UFyJMyksuwVYiRDfXuZEVIQC3T+wJKVGIFdk
pxVglo3UfVVrWpvl9CwcA2K5HSPhcJju6RdCDlvyVY7gzVg9nIDMqvk9qMVVO19a3NYqZKSWVFRJ
c17ocT5NWSmEIiQVPJnAO7fUJwpSDWYDE1PDRccCse1s+/qU3P3gAcEBGDl9qPedNg2kVvwycrsB
t3kM1RpQzHrUeR3RnZQTdyoDWBQLi3j2onPMs439gKaWKl9PcfKJZfS/giMex1uKD/9FbaYQGp7m
T0S6KroBQL5DQF/XOdWMJC9vX6yfGroUcKrTud+sYryXYOkrLcTC5rXxZSIjx/rsOdVMNxoaW4Dc
6MnnHOmtXzOphVnLQr51OsMsoQoZNoWlEcHELccAHy6xoMosmwHSCv1/j0sxY4+pkAvNlCKfu6KM
rx24at24kup//ekrflBfwxL2hVQC6T0O3DUuVdvMHyGNqbIQjj74Ig2Bfhn0txv8U5LtdF+OVemR
bYIxgXRRUXIIm+dJNVFsMRbWjG6qg+oYR4v52WyzwvW1ScgQd0FjnA+gB9jzVzNxU1y92gPkJJ/l
hhboBGuUeBA4cUI+y0Nc2qO6tjNFAUFKxVyLjXjOPAb6ozclzwfpRxDZCGEGy2TnFSHIJu+bnPNe
PGWgkjeL6SGl9IErjlW47tl/nVXfxmVzfryqWGIZ3b2yBqBgIIjn6zUIS1IPUaFtFPL/esL5mCz5
7BAmL+mbOqnNo/zg8MgejhaHTQxYS/UsXC0Sc+KegTXbZ/8ql8Uxl4Oe+PG/7y8p2LLNf9rjCF2O
NiyspCwgQvWp2ScJsBl6rRVpXzXmjvNtAenRjFaB/4mk0AyA21v+ANvMH142FvzT5CnqtjAZg+ev
I+rD/w75xA/iXUpOmG23G1/Oo7lbagoyhRLS0NrdbIo8kvMywlz/uzP6kvJZJAbxoD3bhameNM1c
El2oiyQ+pPCt1Vjpj4RJEaBHXhnQ90IWPaFLGjgl7O1p2fGT5MoDvHM9zL9NG5XnBAOVlW/OF1xS
LRSureRZZROPUm78VoaSvaZsbacU4i2ZN4gxQxWLycbpTIrQtelzmz9oaybF7IpQ8/W3hu3vgfSQ
WZplRmLv4BrnEsjh3ftFDFXbYEdfKGpmvcnUZ2q9XAW2AK1PhaQlh3HodApSMMmkGRkcDj/9j0gJ
D//++R55UXUxY4yuNwXcoLahMTIPWqcXsKOPlrg7w2dwUqmsRU0sHwdEJUYiHRetFrXaKRLh8Sm4
q/Xu6vDPOcbfB329+aUJw/2s9xmLenL3i41FmSYhPLgL0ildro0p9pQqFwG/SCakF9XRWJm0Klnq
vC473e0Bs1PAbchOy7WXml5kQ/tfes4jc2t87z/yaIHDczFdC+r4tv48Ff8NN1Jfs+i1kBal9iwa
zp+ngQVyP8OyJmstIltllIj8RvF5uPaYgmdKzlc/oUWrU82EQJuCucsGZAMDj1RxcXPk/n2F7U8r
jvc6bf8w92VlsJKm8BbaK667m8Iim3FkMdatjXWDxDejE6pxFCa+cu+ZFjKaSx34X7A6RP9SIxx9
3AAJFopp5LH5HucrlUjxfgnmM7/r+mJy5NW76+1PV0Kg0apqLQ++sxmMV5HYoTku74QWIPSv7fhu
RY6WbDYRXWKembO3ycp2tsTv0ZOeVWQxWZqH6e/PEh2YtacNRenktrW6wDkfwiJpr77/N2y59t75
q61fGjb+tVKAa4ezVgfARAlluaOS5UilW+B5j3KzuHXx7UK6nwKBZUazNZ1DSMs2buUn3ZZDcJ9O
gnEDmhl75ljjt54nRIaxlxpAce/9h8KmLCM9WjnG8inNVWT8N9/zQEoxilfSPJL+2IWYDr97Pl35
2ZYBfRSlNlPGj2FMYEaMXW9f1ae6g7mez2ksLD6thl16/w+UtKxMgxlDYzSLV/lRFwro1kgmPrZO
rj/y3fY7gBe6Jdt+rO+YcUv/iFLbI8/PRahqalDR+ZVV9dnqU1xQlb6iftdK/rZ8GLWSQ94ib76L
sqmVpPdvOJ1D6l1bW71YksLOVXsKgJv1DnNAn5HhPzoLARVaeQrZ8k99EyfclzKx8WQyDyCt5Ple
aeVigTRPMEEL6AsC4HwVaEV919dt7a5qjyPrnJ9fNoE7tEhNmPbD2/G8Ubu5Y6Fbfrbviu7TwSNF
5xFZSWaTUI/nKfh1c8Zvh/0ywAlxKA2wY9dHbJvrqzKqgNMwyVO20clCjcucNgwEyLOrgfHyWKa1
dGUV9/MSxKjMkjoNwEmZItAgcsOybU59tYIcp8b1ijG16soZ2IYbaFxtWWOx0vQsFjA9DDXU3ePJ
hCP6dnT1HG8bL4mr5a0v46QlB+4Tp37nvIzlXXQb65YjI4WuI+J+3rdHSHiLJa/cyTt0Dti22Vch
xE6HbYcsOhVV2PqU357YkMUzyBX3nvYOD1kJ1CyaOIJCG+E3Fr3eyGXq8mAg1qA5H3vD0P0NSYU8
pH+VKF/QuyqSSYQVVOUBGt34X4ARxjy2b3D4dF7i8CS7pD6MoN4SsHanHxJ0CwS3VWsP5xeU9uN/
kVojAYd5L4FP4N1uNSgNn35bfLy86M76df5aeS5Xfcu/rgQZFK6AmeBU0QTG8d8cxUxzSz7xefux
qX8IieS9Nbq0kA01dTGFeDOKxJb2DwYIJhfauhLLP52dZP4MvhjQKQa4fDTR1vDGCReWBPQPYn/s
BHsx+tCaICsgPfXhC3j494yygP7u0BReW0wbcjEjQqZX+/1kRN5QznMtdBhWZeAbb88Rg/L7+8Rj
jqJAUEJdqq74imvFU7qViCvyrRouqv3j7frx8F6YYaGsxRTVIsfEyTW9WgruHFGlAEWtG3zk/hxb
IsivpYAAnyxcVSUpNR7vdu3Gjy0bDc8J8VVldKPluNErbXBgwcchc/qe6fglujn7VVKEJgk55PtV
yDFzB8ty8uoVe/xLexw2YYvilSSDAcGpyBWWaLxdit8WV4D7JNM4wPIAQ4JhuOzH7pg+MzxBv/TP
bMTPYwVIggJYVqvi4uen6NrOAD+C5eAW/dqQWVlR241GmBt0CjPDG1PYMXu+OWoxcDquStScdSy1
J562HUFd//qEJb++q9kF+5dche5pqd3fUDdmscrxCgPfIKe07rkOijdBfTFrg7feeu61ofx3+3Qt
1xVa2IdsWMR9Y+q1Bk4+AHR6BXPh0aZiL1fSX4u9+gbNKjbAJ6yjN1CUdw2aoFEju+LPw5bFA+y+
8YIv/mqSnvHekanFrZLazDtNbKnE/BCKMg616t23nhWVeqi4Sz3AQLfZ27HdFXka/WcWnXU08+kf
pfLsk2kOZqo+VlVgWEgVytpaE73vFtyKlVbuLJmLFqj6wCHF84OPbWKPFrz8Dc93GxGmHQJnvlaM
MXrv5KmXsCo/KvqPx6NzozHqdiZyBmliCvNYqHONLSJaMIt66yqKNAZzUcPervFUAA9P7/rc0Fxe
AGT/U/+7y+wq0SzKd9P9k3doOErVbqekpehY08YRFwTdd9GjltDTCECZ03TvROIzJZM13nQ97VxG
K+kmKRXsuJjuE7uQnRk6oBUCVmprbmykcJ7NY5jueh78uC86xjlT0sesduGiRjoA9+3RycM/v0MV
Q+y6GlIMrLgZv9881ftEJl/qDNRUast8UR6F+564MO4V8ONrckKxC1YmicOwnKrapL7M/vXKSy6V
S4nCjJdoYEMkC+EY4jTRPZQsoe6Z8j5V3/LolXRjjG9PlZcJf/T2hGUxgWNvCsAcfFptS1nbMh8t
PGquJ5pkKMyZjFuel38VF/kM8cKV6CYiH56Ao2BNpKMMNUgFFhU6yRnLu8otmFgkyl2jSFveqEr7
9T+Xgtea9LYVjUWtCVK9XN9YU6WKOWmovg8VG+ZbSuCaFTeleBlh1yQJvceGY2Ik+saIpdtAVDMT
ehZarUGkBFlpPIQjUOy+osRiHcycFLd5ArkCkge47xFYFevyNgzha95nEwQFr0vvHlr9J1a5r6QX
taY8b9CoZSMGDyAynGQkVDrVKx5IUpqcSqaBmxJGEsKfHPJSFvr2disMqoL6uJKB4xkr0e1mone/
EFqUUc1M4pVFc1DcdDlPQ+0rBgLDpvuByBBhHsdjkmK4Z+JDdd9pz9UhtuO8ym3Uz5J0szrpS0uW
ISWkV8OKkPGa3Wm9b3cmg+cS1FkcUL1I8sVdR9WoCzaYpmv//W5bWhGaCCKaOhaxBStcjBVLsphm
bEqDHF/XjcNbxvgksnQmOgH1L6cq+WkV+svj8AnPyEaAouAwYk3RVVYikxelNLIyl9c0be7IILrz
qZfuRjzCpbRWfPmcIzm5VMgrkh19vaNBGzKWWHAuB21Iz/JoUOrnEBjeqUu5fXxL/PRPhxU1T+0e
Bm9LNxsQ7fmsp9Da3UDw9H2vk43HqDY2I0aNdQq3406v28MdpPrZ5zHr7xZEgU10BmDH+hBOwWty
h0JyF3fn/FSo6qIhHHkiOnpZklKreNDkCR4A5Es0Vn/BSCNIYExPBHafEFiOb4nLy610J0a6rB1j
zfeBI5XoRs8TveqYl/51z0ecpsHmGWveEOu2j01L+3ZYyOowwzsudsg1z1X3L9C/aLktOpK3o+39
jONwQzD4Z5/ryNPoUbOxUk+X7SOD0WI+QaaR0ltKIyEfvnz6vKp2AiQQi4E9z4Sx/Ogw8jm7hnyR
7Kq3Lh+bVDsgU4CZJPxQ5ylqLbHrUW0o5Wy3HMh/MwNU7PCMOgUt8FMg+N5qLjJTglCi2r54LlIY
LfjT30+nV1h5lBZH0rS4bxG+ozUzLOgOhAumLdekMUmoBhKe0jGFjHlqDLgwdRdUdPQOwFZehtvD
k8wz9IXwITUloJqh8CkTq3kOOSnvTIjsxXGNy0Dt18JdJqh48AvBLXnq7GzUwf+0cFeh/mT2H2MX
t+00Hh4jTJvU2TRFwvkBMtNeqqExK0cTwilWjmnV41GCLD+WhRRrW+xafCa5il377UknvFnSC+6g
rxEGU6ReM25O8EoojbnBvkdQJqCMxT5dFK1BjOlVBWfENz5rFeML/+Mczaizu4s3LPOAAMofaBm/
rUO3ggvEa3uH3pnTAwLtY/Qt79Ro++dMkz1uWWzD2N7JgsyOyz/Hg6q75Fi6VVVODjsbs70Zmmdm
WlhQ8r066ZJKvnNhuUigS1lhdfsZ2Nt30yQahJzokZqr6+goBOVKPl/zXFBa5nBlG/h5oyvwittP
TkoNKOnvKZ2P6DmQAL/B34B6kPZc2UaA0e/da6kUddxPqwUoMP1D33/vOygk/dZ60dVD3LRWWgT7
QHs+v185nZjGjpi1XZr4HJScsCk1F2Rizf1f+ADOsnbG30kOCbdGyi5DEo0Clpvnx2cE4nCe9gev
2b58Myt4357pWHRN2hJHpqVs8ulOutShsxeo472vwp5VSDMEad5MXpenE5SN0YJBssJSQHdw4T+/
jHl0HxOuAtrOE5Ny7dkDQ8lw0cBQFQJ2W0/rtYbHFHvi1+ho17BrKvqh0hH1bPk4XKKgFvt9qAMg
nMEzzgaQST90j/lCBB2HSTG5/CGBAprITxKKfZB0qLXTV6AQb5NmNfZ1Z4FzVagWDjxg9UBJLodE
AlDlQh+uyJOJcbbww9efZ9Vz1sqJlcFJSMTMgbOxcahn8YfFToGSiJOtxUA8maozT7G0kav/qgZ1
p7nC6VTygm93wCNd9ePd6hRSLSHsNBITX493AwrPytbyrY+2Hdukovm8GucaSVP+hLTGQ8H5wfCo
ZgLzZtl/nAmvhddcXh5kaKqFkFqnSqvYqmWdjsjEvvWKwr+t0wupZV3UXmcyrTkF0dWRJCF+We8g
96XI27R1WPTX7BnTOeTzM7AtOlrFvZIxWdmZN953jcC1TcLhEgbLoTbF5jqeEanb7h1R2LKkxqfh
tbKLbeqWwC2k5aDDfSy1I4AfqNli0A28TlJO5l/qtYdhxqwFsGkNVTvyVNdPEPCHmZwZZ2x9XKL8
c/1+bId3cRFFaq7aGJwc/h0MyxPbncg0yIxDxMs1oFt5XnOhMVtQcUKwP8dr1tYD2KXaoKZOPxN1
+5XkYtQGG0IwgKueMC4GnciE48hmvoAGtmOcTD9vG4zT8bUcs6vIuLoUdCqfeU/SDVHPc0GokoA0
h8AI6b95it4sFIEBTJKxkM2tyHAxcN4UHI+1sotqhXyEE4WG8+JUQ8vbUKUFJFjZLCOhkeUpqcs1
4WedMd7gdRml9n+894OrUt4/0RGvpd3gVd0g8m1Ny1lPAXE7HmCRUP1Il5drE4MueJzgNH9XCAVQ
naqM6wMOhpcz+MwLQgt9peJRr+hcnD0eVDvuV45BfJ+O1/WeNgV5mijX5WCvHAvXCEbS1T0Mt4he
Nzy3DshHyLJc/EHntSl0NEKKJdw1AgArfssNjr9vywJev7emkw7Yrh6wRO4Tn9uD/lVXhsU2rPYw
celibpMXq+AHXtF/Zz3hk6O10slZar9V3qhz2+8CY8PrcPTq9hcDjlfgC2OMzacOIsx29cAZ+ZHi
fj4ACaYZp3Z2T/1p7DGneZah5ObeUA+dnCcydh/UG2I+U7KzynnzkWp4i03KJHc9Xe/yMxaIX5H9
xni1J25FDBKvzp2P3la4c2RCN5LpIK2qW9fIFWgYM9gYK1GxgTnCMoBnLY+FTKPULjtiz467efas
M1uLjJJcn1PudDDwopmWOnBMJaXHy3FQoT/zPsdkGQsP7efAPeEF/+6LxoW/m+HqBdUBehyTtBWy
zu6R7YOA1PuPCO9fLaOr8YaEdNgL+sWQI4lZGi4ddH1wDqNuyNcJs54J/rhXqoLBkSNSzkSJlf3e
ksjMb1IWAi6PohT5IiZHel8iECKF4GOp/7BU2ivgnwZiUR7giDsDjlUr8gOGgNC7jyfHYJAPjjn7
1dJtFvhi7Jh2UzzLQTbbISexXX+F2SJh0Yj4mnXlm69Fcn5Fj+mHqiZRFU7kGJ4Hd2I4ZM3rXOJ2
gNJ2bqkInamm4JfkUbrNoYiqIwYRKPS+dOqO4KqjuMucyLTeWsXG3C2YdtTUUQkRNHQdt+hPzgG8
qICU23oCKFdUvIewKY0EZxf1cxxgPiinWQcI0+JD86N1LnLsT6GSyBFKNIb0OriLJOLPtwYLwoZ0
v/fCUJZTXt+eqDa1sJBab2U3aPousM3dPtH2Zhpa6eobGXDwLpjfoKDtxNDf9SbtKdl9Sw0UMU2T
wQPSLS9Bg5iPCwhkBTe2fADT5Huz7hVd/HjvCbUsmsL0I4eixG6yqgDNvbvmiyviGQLS8r+CKTpP
a4KI6m+DVYRb3oGR7Eji7hO31AOQjiilcjOBTmNWlSpEeZtI6fCTqARtCIg1ViwGml1bfQysv5XM
C9QFAxK7YSmidGXCi4CppcqCUGkpouSfOQNAde/7nR5ZGrADAoOrUbHEyljb7sA2QjsZ02Tlpscd
yI/UDYeO8tC1FjxwFAnHWqo+zpy3b7MwqH0/N02UfN5LyxJNOW4HrlZrVRVh0FF1K8Y9uGEOdjM6
BKJAEoB10F8miSxW0D5hxy22aUX7Lb+NF+wXS5Tg7M5Ria9E/yDoU48iNd3VqKNbb+SyS00XFTmZ
mOrIADMWLA4zZkFNhWLmFF2voivsrRm9Ibxd5EuBNtK7IWy6vuFEj+biJDMqKBiyxU2w4vDatLxR
Av39i85oS14jGhO1uUbFRbPz2HDol8x+RrbzAuqcoKSHj2gtuKdqN3uS7dO+0BymeXYtBdoUzQ/Z
9rSGLDPfHQ+K+E2XlPIPSoiV2lTwAJPb12uE6+cRcTZJKO7wnDFOVFNuy/6We1GiCws8l3UK5Sgk
Dkuz+gCMbahbV1/yiH45awc/CpIxNX3yQBPt2zjBAbnZvnCEzPGJuiOeE1W6Uf3cRgFZUR30Elb+
+0FCV5lE+PeXZuc4e9BXO+3gzqyi40WiVuoUWhXgJ85vuU5Illw3BcRr4Ne3iqowaHs1E3JGnRP2
ccJM1VjwW3NxQYdEGSHWnZKPzq78y6MBzslcb5tB0rgyAcVEaAEImOAXrMD2D4Zl24F/MQ+T0iS/
+CWIgnQetYHY1ZsCoyiFWlaJT/ocZH/Pz67O15fwBuvZsCwCht+ZBsIxbg6daGAdhgtGpA9Yp7vZ
mt1SS3PfBTwu5obh0C5VRI199/AH/lOA1naj+La5xtvyq7GBZ1XYR1/GkJ6DDtJ2i3H0CRscSN+Z
cUsSObz0N4wVvSa3nKMon7b6s/4fG9Q0WV30gnd+O6VGFEw8uI8M6tl/uIeC5Vz1mdtAdwT0nS5R
d96dLcPu6Dc/aIHu/yVlEcPzn2Rjsph+fTPYK33iyhqX2xFBfCZLbRgHUD2fl/4YygUAfDxLU45M
6Kc9I+M+z1x8SNJFosXRsfytY29AIZu/310pvpC4wIo4/MrrAdU0Ott2nfKD0aIUnOTUxDX+6XlR
eVnWtZKai3HODuCroDpj34aAn3uv4MHY3NmW/ERTYhyuoArYOUs3i1k1x3NCQ+Hywtgo/P/BKvvR
uCBL1hbpz8sd3fVyBP5ak6kxVBOcqnDcFPvLfGsJfIbK7HoiP2SmTKCitcy8PAkL7HXXbUIl20ch
O6cwdCjbR8iPrtvMBg8lSD3QtTY+oPx24jTGmnsKtdjkeH6zs3wt7cikvdvlnwOpAwUOnHWGdlM4
sJABNnemDj3EBMQHGc2N4nbHotR8peOYeViKgNIX+9TrdwnovqUFhADLU849OfoRKg5g9n2yuIUi
PcxB+Y8ohyjGO5qYTQyP1tSzBo75nq916Dnzd0ZCNGUHErHdJWq82QTjxuLKut4x/HHBEk3A5jKX
WsBnMAVfo1IHN9pLw1rd4UBrKc3NNpJA6vVq46w9jJBiVR/DiiQ81crJysvr8ApTE3/dKer8F034
/1lZh6J+legVeBcq9t/GxG5LgOfk0yiIe+CAtWXeIeNnd+CxXfib2+D/gd4JRZp2u9Cqqk58mx0D
/yd6mi4OKAbgcjJbw8VYuqwav5h2+U+lPHSY/sAor2evy11gWj5rZuqpmKQUUk9pt1xsBA2o7SVS
zpf+MehA6yuBOq1MvUFyfLvcVd/SMgQPDOqnE0TST/DMS/pxg031oD1ukhvIZVxCy1sFzwB/rWnu
oabm7iPIkoMoJQ7vL87vh5zN6eOhy5A8AAYqLiKRW5OAnZkweZ32BPlbP8WNYm+KtIGGUpiO3xK3
anL3jarrFUlv55Fcsj3MNO42pJQE54eXiZ9KjxkshwYYmxjGt7sA1WNM2/dX7X6Mq7eLbICYJXcT
aFhYmLnoIqRTh0sQfAjqjGJu7h3jsPb55aGNyjovqu41lXMpMEAIzNGBE6y4bT7FnihgiMyNKHVg
XyGnPGciT7IeVUprn1U0ppDKWZjfBb3xOJX/hwuILpD8cQobiA72VbZjQrowD5BExIzpe9g6psGr
wzLC3oSbzWM45+QCULhrh/gq8dCTPdwlKTQ/hBzveqgP1FisawTzuLwe7It5l/zzVDTVNb7YrNeA
5Xr9cyaJ6oh3oI1Ht9xeRzJ1k2gCUuM7gkOs2FFpZDPenU/Rhk/jQG5yhOV3gKElvGIZjeJZD+qD
2tXoEFfzQjjCV8cKQ7JxDUXNt+GNL93sSyv63q88JzFkS/wHgj+F1i/GiHl9ZgGoUcRH4fhTEjLP
QdXg2n23MBWPcTCQERJ97A9fRZGY2fHXmD0hvjdrmw/dczzPYItB50R005Kt75nWReKEVgU8sYlK
SfcEO+xX2BOenyvULwnuX3hUP7GChFz9/c6W7mW+JzDPeyzW52IvEIXrDkgZneNB95m9dMSPwk1o
wvYVbOA6OcVBBGM8DDkINwi2LpNgjppxjHBScwynalgJHVzc0710fJvtb7bq2BO4UcMLMouvqd52
3TrINRS/yI5pXt1ry/ag7QB8sRP0iEtDSTRC2hSHR5ZrSSQ8n+oXNl5GM+4LuoL678qjmiamYYi5
AnP4fZAkDyo6VmYZdskZO8z8R1zjWFpSYvKbKplkrU7h6Khycg8/ZUddiyUtIhpGGUGwYvRI7gIv
9qZg/5/vEzrmI9kSQmjwGd/fh2pSpkG4AFNioToK+/LpmBjyrQPRT+zfsnCpgyj1m2a/fa7Kmyda
/ht1rPEUCT5bsyI+IDn5XmVlPjUHiCmqZen3iMdQFeQNLWYJSU3yJntTEvmbmIFaPtoxboxee6gQ
LA38o1H2swW2MHwrilGZz3NQBUmlzYG1Pw2XW/sNNABP0+K+ptDOcTlS3AIw/jdJihKh6jeJOims
A/KXqqisw2vQ0cvQqAho28XDNveqWIxhAourkhAL2D2A5xAtNnuCmy15fXQEKY7WUw1xrX5Fz/19
DKxJCqooI1p+p+tbSO/97qtgGJCc1QuF0saCcI+x3Ug7WTm0j8SJrrAgLVxyQgzOMmN/bGxnXDHH
yYmPT0daNSCrrWYYDL0z5NRMCUohbwOL5GWEkvwD9RcaL+r5oGSTvjd6CmUcPvQkpL7odZHbEMBv
8I5uWQDwlNMxg2w/mn6xDH1VT+s2PH094VkhembyNHpKjPSgAKJBKVWDwzS/3iLmOSI06DXq9Cly
UIv07kJFj1RNmnV6YHWAHc+bYMZs4CuGqzGePfMuLse3pAiB0For6An7jNHvUeg/IX7Poy4cYzmk
kax13DwYuk4q1BQC4ZEwyxHVZRce2SUCTno6Ph+bAQQwc5PHErqzt64AgM5TeALQ2DX3BYHArEKv
qJpaIMRuNkGK21PyS17u9j7i+FNJmL/h3Y92fDuNE94N4sN5zAVYb1TNIAdDJrjBvLYq+mj/fUbp
N4bh8GTNBGQ4fRfvdR+v6fgLJxfIPn2Pdzb/TXNAAOmKDLsThFpJyXcmbRuU7+5k9gROL7867bB2
5w08ieTvTNNZgIyQrhiZFqWx5TPhGbSLpj7HhsW6DXRdDLMn9D9M1GCraaV6bi+sJgf/t0o7VoaO
VkUJmUy3q9cdxG+blJpPwlqxtSbMn/gV1opbb+JcIO68XXjvhV4IrRH4tjDsvhOe27mF+BquuAb0
ncNPxOALhpOsRPwfQqOoB+sZ7IthBwi0zt0o/DoJWRLiVwI/uCr/1q4OZbPTETIKCua+Hl5OZliV
HAdXHU5PGO1dKeIecDatdRoQGJJ5WoVpOoGb5d0wP/T+3gbb+Bia6fKizH0ZhqshDiLP/GdQG4x3
gP8bwml8OU4eQ9IWBX/hxKu0WlyhO7MjcvRvdPlwyWJDNHRJszRK5zEZjMsh67lYqzmObc49k3Mw
bCEMxb/U98XrVOKjj/t48GEK16bTis4ZtaK2vAaicmG3OEK7COd/u7g22rjGFaEC68oQ8WWLRkX9
LtAyrmhZfh0f+9ClZ/Dw2fo0iXypEhBIP24OlaJayd4jxvM0X3iQSLZi1UGNG05j0R1dfs85uiU4
Fv0O5PuUHGsN5yzqV3EF/5kSyuyDV1Z7CXCf4q9vsGyqh9CXlUK9RpEKTaId50fZToFhAeYXK0EZ
DDOnMUlYvzywELi/cBLtmnYqp/x5qikyRjqhflWQZfoA8ODJOUVeNmE1BQEnoIo1U7l1D1Z1c3lH
vqVy8BIqCFLrejDEB8uOVAgeLteJTIbd3eRvm4Xg47Z92UJCryulCFwhbJUij9qvpUNeAS+aZdWR
JGFtxwjYMyNUPaquI67FqXZFZoUb4GkPM+DwhegYfA/+c2G4vus7qTySMjDgbLvRBWC+F1/MhDCI
E+eEv0YqZSCpZOP12BMeeZmlg+3sefatHTwgYqJGWqvAgf62mBFreh0b7m7UA1msrqdePdIBxoD0
5gyx1O7wKUisieNEHOHzwBSXRbMs7F9FzXVb1Fi5xdGFjeuz+YkCWa5QAQSaGaVikgXPDOqWVQ6m
kZTU3n+N0LGxYPdRfxeYInwomyQRK7EGHj62iRtcQjxl3nxB+x3zdiIDeXbaHxLSCtV30zV4YvSm
3AVHbCHo483cpwQx0QnHzISqWldZ179f89qtWG1avTVhO49ANQvTg13qFZAlollNwDktcXFtuYXp
IhzKIblAMC4mihCxp2mxV3o8I9weRZMGj0zaReEnIJw50JxWysA2MN2SfOWnMgB4/cDLeZGuZN3q
8OhTrbKlE+FqYstD4PkX6U5WumVVu3oHy+1ikQilAYDWr3xaOwb9pZHYtg/tyVXd0veKqsS01qjS
rY7OheHehE2VVm/ix1C1rd8mGl6MTj/WD4gY+PgH7qN7qgDXjQrP1noOPGTF35nhfFTAGgT9w6Qv
Xx8hgC2suu++zsQmu+v68i9RrEVOa83DN9mRgcS4zsNTYgzg40W1Ya1PHQ7rrG7MBQAIAxL22eqj
T/VR1ZQ6L/AyBuIJmnWE3yzXnppMSMURTecOZ7FidaiBHdHePcYlpoYVc1A4kn1bVitSrOOcW2Sx
IVqPdXZYicuKlleSqVsQHEMaVf8S6PBThWHMdXHz5Cj1AGxYn1e/0/WMKo5jtnz86KirG7Sf8IgR
3yRnYep43kKsyFYp4MTud/gJPgte10vPBYcNRTW0mR0xg2+sjaOiNKtRHVIU95O5viTezfPtWMvc
O0Q3Tmv6/zx3h5RTVaFfwvgagmnH75JSrvfEL/lzWwDzMp/SXPrSYPUNA8LqRenXAZlcMK85+JhV
tPMTSlxE+Qo3vuq1M7v5aZQiDMB1TB8/DpIBXGPvNGeLziR2B7axyW2Jy06sU4wCCJDRey2FB9nF
ZWOS71w8/YrVZYwgFv2RNawW3k7+W0HS/db+7SKE6RZHG152tHChpspjhoT9pZEdm9/CH8UBS6vT
WvekrCRwDqWRllTyetToG8zqPTdiYxJMH17fi8HxNnN0nzUO3y9z9MpKMTJdEyF2kyxmbZANtWeH
Ny74fDPZRlhKSva/DEOh+voXdQycKqPvnLSNmaXvF2QAucZrLN4x6TASoEnAp9mBNL57RUBh2r6m
adWYjpzIp4DaCISz82p/LazINR7U2vgr5yrRJ31ZvRDBugjfcGnQVuwVyHqetXs12PXTm7ee3ovo
AbjF+Zbznt0nGDVaMJuXat/ovjmY37ZO4TIFXC7/q0S6ANT6ySRkowz7y2tpcFxl7tBI2I9EUK60
bGbL3f8pcbelwQcUmx6lVN3CXTkYoWRT+oaNhpfqF8zPFNHgOB/fhHYCNPYU1DNmhbxRiUireQaY
fl3VJ6jkvvP7WV60RMiXKOfCH+OhF3u33qXNR5ZieXstauvtrmNrL8zZQ8H97/saTO33Cuher3T4
RXceCTpdMZ60x5sPXHFLWfjRSbcPgT8wH+j6aIXqZLO6blkSRmn2aPWBccvkBHcPxfhI5nu+jPvQ
1LDx4y7PRMx88E4Sa2ysfKO91SZ7/tghPI3RwgRTAL+m72xyzpmnvPIGX6oSIBaSTY82C0rJ3Wbe
Wd9GGsGROHXB167FghRCPBsWQOupcilo3zvP5oxDV1Gaa2/itiPy8Bhq0WqwBX4smYbgrB5Vhwxz
FppidcCCt/jtzw1QLvCvYzZRGglGKc0QpWlyBJJKGHMhNqnyBw+kShOM33kkSLk5Oipvl5j8c52i
gT7RSiptL1DytrxlwyBNLyVeU1aZOTD3QWXCJj/Ws0H1BLfDOio8eA46deBnHhkm6ew2XLcb4iTa
2/+JD7CAgNGBDiH4KlbiCQ6RryVd0Mkk44K8mRo38eQI8qeOMm7jpOT+xuTyP2Hwhot8NuyNY0ST
CftqvepkiOaj/y863VDdcaX6wjwAlpJEwi8HETkrbKixIhyVFYSLI4sw+FqZvAWXGfax7NeGNrIo
NaOn/rJ4U0bXGl3cZvyLUuadi/DmaLPaRYGL82PGDNM3Ggsfnd6yt6QLmPotNju+uIJsgvoVJeu3
psDl+XyyRgzAMAWHyRL97dseu+atOV6MFG70du+bPwVmMrStyOgXsgTKYukmfDBpdjVp4HfdIXRo
r7PicT4V3gCA19Q3tc6cfcJN7u03jgFMZPY6zWN56Wt8Dig87N0XrR7N7I2GYrTeD5FasALF4K+i
A74cnHJC/Gcjb5wcGz+0X1YmBnMTotUxlvoq1s2PL1bmRyvV3qNDOSK0TznnDE+SdfsPRjqi1LzM
jbOZe5o7VMFAFtDM8DilhQ2lFBM5Pl8c5+tge+lBkJv6Ya0i50k1WGUU+S+on5OMz2W7YRbHbMl6
j4Y49/+OprE6iwo+2efAeM3qFgSONIaP+4QOS5nCukdpnTFggi0m7P18pfcgiDf05nefQK79OmIu
bYhCzJxB9jJZNau/gUYSQLHmyybyP6P4U0c7NQTT1wu49P8zflty1fDikVw5+Cnu9M3whaL0eJvi
zujPkr3vdfYpqpGCfUmIPsOsBdbeDSJDdcC3KxcZs4FleW2Q/joW72sd+wVAgGOiUeyW/uRDYxZY
GcsfcxxlVs94tv49krW6w5Hv175N/eUwlpjy2fYn9yVC1gDcH4MUSt/ZML7djqAB/Xj0aH5OPLsy
0/1/uiYKjZA4CPDl/O0hJs0sTUq8rOghp+95l2koaquUh60v4bIxBUREJ/4ciOScWosPdqdvPJCh
4enzm8l3zp+8UTWXW7YPEsYCCuRQcOKMvdknUbbTZt7cjHWUMcgyGp6LnNgG6ZxmO4tgtMeOHi3i
o59YMWlQVX6vrypuSxe/L26wEyM6PkBlM29qzfC29jC6CumTBEgWaxGslMOdej3Iz8JYMDVSPCFl
/Bs3dCn+zTUEsPGYI1qh2NNqtjnY0in9TWKXPtc8u1B8dPNa/zkLqhFcwlCj1yca9hXDZcQxaMaO
o79Q4n/Dk8cb44r2BB9AJW5y/RwQ+vrx3MpnKWXAwvepB33z5RBS2LJ/U1XQgcjtbKJ2CS8dvUO/
mt4yQ9D1wfwtJ5WUPj7YF9QaxjUA3HgY+UmWRYChxQDQVLJDxbgENmRTD+4VFaw6EgGX7PNpA5hX
pUL9lt+ITy2mxvK0TGX3Wr+jiUS40tVa7KjofhlLEgdkrTWoE3P8U/NM+dpVAduOX98DcpGykpd8
8UEu/8X9EHd9cLRaN1jGZpfRxTINiuvcL0plhOxg420XG2rHli7Z+x+MPpJLmulv2sY14PkNs8G0
1DsDYcH8Tp0QazqFebgKmDk4/ZJ8Aok6BJzNqei0840S2b86PGQvkknBIMtVwqnQ8dVjE1TlqqaF
3p7TkYqSZNMwECedALBS1sZ0//8Qz107sYvWSZZ/PYOFEDNMPipWdrpEiyqeMe/6dz7M1Wms6hQ1
IRaB9t3XNkuv84WHi1BpYJzySUntP4shahJ3Yd0nV1YnqimcL+YINpBol0UIF5rBeAC9+zziJD4Q
Fy/fosDtOBOjQvu1enry7VqEnGcqypXXxBBcCPYpp36LdIjzm5xPSdRDCzRI1xnpaftxbI5UbmcX
VyyPJ1lFzjCDZQYRqPcVH9ZtwTHdxQ1PXt5t4WDQm1lcWT/OhEiQm53hQ1HlUf4ESmm5eQirVwvZ
fMe/disTA9L7m0yOQpFUcgHXZVpVjpTEuO7hOnNSsiqAfVa7Kt4oURx3cUx6E0nkIdbhL94UBG0N
YKgbjn4YBJxIoR5Hw+0PdULXBLIPJd6j7BcJ1p2WpNuyBqefBFkdQ7+FNHF33dMyV61RA3ndTFgb
0uvISAGtW5stXmEOUi+WYdlvMWDrZOAk+8mmFutHe3U8/XpmQgFj85GgF3BqJcy+/RWKug3Besmw
k0TZ+bPdh3nWpCxZ3WvNvxRf0yKuSTQS4MfRE0LA7SVOoOkctODMyMnlr9rm6HqLhl6eUI1JhOCk
+YXOI4Fzcpzxn6Y2qCjH6JRGhX/bziNiKYe6NPtzqX4bQL3ZJm7cPmefACVC6qedcIQZiXVBQ5ix
a+me4zDLhurAEZz2L2WbgKb4B9LdogcUj0SUBBj1+rd2Hrm0Dt/8huNXDgWR1QKr3Jj0Dvwuxw/k
pUaJGEPIqeHt1bQXBCRQbIY39/84ESBm/y7zz4ytADoxxbNJoC7M+C6lVJEIQCgwUNbztu+LY/VJ
EbolBz4Z9RtoZ6Ylje0pYlDiYessae5oEg3ocT1Rjzkp2jsgEJ27X9dSIDamSPEmtji45WqMGDPj
EB7jk8NgWhCPjZCqwjK3kkKNKEMKbtJ1sRhQWUIZGdeBFWy0tXpfu9ZOZmPSouKY0f6gCjvT8C+E
q6nPnvOjQMLl4TMLXOenblXfhywrkqr3PRcJOAeWGbqtN40j4+XAveTkPclMPAldpIy4QrV0oA04
ArwNGFTBw+TcDUm1iM/YwqPaDAl8PzU7EcA3M4E3U9FGF+ZRqVULnabtf+5D3rdkkpflS6pndjQL
kPcf7Y2F1ssn2ZHqUYa34x1haN1X4/XvTDrQvakGYysG3mNxYil0JnrmFGb9V/hvr0ddY3CWKL4z
a1rXb7J+X8IDCB3OB0v6VHxwkz/Sn/0uFDS7aWHzaubuBQH5x0IGva+p0ahZmWzyeLgG0ZoT0zH3
dJ6A7Hgx50+g/zEXGv2PhBcs46vAT9fxRjTOyQrd/WjuCiBmhYgN9JGylkqOdpmVLIQVEIrCS5Yz
9AI1InnIluspgQ/TFV/T1KjJzWHqHF/rvmibKzrq0wGhxlgokJPQYwiKo63QBWLTMUWDWKLgkIf9
KIG6UmGQfzx9BsC9EbTPwsrLWECKZfcD0tZMutHtcBFPHSW5NwbEHGH8iJPfdhnA5hlAoCEObSj5
yaQGvgWuof6aXn2vkBIywhHIX8pe9kK4pHxo/UPO6xptwPBlBr0Prfm34EjNF7iY6gfGMC/Wa0Ip
BjmJbq8fIk4hW76F29uAk8066A7eAa7IEBNFcMIL/zZUQzBwvyS0HMrVWE2k0zS0ZwzikK8oX1r0
mzP6+5/lExQDQqUPqO3C9VdtGi5BPM8/Q5e0iGw7uCjXJ5aRP3z85P/rb3sQu9gcpS+a0FkJR4I0
2Z7ohEMZkUlr2i2ekdaT4bdhz1Snc3UkiI9d8AB/ItooYhGgVUny71JCj0MiATIf1VTKYpS6zbNN
kCrgfix1VYh9VHrJBPQxeBxbivtwkwUnaZia8yE9lWM+nUvscyDbhhT/FeGdYI+/0z1KabmWA6C6
qh8otXM/y8pNm1q74tZ2wMVJEEIJ+mSAiXrn0JJ3D+JIjUow1xu4JqgSrDNJ21TbKcpkITDwo00/
+6o+C35JyvSNkVvziLuB21H+J2y9/SnCJ5tF9iYWCBjoCFAbDb+6tn4LCi+seSf+a6/ZFE4HjMcG
KjsPVSw0qLSGZiHchfbxtzoxt0RalWReIXc5mPWtn7wPBEwx8FumR106WCGjWO2PyQdFUPi7uJic
VeKv1cbvZMY8tUhnoZZD8teS1NhqdDElPVkzVG+n3jX4X33etZFSTz6Fl1tgmpicxpUvqegKi+Ww
/qNl7qYcKKPvlnm1tA8byZYWh3f2tvGRQBXgzEs14DQ+zweofo1rdKmiXPlS3a9cZZQCaYP4oGIk
w4ZUVBZzXvGfZRC1a2elCknjvRPVdaVouhWmhvnSkNF18tsJLUNVIR5OaoUaEBDBehJrsmZfF9gF
ikDhKkqpWnqPkRlUyK3x3Y0ZX5PPG/Jv48FA3OmFkBx+AtLWynl6cCK7oprnxDy6yY4glgx5H0Px
BbXj+fpVmru0Du/3UNkaFQPRp70jWt6dufWtfQkyIslzWlnQKv3gyg44fkx08V6kTH0vjOu46AjV
Gy3QUXbDXtjUrpUt2IU30pBSnHouwCgWTDT6hbOfQxwvlk850MUz/WeVCm6gwVpFvTk2gMMQSIAl
Z928Q158hbrLFsc3EwsYybOxGl21qbF+JOp8Bs9cmpmVJ4rpbaIHOkbe+lNNBbSlHLaDaCOBnbuQ
cYZnf9CeelE4gUmbmjp/jci2kisPuE0GyrcSANm3QXy8iPNXN6IwUg3zs8GlTJuT63YEuTsfwnHG
iL1dqdO+gzWebObGxA27YoUKKVEyyBOwXFgKmpwP1sGiVOjAAlwboi6IxTlCgWFC7UHt9QebKFw4
KiOLjOGpP2EeFNikWRm60bOjRX/9NgjmikCb0Zq6+HFu/hX3Cz6fWvKHbpyyMeKBrIrk5Ldarpgl
WZAeEgZQxs/dwCiPlisHzjZpgAOPASIOYNLSn9545OYy9hoVx2ZSX4DkovE4ylQlKruWQlYz0ooO
KmGXMRI9x1SeMl+QQQFXnYLrLIvc4ys6NMuFimZcD8jqJ3z8/gj4jFeeCQHTTNzAj+zb1Q+hFxCE
uv1jGw2QEqg9ogEWiBOgjjUwqioJF/VVR7qILGUNS7YK2GGkeVD1ktT3LNP1Zy1xzT+SGfHmms78
xaogYXxAUV1QV+CrFGlT2hekl6ZYWvF+FZNf9WQF1wSqLtElFFJN1P4z6gv2XTYNXgEQCAoh7NgN
LvYTNPywlwnmp1TkodsfE+T/SgbxSqMyJRiym9t+cZYqbDfBpRpuK4tR38EM7HiWZ4kWfBK2EtUm
dhRiWjXvg2mRBEJD65w1hQapicZ4w2fwci6+e2ZagY5yVcz/d6XguY6fRMCHzNq5bXy7Imb8uuuO
twjoTzO8z4B5+1n6SqY2E+NpXjQTJyyeMpo8WyD44W7ICKnjkOPDbu+UsQyVLwXKIRnKIdAtiDI4
tb1xM9df7QKQAxjWg2jqz/trUquMwjAKUX0uRk3peFoOqv9s9B516kWCIY4a3bpkh3y+mgi7ocpl
syi5qXGMb37xrDQX/L6LecCsISgjCUTaj98oJX42r5DYFKQ+Ni0x39JgNp7YyzJsbkaIvA7n23cK
uiI0o7+zwxk4WanKHTMqHKbCVrvpPVOGEREyWpcHFY5bpIHU2aBySgaaLMbIu6U9r8zCJYnot9f4
TxeiiJYiw7mPT2gMeVDnS3Q6rPE6JXvhYV2383bsGeUChJH/gliuMCQAA3TJXlZC5NO9XCmRUEFz
IGfYErFUd2rPxzu/jTjZ1oh02K7BbDeTmfNH+twAmzBE+6RGXD4pNlNE36W81+GceD8RgWNiDj7S
uz3UpX4Z+HYQI6k6yvb+LSB0MUELeaFMu3/RrX26ZlYVGnK3jPFY3EEDI8OnEWtG4bFGST6d7hDR
8Do5flX3m5XTLYYRST3emCczfKMIkuopzTINm5J9vEqZkvCdfH6VPdDbZQsfRaFVz+quOdCIMsM2
gZfT8lVIOW3wTfQ3rbRlCizqdKuAFlmC5d/utM9NPdR6LlzwTKhA2r3+L9J6e5tvxuKTMW0w/AWo
W5KbaOP/UNkkSiRD1ZkoUKJJp36b+4WpmCKqXTpp24yBD0WvKqtfLikTx5nYCW0YJPcAbbj6FwpU
bJpX6p0/6xKpTNfUnZkazD2ptOioSIFD2XP2OP/hoKZdMNx+HUI2lcVG7M6lVWuvWbwl1RWZ1k/l
Zyg0rG84mOZncISvkI2gmg1/jTy9XP/HKJielzgxo2Ar3n2lnkmSYgnsbMD3VLOrtWTaqoyyatkt
8vroEJ3PzLKH2C+VriLte2rIeIqLPFwuu5scyata8eUFktpQizEXuBVOasIpofG4kepkC63JU2jU
X4MwymRpGBh1Mvi61gpRS5vZo5tzqArD5pooCusCioifVdHYi2vyj+RB1r6BlF32htZh1RmR9dKu
UODUFfY1quP+8EkmPb3BAmU7hxOlnt96WQuzCiKH6nIGwmrg35Y/A1CMbug16MfuzLXLZ2o75vVR
gKOk8TvDMF5XvDX8iuFOfXY7AJSDsuWofNyf8JZE2tSqwI4Ba44o1kkij3S/XP9PELo929OQY2e5
uzE2zipwQQp80GCS26YT8CX2dEQ0jaKoKG8ojEqxoLH4POeNhPqbm6oX9x3W63dbWC1KnfRJPy+q
lrtbamlK6p+98InVsAjOwWYzarnZChjbP+n40oM2Z5xUkbgrOMLmPwA6kjjq/o0Ma2tcF0T4itv+
TovKwrKqhtnBONLz7hoOwSKYYU+rx+G8P1W67fbfg/Pv4XesDr8Sh3hBSpfHCcSexP3LHkpuHzF2
wfeYQLWARRErcU4+pHxPP8VesbQl2WXNToLswsqtyDC3tuuPxg2FdNd24Bx8QC7fUmXlIV2WNeu8
cIdIKu5m/0fNyQyNvz8XNVjrkGhUTrSJ6mqDG0KlqzmeJEO4MgV+m/kAIFlHCUD3vEPnmaIVzUvb
w9CefHCzpKej43f/Oo4lWoYfTfHImxGwRfyL5oXEKXo0DFZSCnJy2i/6/tdVLDE0B4FTa10umrfY
7Aut6XxHmiPytWKuxoLBFQgJOOzGkA9uEpkBoKLIfhIZegKLpBfwKp7dHYdZzs+/3wiVS5RfCdgy
Sc8h0Tl6T13Hrys4jN4hqSxomfZRU2xgJKH+nGOB1N5xKDMdAMBrgTteAEYrKclbex4JjVYC571g
0hMvrqMxVKYIzdXMHt8fMSXRA+vFgnsFoWMinZRQGC08EdpAGPFYgu/15HS5KsXR/tQys0aTnP6f
nnVPK1JcWms4Tm0KS7I/eL5L0eF99ZGebze9kLAxYleGOkA7NM4MgXUaIYOSKYjm7VcN0qE81Z8B
Mknu0jLD+ZCJYj7IitnyVP9E222qOQW00DGnLyxQ26cyPVaglwPo9Wh0gnldTBuRlC28G05Rrxdz
4GV10YCdCaHXTqZhg9xluOWv3lOazthkwkDtnERFho/TqlDTkFLWnAlMZDlfQp5BP7rCUBM9Uhsl
piEzkBt12OcuyeEcOITE5JPaixh3NrhZrIxy/V0XNTRM/ZMR5hlioEf13Ocvy3y5StNEaTP8ux6b
pEM1Viyc02BlwKJ1KYdmxoBSWgUDRRFcEY7a3sypQ6cnnfYNKnXpNZroO6OOcC+9nCq26Y9UOJZ3
79JIPly0YUoDC/AgNYQcpuYmGYEPuoxqtKQD1FOo2u4C7zpUUISNnwC9MKJ75iBwxaJ2WqiD3WAk
78WT1o+nHpDOVYnjioZfQF4fSw2/PgbI9XvQU8y11VCQ6ih7UBpzm43A4h5HOCq2eUWGEvzUDyx+
ZALmVlGD4J5sMv363uFED+8OtkDWwvMNkpwYRyNeHYEu0CvN6uRYfWs6oBuQ06Ugz3Pft2nDth2x
TffhAsGuXi1z4JfPz0w+vlefh0WXC56G1UGEP2krjRDl5PghvjaWovJoGZPe7rfrHzg8X3AezilQ
WNM6ZcO58zP77pg1+D8krv1B71uxbOsh/xjYICxojz8qRXOQAFK5iJx3v97wfezpR8l5cG4h+Dew
ckR9EMvbceNlYdlN2r6+ZhjEh6kRh3MP+V8HYOyt4EL5HQ2ZxJIEm9VxzW5EPCOX6EllWpvfZtOM
4ZWPK82qqDWzA+NU2TLW1uMQ5dxHo/u16TRfhHi9nholyMe50KuM98SDFIH0OC9pwRmIOy9BwGBg
Rk12j/rUTtmiL2KhXzp/567zMEbrMXeVrW5admFKnA1/GJisYC5A83sY4a+D+oVkj118YPWw5arJ
+2omlxQPLawpzVYzqLa7RVp+8F4P8TUG3oYipr970aqu2cEXU7B4QecPmcaBHSm3k5qWWjMinTnk
lkJzKfy0tAsrTw7b+e7ILaDGxStiMWSZ6YmRdpdBWSvmqy3f1WdtNHWrSNemTaCVDsH1geQ5lyk6
dG7pwt5PCTtvAcFOZPmnZDd1LllsOLU6Xn6teL2a/e3L85EK5oql+ic+D/Mr531ZsOExHbSxFubZ
hwTt0JRVXIddmzn4ypZ10rV6I0NlEfzChGMykvqh1JCIyoc2ywcwJKtCmB4fjYmiUt+KFxrOhA5R
P4DJun0FpJfwr32fUdixyELK7cNCgKSwuS7dKvHkru2F6QQKjq5/JZrb6Kttm4+LaxwFvqVr15Sb
R1POw07dYq7dyOm6bIFyYe/aRWg3vxJXEfmGMvM2Jgr0Go68TKnPuOXcePJ45YNgUaqnnilCzVju
0IPAw/HQpL7rskmIIOUEKou/VUjC+s3BOwECSDF0i2a5wv/P+btkeaxhKXASGmN6TVYHernqBzUB
2TCkqqiASUs0zaRe844sZ4K6eCyGfKgy2ACGmUoHKYS3E9+s3tiWeGU0c967a5hPdGaoc64VcPdr
2WSho86kEXui2762eCtW1+nBYolSIyDuB5qbouFOyA5ejueD4UW0JBkOJKlQ8cmGHXrM4dIbcNC6
IvFxkepJD5A0c2dLLAx9ttGk462YihWCllLO5HMBRqh85U3QnfmGm9NEnKLxwcouh/VGemkELkMw
HJZu/tnxnfE8OJBSpoM3O5sAiK/yMov87EVRixFoYTQWL6c1Uhehc1Y49SfMonG6/v49h9PiBEYi
T2SRhVOW3zzmRYNNNo8S4b8n0MlB6mHRJegEHTxHKFjB0Cpcmg/rFF+QS234vXKemGVSmIvZPnK/
L5f47TK0omb356FZXZ8baRf1tskDfBS/o412s8rjTZ9TVAQy+3XE753a98/aK/qrAVx0d0qKV085
lC99in9AFWyjWfFG1acIzPaRrubxslBWy1ZpotQh9dhKmjY8MnGSgQm1r0yp6naUy6+OOz6Y2yg/
62bzr3f0IOjHSSn07RhCfWl+Kr0R7dXU06d31ChDStDagmw7CZwIRr9mODeXOa1+qw0bVVVqrih0
C2Ma1a6GHrKeB7rNq7pJZ0Tce6krBz+v0CfzwIqw6spJySQHBUoXWUVRHzibYXMMjsVFD8l1ab50
m5SrhG+TYefKrF6dzUWZAISqOZGD17wAvGIt07qj0Mvh5yN2JB4Me4PP7leG3CF+cTLNdDbChpP4
qM0SGDRsunjEMP4P9TxXf4+pNiC1twH06BHgz44KnnK6GtYKUFOP1WcTTJLLo8YFNBExyVh8YFFQ
n42MwXTk/SI+jrGhCXzAtC4xRCDfXM6Txl987DnDrlDLtn23DqVsAL7se13nA0D1PQUC8PJ4Hi82
TBdba0yRfvLcc5mAHGZRbpmHccxkpigTdZnI1IiDdSWNkmu1zoAPEWBxjIlSyhD+2Bjl0Rbm6ykT
bApxKcEW1+tfD9+nnM9JM/0KGyxIPo2eux9BUl9OjvwYoXTjURHS2GBi89H95iAEOS5LJIKyKVCc
LYG3KwwdA2xaEv4V+bCCu7JEL3LQMg7ydfoSphsEzJ9TfrDvmi9mdVp4Tg0arVcse9L/W7/Pwpav
csDL28PKaFmseCKQhfdhTjSAgrDVRY30uLR9C3KaVU8C5/Gx80XLwTNxpjg4FFRMuG89PV9zoMv6
i68YYY6bHODsaHZ3mih+cSx1AK7suj7Q5Wu9i/28mbjJ+fmkOsc4hGW1sCr4OfL6H4OXrpoSlKTX
yG8Nbqn17rkeS3HbIl3HJUAo0y+oCnLwmrjX5Kb9UwrvsTOVn6j9Oe7ss1x1YlXmG/sVn/vHKyOJ
NpKg2nUA2O+bOFM4/HOIKCZp6WKJvBSNfxDjNW1atXzBTjhdxkql/bu4QGxkZZy8S/b2mIyGwXpV
4zC6k9hG5zPo2MLmUOcEP5hFMMnZzRH+Gp7nhOgiWfs+tETBc3UsxBBj8gaK5laMAc5DXG5wyzIb
GVxHkDbLCtOmbkodhtmHJuPBWqmHtXWZLAgiPeesjnPOZzVdd4t8BzndctJC6DiOIppfWKdKDn69
UlWVR5/3N9ZtMcLbKj2NjirAvPMVu32mjM0jj77xiGlZtst0ATEz+tg+EW7a0xUpjjJIyomM73RW
vcCfNrYnPgYOttxUhVT2u3Thsvlm4VNiMogmbo7QiEW76qLz/qiDGAUMnbXsmSw8hQ40dsVBzKDX
Gwb4QqU2mvW4h/iRhLdEGPr70KDi5LWYJwCYjK3rRnlAOUqOjjlbd8PVhmxn/TIJe2sUJ43Irq8C
YyCAFEocps8KvWyughtfTSqQaX7W2SbGHu6u59DlG9YcNnmveBQTGSeed5no5gCWxNxLElA48GHA
85+gmg01m7dBpLK4EmnfaL56SAKTpgBL3dntA2xtV5+WaGukfaimoLC1VnMmdKo3WjipO5KTW/yz
sglaoOBQ4kfktMqOnaqg8G0fp7hMxOzVP/Gf8nnUR/gAgLnjNJ90MYWdUiGf8Z8mXLBborsEjrCN
cmNpTeoxraPZBvFLmwSAMCe9nZEgKq2Kn0gJ/oYVia1i9OQAclWFvD4CsRP1crH6ZYKBEzazihSA
uua16Jm8JDzl2rKqTaruXDBUooOrsA7sAnDiRZeG0gV0A00M2CSEbLKPPMTLlAS3W7DVlyYoyDt+
H4vw3liMgIjRjrc8BWp5pyLFjH0FvWLGldM/cWChFSY+2mmdZdbk9H0bpl34MtokS33ultAWJPAv
n99OEd+mbWkbQbs/XHp3jWtqZFyfvVpIyIUUtsvMTyrOi40Uew7myA4/SmQ2DOKehDk29bcz4DFH
0wF3Y2KZAiu7URQsewUOzis3xf/6TPP+fcoII/iognUb50WGmEDCK5OtzXywB30VUh5BUx1b8Hwm
W/VpXN/cx7PIZod7f7KlV6L80urS4YcyAdwZgofgBzYubfjuNPvfg5GPikzOTKT3YVBAMqKBYULc
TDItUsASZ7ZkZwLSJHmn63ssNGiDA5rHin+09MTBDauDN2KYiIJLIWpS6nWXj0iaTkn1PTkNaLGk
I3HiMsAv2wyIyI1IcmUvbnWd/v4mRK6rQ5sKC3gOr0rgXgUt6ePhODIoXyBy14HXgfMwRTSUbpN+
3sAugkAWFJ+qCE5jyxc24dys3WtCAEBBlcK/2LknAuWk9XYbqcdQq0odUhRU5K8imDPCsTJ0toxO
ufq6J6y7Dcdy5thnW/rGxkvjTU6jx1W90nHCMFulgABNA90M8ln+nud+GV+NdGCTHKEyxtWKbzrJ
iLYXcOpvlqbC15SsBIZc+ajOA3AzIPk0Eb2HHY+CWHOmoYgZqnvB/DAUfJY5/A8zvuHYi5wK99pN
+vwabDYuS2dfDtAl/XO/SCO+hfdeOjfxFZEM5NVlGfqYwng5SHasSVeO347XQc6/ux81Nw5fWmog
4PA09ilF2ZNMn3y0vO2bZn0igxZrhFJczUeHKrLk9im507wFV09+62ub8xrb4P6o+js5gKNfIMyX
6ZwAboytD0llCo/I4DEaK41NPBvxJSDKUc+Vtn0bqZf/2d5bxNREZ00LTdDhjtFtLATcHFY97ZvT
546WYvj6HZeFM7AytLIcvuPsKpQkGMaqoqRL/BXNQ8Mig1pvLa0658ur7hKzcfGWpTuFFD9p7zjw
qg33A+vtvvQ3Z3DvdX/qarth+YazjlGTRwcntMVt/hYV44HoEU8EAy87Z5sjAMpbyslFnv7R+cDR
WDmD2/DGKL+ilhn7pMRq4zPi0PhSdfVbH1B306PoJ2bEi1/H/ggGCDstHJS9DwkDDFmJZLQ4S72q
j4Ku4UtjToH0+sIE6BSgqJO55T05rsLqju8j32VpfVohUoMwdToJajbU66rlFfljOfG8Ma+tBRtL
Lg9qRsANZWWmzQYnfrm0C36PESsPsYR55x6tK92eZ/3Ywo2WKXzjmB3EwT3vhfaroKL72JUOhrMK
65pU94273Fb36S28Zcgb6PyYWcgGA/BMXktHTGfUyZanvI9cfjx2K7N8WyfZ+UQ10IozvDaR0FEI
UmKSSN4ZAtXIrYiMxML/FY/Auwmvt7bTZ20iwn02Y0rGWriF4K7l22uVw9zSRnq+HRb+6sRsejzo
gP+PZBj9JV6yofvE8sm6e0TzAmQe6H0nY0H29TJKZg8kNA7ww4/0j0yEwqpReW6ekh3NoxVUx92M
QER0gOAb1kCZhlrP3SkgqvJlxoyD0TNTdci43BFha4VsKtahtYmATU693IUFbEDU0TFY5sScfvXo
AslagJiMHJ21PXtyUTqJNk9xT74wsAVItXVufhYkGbLSNZ/f2pOySsMT6czPzD3i7Y52lztEJ8b4
99RPVbHMAikCeaGeWCcN/EI+W+lGNhuLgWN0g9kCrLITM8mCZR4ImJNcZIL2Pf6yXwjXp7Im3qqn
28piPJ1sGnniO4Wank+peNn6LVkJgzVTSGqSsGO6WPWUqHuHYUNZWggvMZ9F/vhGWeSnZ2qXOdXz
tWZGauf/EwbOaulh1A7JNNUz35AyJ+RQyuhNnr1EjhF0uKgPU+nOcugjNVN4IEhCzvEajLvoMIbn
IsM1pYz4aCXhGuQ/IqwF/mGEaia6BE/oJ2QuZHe6Gnsn2haeoijSS9om4oV+xA4AbqWHQV7iNiTH
puax+j5NoafOYMD6yjWR+PDMxT6vohevTWrgVa7lM1l1nS4gMWAarMXpto2zX07OLKTNWptdegSu
RvPH6RryhEZpjUJ8YyEcmXIPHr/575176/cZng8VWiKO2PP1C70Nka5kmE1fjxBUvopxC3AsSChl
KvCYPHqMc2nK/z8Ycbk1YD2p3keF9kGAoVyQtt6KYEZVHZcxfr1s6ScS4na73SAom8XU0nWh0LyP
aPGP3gO0T7v2y38cg4odWJTVQtkwkO5E7kZLlHi6mUSzCYElEbtTiM8SscSw1nLlVUPQ1n0Tp33/
euKhd0RYGqhiYKnlpWo0BMWiRepw1r+AKEqPLOaqaK+tulhROH2cjY70RDMv4oF9FT0bJoBEJBiu
usMlfiTKVt/948T+qC4DoFf3B7I+P8suHfUElZY1EOTy3Wa3bEtOMKWSW8J8rc9H0msakWeYtKph
RGG794igtH/kmSF8wF8iPLK1cGdskMzhfs5FvvAq3F4iKqh4nZyIIe2Vm08UQhRJxoX9L7Lo1ANg
T3Ij86eHpp0fvfFWaD1J1RXYgubOIXckBfdwESPdIUD8WsDiG5Ii82aD4XQDF44UzQUAkHFFjgJT
Oxu91rmtPiZx5iEyJsbQuFWDrKv99W3nyq+/S4aHkCsbX/XH7YGUhq7VhBDnhP4DvSWt9eSHVsJr
6GYDYrOCDFshG8pGWvtU271FbOQ+yEMLv4jBO6EY3DANVEWnX+pfrR+jbgul59WJCAAG28+hbg+E
Cy9UlFAN3Zo9AoyWAHvqqlNdXPaUm9hlvFm0JmUTNcWANAo4HHB69qyD74jXhp9DWqanA4wbyCNh
zoMyOhtIbkO1ZG6p2MRWaa98z3cS1iSjnOUtUq7aJ53b9P8kvdMOE+fUeSOdRFQLqErH1xluUrLV
DllDNlU5qrBUsfTPV+t7XLbtdBmW+gQEtD2zD2jnm2mA/OsvCUELvVULxtHsMGPPbKAkW3OWPcMo
3UiotjoWYB4roMbFTq0IPThIOIBAIHQ5StaL6tK0ijSrIFhx8IP1Gl4OcS/oQZ+QrqScOo3qP3SO
MCg3O0jNH4wpMYpDmB/nkLaWKvIVMr8g77j6KFHg4N22STUBeon5CUjX5dMbnAb8r2fF7CS4iECj
9CU7HIh1udW/bYoybQBo0Szoz05w6tAwHzgvgRYylsjKbVZcKY+3kyJG+bJXo3CdRTknRngDhvkM
eMetcdIWqp8UFTrvSkYtWXd1LBSP8g1W2Dd+aSmVXFDYP4IqWpp+6ugHJFczcIDBhVAd4KeoCx21
sIHP6XtUcde4b4VNAhrAVUR0Kf+TqCj+jkUUsPjYGtSro/8YVywxgTziDNOltNHk619FtiXWwynB
tGfbFVfWhnPDUVLcAjv9fmWPJ1JW4gUcOA2Xo2lkycRBYpbMCFFL3tXX7Dk2GLi5+MteQSu1lk3Y
uNnutAewfOQWKyfE3VO9ZrF013rswnSmoKvb+dR0JSuafrqmJJHC9a8fJSBEwklQbo7FAa/LX2Wx
fy0Fnn6His7FBRskq+vmIdvdcd94dGCPyRWOfX3g5nC6z0cZYfLty6AMBrfPJJA+wbJWDWhaX5Fo
5ICmec/Xn0cpoaEC6+Ue9MIm8mqY+W+pHD60culuz77OXk3mE5Q90/mFbX2DH6F/AYQeirGS8jmF
AL/wsYIX68DkrWQRaO2EYtEj0bdaAavxJC2hfPPDvtlQJJwMNiT/7CweOSZenMsiAsNCSoRjR0vy
JbCos2e2MdGtrlc21lf+l8joe7kDuAdS9znoco9MFqqCI/2YeQSDj9fHTVGWHANecK1HhioZeG7n
anQqKUTpZ633sQ8Jfigb+Bp9z1rwQBj6AgxIwgIUiROdRPRTBmsmN/9+oTG1AEq+tRI8IJQ+Axxl
pua86HUGlAnFXL3Ep3Ew1yQalZ11ObdqvjMy0dK/NdH8PW+BLAo0sz4zKif8JzPxHAb/PlMFoMPG
2R+I+Xy1SAa8m8+EWDqu8/R4+B6Q5LGxVb2lBe0wa/Hi0ss4P1tsCXZ/wxvOBD2W+LWi8sR5lOQH
vB44bEcXybSJ3+4AOoQJIFQ+UfJcCsOwtxBus1u8FhJ/2NLS/AJu3R7ZGSTxiymzcHan89rgSaAj
TfbzolpYVXImOFkkia/D12EAeCSVX+3U412OHuvSphXhwGrwirFG9AvZFVILgI/eBYMAkrRYMRL0
EMMfV7s62rbsnGzOEZPel2fsqXmcWRBMfqqEHAYCWSyFlLz3hYkclGX/pvAzHxqj+5/I1+160O8y
cdv2hpvTg3vrmJ41J1AxigdN22GCiyMkye0GNo8o3WIhXBXLl7LdMmhs28kkBK8MVHp7h95CidO8
deGcrN8UiK6G1pB/+NumdHa0O1X5ylCmnQUN6dkZxx433t/QStAHKBfIzcMIIglkqU3AGgQZV5oL
B3jRp1IT13y6qRBOfdeTMf+LV7+9gLkPZ98Pu0nQSpGIQMAjDfnFqUa3IwfJTnvOLYnLnANfQWE5
feRsgd2piLeUWc7x3DT9I6xIxvJSdFTf/k18BCCzbA3kglxJeTo539ld7jdN5EsFFsXGpKci9clE
AJn5WEHEqI68xQaWXnWuz/bTv/H356/zz746XgbV7QkDYz4uH5gJo6TwgAnruqqJxvCFVQSQvrH3
M1Vs0xVe6IySOasiIJ4jvhLTSRpQji5MJ5cshWiU1coEyHArujy83XDZJHs9K63kyqQmSwaTHJzL
Hs0L5TmqKH5iwsEfi+F8mMXpNE7gagM7VcCEqPFRqD7f3AXoF0isslOBTvZouzvDA68TdPf/78we
InYDmLDLjK6GbpgOLJ34wQZ3PFrJEP4vGhGXioPoeFEdJBYuU3iYWeLDCnJCQXQIfOXqA4sanvO4
Q3T+ISRrZBRaA8VtMD2Q3caCpgHIsWb3OI1j1WMeLj8Usn0kKRgqYAKX+dW5lj4bwbjv9txGi8xR
sV+m1iqUyb9WDD4TbCSIJXFPJtNfbHn/23fFYOl/FoIBDdpmRZzHodje3UH2gV39Tt3xWM9/U1t4
q0xEiwq20CkEN/TLhJGqxyeeu4qZmtggX/XvVAM1gJvJulvnzFGU+D9udljA3iS8qnKpLq60ST1i
WENVHmrFGRUAiIKiVqdcttaFosBAxWWlbCWVFhTYqnj2DFDbWifqEdeIGWgAyNItCuRxQ0Zccssd
Bqg1+Sdu1AN2xtSwTkqaSaF1WiWlva6FhK2vKLOgEo9A/9DDP0cKNXWhWaAzSxj/opFNN/N+Pd8Z
2uHnez5pksYwAc4uzthL7HuDojNMxIW2qRpENivC27oOhqJnE65AKoUwFK1R/i7Xt2wp6NsMGbR7
EDC/lvGk1YMhlOQptF+zKvaecnAvImun+l1RraEwDZCQbHVgZNXfdP5pZdqkL94j7B9tdoXsHNa7
7UFiX5hsooOYbJfcSbnKFCA6cjLm0IRCoBtqFBv/92i9zqu+KNURY1x4iWyBuvpTDBhXxI2HnOxw
I/4vXGFf7qC8oYA9Zr1ZDqcJWsXo87nCCWZZcQkp6MePLBflucweV7apssbH6vMg0MuuzdEO6FiB
7kFTsUOT8efYOR9vV8PQLd4LI7EQSNM5vNAnn+F+WH2RftNpKsuR+DjxZtFAuQzvyLfYk52owq0r
BBsSh0h9PdJm2S9VV5EVx5QQ+34fcwT+Y5ihE+1JWKqeQ4MMNy7wruQ9DMxlavYkll8YN2fRyoUG
3zAeVi0S3X3umC3SgHqcyQXWpIKtv0RhOsuya9yFk4aAiPOMFmTe1FVj9lP+6dpk/vmF+6OlSSb2
BjUSdt/eVTykTPhs8j29llvc1wmpfXE3bJLPXM1sCN+DvK0Z749stD8/RjBiwPPWbAgmaNE0ZxIN
cc3PtUFSWfXGNkV3M0VTK+TWkPrIikKlsYK42QVKbPGlFWkLPH/w5rYyBifMZYPJ+M7B6Tt/wjCn
+ZU9c8luhOraNh1gUOJ3EiipYYWnc5AR+TifbJAeDZStQn4MxJFEcse22iXgPVT1EGbZLTRlDCwK
kswSYfVyb78o9bBrhlR7yNJBUY/TFuXkr0h3IigxhVd2ZWN3NK13/njZ6AtydZ88jGJEsRUfCcWy
oyJN+VP1UvUTT45ODIbzvTvRZPmnFXK90KaBzViJLzFK+5W1vt91M47tQI1dLMcx8J9X2eFogW0m
lZb8so2uDGiX9SMff/jOKu8ti4IlnYC2WAQ1Dx7UqXfFs89L/FWvZScNuD4hRspXAs+F+ZsNdp87
0GLEfOCloanK/TeR8/4T7yMrpuEMvOs6zcFOZgcug5sgNRISqWEIJvho0pLVNbQVtC/PFleFGz1U
bDNejMFOUFmLj/jPTuVxeIfZs0XbMaVOWOOGm1GMNs2ckoK6gNli9TL46/AlsTMpoEVT2K5L1f3r
qyRrqYHAvSVhjfSPpIJ1u5F/bdSM67DMeb+NvSJKi+UwVrNkhnliTufo83L8BzKWlt77g+tVrK7c
8haHIVYjOxhiJdgxngrWE9o/z7XjhhbZDNnguakiBimOfrQd1454G7bdQf0SJLr20UabcihJ3Q+F
4ZgtYH/uyg240jMDbOOMYYfdnZk3kPNPDWBHKfkwwJTxmJoByg7EXsX4ERRqnmZfcbhatETn36yO
FXKf3VvcQHDatgwCYHR3n1QcV5mD05q4SNfpu8tNBajYkCxQ5SBf27qMIa+pBFeogGWXUcvsIE4k
rhcfJGAAVjbthDRCZgwNvRpZ7aVsDWVeQQM3EjuplX8MrECPJcm2UaTYfjhBU1/27K3VOmKksswP
rXFpY2q/DE6wt+1KRajwrHjdVTyOFWUWWEN2//jR7JixPw/wlW6UVAqc30OwJDPAKUqSFTDR1IRK
4u8fP9G5tpkY99YgqBBb65Ri7v7a+HAOlrP181p4EuFouJGSVdSJj9ofe5V7P/brBElVJFdOjkkw
XZPsXWwwPUHa18rndch0mF01ZJllFmaJW3ygq8iTIdqjMuH8yepMwPxQrLr9fvDTRCQLuXbXzAg4
GHjnLl4DTysFqS2Ktqfgykm7r0HU14FHkkieLvMULdP/BTJ1vJGYyk4ibtdPFS8QtsmNXY6Xld0v
aOFZ3uaF2Uth9DkyLjO70c3xQwufZ0vZIVGULGuGxB0sQzF038RhphRDW/+myWij+cs95KxHsSIR
AARW4JCExBoVbPSa+QDdXqx47u0XzQkCCQTd0L2YTAedxrMZJCOhWyf9HBsIEiUF383sOywsI8hr
8/cPi6PlpoD8t2ZtVM3y2zLdvacNtC73uRguEl3/T9IiFLtIH0r1mxVpGA5ZkHYuHj1qnBiFHQ9x
I3Hnae3H2LExFVIpHGkNjWGld7Y+wmBJBcxVhbzHBK36n6n/7buYPhC1iDt89DJ5A2NUCRTZ8ElK
U2+bJos+t0G4jKXsofkN2jaLWL60dMGea/gE6rlGds43hhriPMnrrT/fp1guTzW1v6UNOL+Mu7lR
wL1cvOvYyc04tt1spBmJKP9u3mLkLgYTKOKUBS7Ngh7X5OW+mcMKAC8L+mlAwITbzXKwjV2jPJGx
pViCRarz/VjTuQ30i8m1GcZfvV28rwZl/x/qJvmAzIvwJsT0jP4jLn0gRiLUxSvmsZU/9OXF0Vtj
QlEZQW9dTr92Kj8vfNXyFSQEIQA0oEttNuiQnIYqNrStWn6sR2IV69G0xPoKCDDPXK5At/viyW7B
4klV2UYel7ImAOChCZKOq8ZZBtfXoxOa3JGw3Ecbcx1a4dN/RPdzu3763o2QZzrUHuibPfylaCT6
pkL2VGhEPr/f9CAbOvV2bg/LrXt6cLBRbHu9Y6w2X/z012/K2r2OL43RyKCjbesNtOCGCMIRzLhz
Uurav6rpliQub4SoZdX/kl2q+NhtnyVkxLUaPkCJ+0UavzMSF6UA2hAlAV6vdLmb5Bl+L4tgvAJX
xHSizQ0O83jdisxVa8ut6E/fCyeuSD7oHo87pUMLNmyC53dI8P4w5EsgpvBN/7M7XG5q8bRnNimb
gSvYBfs+z2S2uCG82KgV/knoyoNVWn2QwJo/zBwp9p1e/V2gdtNZlJA1nwP9aT/Ty3o6U/XMxEL/
otV9fKph4Cvh5MUMAjADy4VUsPAcw9RivOW2ROgs71ygeV/ttCYumP2gDy1vRxPI96oy1bf0SLUv
2sIqJroEOpmJw4q5CplU1xyZA+pF5+/bzy+QvyVs7/Uiil9RTO8Pcf/QVPxe4hD+K1N7yRc2EfXg
NItbJRwJqUUjdzb2Eha08S2eD046wsJMuDm/bjCUKJH6A79scUb/fUXDyu/PFCtMcakweKAE+p1s
Vq4K4eFrAM9FEaxOWvRT1MaGXpq5CdFL14YaFSblj4rKx0V6JsHW3xji2VUl4Dyk53EQMrgwE2RS
K4GN8nbJG3nfgqZxM/LMRYuzsOtlMegA/FiLOAoVPHAetu24m3ZIIy5x8OjRKgm+96tP96ziQY7v
WTXKmNy9Ug0zvbna5uPP6cHUxRugShykN2LweWIpXbzXJReA8kwP1uaUaiZ62W9yOeIxvTBirkTQ
Ce7fCqUdYOiuJK2IFVYwuMRbRxOLAzw83BNeQzHIId3LrdXPvhO9R9aYTQhJphpKQn/ZKu91NaqQ
Vw1UmWkFXq/WcelOotTFVf1kyeYOUkXO8PAJVlQ+2V/Jm7xEsTBGjZGonjjo0HJwipu4cnYAiybT
Cw86Hk4deO4BMbhKU6NweTkJOh13404ZfRF3OUVv8Iu6017JAMW74nhzTn3L45/N3VzqYFdmMQoq
h/DFjBnGuqzesRVY6nnK3/b0B9cbbo00BOPRv4ubPak62zOtBfpHBzJFkUX+t79L9/Ti1OwHFCWb
c4u5flGm6E01q4CqNunlf5XxN7Pgrl8grjL5Rt3YSIe5SAfk4/qj+n0LF/MPwPARd4Mma2ygSXP3
NIP+9vpMZWsYaE8D1gSyBXA/ZkCRu+MZUecVzRgRuAz2MkXID1bH1iRUpSd8vjWk+VqpviB+nIuL
yA+SK5EluDl94pKuLHeuj3tjY3TZH9W8jdszIjcGSY729TpIXkwrzdrcYx/94TOotJrelYiLQuGx
sLzuc10VgdQ1QQ1+duJJ6WD5INd9irJNcqUS1PX3bwgJLEmkov1GEQ3/QaWP1ehuvry9SrnYg6UQ
6FrU65CCi3+QgQiV3pnfbs1mgYYxAh5zCnbLKbyfn1VbYtUfYynqTykmbqHzDjJnJkTO3eNDqwPb
8bCyrt2rOVmUHBRWAmqwsyWJ87dpHhCX3ALbJ9lP1Dz+9PUHZatLxG2CTED8ua8MLjZmFJM87epv
T9+uDfWrE++NoHeHNzFWYM0Nrrt/+DXceKgTSs8gCGT25OfhSROtPDvEEr8UUAr45QxWixRmYNZN
AFG1eyTusvJhchbwy0KNJvYGixKbQlSnQ5nbidY1WYBaTLf6YjODZj2YLJEgLFzFh/dtGAa65I2V
KNoqZ9Di7kftfnHSGh1svmC004IEiNDAYhKu4qdyK4Ad7SvV6GMZlQ6UflMetXJWqNShT2ZQkeuk
3o0/QTx+Un4vzlgz57Kya1ADVN+QF8XEdWl9tmG02uSiwSR0gd+5z12ugkLQZUthVngT8kuMDiVB
CggmBkqjmfFV1I7goGZwsbng7yySXMOsMlL4AYg2chF+Bq+iNlJoylzGqbZ+EvZZRM45TuyvIvrI
4iPsrmL8wGCuqSyxi4e0cWAL87lWAkBxjFc125q1SFJMFzK3q/kUdiKkzWwMHw2+LdwpwN+uMw10
E7xeDpvZjVADayIO5pz28xZZXfjhIElbs12jhUyZHHgF5yqpZK0n4Iw7efr7uZit8rBwVegtjHam
lxdDop0qa4bGPdVtQIELXhcYSyUzEuT/ZrMWOAB7cu4BFCrcmPxmmpVWIWH6oaus+ZeHZUckdIpp
UX+VoL3Ov8E8TnS7EmBSzMW+8qEGaNuD0zp6E4FM8NYuHWo2Q/+D7YmMqG94nP8o50M2RphvwFna
MN4NoVQwAzIJu8HePChIkkw0A1G1i15DxywSbws8vqdETscZEnSW+Ns6nJENVrBhPJaXs+N5jrxm
kxu+j9mdEL6ddJqSZiRVV5LB24jO8ZfXE4Zh4F21tGFN9D0y/7gLid/+hl5Q+Ew2RZzYY2zUW+7d
t8rhx91MCBJjWybhRuN71fZYNE2pBh/GAJ6ooi+9tSjS0GyORuipo4ulXiRRLOBjOFdZripOW68o
E9Q6baGG6gKtNnvhpKoecZh89LJVeYvwrg13euPpcHsCm+ZggBGNqp7OYpQlnULUSM0KBT5xNW2o
OUGK0QPMUGbQDDunWKvMVyi2wv7yycAgjq/E0el7fnMk9QJ2TK0c5unTTPw6c/mCxQXKNR+sFJ/N
AtCcyxNFFvlnw15D9a4zurqQJxf98Dt4OysKPFNj5tLw97yDtCswSM3d4YpxGpb7NAzCkkMXOrpf
FAALp/exRs0L7ttN8PPFc3jqnIVd/2+yx0qnMfuWIcvTd9NyyTKuWIH15Wywn0Z8FTndID1KNqPi
Mu43sXB1iayXZk9U8Ne97VBIMVHUkZr+PW8qTA/vVXe1NWelzruC1SCEIo1mXy/99wuDeQ7XcVzC
gL++Lly14PWNu3Uv/Shj1VAWBAANFWUpGrnNaQmFiID1LBKDFyOMh6iDviCnndMsLiVqAhs1ynDN
hXmmUNbbu6NHcZddf+3c4YOF6ANLOPdUArZCxUerRHd/hvlm5VmZJ10ZujfbBQ9VPaOfOLJ4i45H
nJlEIfjgtYDSblRCeoL/jtannyMw7SunghEkUNUkAE4TgiD0lSpIcXre0xX6oaJZVQP/crCD22RA
uBMrz5vpCK9W5krRJIAEw6KeqpibiK4MOKPiLKwjyYRSHZxcBU5ftHbVoAPYICFEU4RC8MeMDrjL
deYwZTFUuivNaN1SDt9T6Rxqdkq68LBYeMTWNFMOkxfpDlzhIf3ptR4ohrRkODyO7T12NPnr/LRe
7Hq/frTPbbk8KDlMwebZrLosw8koIWW/jbN+Uw43vAS9k6ffRVNgD1TFYZZTgqGnhKXmzwJUEUXM
t6UmtewH2kBnkQk7BQwmZuBEJ2Jp5F5U13BHwdT5+K4wGNNRSjITWNL2zO5Kmr90yic+LNEs/MFF
ac/nxhdTfGpKYaEjnI/EUNKlupV0WKKrxxvArqbfJgt6CuFg/wtfAx6Cknr+2moTDX73lMZrb6Q/
UAwg0SZ7eHulZGhNojHfIhr2PsoPg+lbOSxnsGwGDlPgUCUtdgewSI1amqYM7oi84yX/AeVfSd/m
zLAswQObl0XWTtPJ4ilNsYFiXAD26WNL3UeBQknryWhIblv9zQYKWSt6L7Xe4aWRphGNTpNSzc60
PHghdwpfd5lxK7qCMVuGp/v16mgxVq6L9KNHWJaYp9EIGdK2daLaaw6PUUBPZnSDXguY4xWmGRFe
MK7UhOAcnF5N9RVx376F4IpIOoim4pq8KUSLBeH7NaoqhlY5U7WCyIKOWSTcPxV8W5B5/ig8KPpN
9gwrEsqAyAtNOGMvYKrd2fedZmpN6QuEWCHFng1Ci0r4Phmc0POPUwG3qyK5wikiiaVK+EO2B63d
R70LJp8Ek0nqKImw5kkKBDq0HEvANHjR6YFhiSAnN3mxpX3HXfvGKNF/jNd6Aw+yJdrd+lYAMCyb
jSTSchOCaEwjyP1pB+4IN+c2lUxdYh3l1A7xLPyTSeLRK0EIAaPMO1VwUFd05BxDpQS/N4uRrILz
gsyEzNbef5MAPD1RiNMpk+FZ1ljyBEWqhzf8GOWBUxKvRqyI2/d27Wx6gnEJVl0oxYcsbFnwt6XR
5nm7qPgjM6z5CxoxhfdBW0zND5nSGGI+WH+4u1rnBPoHgR5Pa5eBCb4S6dcuvisSUbHq/+UkEeLb
6iBca3gvIiiIPnw27X7lqQc+A1ujOs5VnFZrZS977Zs1smoOid17fSPy+rs3kQduyvX4vmMSeBoz
rxCxpzWZCnPaekK1DrTaWboZzCK5MqgRNx0NismeP45sW3paewbeiA7ZBfKSRcR0lPE/B/mv/gIo
f1GfBd7ZzqOU1cooZ4JSGcJpToPRrO3soz4EnurG01ySGw05nRwYt4j4p/dKz1HV4/wxcfB2eO1Q
U1mylwEQvDEgsQhCEZFIStBKlPRtwZddw37mGz3MPTcIbFJtmNrCXI95hVR2cekjEnrAFiDO98ZP
lFCK0BV04b8UWH5C2x0cXS0r60Oiu9MUjC70IDU6Em72ljOmNhZY1pF9okjWod5o4YwXuf41s1pL
a13f0gX+H/+G1jdcUF5t+RYrUvp8UN8LigUOea66fOmm5dpPlYYvO/sGJ6hIvAlwBv2S6sMxGyp1
6c7c3nqiGx179naWKsQbxeNuS07GZpnTFv+goV0Hv3CRl2MVpy4Oso7Q3lu8X+6u/rOP/TN6dUHA
oDY84sA489m48Ui/vPb/CEcMsHfFOgARQdrrBulEJJjEBy1pF+S5UNzdG2Isd19MXXV8nhz69IoG
N05uLHmxQsKhQT5jr8pdr2nCaTeYZn2ejrD+0xWkhoJuk2VmYQBGDDQxjNAyj81CZuWPxBrVEnSR
Cf5wZeybDJw0HmUvYC8K3Rb5NcPmXcY8rZExGlQNX1ARJ417HBjbEkDixKJCrMM6hNrCzQkPCBpU
2OZpARwM3qJJCG/lOGWLxQVWQQ+ZCjC278jjmih79UzHO5aokD91H1x4jSXuC69RXL2vwTn06GtU
yfidvpqm57hKb3xRJWHueJNpb0BQDnE0zg7FfoZy6Ds6KFTYS3uBdGc0sacv+Qc7E3Zng3+UH6+q
e/w5d30KyxkBzpI0j+pGpfKRxC95j62QnAi5v9xsf3sz1mckyE2M3wAik8Qxm/NVD3zdfCktSZsP
EDXsRDtSP6lJghLksdJEa+eqtm73P9Ith6NxI1Ds9+gG26HZsOZc42lZUfcHeQYLohvwKvurYehl
zKU8uNPsXvxy91QNOldJdfvDJ4s8cHigOZjQm3Ef0NkzcrccJolh+fo1m1HR/54m7JnmgdrOFV42
KWqcyhgTHnoEgkuFbVS3LGUmWMpUoUrvAunQZ+p1eevynj43mWws613NISJ+TyevuGnwtN0DKe+7
j59Mo6K5LcgdfyNKWxz29U3/Cgvwt5MA8XedWffgyFZfwVSzZART4xfDBnVTLQMX0gagWBiT2rD1
S726sNzntRcM+KKUoj29lIMUi6K7ihaaqarrGrl9BsOFTkoqEIbaFs5AAlcoH0mzd6t/u7rAlcho
D76f1h479HBxLsrPhZUntnHfVNBmA44OJdlvib5nTTh9zOzrTpRUQSr9zl0CUttqFEp/k2uG9/Jp
6AxBi5F/JxvlFD5gWS23yJ9yyE+vmrp71z25JFz0x139uYKBEw+RJ+gn4jlsm4GYJ0k9oNJEPpCl
CiagrOPCCUDAXzM2zfDAxwYWxPbzYZbcDiD2FMrueUQ1ZzTwuJ7AuPiQWJutDx2HgQ02w8SRX33k
qYMTIQLp5AVj8j92VO7CqETks7iWKcwJfSXzKrOHlUJxthGPm+p1Hd/jQ0tIHmiaU8bRMf5utgzU
wwxJq9e1Ec8xol/j6RgiuvCTnHW8kFgwMp2DwdtA5otxoiKD67RwwxnpN7bRnxbN9VxCHy1aD51c
DNKNQqRD9d/Le30ad1BMb0afjr3ffXgwuJCo/4MvR5B69odjPJ5MUDQtElwoMDGKsMaKTRL9q7Ev
4rdiMR2RVe+J9XWsNXUtw7tKpK8CrUYNHE1OPx1Mr4u2HnNcJ21kivPVvyZJMyYY2DrSEbYTGGsu
XO/2xa66m0KqvWfpK4s67Cu4FppB2BY1lkW9VwaN5CyH2IT6VIooiDRT+KWqvgBWVS28ACdnRuGm
/+oveAHJdrm2Daytae0f33h8AcWh89OrAtNWLjI0/+KGFel0ylzyCGfV1bxdmxXys6TxTVvW1bKL
+IQktxsqhxMUu2Gd2hx6CGyUZgF/cSKPWog9FZcryC6HcXi5S+9SFwuj3Y02j+gOgbToeYGQXHNO
N+LPrPQsvi13nsnHgP26EDo2SloWSvO80yp/fR9wFk7e+vbYjp/u2R2BhZYNPQlIFk5jwgN426Ep
zvgvjjarzmjI17xzFNGkWUlQVbzGPoMv1rwy8FwVMKWhoE/mDzhZBeXUjFU3lRr6JhPeL1bIwWbh
xtKUyKl90Y4d2hRIk9xjo4HY+h4yohwQpqXNCaYKtq9JKEgM7HAe+QoaqFpIOlPcF110NfJgeJs+
qudXGUkbSAcQK3ry4GdETS+FeeDVBYaWoLpfd+3rXIh/sA/O2JU//TEgkLbKKwWAVGXWzAUh3giH
/vdHHlyijw/8A9BQf6A0smO+q+SbYSd/cfhLKWsjh8a0EUVZHwuwmgyhfEnNltmE9Wn3H1SBsSU4
lXooXF6TYc3qbFIU6lXI3RgY274OsiE9QNDo/r5kiDQBsgX8vl+Te42hiqJPmvP6N/S68S3r4RTO
tHWo7UpFkpEUDOi/Dz9R6UMdtHbp9T9MVreaza3nERcWCanMfoirdCYbFrS92v8a3zAM4qa61Cuf
LkFo6nypHQWFiVkBSzsX/VahK+UMwRQpuPnO73SR/nC/kXwNYfI7/JgXLkc4xnNNUEgTbt3cZDFo
tblCFgeaE0h6AftEgAfvdK+ediXGluY1LdcybJ7U9BmoJBjIkPBNgpmG7otbW9ZeO9IO7xBdJ9dG
B02Fjur7GiDwInmatsXwbrEMBCF7aasEQ7e4/rIXIMPFzWDR21Vg8IFETjjHOGiNj5ofUqh75OEa
KG0v4Kg36aSlEmEOQfxureAm7d/xPJeHoVOnZRh8ombV30jxyHEL+WLjkClV8enm1r6/gvSl0T6o
Ym244oYJvW4NeXo7VbMa8iEggZAOLwChG9tGS5wDtUa+cQRRLXKk3c1+3br1p+IjW5o6AXU6uEbD
/rToExWsQbC1aBRzjs2Zsb9k0YbeTc9qTiWKgmnvzJ96BcvIAHl9Tjt3/zQLxjiD0Zychvnv4EB3
ZOAqkFKL/F3oUyLGT8xkOfLaImM7K6ud4Gs6UOqgo5EPylQS6fmzotmT0GyrvC/IS9mhvYQDEcg5
LZNs73jzFCMjGN5FpBL9kaP/0Q5f3IqCWsakAwV5zaqv+ZYeht1dJK+Wi2q1OJ01wa9Oad25NRzT
UF61aMSOIcoYE05xJa5M6vnFY/7fEOmVDo+A25xyqESV6DegnCsyQv+yKC6qHlG1Q+GcCQE0OqQm
hOvfHQP27BKMCu7CM8oyG2VAqdce6/l4GeUnXIs+6ukWa5p3EMvVcHIYRvEGNuiPfU9o0FMDSdIF
tOlM8GPJR5qxaBhT0FxsE/aDSpLKsy6TcNNHROx5wRHZg3AtMGCne2dvJDYH7cktdbdEkxzsCqdm
49CWq1t5jdULelQQzY02Fi2Lv6hAQUjf0RKzRaZ2BtXTX0j46budHma+BiLl7Fb+YYd9lhezXvk7
JhX/ZZYqhFh95LCy6eNU0VGhCkVanZ+xTmXi+xBGbR+CaKw1EMQl5rCGHPlCWMpfUt+eDYhgGHu3
dD7qmar32rM5+yv4+L+RPzd/K+sLzr9acXOPqzzLstvO679fzWp61n348pVWa4JQDUf0jSyyBagT
A9yENygeo/JwJpee0RiiBAZ6C3lo/IWTTqNZDrE9oh3NeySrN1/GGvEsS++J+vacdw1Cq1HQoSCc
2EgY/hVWc8uMzcLRofzpld/VLZJXZwTIxfoXlRHp0CdhHhfJuSQd4UaMX2TuX2q+VL5FGYMvZ8ni
jNqzsaAHRTwUsMeW3zJOvSqRT45TzpwED4bYkbXNcy5KcLNxv0ipsQHXdnLZReqRUWpmUgvWeI3W
h6kJYnMFHKsmdsCz7EZ7Kuz3Rl+I2/x+4Mck4P9ayqma2qJ2iE+hiKasQ2630VoiI3ifofQYjAeD
Id+sJQKbbLq5B8OrYSv8wNnweli1FJ3rhy3E1Fx4VkIx23YlHjHfh+lDGNKcGPEcpRGvIRGEreUa
WL3XOecqBxvwPMBFL/wetJybOXXNR6Jhb48ovbMtUuRZqWoXbQLUXjWGK1FUF3jaWLLSdBWHcEYi
ybPIvU0kZ/pbIuYz6VFh+FIxdXr+uJ6A7FxUZorKSGtccCz0aajA//oyop2zaQdvBTTNH5MXaybL
tqoYAabC2pJEvhkBRX8I0b7rxeOCg7bXAbOPkkntZiF6OVzyiWbEH6KoG1rQymRkN/bAYRmyXayi
9u8e68bAiCqdtkg3j89KjU4jdtgibzIqlyQ0ILF25do1zwnGtXZcKeQ8/V4Aitxt2tSlqFJDEjoF
FhGlXWtfUyH7mYRdxwIiHDoVF4nlft3JlRAL86R7nOemMYr6fQ6XqTCUDcBAYtdTKD39pQMd9r/U
a+0xkpNE//fOyaWfIACxGgrpCBwAZEL2OY1Dqu2N10N6su6H5JCS3j99X5SYGSNRQDBfZBayigv/
gGSmLwVHMKqw4NVI4YFiaTK1c8j07uJ0lolLW+l3tz6OVifNBOC6LS+DdpPtoiaAWQjkNehJe5De
VjNAVjgrOHIYHkRKvgVfDYMpPiU34Yi2/mD7lvXdZEk/hYpkhpb4joNra3WqpHslbjYY/ivXv9nI
F5u7hp48qZqOsO/Z30b7UlvPgMGkG1vNwqQf6FFD2/X9FLpJnom+FL3pkG36SCM/UKWV/d63Txci
Rwi2ZhboIy8ieraF+EdCZ5ShxelpS0Rc9dlUhIYtWZ0Xrnc2GhJwCBhdnwxOX6mYkMJZlZ+6OZIe
g5G5nQYww25ni5CK92T5fMIArQYhgA/Vr8UQb6Jbv8J7UYglQfmkkzXmLDRZ4o6G+gLoYGF+I9AK
J5XUToGoxeSyszT0B9GNLBmtGq+L5bkLSbvQy7hc2qICPw5yrJ6VhF1iEmFLo2nZu9l+fvg3JcaN
lxr9TRIvRR9bsglCXiiEyzuOsZQ/XH65Uk76xJZAMB8bo1+dUnrA2PjcrN9FeGKEg3J1a+SLiOCk
b/Yf2QicP5Af0We6aSi1Uhb4bQnaytaRD8fAtnRiv8Lots5O8J5iy7V2sarQV0wRZDpKXPov3dpJ
Aew9ccq91ryUud3uO1EVgSCle2WkBjbHORcn65Xp4wjNdKGw+fOpITZ2knIfbnBd1O6JWXAb7s3r
O8p1GWvMRmDsBiZ4F8xjD8cjb4qaGf50h3D/rFKkh8Eif0IJos4+3ihoerm5b8pyaIDFq60n6mP7
Edx27xFM6jGf4gk8B31OI3Un37ErplKZwOMFhFnK4ostlZXEr1y2PqxeDHcIASiTs6RacBclD+OS
41Eooqt2gshOdFgdHAd18wQ8w5J5tnFkZta1VqCoBEPVxZbTRlGTJW1LrF52+wlcSza4ZcngIiZZ
dggQj+az7wdi3W55RgTLxS4ha4fopq3YfVxNvmCVADvmtJOA+/y9MAmAziVeKe25OFxpyr0ZeWhC
QEUOmWjUr1Ick+m20tJ/DXuCX6iKFgrzubTXmgZwcEQShA/f6jVFKxz8dy6K/hmeTfr4hptnKGqo
9w6PdMNGjSY3Xb04Ur+wIlFC2drrzJRYroansfP8hO8tkhAbQ4nd0nPvGl1VbDpSzDn40cBMsQ+7
2TD2hpjttK1yKgv4JoHhA2kAP4I/99gyF/Of0OrmgcKsXtcgRAIVZm3LM6b8A9RW3LJDUb24Xlyl
fSDMg9O9r+UKuu8uaLKLWpacrvwoNso4HDM1Fl1bfPI21gjz0Wfi3LTMT1F+5d9a51row8BcIZI6
ZoIhaFxrnIeCOUMRCOUK95DqYZyTla2UFqCx1BmqxMUQY8tFW0rp+CDxI4e5wQ08hQwvlMeXXmBy
rUiT4Vc0mYxsc01dbUTS62DsdS/IE6s26OqMYmdYHDrRmKlRiE+2EsjFkNoMrFXXxMrTBHmKsf3t
Eh/0DZ4G3C8IKNrOMakW06snAH1Li3FvU/zLWRz+Ec9dd5DEztMZxy89yYmeLy/Jisswzc1qiKFy
ePlALZGUSUnqUQIS6vnYq6e5DX4PP/E2WQAwTd1g59GAhKvAuRtK0613+l6cnJkZoVRb6rm0QDv1
OsmWhpVmtqHtdRKrrbAIt5jBKxLYoOWekaN5Q8n8mDxSwgSvugGSsHpkyLg3l5PHN+7phw2HCqZs
aEg8/46XRzV3bQgzw8C32Uu6sx0V9jCIkDKSLWzbKh4/uUUAdYCujUQf1d1LhQkDFLqKgQ5UtZjG
wYB5DNAYVWgjPZdwMeg9khVM8VFGQ6N7exsqzJOhpMexoLsTPP5ZSKAp643+IKWYZIVPhStLqjfR
BtdNrctm9mjzOoKjv7dKetggkMvCHISi6Mn4ZvVj6ycyvlUnqDz/lEZiz3Lo7ZRrem55ZyX4y4jp
KrLZDgViDq0F3I044NuUOOvHs+VgyDgAb6kViSFeBfY2HteE0QjZb2ujXWTmZtFEKVoIZsPNwJla
JSYVXKP8rTdU9YOo6HAb7UYGaw1iJ9P/8OLtcV0gOR8NWRrXvJiILTHmQA81oEBoKcmmgh2gZh0P
XrC33t442PQbPGBJYVDqpL0V5qWhRSbcVvAaaoPqdKw884giKFkVWz/mF2NZ3+j1LyVUnQQhTXuy
drr4LxvJ3f8ad0/XVWZ35ScKCTNsVeZb5J4pZNnbKgeE0/mKFdVBbtnK1HP5imDgIsVbcOc+GvVE
GIGpXMmoCzrcEB4iLltWvBX0+MvVINqTRDcDrR0/6vxWgjmaAVrjST+/Vxk6Ct+v5Fh7zCIatCYU
DQExd/nLqDyIDIp7TmMDtkxm4qmUzQCB2aUNfRT/Fg3gIQTW9fguUFRFDce556CWG8osN00RBBzn
oHZ8rnyQP1ObUmPPUYa3M85ZGuO67RmIBW4vV5OI/+p/nCeOw1BPKlw+uhxpa96wiX8BXglihuy1
lVpGItsrl3STfrgBf/fyyu8CAqSCBzUknVVzcAIouTDN/odbHbNpCNxcxt74BtI4uQG2NuwMnKuK
Wl7xV++UE2JpIQCiiAsUvYXkiPmMTYzLm6um+O8Y24jwiHqmf7Q015T+7wcvzaLV2gZCzjETb/8A
X63Ab4IAEcbGeiAa6Mef1WH9BK2JwDZuGdM/l3Nk538Knysr+LMFGrtVQNPWbtMlnjC7YeYX2+w1
R9nsTBL/skIJaFPpl3cXfE1w9FnIWSAuLlCbvyJjI5ikQ9c4nfCpoUXeFzcicTKKh6JA2OQqHatP
bAtNy6Kqr7uAkYvaCZ2mzf05NrwTd+pVkDTBlMKaayCh++27jfmUE2pScDdxXae9wiQfD/IxSNWJ
1esasxb8HGFp0aQzBScPnxHjl1N99N8qgT3ok7i4eOnzHYbetlIToyRBdrdiXV8o0xM3FOETr38i
u93UZtG0rvQhYQOspxo8wmUd4cNmUWyga7Q7qul/I1TU3K6P6gz2w5bmCYg5VU6p8KEo0CvS/XPi
G4/gOttcAiaiuhq1M1pCJgG8v4ljTpIVDQX5tQPe/2oAK1ho5uxGXLZbN1J4vdH9QFoQ0vWxOdKL
JqZabWL456zKBmQ9+wsadjrgwj2m3yrKCGN+KjCtdLysFShlb345YLfFTVMDxYGlOw8LldcbtARa
lriANR1sVBQo+Vi2te/yNCNSvEyMC8ieCdwGAkLyneDhQ6KuTVz5nyoCHW7VMRbkG3jcG00HsAvE
4UTK3l5xSvoyqAjyiQB9taBwmHldFshBx9Rs+EFthLp76Y2wDUMx3lBJcmmvw8sMJ0jxhDBBOoEP
t/bTN537QUJ9BgbnjCPTusPBQuT0Gl62O9PZ88rKVlO1dn5nsHRozxrap0aPn+8MvUsCVxGZOobR
xGdslqvflRELoQGIBlubyxSBMyNO84Uw8d7J/ZvtuZ3Jt59j/4lNZWHj2CWSzPPNKVtvHeaH9WaJ
QtWoWKk+tY+87AVAQQ4/Cy9EkExfpQDKaVKxugk44tQ2TJH4LyqpIRDxUSITWoWcTh+BWWrzRVdv
hsbM60tcEsT+IHdD3lFbvNCqwUqpSlAgm9TaGqhViXDM1JSctvyCOBHDlLCFjvq0YhVKrhbPaiR4
OQLcb9SvwAtqvA4eyhEqsK5NgwxSXeYcGu95v7fYk/Ugi8XvDtMgdy672yUpezRR3bQ4LzDqUG34
uAqW6GgTdJ5wtZ7ZJ2HGqmbZxHTmQEV9CGVy/KaPkdMYbPeulL6c+SX+zOExcOf6TmLe5P9dNb2A
hv66k5xgWp+6Z464GxzfmXNgle7asS8IRvR3dpV9nH4kDffP9Kyq1fSQgj0Jougtrpxi6Q2vlqQs
rj+umkA5WN2tG2vgW69OCVgsJRtV5BsgA6CxzrDC9IFBcpqQROSn94IP0hnd3fAVSM/WrUF7IhkD
LNJOOvntHuWNAao8DjnR5UgJ+482f/3LRVy/YlWvMjYLa/xOsIrloxKevv5CfGg/iGgNCwN2vwz3
9otN+Re6SIiMCmne0e0/D3ftRqPWF1Zft6O1I5pJLdyu0SuDBb48LK4z7cLEirN6kKsTKOtCzPwA
yw/KvpCBZsM5huCZYXw7s/kXmU+H03rs5leiyx6FUBdB1VTkdJT/5prMPzXydhXyIcaFjn/HSW/Z
O8dhQiqWHyx855QIfies/Uc6kvarTRZbTg6MFIICo4VYNIBAsRf/fFfTgDnruvcRsd7YNyG/UI7l
v5h0ycNP9w8i3IGz5HAmpR/gKhk3nAuHNnrxj4QkZI57licNW0LkF3MFAW1biAZ7Scyyf2c3/jFh
y6x2Td4h7N3bAqrK2OkrbXDDkCdMZgfrV/QjpowHvpORXnIdH0ss+T2Mm+E/QW0AjUt9EyCLDHjB
ddZb1p+ZNxHumlWCReVl7CMjPg+fhxrkEpvCvac4Tr1qlzY0J4WKFUepL9ouGth0Ex2q+XJLExI8
6lrayWvHTnyWYA8aRHf333ZJiGPsH+U7vAarOWqQ6Q25i/MuNYfBOm4bBNp7Czj5pyc5t3hNX+8d
k+17iKZpSHd92DkRRro/3gayveyFBXOKX9j9kKIh4d6M49W+9Tm3EZHR/Gncf0AMv1l1SHYVgWPB
Gp1x4NB5//88IZxmIHyW/LKseQbf5lvFYQ9+CIjIWM+PFO03lyg2Gpxw86F7uzt9pMEBqTeaWhW7
WdYTfiuA5zXzSPTeM0K0lKnZqKFoPgWVDQRAJqQ4DSK7hgH2bowa3Dyw2oY1tZypbq3jhwvttX5u
U95Ad6UPzxjJlbuX+7VdAAOKT15hTlSIX4lOJZFc1LWkogLmjhfqJUDMm0QaFcNyj0wN0zs6z9nx
ohjljnr0YziEhzcuFdNmnH67zCsUhxpm2LW4k9ZB+FZw6k9YzlxO7B7sdm/IGpvcddBW5eoe3Hr2
pm3CwUBaSq3oB2IskoH8HSu0Uo9+7vKg9bCFzzmSQV+dOpSsK+PG0/RWsFUQfX6gMZm4GbjfyO8c
HOOALDM94uvSK0NE7bcGQy6J77/AjXFzOCdmsfnw9qooetrIOIH2OiLK0zcDt6KPh7gMzEkngb+B
74dBMbWmKSmLTPzHxuxQh5VjxkQz9kf+JNz+4WS4bF8yqxqQZRHQuFDEuxypkjcKY/XH6W+CK/+6
tk25IRx0XkbnJFfM+hrJZLeWw9WziZa4PCgJ8elGN0I7zf533jjNL/DNq3jT1YjeINjSVPUlw26q
gQMgA9TJI+c9wXPbAOdbsFoP2COFKDQCDDEQDvMTP+9E19T87T5XIYrQQZphhQmzU6ew5LR4M4Qn
4OdJ1kRsg+jDFJFolP0rRvC1q8/DuF8WeeFt0ifrJdKxMa39i7g8p+9rcW0hW+Fxve1yFZrFKTiQ
F49PYc1uWZtEzSjGfAFSayCfRJfX5OIAFX6PZf4XFaS+XyPflzFcW1DbcHW89TPiHSq0r4eHOOZe
l9TcNhca/ItS5M/W+AijdpQnPRgfpapmBU+5oXLY108OEJjVM02JCZr3g1dVf57mp8gTZBxdjrlG
HcLDMNDuusowfd3RkdcDz0ORgb8s+HEo772fuMDd19qBYOXymJhMx+vNUi0/N4vJcxlnscxk5HQR
62Cci+oEOw1xiQekYbXOc4GRq95nBn/Nh25kMci/bFbSlRQuF1muOz9iZhV0xFba0PQfkSA7Rcc8
tGkON5xKD4xTkj208CHQ1ZYbd+DdlkyyvkLjr3fvYx+64+taCTqacWO2slhXQDv6tRmNqWNILif+
Kz6d+duTcIS+HtTVpcn47+uXZsgP/IvBnh+9ILSGhryfBiFRmpzPkfzbxBfPzxcfElGA2Xp+v1lQ
Bhibtjs628OCL7IDjXwhFkeXajZqFFLcdcnzxPhu3TGnnnO8gQiiPNyl0Hsu2TN2ho9duHKsxwV8
vIFL60IxzbUb/jfKgdOlJ/yqAciiVIqUBY9SvjAubDBVRcjpLralCm2m1H9dteeQxLG4CnyX5uPO
TOzq1IUY2GGWngNJEnMHkAjoMth9r8jblIkFZZPHrypgFIQsV0fvVQTiR/5nEQgRQCYE9jKYS08z
MZ82Hahs/Tynwi64aTfkeMd2I/HrNqyYUdSZvJt61upCwZEw258UFFo3JI9MuDLMCB2Wy/JafRWg
sh0za4o0qzqTVhc3ah4eFb0/xbdN/bZjXqGT8di+n79UQ21T9RJHCJm7chHq4cxU5+xxm7tKuFJb
HBu/ZIzk2iAEfhV/sbPBvT8Z48Q1w2kuJQI4hxpPc5lFaYxRk2Q8nS0YWMKSAyzmyH8dRLv9UjEo
VSHDpv7DuGSWNQE1yndg+dJ8Tr5QxGYuZlB/G3Nx0vLGgj6ooxzohInV31JMUdAHqyuT8mmG2GiD
VNQ4FJOF4tPdj1vwox90nQnMe110mHeAMhMAcCg0X+v/EnyhR6M5beOWEejjkc6Bj0MTPZtm3yqT
pnD+Qq3DM5dqNOl/dj2LCLQXQ+H2+z/8/AJQ6ggm6MGla3dEtztDyjI6uJL3tbY1abM0pBEqynPN
bjsiBia5/A3Bqx2YS4mofrItqp27j7TKfcfgDsEWhsN1GDgOJSIkOGc5xi/iF3cxuWWpzHXzhiFZ
ic7MGic/W/1wlBGystrAA1uEPkgjlSXpWIhw9X76bnPYqj3oG+qu5MEYop+z28LIOY7XcFTZIhHx
9/bZh65MgqqOVUHGiWv+vnfmpStoFHI0nun5R9Oed85+GMVXSaZ37bb7HmmTZLvj8pxKwocNQuNa
uis685Av+saBDr00Nu65nNq7gVhfH/hd1LFX+Tu7GngCVov5ZgkPCPom9CDJFgz2USeFQEJdepdE
VAdhcHyYCI0AQnd3FC3ytFkXU7Hng6y+ogIGN1Jj8AchthanQ3Tpzjug2eWBX2EqMs5POsBNuk7T
b80bYRwnlfF66OEQASzN3QWkZEh+qCbl4m5g7139DbzC+17VEKr5gIiDw1BcIFnTu91yi6ggIa+5
kPNNrLcKNYDqOnYXCJBJsrozhpMn6AKP39IqWUfEhjrFmMdB3bh7dSO2OcQUxqOwR1x6YP5OoAkM
3putEQsDM24dlGA0Fb9lUFtn6N/rHAMWbWam2oGMSoqSrwiQdWkvYDyuLIS0tA23iNoTGAXMstK8
tJByfjabOGEi8CTua8q9hyMgemVLQlQa+wVv3yeDawayBpIhRV3KmT0JmB1EMTDQjyQrugOdokbb
9ve1w10jYgEEwU7sbbym8/kuNXszggb4eIebRaOkCXaz2TXZDHvEx9PXG3ZPEDToBT+WwhQus9a6
LIlTbjQ2nCn57IKmPsuR40yhVxyTEf7n4UYld038l7NQVoHE7UhYK8fpdkbhHYZ2PFqM18IIcBwt
qUS2sygJSTQ08pxD/sIBZjHkGKs8FdmRCp2AguJGSkicIsuhs3WJ6JCBw7X8uCmX6xIOcjOFUC5z
N5ZYEQ+on81s1oJiCD577v/0bNyvfC8nV5aJTdHltaCmaY7ke/RQnZXQgZyoIEcPw+VsRipizQZr
H6Rnq3B2FATxa7S4RXnXiAwsZqpHzUiclmVJ33xtzzyDdPBgRPSkv7aGo97j2s01hMzC9olegvW2
mupLYPYtoqb/45HqQMoE1k0T/viS3u5oIXTqtg85c5moMH6Iyem9bqnfqwcQTJlGH/lM+ZmkCb5A
Z4J0P4opgQTs4w57XXe3iCJYiHVdb1lwHBp2DD0xcK8uCHtPMjfjwR0JCb6KDpC4P3XBbY84MwgP
m+mDSrmYtDR8JbmSWdLeW9BXyDtocsqPtA7SN5EXT4dxUXuEbbPjz3FtsgwGXb8yV1+9GDi9j5in
lXiUYvy2j49xx4RFQs31zoauIdtdCJpAr03Qzc9JNf7tJja3G18EdatWwMkmvB12+K8KKH61bFQQ
xY7bNbbZcdw5GAVMG5oyhGMj9+LW/9j5qIBAl8LVohk4jml8o5ah+XHtJkkNhe5XfU+4UHVkABjE
Bv/1JS8GfP/MAaF+9ewqGG7kw86dSlYbgg/qqS6r0MnkypuqDmdYnhAFDOWDWBDKvvV3X+TkpFzx
9CYU5ss3qxVKpqNuzx5ZrnreEs6Tzwh5JQqVtmTXQOsxCT9jwwCD6+fCl87WXrt0mV6v4rK5eF3f
tY6/vjB5oe58uIfVh2DEIGVsDzgodkdMZyZ0HFRNFEuJh+LuzqYLCDl8uKh2fVJzXozZRly8jHXt
tKNNvKDCiFHPF/oZL+Tuuk4+OjHXp7ks01h+c6VLIqXpjAbqgHdLlNu3ww73sinYSLUfClFs1LNI
sDuJdInVZT6ysLnd1ul8M4XSiC9VSSMAjBa7thk85kbgzbqxbw3mL+B+BJxcUIQkBidk7FmF6vOD
mC+Nx6qGk9+50Td6jUF6qCjsgNa7XuBjCsPZ6YGbwS38Fng+8nh4s5pvQ06keDQIhem4o89H5621
JhPbgXTFWzUsj5O2w0Y4K6Im0F10AshZ0+RDa6SJVlK6JR7nX6xp4cTTo9m6OZwzL9CFI1xLVSiK
nPx1P21+LelxTKb7gmV2yqeOFtDXpcx16uokLHVbW7bvMLce5MSD0fEen5NmzsfhqgaKXCDFTATm
X4k+zqxbDxao2Q2wu1tqMRinSoJJ/01upWK47kspLc5mBhl5uo2jBpaB7nk4ywAfNGW/cuYAzRt1
m0cQ1qE70zNWu4ii+xPKxszslSRxbdJ2qT4ME0tJYTc908B5rjGfYvgnjBbQh6FqDnMW2MMvjsVD
KYCx0GRIK9AV8mV992edegIfV3vVOLaGfYJ4VAyhg9V73vm/N4gnYDJuwBtM1ya8C7Nijvi7jbQj
yERUQRr4hEZtfQ8r6gWZd4wHwyBu1+IXBRtOhaGWQ1kQRiUhNbUZ7BlhbnQOr+e3NKZFgHnTtAj5
U6S8LUYCYvguwKHTwVCaccq1lbSmM/WBCFWrqzphIG8c7HmEaU3vde+6HnYhwdOoHjzMEz28HG4P
DP0dLGyJ9TePwoixy2fWK2Oy6iE8TMM4dM283u2zwP3YCh0BtB6HaQkA6EyhwTQWPT7q7rttN1QS
CdWXOt9XPOetCdfjljEtYmDhz6pnW/EDPJilCe7/2xXaWXoF9kOVRbipM43UdGpAYFUvAB+KEGnn
TtmBn/FNZFB61ddCg9xamDUyqkXajDShweI6cPvy/v9Wg8cXrm6JoksusxjhSrU15FKVI7pBn8pv
eynalj5/jUwE/fxQnIVWt70VnmyVKwq5rrdhntL/46gbzalcini0ylPYhIFj3FQjxQuiVzlCvUBR
/qXcbzbxqk7lxWRB+VehsDcHsspn2DtWsRSB6L/Hc/F7xTPVtq430gYUc1+qg431sPXjrcWu/7Es
P9+aw4Ji7LXWgKl3QBgtsTEYH3SkgXfOlV8ZVdb3QqIvAgpjddY0gjIvgiwWjDkXSaq0Dslync5m
Ir7d4i0h00b5g6QOeFi+SPFm912AVn/TXpq3u7DPi485iDFzRHwLp+LXe48mIYl9SawbGjOZV8NO
LOhfOhjAk2q6Laq8LoDmDIQwe1bumQa2svyMAtS7ElVe8ApqLWelElET86uzGA140WZwwXAPjanQ
fn0R6dg/0cb5oD92Retv+hoggPEtWJNqfOeXxy69vDFByKv4eTE8WJ4nFun5kwC9PybPxu6n3eHQ
pD6MkZjFW/c30o3U7lsxwNm90b4QDgHWXqYhb/0ir7qkiPY3Xz8MvQ5O2OisuKFvk5KIeTsaXH2T
oOmEpgg2aHg17Hs46DjeaaqVoipv/0nFV0nxZ2VCRaUnLaHTFVSy8Eli+0gydTXGG2D6bVce6B1b
CiUfZcjtwSqOgO6xAxBWgSS+5a2SLVz+A/rEFVEWiRhXyLdFz6xDbnrYEWJnKT9NPoPcMWr2j9Ng
9UEjCSngSyfDsIKIAR/fLZqQ5GlvwT8bvL8MBVSTA3qG4SElof9xvUmTfuutDkTDultLSU7QzsNY
FCi23KK7eCKUolvV/ON8uoXlG3bOcC1rEURB1X6/cUAvDhc5BWoYuY6Hdpy2Kt9z/GAHMtVj7gMU
Qcuw4ARtewgp7EdN5t884VDgftLfbticfJ1m9hlIMGW9itnhIk8BnQSv6ez3oQH67sEcGmsq//Ue
f8cgMwwwhSW2EfPWqtcoCvxfsYjIO0bUfcWpVRTkLyZ2a5stfgS5dnF1GlketBiG1+pthxHhZrc+
oA3F4los6xwfRuMdDBqTxpfB23iZXIabrzdyDMbTLiOku7VDcuFB5NVJXBEYBGrNbDcyig7GTHcM
gjxlN/TMtswHtLrH5wW1Wjn9zOGifWPsXw/cgL9qqPWfXiqi5DAutk9majiFXt7Dvhqsj89zYNYg
5QSgU/imJ/M1/CLiQkI1BJYySmOuUkxWNdyCaUNJmH9yoTvGG/4QTa8Cv/pghDGC84Y5U7njxAOU
V7DPtdVu0xB4atDo+LAEJj55alZQIYsL59PXY3rxQE8v+ZTP+l6kI1KNTjopo1hKraFbi6xlakwD
JGVAIg26oogLvpOfx7oBvPkN/18krh9A5V3GrL+jbNkDL1hmmNjsCXOM7nA3kTr0YeEaWJawemzA
0RyhGtlRbI+lrnD+xNuWVV11Ye953vILFe8xZ8N4sAR3XSuQP4BO4EtwO6bm/9uzw0fEhECC40PQ
tKLhPBWN6uRWCWeGpeAz4RVO9bVvvPnnX53qQ+jHON7dwXlGjkR/INJk2HDVZJ3VCJNXxkorACSn
usNmQcjvY3voMWAlFFNxVmvoAxQyfrihfcTHf15CY2ScTfIvsMDdSq2JJ2eh6hJC4b5objTgiLxX
Gy736g54A4nkuCmj5VgpWF7XqkHoSLtNmv7O+uZd2PYV0T9iuTUjqNjoEWxxFKOF9nDyj5oA1Q/R
uPhRm81NU5wgQYF5Mk3qQLbgyv28mnWk/VYA/nowcco0/t06dzHgp1prjsDzicOnfr6cNgyIqPby
NavzD0jHIJ9a6y5QPoBtelZGv6ULp+7Xqun603snIkRdHJWussgpTZrp7+AMyvrzVI1laCkcP+Sa
/K7G5TvdGaZ+hlYTJQpjY6SL1ZqpIYA8gD7HJRtG4LikrF30wRou6zWB3orQZIvl2jpKtJxfnNKz
SQvUPTn0g5WS2a3C6RdIKDyVHgVfSnM7hYP7YCR5W6JV6hn36dYOFjrwmt0SmpLEfjIouSVUbJyD
FDW5uZymaRa6aofOWGZ7I0WgzXgs/8mfYBirqO1kC1zRKH9uQYZV6TApAQNYLi8B0SydrIAQFFir
4nFxTtwLFkSfk302tjhiKaOuW5G9xim3Rjl/GJLH+AkloIpa52ZhZVMuxPmJ4HeTbVpEPjgd30OQ
w16BW8h2ZZ+rciv1EPO7xNWfi3JmyEkeYFkJ5DSeu5q2xYPJXO+cc+ANoBNW8Uvy7VovL/gSTjmE
G3VwNOrGYFC89ki8HaKqt8s0Lj1i4MQmivFmqJd2TGz8INN6nJ616NE9otnt+AZFgxcMIpAerE5X
TeXQu8VM9fVu32UgKoLYnYrmqTCkE9/ON9a3/ZKuwMpDD+cdBXQ3DRRsQlBGpJZ1GC8Hsv65G3A4
QVDQhTi+PJ+J0yz4sLWVsR/1Kbp//Q9N62/5TUB9Do/Hn6yYqmIXiMHsTvIBxfCsgypuWp/iYs2r
0sQ3MFoYwYGCFMrpESKc55SUIPq2K7Mt0I80yM54Z1ffFHPXo2aEWpTRK6QdJ/0fS5cbHsuqSa5R
PIzHX78xxGWT+3hEjVqfrgBj0HTA1LvpFFfzKKnBkxp7S7D2NfhIVJ03RDCLlfF7Q9saPZxl5EjX
FdkxBx65jW7yxrDA+GkbECUqDAxt7Iz+l6miNkIpEeWUbJr45M6IW4LTCiKJBWiRPu7IaAW5sQ6m
RLOI4EWQ0u25YIu6P7k/Zwh2+R+yA59C8+a5brrT0SrUwPnag0EQZkXn0ZTfT8U4y9moAvsU0gKb
zi598lhqINtu8CqtYpShUD2aCK49qC62q51hUTsbj94dTM4Ld1P5kjUiSk08Cbae7VgwOKn3eXBG
XOvnEWZ+EbULj3tfFTHnlX3c8JOCKrjqz7Ptti7HlxIuijFW5j9DvpClv/j3RukwY6ycXTn5MWKH
8mG5WVfkuf0Gpu+ajksgh4qLxCvrdlD7OVxTnKcas3SHXeXqRC99STYsNJQDosbKVxHTrgkdvySD
eNsxEUkFKjMQBRDSIYa+uBubHeBPhswiDZaLqRBREFBS5Fqy+sndMpyVDU0MwKQOot3EA+ViriZe
go9z4KewUT75s9S+CPV5eXeBqO3D8hAYCD0VLDpq5tWzPfSWb9bc09BKwtVN/YL1JOsrmaSYsLF+
l3xHj+aFhfyXeTP7XKaqALRs95rIegYs+yLhiVSnGeq5S8uO61bo4vpRpkUcWLdS2iE+Hre4OdSA
EtVU5iPzOrfOuRtuYIfz3ZmW7vkAnpwUS7wxV7IFvMIEa5Hod5N92kg/EnjIIorhJUqRPqb4TDB8
5DaZMEpH1g1yqVuOW+RXxylG6Z9bOLfgNCDg1isiHmiFT7OnuVCCIfv+QJ2FahsT7mA144Kz5hNJ
7T0KPQTL6+2Z02aNuxoMODc7V/ZfR4r2RXUsuGk+EkuiRQFto8MHHUURTqhqRYc+DYk2ZGhvPjth
J7+S8CSFBZbeEXT4A3u8N0FoHu57478Sa4YosSX3DdHl+UiET1Ut8dmOd4HmQiNRfzJOw+iKQmRu
o6OHglF49WfxQ1cUmVoABX0vFKPnyCT2HblFurVApIqnvvyX4x2TcHCZ/CsDT3r/rbMwy9wcDHYL
NRDSilQ22LCMIoaVbXW9ESub/Id+0zN0+9lnlGa7S0nl6bKHKxqsaWX+HW/gqot1qgKic2YMXF7I
GNjucympvlESU/JxT2u4iXSMkhnwHY+2bjqhezOu49JHAuaudlysxDTTyWo3ZGznSfRIvob2D0Nd
W6SnfOqlF5QIvK3ylPMF90QghROBrqrgpSi9th1N8o6qb05NG3/eGX2rcZiDL4NqTIthKM7ISUVE
l9GG7q55vOlVnlP9uv824a6oxGKEXVeuFxnJn08MalfMvrBYHPBsAczVQa94BZKZWry3KjZAuK5E
IKC8uCxaPDi/63Auzp2MJS9i3Il/8uHPZIGMHviFrSxPqZWbJxX4Bo389ncHV4TW2dMImxJSda02
LICFXI3FT1DSHH7bxmk8UUTqld5Z93PrQawpL+xFJuZMo9s3anE8vHcAbCbe3kOVIFskNEX4G7Ci
nIz3WiPhc+sXgC3ThbP1ujfnYu5UQjVOLwR0CH+z74/QE3Hov1TqG4Ngo49VnTzmOQozIa2UjFCM
Z60mZzxZDnRfPDsIJkjMowVW0N8gLStXZmwwqgWslZSnXTCkx3u3euM0re1VFaYkT8pq4p7HO3+6
s5UXfmxz21oT2DOMNvs2/Ad2K4deSKpvoCuUD3ehg61qHMV1UZrsT0OexrPkji/wXoFIWvdzC1uJ
I3mSIiolynbTXhX6V15yVLGaF4U+Mm3xWsCeCyvLwrwrQDoH2GuxfQrUcWmpGK9QTsCCikoidpst
cvM7rG8wyAfDtQUR9j4CYsAW2gQblUlXbiyVDiHSaLcMwO/+jzfjVWopPq2JAtWR8/W5y5n/Ftx4
yJ2CxR5aypXkD8bVhedXBlg2u+mki94yvVjk5eXP2fC0/AjBGuFMMPcW4R34C3ggOQgESr524CpY
kkeDO1EpRfNJDhBaKK8gTJlYmScAncauYdOxDkypg40gAXVzPPBS1TyTD6xbzZcPv5KPQlpQdsgl
WKh+U3NrQl6oYArLCCrBITksshBtWN8sKIytg+lbSSRSEVPfZ6PEVaqB6e9RpM2kOwytkpHx/Rnn
Np8waZ4fUA6j9wpV9QrLBxG7lAziXEh1sh3Gsa7e5oL5Uf7tarNGIif3gK0EchQ2wZJGWfyNJusX
HPbq6D5r3KwjsKxr9P4bkG+OBTZWU4JxIgdu+kEclFKgWJUG2CKgHx6dfUz1MT6r0gx09sS0/uSK
Ikj3nnuGOdMneMVrU3U/4eQJ/8x6Pg4lmPdV3+e/KEl+8VPzcRv+oiqiUZhVIzBgtxhnI3zLxpCk
cv2OtZfvFQ/vdcv7A6kxu1CYMLhYWgeOpAM/DOYC0BJMkzkr6Iw3LOtdpVk6xUucIc2Qi5sIhHQO
xx9PqdOzDVrG0qI0YJ7quvhRw3vw3i/CusZ7JdW9AaCopgJoq+ahBE/3YTqeVVUJNh8hEsPZES5n
CE/V351W4iks+mfZb+y6+7WuMJciXIbv3YjPNeaSzsrZBXe/nvPFpQQuJfEXUywCKlmkZ88A3Kus
Na1GMoIZtZHPERD7PpUrBgbRzSwOdFghSCF/9FhBmtYQmN1rzjVLfpv1b8hXC/l8C38wIvMcerL9
w2JoztYgy/OnmvG3FjP2HHwc0V5VVj06f4j0aBji6ieUM3yB0kEmn1F9P1nWOChW9YWbODjckkni
2m6Z6baDn0wxghsUnVeiHT1VAcYGG8m3569KoImfIPUVAsFha3W7V4Wcq1JEny0+qzO+gtksY7MX
wQwBDudjCk2Ou9v9rv4aK74HZSLsXn4G4nkR5Rfey1dNsAX+HObAafApxc+2MvyuQo4LkQIkJwPA
Jdm1NarT6c9ZK61qu7nYJvCxnSE9ovJ5i73fcXgTSuuy4fz1YeHfHQBCnb7IzQET5HlwaI9v8dYp
V4pUPP8BnPYGs0oKZx+xAAHIFtgYsHj6kGLyM1yiev5SnoK+9NENIDS1/y/cc+gl2Q1fgbGBFrkG
pp1aznUJiJSu1syMqjcObrIT7FoTA27zf7ZtLKMWJDJZD1sXjgZSN8xKaDJzIV+8QO3W5b/VBRwz
V+XJ8HMmpv+jySKu2tZ4+cn95btrffnciLnvHT2YrNeONEJABRvMCIAuKjC1Nc1NYDlxi4HVeruZ
crgPwtjwXwvsVqIRTnoBf8sJdz2uyh92/xwD3fldG5Y3DKgcx9iqq/cjVixUYrgh+cG/wMtu5z00
6DdxxA6WNtzfZC1ndjJDOmotR4cQmQoLV9saY4Uf4U42O6BBcASfr+21Mow/ykD5B8BpBT8vB2Sd
csXQHMZqHKrrgeqfeOu6NPNkw5XoPkmSHrj+CddXvZa0ZoQis1LfkPmAyDtfCsHHiQUAOTTJeUjK
fZf/stkv/cCpva9r0HkwhMneZgxcwh4+/hLICRQtbj1k05Zm941Ogo0ZEOXjwYPV0giZC8tuMp+C
iSM/W42C9dh6Ep0A+JmRKggg1/UeKivHppmEL2ky7HwowiN0PMzWNdzGQnUX3uiwwaBbR2oOSak5
H9hSFRRoEvAhKIeeIXUsjz88f7dcIo9hmSfbdDuvZyBP0v5mRVcb11jn5fprjkNSBy4XVO/NUnfQ
IJniaypvVChCGZ330V/SQKga73BYyf378GKZ8Hse663VeZtOEtub/PxKOKO95JE+eE0azictbDsG
IftM5gz8vr61/+oloVgxvntPx6NP+NIoIiVzWfxM+E0DEZP60WyIxrh8vsG3ggl1nhLyLPAT94Z5
Pd+iKov8+3TlQEVDZpGcz0dJ6bTd4Bki+Kj+TkChjxCXjFuOnuOQNQcFiE9uZuybE+H0/8nPfr7T
6dmANlG3WuhPZLtymwCsgP209XoU2Tw1xjdXnmx0H7kgNBkYlX8VLJkwX+wMleMXpWeQKDEChnwo
4OF2w8WQJv34NYms/9szGKV5bLrt/0Hj8KmGXGMOHxNsmqB0eEEgqmzhDW4bTeaq+jc+Bv0ERQym
aawaHkyaU7oQ3jAoLB4oltc9CRagzJi/dJRQWXwtbCbzZt94A3n/9rk/z2RvJeJW0qvuEVlOK2MX
U3hXngvNhIatdAjOmqoT2OYln89WD+5lIINQLEhMo8NPSXGh7ZCBZpxSVbK2oan5WRT2wq4VD7r8
hUwELsUX+GBc55dns9eMHuGiyjAXzyEnAopx6UvF1m50yL2998nmmNBh735I97tSWvUkPEogO3pP
O85DxiwquZdbcmGnba6xTjFLZQafVX72xnK5EJiVIrFUaSw1xMnFIElwd2X2ns2Dt2CF3RS7Y47k
8+HjA/WpioHeaM6ahKdGE+Xlwe0M7EIphah+LRqorEMPdNNdV59JZ/Bk8jlgjSL27Q5/PcnG8gAd
D8TAPHgntT6mSuqOqt7rwxWPOaoG2eqxszdSsoqtwhOlJrlzmR5SwMaF+PSV+WUq0So5Dzv6YCsD
FNMsRpABalvLWotlYaHj8ynW4gGeLB6Oo6Rw13vi5DHrEIeX3KdQFlHxwZERIspOcviRBebdVk7Q
18pr5hvF/4M5qlmS1/6eYtWtHF38vWz9DmnWu8SvIhg01IHk0pcWjNCHQebLYCzWN9L/LYP3B36w
qLBg8PA7FWZ5XWd3XN6xi52GZefHF+Zo4FKXK3A0yLZyLzoV4B33oXrtRbOfy6sfR3KH56+zvdNU
OLQc/q03gdKsOYV60WLqQTAKWGJh3gi8eQZn9WqsWmZ8GNMC3DzSXO5pbxJWjz0a71nofQrxpe+m
WItk9z8SCrPSlgvitDR9HNuHiHMm/O/kI53Ou8OCsH1soLGhwKTvXGpLzDeOI3tOBHTwl0NUB++9
tCCj1fKGZew3QKltewHUtWklUwiesocZ7QGmox9mjv9zaZFL2DUXyl+BQtUcA3cBxWmgqqPqczpg
TIRV2eCZknx0MgQHabfRSdL6dfDeE1snDZEuuIYZdu4uZhaK8fnsPjVe6UHvnT5Uk0rqW6pPgxo7
L47jjA2JZ7qShaHWuAPPtAuf/AhhG6dxsY0/SNl/sPOE9aQsSGdb6uTja4bsNdAn1mMuMkBQqIdQ
/V6GVkumdYkktPywNNBRoMFDAdc8DZsLV8JODlzckl5MF3urjx2KMxKmknLIQP4b/zhUn3OLc6Pm
oyZJDmW4ki2yyQAWiBVgJnXaGskkraj3BrWUPepencPzh8AjVUOAzNEVd67UFsFQ6pg5tPHDilR0
2BET3KcEJBohdI+8afTyUr8RbZuiZMXVWsxArPMbOeq+AzV83LaA07btxWkGXVuWtqANYwb5lvV8
43pXvYFLBl/DzVzRA8rOerWuvDy4dvkOTXDLmr1PPWArmyCnVhS521O5h7TeFn/TIdHRxbN8mUYt
tS8mHgyJiCCnQnJuK3dic6wTbajyOup1oyPP/nKtNmcplukRsLJKaySyr4enxt4TUQZyJTHFqalO
TGOi/FlHdhwpmmn2Mu1gc5USW/qJzI4LWAvlfgt3HlxO0F1cTAHc23qUzT78x0yT4x4a5dL4/0V/
0yJs5z6zb+Zd+tfr2+AmLOJpV3PPiPCYJKocKhy7y4CMCzXZ3n5Ak+FpnsJq25s4KZnjk+b4iqUr
R2R2XJWkSw9rexvswVwlUO5Wi8upWSHlUqgk0aleKKj5xMDaOZLWhFtEu1/UbSAxGQCm97SYPMCU
NqbpmL/3kXPfi5q/yov17MFOzopKYOnlsaMUe3B/LPIfsuBicd3g6fcCH9j/a2Smr+5EuGqAEVBU
9J3BijlcWHjLsNiyEE2r0peQrElmu9ISimzxBsvDMSQZgND5IboN8VCVpJI5TJnwkS6km/OM0IQR
CesIeUqu41nu5LBxFZkZobpktBPDmO7zf31jDEwrZwcxF6fIKTat7VpydNT6lYl9O4UnewxCiY2f
ebhFazvhVmIZa2StwqX+1y43T2jVoV3CIXmlPdu6pkXAWWZvJI5Tl2cNSum/ZUkwCmjJ6O0u8PNE
e3smevx0RV6oNitlg4PFuqgroxdGuBNiDaLp6rrHpCSuRxQjE8q14pLM+qeKOn4O86BpiKmF4GUP
Wxm+gjMbN2YBPz8iY56VCiHSyevrJLBTLpk6gTWCKULdOb73rnGIUinPr6zya2YUxscGZVeKxkUu
lxUwHBnD6c4m4axvsM+O+eQGOq/AnfcxjZ0100y449L6iAAJcPIcuJezOs/RRV0yDVXDtbYgszUx
Mgx/KSWsAINqZOGzSUEYtgp7nQ1jx/40Zkj+Vy1KuWqmAcFIUwmJHbUjjB00DPndnd+4dRx3PCHH
lbzpdbEMYep37spSdzGSzRdismZNN/pxG/H+B2CBdjMdQ7HxTdC9MO2qLQSX8/QZX6MIIl+HQT/3
lo3HlrTzQlvLlK9O4Da+WEDSU9NSoA+Bxw+uhOt/3flktPwIfUl+2UYdNCcvgIyueUwmHHp+mrWZ
oMe/ZPq+aMPqjXgMXutP/nVD55NMD0stTWmP5voge3EkonlvxOKPb0nMpue7SxAcBTxXQN9Y6UUy
PR3LLDYCQmYOmi9bAGlKN9f2fn2wpCd82ivcHUuYzdq2Vaw3YWvDYj21Ian6H0uZ0jKmRIv9D/OB
j/yCu3+vgd5NJFucclzSxQyANUji5hGRDj4mCwVvrZR4reTm2bcA6s2KEw4ZsveOLAQejyl5xzt7
QD8DsRFq1AJDmQ03HPIwULf+fRTQ3uP0KbLAgHAUlxIXLxOoBEWyv2d2WUHefyzM8rZZFQev+2VD
w42Emde/ZAklALCRU/2/p80n2RHyDspeiMqwB3Yt5lOMrANdvkwClsUg5BfVnvYcaILw9wV2Vhrz
CQvkdTfamc21scvBTet51gBTKZMtgbY/31WjqyVqbZR4+9tdp3p+7jbwT5mWmwO1Yb0Pkw89vvgt
MTraKQIZlbeY7bAAVFiizYmbMYaSuZD/IzpVKNiuuFnlhcmsoD8wc+I4YBhuFLsqKKD5Wnf1kecA
JUhoRY03QIZVRh4PlTc8L3v9k0j9SMxZ3mxe5oVUDJPeNxoGx1oe7ym0DSQLStJnPffdOkFFwXEh
mj70RVNfNB0Dr633zchRcMa5/24MQZz4rwB1/9yxf2lrHmGmAmKUg3mb6CCw45gxG41etb4XmKCg
hoJ8j4zm57KGU8TonEWIvCAtOAT7J+YbJJsCVItmaqA3aR/+9qcOxgA+4VOlO0Ck/QY/jxaD87J9
xMRh7oE4l9FJq8q24RuCKcQRPJ+XL/YTjbMdlkqeY2qfEJ+Z2GcAlEQ65Y8DltxZYEIEvWbXZEZy
+D0lVywCWLDZxr1+EaZATxDaKO7sBTyYmtiBKU1yz12Vq7a6tI+ad2vyRF0pd0rmg5UQjxVgyGV8
aJyI+y2MG74r1Ucwkb09xSkOUQ1Q8ypo7OOXdbtXDL5MFOr6X0c/HPBY4QwBZKXR1kaO7lUQeNXu
XUIp9ew7d+FkT0t4a8ANPg3lJfOCBGpqNzp4AyKnYSm1wpIj3dpKuyW/6WF/pbDQ7FFSwIs7UU9t
r41Ed4+KY5c1/SxoEXxEebAK+xv8+iWXlDoVj+oPu0PC51K7RxATYPw+IgC0Hzxb17otS/yDXZ5D
pibh09gUN+FIj6B1VoGA4PLljAzide1TQGflv2bzu1zBg6YxSCd19ddPeoI1X6GQ4SdryIWpGIk5
hkOEfbp/rlxQVPuheJuSSUeFPVrcIwVURLhZRCDPY8d/pb+64N1oMjrCvHdefQLS9/kfWjbuBWtW
a4o4FEa3x2Tyl7QnPY23YE1BMzdz4ubTC9gGFNKaJ3098fZULYJgGrlDTWC66Wr9m/UwpXlINEZc
gb1+jDp8VDEUnpK6KwKAAF06HxXaGEca2HedMjmZKevCh/a4I19u88Bkbee/kuFQVKOGgDOAfUUM
F3ZMyB4uVW9ja9HSQHM7MrSMoGJMfr5hlacEcxvuCwhvPA94coeJtomVn3fh9gQOjz6oX02uXb+O
Vc4CKDXeKcCkwtTrqmzf0q91oDJ6iI4ozyHQDDTgGIckUKFsL00wXIpM6E0FYO35x9PBmPIJ6jag
kxjaLt7GlU3wkLyO706abq/SRpo77v2DDEucTKpU2K0c5fIUNOwuCkT8lvMpvBjmTdGURX88np2j
Jve54JsagjkhTQ6D+x4qxm4HXxEckDkGGlKRu/bSj0ud8HYkt+uzO7qaU4DFDceov5tATT38//mK
zAIOxjjUZgSu+Bp5YEcRRJsthv+t68R9sqVGb57KPiCXCD7R0SChUVtWi7T+qaLS34s50t519xmX
FnNlPOvfxN+p/wUlenbt8gYz1211Kw6YACEeHFlUoXy+D5ueDgVKfujiL00DF61Q3L9s/XnDqydm
oFqw9b/A013+oBRa/spC6NacKQsEmRyDKFHRHesPAOptYG0vkpZE5W0pUi5F/8U88sel2gVk+Pds
j5PL8cAB9g6vZCDxzg0UZyqRyLGinMP2ln+Rw6ipqWKN0YcDAPXtJf39Bj/igbbY5T58/8Qe/u9N
zgazx/caI0FqYkwC2WNAx4/s4ARi6nVoSmcFK+p9TK/Dk9ryEpp1tnnM6y/3PBpjW4gKkw+3BvUx
pgg7Zcke0scZ3ymyqnTuQRrXM05+srpNh4MLNY2uH0vqsBfTgDV7a2nmzSKyVCaT1eMcoyHzj6Uk
02VYFrtaj3xCNC+0mXQghfv1dpIKrZETFNuDT6y/p9zc54vweLo8dAteeLjHWVEryB8oJkuBeYLz
OTaOP16yFM96rje+DMz2V+UceGn6u0u+mKLxfjRcrzChMoB+GRp9sQWazb5aKuzBbUgfzC1DEAFT
X6nEUc/1qye3tBsJbj79U3QpOVzht8cA+VxepuBkPp3vvvkiQtufZvY31aioMNX9llXIkvmsyAJ8
Db5+xKUdaNN2ePJiZqPgiwjuuDxY3Acnjlm6aUm9A1jNKUBLz0H/qmJqpF9G3CbftXcvRmdt8fVq
V7TmK8eteRiffigjpXrTA2KeJZniELDxxa+5Hnwk04yHr+0jKLO7//H1FhDEb6ySwv3THDUchSQ9
2Mek96jPWmVJhrys5RVq6sBinisOFuTGPAcZ6ZsKpEDPfOnNpzxult8/SarkEf5HPNy5M2aMEXw+
Pii6wWsmqtrwu2MTyFw5glCetrr8t+8zk2tat7OQ7Pj/fMVQCIJh0husmwkSh25c280ZDmqb4ZBT
SsrcLjk7SwMk4yqYfmEBla8nuxVthlzfhA7bKHMZWNCV/j9k4cABdx0LBkzz47wWyrfhuGKJ0N1v
E6UGykpHInd2NRtT879FaEhEWks62VlAV6hjSpvehQTAilUzLXbkCjWoifFxSUdKgTnQxdx453IN
uFVL/9hqBPUq6uaIV0ByFAw9fHOA2FrsCcVdipUrkF5lCzQk0iF4i6I+BrVAnnORf2R7P1pYtfnF
coORqfdt/K2hhtep+o+xq5xNeyLPKPGLWGTl3LN1nq8WQ005eNq/tSrZwHUm4q8BHEgyKWQKCdpG
9BnCrTgslt++W+/k4ywbFrdBs+WpuHEH2GxAnNBHzj9iY7nGn+NvYkrLCxrdAioWZzfLV6kj7IZn
BQ8zUSZctaxA3LdEy4SNVl7eqxznZL/nIuwAozQX7WQXKtr1Z8NbPZpsIuFUEbAxeA+DfoyR0STo
pJo9npsjimkfPWo2kHZzEyC52L8z69AjEuq/uqM2cS4bCrr2xf9ovtMEsoC/qb7cg7QaKsIGt4bD
qBClx+PosbtzmGcBGwfbDw+iUHa0MRxnNoPg/KvLMj/aQQUiE/Mi6EWNBHyp+zigJwvxeFU9yZKg
9lPv2DCBbuabJe7SIuxO1k/dOCnBkR6NCBJBimOsf1ICagVZtsoyGgWkXDiwceiKZWu0BbUbKh1a
lzswpAYmMM6hWJJ5nM0PuQJ4nvhgyFx5XwnKAk73779gNrAN+MGcdO97iEnc0c9CaU5oVIrPi8s6
Kg6nkGkh8oXYhbtE2q4DHelbUxXz2n1CBP76GyhBgIJNYaSbV7ien5nupQZGB4N7cW+obdjyzR+M
0S4qj/hXQU1bH8pJQJuRIJNo8RXLNKJCzxnH5zpfGzjjL+PBvClSxYk/M+S+CF6DWYfSPZBQLQe/
JOnk6rBB1G/mSGra5K+Dj/hJnWxKQl4lYgos7OZZTtszfaMbgaS/LGIym0IiKBpcIQNYUItIjZJF
FKwdY4fvX33wDC7QTOY6StVbD8cEwno20CUeV4JWNFtyGX9+bOJDAyB9UwUzySu5lfeMfbGb+RHP
Wcny7GBEqwiFrOZ2IovJdpxJnOci1OvdKtnR8XQj5x7rMJWzZmwePwNeAkqKNj46UYd+YtvIz6jG
irgoObsyHFzt/WKdjbilSPadslEBJsPaZW9NVkTouaoimKJz8siIgkY0PJLOXVDA5QqzJHga8rJD
qmHSpXbyU11H55BvUTkhQTjV/Vv7r41JhAEkAp5dUf37PaK+SEEi1OGl4XlHqytljsfEyTIV3NxP
Qen0ww0E1vvFsrlZvUrKFsRuede7jA3qQz548JuOnZcZ27fomFjr53lxlEDFOEQ8nkWjFFkh8zV0
GfKxx6Hzf03PHxUdQanbD14K/Bhct5CLUS0Q0bLVhK9p1eWwjOQKHeZ//EImDuwOpSCcssqazKgX
abMnXAiJVrzxEnYwB4P4Q8pBBWju9HlMi53sdgI+yxeKahW5xCT1ZCbpi3jcwcz9tBEeIUxnDam3
GsgBX8fJdLoQVfXxbHnJA1uiaMxidm3CB1RtWsXCcCxwLzRlFPABbBOIDFDhFpjgF2YLEJZVcMDF
YXt+CfyqXw+YKBWjy3jhTgS5DBVBGo4ZRI+gm7jlh5f7UDLDwh00QW/FRYIAuYdj2jISnl/ltoqr
VpZw0MHPlPjhZW8ZLiNleQ7mAchI/3B3p4ztZrndlTxPbKrE0TQJSRQaMGRW4EcXSKVzQyyMMubO
Ey3lLBuNOfJ2gSjVdv+r+mxIHXWiECUdyFgbQK8SuMghZZ79HUz3ZLFequ+q9UO0kj8Bj8zDSZ8Y
lQz5SZorZWzL6zzXMU+lquc+tWBPP0TjRAPbgn9bhpw4u90Y55BKwTbigLHhj8hvdcLCfGB/O1eh
m/E4IO4a2c898tLaKw+KfpLUFyDaDcx3xpYKDPVg1si+QE7BiUki3p2quv3WE304Phmxq6iqqNSI
6l3mO62z0/DDJ2Yr/gtTzzcw8RQqwR1Jb57U2gsrHdvFDtCux8IG4dCmnLb4kCaXaHw0X43sVU8l
lS1MKTGgRNDk/QjHr3D7rkHws1gXZiKz1NU2PmaXJwMqVYnMfJTLyeES9x9h8dv+3Pjhh/+3BQZI
zdlKkvowf5gjYHCa7GFXFW6fXSkEky6Ift0l1Vr5gAChxh9eIRyRVJqJGIw8lKDOK3D6bgLEPauR
d+sqH3+4SYDoW4+bPC5jzs9OY5lXNHPZxWA7BQg/cueddUszgnOrS40hvfayYYF2W0yYOYcWcTq/
oG990DFmKx2Z91PXEsKaG1cLMwQPyU6T39ufLGYlpNIyQWZT+PgSa1zbdsYR6f5D0ye1kjbWGB1i
cJSCyujumba8HvhTPnQP+i5CpF6Ev71Y9PYvU3yO3YBVoVa4y2VrHqb1Hy+z4X9RfgKCDUman4S9
UjN5igTRqRuDYkBxiw5VJDkIZkUDaNaQothVuIpgmXr898974o+X1ZSsxgwrtB/pqblciKUGb1sC
sIjF/XJdc/Yb0wod3D21XjkfwbRSn6tLcBsfEvKjh7TqL41uRr+oOIWFFghdtPWWEOe/57pxFogU
vjran2mzYFUejL3eIRsbSQHXiT4+le9Z80gZ4cy9CN2KkyoO+g6C95TkEsfxTrUvI6PR52zfrIbc
6z0uBFNFjMIwxZAEEpxmJCRUfGnXtKErUX9oz1dkYE9v4MhSbPCYJ/20q/vr6XP0nkigsh6iGatD
/1YrEA/ZeKyDJnr0ovGrrc1MlJLARqvtXHcL7aDJI5mC98Xoy9T+XPYoAWoFsBScIH3j9hgx7EPB
OpiKqfac7mx+wajg+KssmF/2u4BX5XLSEFD6B5aAp0bJbdz9eH06uaxVvN0iBbU3VIC7DDlCsvm8
NvAe/2z31YJ1Cm0iozN6sFKVBWxd95LBNdae+FjIjxLfjmrLW3CWHDSxEnO8BQ8LUQ2WemhZniLu
2oW2/RgzQHbGDygliYQYrpkquo+SVMtuLEK4JZ4dhlryJYWvfOCl/w/WetLc5Tof6J9GtbCXThcD
fjciUJ5zm45u9oieJMdHbr1ySyQITkEjKZ3ihz8UqgU4cwg4IbhwwJibZNh17kS86eTJq5naqHr0
aiFqdbJ1BYUP1hfOQvCuHS+pcDoAljXT+sXSTmZCk816ajzHECmNyQgMvZX5T5Rxj/Kr6B6IRi4D
vyNq6BDdYcyEsbYGg52YY4JmpTAMoBgknz0ep5nSmOUqghWeFG09i1v2JVnEZdNyWGHH0gec8YK/
MKn4oXaAmphN9h0zFIsGAuSOBhE0KkpWztCIF/N3FkJgjbfjg1vlhDTnkA5V8Y4qvVs/x61q5Twe
f4Ilcv5TeBlR4BuzrF0NiXsGh+nC8uLWhVPJ7imy1RZ2N43pmyo1eJG7Dm5tD68BbKn9fuh81dAD
/vclLgHh9jVtQDG4tH0EP4S2Q+4JPrV0sJcQwOCP+XM68CyM66czUH2fUAoU6tmV8fBhy3vpjrs4
EmTOgzX9bv60+/dBNpyzMdsWtQ/oJvmZB0VDq0HppLTIDnzQXvpyqHm4h9/nVK7ziFCKV1YjwsCw
XB3flUWjiTZEUAbLMk4KVVEaxVrMIf3Qi/o8K6+WrA46qQfnqwSohpRJ0pJODu8l/3zc21nTkcjq
DjwlwywRMN0kUErPcYtYhqoA2a3a55UFPgU9eruLN+lJKdzKzbqY9AICKZrEN6QqkTBK7sdv3H93
d3t0FujD0zycDUEOkQvuym+rJeVsyCEGdXVVjnU5cHSqkXvHXiYDhnfmJ9oQPvzb58LCZb5WvbPi
hsCo5i/uFDJubLPj+YMkiyDTlm4W0ax1su4tw0hN+KFPMk7pVhP2yJLjT4jIee13+cu3Sh7+2d7m
ffnyvg4sejHL6XaK8IIm+K/8nuLKRvS1qI45pAqZnNLFKQhRaTjNZkZMATh49bki1NbVh3/E5kYh
hS6r0cA30KcqWFE887y4qk2sSD1Vt6POTiczk0cfWWCl0KIYNj8sJBzSsLkiYNGiNXdaz+ppqgjU
Z5qKDdusVK2inYpp6DOxcgOTJBovjSDr1NkAFZHdNa5mGoWtwGjuI64aWqGCo21UQSyPf4qPfpr0
Ueun9EqhppzMqww1RPwTWKAmI+iNFrUP1pBnbDxyuPtHFabAVq434u9h5ErVH/N7JhZ4NBG3XJ4R
DaTS4O7TOmnOD2RONxFIMc0W6pBGDfstpjMxP7VG3nDx1CdbkdN4foEuTTXgsTRWY1YVFB4JB4e6
bSqcugO4JEfyGs0Nf7B2WZK7mJnwhwBLjcM0F8KA8zQteoyZtz2DH8qfP9Kb2xp8dU48gSfr/0FC
grKIy3xHUNv4vtZzPXYzPUQ0kciq6l3p5+zLIaZH/HUzaddhYFvKVGyH1mu2uhPnctAiAVp30IAH
9D7Emh31EW5V7drTWe2hu98pt347/s30JRMmA9nVUtyqCYr2nYVEoLUDSIhlqot4Hu+z5Rh5EUII
L6CQGYo5Hh3JTRGptJQUA+E7wVEouJMmTZz2G0LeDjM2ym0SiEAaiQqgBrkxgn57OJvBzsRtMsB1
6geun7PnLkS1g6ChgDh2L6HsGMacUaIYPPSthw3GpmEZfxhrLeYdFUq8g+oyo0FrjmV87BZLU8fO
iPV303BW5CyVuL9R5G0qIyRYQ9PKHfhqnt+46WYFJJ+u4beGzMFG+AyJf1lYW+cDFgRLIhzfP/SB
fNEFwpsQc4aDXZ6BT9EIbwySgluj6EHxWpmj0XLFM9x9d5C2hSgaL4g3gcUMZ0V+u13jQMQZ8+pD
nfwPGLQhWnQfulVY2nqpdRtsDz/TaYBhC9rDBX6E0znTDx8lzadIwT1yxwc3B4oW65kMUgSttZny
KF4ND2tqwJEkwTfNDmcHscf61Bc7NQ0ysm7zZ9peDm1lrHVtBP89K3P7i56HXkUduMaAqQ0q1LGL
zXeqkl7dbBiGciEIm9yrU/2hk/2BQX0XO3lSkZ0R5fKB40yDLbzLxycXGDmg7lkGxmYDYrl+MOZT
MGWPydSVHfctCU0JbCKbZ9ap/AHkUTJ+Co7W6X3uESZ3UNCxGK/vbirDscU3XNbW1UbZKDHX4sI9
CqugWa44UZtRwOSsJVqyw6t9LjFznZZoECLI5sXjtZXaws3naE/mvkrFCAqECRCGNlRTnsp4BIot
mdHK61wPbvE0pJuiQ1M2+2fXixb18PV/YPrig7uzYu8o6dVWR1s38Mpu7xxw8cwfKAOfFk3dSwE0
O3C7ztlhTo5pF5AxfEWybFsA0lutQ+5K9CIONJneoT24AbohyDuGadY1pc192A5HzPC7ls8zIZ5G
5dJ3WuhkqnIOXBvQz9z/ur9cjyQnMnVHBJVjaYszGyBdRuOBPmRTg3ZNJNZ31dH9EDgZFgpglfY5
iWS5JFwOMNa8SAbKxrMWY7WH2hoESijIH9WXumYFnhSwrdBj6gGRcMJ93LWT1sm1lmwwuLu6fXTZ
wJPW545aW+jDHlj0u/3lQa9hBFa8EbaTgqkz9yI3JrgZtE81wD0G016HccQLoYhfrxeDvKuHbPuZ
vyJer+D93Uuu1h9SbQ2z2fqzYlqMxNo08BW4w9ffuydcg/f5l+q5JoeKPap2qzJQNnXE+v0IMq6r
WuFFiCEQBsLbF3GFg47lFt/m4lcuBlFxyT8p3FPjl+8gY4kyfefvCbQDRnXzd3nI10BKrLypNoru
7TivQvMeD/OnYKQI1HbJfxfjuEGUQIIN41nhpluGL3VFSt6hsUz8Tb3+OKHlGbUjSpjxM7h3sVTY
VuKmXu4kJ8a41XDJFf2ByIEAFMmxdkL+GgIQvrF70rA3cLMtWbnvMV4JybIZz6jfnL1GoXa91Jla
yir01uTx8mepHsyQ/njoMfVw65f2X++fJjkDoEIK5pzreoyCGD060ufn3vfZXx1F801Zh7ujeXrI
KnFcjn3E2JERuHBqK9QmLcdK7IoS3Fe6AoRQB76ZoogjtC/2EqckxmUPp3pCLO+lZtiqoP92kLdL
UpaJBnOkxC4gxfnkrf582VZp2MUkbQ5LJM+nW9yhqBN0tONrirxSzMSroDbOEnrxlzqHGu/IRZpV
Gc6L5AbTKX4bZszmlYv9kCINnH0ppdP9lzai8X8GkNnglruSrAxtGlH5Y0eHE8+0jEU+xO0zaNXH
qQLRilqrDc6gGObl/7A2s6Py/cQDLiRIJTPyWeI3EpfNtlWtnflKmzHG57XZil/2oKnjKoSwTn8K
dmvO7BX+jNYwStvGVyolhEQhTyqF2NxD0E0ou8X4xYednYJFp57XARxN3VW6n2xrw+Kfb6Q8bo+Y
PQImdhzkwXoYHVyDyevG9OyFRYHEtxJyE6LoQKcSjAn59JUEXwps4kj9ougeeFWrXZJYtDy7KQ5y
2Sy5pi3/seeNibDz9OgdiRTVfHeOg3f6wk9UfnWkgkSmVF/EGdmdwyyDwoFABEfj+BRXXHbZ8kys
QsDgs+TckcmrIL5BfjtPjXjA/Np4XiiXVqxJjO/OfYVhjV+eiEnC6QT39ElQbPJ352rgM10TMPME
GHu7ZySFbEU0cyGPwAbTt/l0CMq4yadU+XoMyE/l/vTILHFG4Rg4g7nOtTnSpYIsb2CkOeeqJ+kz
jN64d6FwnC6/A40uO9wpGcl9KbRULAIDBGFa2nUNY0zSlaPwiiVIx9wXPBk11eqcXOLbY/kv7T8/
qYlZjtpqPZzC54dbxTOXBsfu+E53Sw6JUPdd8VKeTakMfgR3RExCXPTN4Yhy9nFEcnaT2+y4b3jF
Wa+ECwWNYux/djXCA+kkVv9DWZa/u4Q9lVqjR3a9uiRbGuFg9PWklXkYClo4RALruP/67EIyeb1z
CSzdXwxO8Cv0MUUxLmfF0g2uI1Brp0/7ydMyy95GDAPpT4m//nzfXal9uRb84cMmfC/4jueSucev
rb7mWg/PCY7+BnvwsY9JIp/qdw6wiGaYHGaSVqQf/nd6z5o4Uz9DNpl1g/5OYRttLfnOOWkOTZQQ
s8govqv/83RgQ+pEWKm6PkV4NCeLKKvasStXZTUYJlx53OnQMiEZaIT8tg79KOLErCQ6PgFvmaYu
If/rwYyMqmkQvnd8HZ6isGk366ZjnWHDrzEmyFbq7GTyoRt9y9seMbOnjV8cbLr9U7mUlNdEmmKb
lkCiQ/IvexhmmKAaOrgYn+WBrWq35q0T4rLxP1Kl8hE1JBymuLDRJve+vNEWBHB+EEsmlcPgWaaZ
k5nDYKwVDR4YVagiearEx2D23cCRSYBp+TtWYRE1TwQQuWZIYFyBDertSFU1BfVugas7RGhepU1V
DSh5u0RIxyeT57Rg7OpLaTnI4WoujtYxVqOoBNC23nFn4xjHWxml2iLd+fm+UGCjHQxpDRFIj1TF
mZshKqci8eiP/iPXB0xHs/GXQ0XVPqBc8QHKZ8eGzvu531Mffw6qRK5rzvDq7uEqDcvPlB0iffCK
WenMr6btjpyk+sWLkya7tACh3PJrMGPdoajjrl7Nm+1ChY4rT0yLFbdux/eHnTjvQ5KBR25TbeS9
VPHbVyNjWiEsy3TtIdjJsMaTr+9L678i2S+CtjayWVxH0oxvpQHiaByZ+uhQlsiEJQddXHBuNmEv
OXv180LlnT/jkwwNx2Bo5Sb4oVJzJKOytAQsNFrwVe0oWpVsRT+DdNqcpTF5TEpa3Go6WXX+L7IX
wjrJvdOpIl2fCDiiWC/At+L549jOktkJw8eGD1g0EpFbEHifre/vvJz6ePoVJvt4kscEXKUHXEcs
5ZYyWJfQexdCNRoa7CK8R0COu7vpufeZbf1UOfNzsGhWK2f06lxhRWA5Z9hhXiQCqgdlqnuI+y9T
DZTdgLriDpd4znfC7REOdf62prsaIc6ziDWwhU1KoIsupnGkdjYLFzNriSzw4psfjCqDtNGuIp4b
mN8XSqxmgQDfR+Qf/Zqs2KNzvvP1QIrbeAej3P28gOUMg7PX09Ye9ns/BSopFzIjWtFPr0fOZwSI
QZMpM33lt3myrkCneZz4fFcRPlVQnmfqjIOsiLUiRsuzyjVovqRA7rf5digSl0FiAm5VXb5wmaG9
J6DO2aYM9zSDkMJKGW3BTog2jzP03Wea2rx72zKB10flYl7zhCRHVv07BqiXsg8DDCzx7k/wwiql
e07rzAq26pNG1OEoU3TEwcEF44NLE7e8NrCq1YTlNo0calAgNxTjgmyqKhfV/kvM3jV0lQEIJB6Y
tc293ma9k++KR07c+4iXaOEpQQf/fbBrK/cmZo0wQXlgKr4XRoHkjSsPCUNGoPmAfBm8u49tTgaq
sIrBORa72CpvnDjxxsg/9KpP9Hw1fvkmIBazOL4sRyvTDZFgCR7Z91llUD26wuFQOuG8exCvk3Zi
YdaT6j4Hrijcv6E6HociJ1/zg3xNLJCP4HGSuVz8LLLoiVzaLogdhRtTUHnHwzKin6F0Dh9YJG7Y
ld8r5lBsRT0zt71E+Dwwp8oqatYCa/5lln3vNs7gNZLEItmr0GAX45a3TdGWrGu3j2rwmkNEiRGw
wrH6TiqkJ5Z1NuBVWjT2UWhBGS9a8mCgM3excYdIIItAXcG7PqgoCmtedAGI1Bkx8MPP4ITuWW/+
YhAo/entbODFxXUhg0N7imTf9OxnhnsSX+UM10+Q5WYJ01A/NG0UXSn1FRQujAshB5h398h/hvpY
CTrZ34fPplXPASo0CCNv4pByC/WceOscD94jFOigbO5H32gmm0tX9KxOLs9TtUnNXnaBTYjFmUic
q8zfL7XaJJlmxYbMcKr40atjZSpbKxevsgDY6BFEELq1tp2Hj26OkEESZA1dizJFfpgklgRU1lS5
qcQXtTUJIMrRA1DNVZNA/k1M/aTkKviRHsk1YOa9VKn/p6yWwmXGQM4fLjJuevL5wJTF3XilVvV2
XgvnSkwpNmmG2ZURlffk8HXiT3wLeMwIjDg0pnBVqGBAqYXZOPP0BoEnGMnUoWgop8gGsOAHavZS
CAi+qdVe1N1Ob96qxAEuUmVv0emmQI06O4dNYkbVu8vyfzkeLGw9WGp+C/HmeFkp0Qkrcnq7N2tA
2dXbsPHGW/reJMhVQFLp3cegnTccQoXjxJWNR4rOf2cMuM96ZiruLPtoBV+rY0ZJMC6Cq+G9W+wG
JlUqsPiysn+6Nx6UUKYsvcxjfIoGaPDFHUIuZ0aTirfUVxtrla2NjHZTMHdeR2eJ9zdJ6BH3A5QE
k9lRUQTpgy73GApRGq3n3HwqrLmwuTAWYXJvq5d2pAlOt2Eg7PfwMyVXAEl7/n5zDfBVYYjvElmn
js231vCs7aqOibrv3YFUk7bbiGD7MVlUoUrD3I+COItIVTnJlHuhOr++mQS91TiFhR54yiqlhmji
ASRd+0wc5Gu4T6Gdh1A/k6eKbpQ1bhWPnk+y/71gKkbyTX8AEmOiXr36Xw5VtzVbzBGY2kP2Ex5C
aPWk/dMqvguAacwHmg0Vn5nlvO/g5JU2UUMPg4kdmAP88q9yUsx0jBkkgRp04oJlotIjvUmQUiV0
0VJ/eVyjhCuZTXzaImFKPWIyfpbCc6G1y/71DmERIQhqcIPNuKeOmT35CL0zdQREhG68UDpTZQB/
PF0K9c/KEcUkiBh7fOy2wyB3HhWu5H67FifXfXj0dxEx5IQuHSBKakjayEik/CUR5CXvrRGXNks8
gowRUltzizLLV8pwcwRC1m6yHwWaCFirjBy4svsuCYgozldJjJLY0XmNILNXXzsfBz+8yP+qJdhH
lvGjgEPj7RtTyHktz/ebPTsnR3TRV87i80tOaBrqY1fp9W6g3kS4ecUO6WjO1wQ4KZ83JFCcfo1a
qylQtvvQhPi92UqVSJojAULd9ijK5uzjljLSo3YGBOYpjbLzLNliIA6gSS3pQs4gx5HlQ0JuBARk
/AMaCBIyMLpchETFp4pAX9regzp/6oy8NA635C5v/z7dRUMBpRegwRj3ETmtS2jAwq1pp8NhWSVO
fkvNupU7MdzHHrIuE0jn/hGMyBgpP6HMyzzrzAuVNDG6FIEIYBVaIzTHp6o7wV5BxoXVBwnNKlqL
w/NZAOZIT1x0OOieY42m1RpAOYymaksOif4Iya5HjGIcbnmdPzw2W6U7QM5AagG/zfsdRrGqsmOe
i7OsNJCd0jCCZm6FL5yaRDn+JR4+Q3cICZVpUZJy/bZeZkWpDYQBVF3eUWhhFzCbCKvSFmpNzakU
0vUL1TulRxopa6rfOY95v6M0KQo1aUmbWEYPOIqtWdyVXVSITbQTffOw6/3ix/6v2py4Qc42VFBJ
Lrp/Df1tLiiHXYNV07GTPSnOsRaQQe5Cy+17zIVhAcMIe0YMmdXQLR71CvPoDQNPoD/Kk3bopMYV
2akbocFFLs8b/y0LBiRzKoT+MTWCv1tkJDBMIEFNbOgkfdyYl2FNyeLCanuBKtgOnZhL+T6XxACo
ezmffAKzY1aOJ+A5cjfJ1ARjzvNO00AkTfOuFcXr03nR6AUk3iEjKZHkGRBrnEKhikYocrZXvDhk
2A29kyrBkAYwQ/SKDNf+FT3xEuRUM8GG49EroIcB864rJTO9nPLykcoas289iEmeW5xi4tRsnGTg
HuNSuJPvSvARwbqoh9/g8IRPmSmLJoFQfyrOZptHS6MYnow9Bz2weWW+KjGVS4fZ17aoQvuWCyAa
7/S/P/z/f3k+sKq0+8/91AND2yPZW0o+gKa5q4AAkeqH2KoxLM2UZfIdy0Nl55JgQl/GXEwqYq++
B1LDmzuy8lVEESduuJNsPv4pD1Ri9uTcDsNu4CPBl6EWyQjT5NI67QrzzOZnr/IUth8qYg7zLRG2
pLUvzWsgv23AdXNOOleuuSVTukxqg40nLX/K9wZSH7zNU37gTF8MpVgUalRIb65fX6pXaa6DvcCy
jdr0SAphcySnHcTRNMcpg1yI2XGM3Rv6YqpbAeeDfPtbniYW/qymXOz6Wi4suapHIAi+hS5p1kwd
n3nke76oSDkWmYBUklTF8wuH3BCzJkR8ysJWmD0EHAIF/4o/o67itUnsITcm3a1iOBghr+DYTsFT
7VifD35sTC7ts1+HOnxOpxCgnekC7S1956LwTvrsXwFEkVbCagxVEtFq69L2AR9xWVkMDQY5Uu0c
4XuRRg3E4xPEHqyofHoPhfNECH+u4HECSn/eeyHV0dY0Iv9E8L5zwX2jLK7Tq6GC/L3iCNwDXGrr
yF9j/c137isCLE5VMosc6nAh3bL7nljmB0JcAsUaQZ9h9MlWch45d3HegFgnvvfx+/ywhcBtfVSA
O9fg+OIKbYM7HHlT6uq6APirWN4/lL+I61tZ53s0gq18zU0kmalf8rMUBSwl4SoKnCK+BfjHzUbg
1SA0GZ2jbNgawnfm8ayAjDlmgv5HTrKdYWEy4luBmtg4x+b9r1BQ18i6+MXkC5H7ABpM7MhR5XVO
aQa5lY/n3Dc+JJb0PFHQsYOl2Hm3mmQnKt0dyO/zjwusPEJL70B5EXrgYi5K6QnwUDB3ZuePZDcz
9hroKhMifZ1Gz63ImTlRt/r6COAjQGhIMi+eWAIrSXpZssa+SHbCyww3CAx4bSVf+GHV1LrV2P1j
Ja9eQO80JZklp8dHHLT1JL9Kmj7xRmpRMLkvzfpYSncp9j9LdhX6SCJzMsjGDU5/TGYmKSbgBs98
KWlw1AA5Vc+AhocNq4GrltyxcWA9fOIQbvcYKIjTOXgHH8y7uom1Pd9xTex1ugrOQPXf58gJO4X0
S7+xZAcTia0XTU5WH7UR06bA28zXl29UwDRvs6/QzIVZldcjFp2OO1sBeISdMISqfIABmUtlxgnz
KXzahNjaTI9DEOw54s0IY4UqKqJxPJe8oIREAzd74Es8n+H/t9lfBV5Zmow1RUPF9P4BDyI8uGC7
3GI4fnv1rR16XGAdiT/7vDk5snstSUBdVUNf/ujWm0Axf109uBg/5F53A3aNbC9G4hV3OvNKdRTk
aBToEyqlSnpw56aTSRDAhqmV1mUgDPX1cZugOIJ1uD+ufMqLamO7nda6sWIRMmqyQST6o4KbMKOb
X3kSAIkZmiZe5IzqWCLwOMWoWXWHK++W8unOo35/r7EcSwSx2SiHSGEuwXKyT6/vWskX8S9Q5R5k
hW9Jp7c1Lwv9QMumL9HYx3/G2zQkFdQzdFqvPGv32EyRs/TBNW7XHtA1UkgYHqnnrl/K9/q6wGFY
aeANjX572i5mswz7L6ozpiZsfM6KXK04I3pxtQ9U6EJJbHI+rzTzPTBxa84ExoSpA8w2B8iYxp1D
NxtxvMx+4NxGgCai00LPVpGL4qZ6s4JFQ6xe4dr2l6fYnQQJGsRL1Kx7symziYciwejBPhyxob17
b0X+OrHLd7Mm551dgxQomSko2BPcAppzh9psJkPRUdX9jUFodZuqruLs/I4bop4iK82XOcKJg6g9
yAv/eLFYL1K+imR0fd+bwopHYdT7JISz0ssBBT47fTX6O+xLpGyY+nF5aFYG/IaOIZL9slr5vlo+
tqKhqem69sTyAPKDUqx39+GlVxrJAN0PVR8nJYrJMs48bSLQ2xssQVVHN1qbwsb+aonNdLbYtNI5
8vnST1IoSFUUONyeVyXCN34TuYRvwEoloP7XBTumWYbzTsSfwdwh8p2KNC2QS3JrnliQbY8lM8w0
gWjToTfr+l23ZKvGn4kuu9WTF0wo9b08APkVM36oTMPyyNOn+0gg6KKTJtTxgcZ7CjAbYc0HfE2E
ZbJ7RwO5Tbyg4kqeoWi5fN6nbxTjh/NzPFm+tY3Z40OOBHcd46D8WIVAKHFMDesoHmqWk7h0ilHO
uXdhk4+fLCmNrnQt0x+4uA+AQXa7mRL78E0uuRzw6gqXbyzep6HFOIvERe4kgjcz50uPtEBVXE7H
Vl5QBoO2K/iuRM06oIc7VvjmBr2vvECTxSot5qEmFKWnEnBRfD8rZEwZxAevAoG0iuG46KhhoQq+
zG4Jx7RJTpOea2Ef6nB3mTLVKPldQTo3l0xaXPWe0Pgk18v8BpM0i6SCwG1VnuYP3bizXpPIoh76
KKQKM5tAfwJcCS2DcO1Oj0mRe1fwMzvLpmzU+HjZOnuP64tQhUTM4Jl8kKAsTuEV7puh0vHvLfqI
vMrg9D1KfIsVW6gsbqDqbtMqQZ0DHiVoipNinTpLwznQTxfNKvCECX8y3d68MVFE2o/VtFD4XoUW
U6++J58x+9knlG4v6CSgGNUZaTcVRzMsQqiQzXG6MQa3iSiDAkdet/E7Yet9doZ/+7YIR65nAw9z
AJV3L0tbHj2Yh3y9NqfndDvKpeZLWKfY0l82HiLpFXbxrLHoYAaf2LToUNfvWufK19RSdK4lPLIO
uxCV3OyZxVf9c4/X7OJwkeWTnkfPKAazJmt75B8mZKiAkaF/eaJudtkUFx0woWgSQ2GUSP3hlv9j
yL+d+olMPW/yj/xTyI6DjR2DoK37uCPUd44HJkwq16o2omJA1w43+WVRj5VOc1p9kGhOChqF0iA8
id4paIb/6wwvSqKjO+XASQBot1A+1/5QbS0VDP9PtCfE1JjKdDG8/bqQVglAYQ9vd4aMt/P3ASs0
03bIaPiMJ529LHlzUQAUApe8HEGU01LUj6Q0JkdywSzI7uw/Pa6bsiY/ELH9SRYztKqBtsGCD4+i
m60s6n7bV/QaTNOt89uVjoDuiq4T4+9yXiJE44Q47tUAx5GcEb4U9gJrsCMymVXGL+GMtV12aS57
pJwHRtAMSWjZpoIrtF3P0EcujNtn/NSJy30jimapHmOcrqUev1jqngyHV7DJ0RYzenUY+kZiS5hw
j2/MNBxCH43uyGSjhWwBz25lp+TCJeJxawoBY2JDmpxOQ6kvnMBPmKHMpC43lhIiwUgmeLyNH87H
AYCSH7uXB5Iqk9LMV2Z9LqQ0vpBrNChWFLZ89cmcyYk0NtLEXQMaHqYGuu7muoccjfPjyfkBUIj3
Ew2CMP3xBBx7+jQWSGwTW+uEpnpuUW94vGwaOy4SCkKg5k0Ext795vMDCgxM6jp1hfsco/+iujlK
Kz5ivRPN8oOA3Xe+o5IngkMkD+JYLpZ7Vl93SIkpK1od+bUzVSLKZc1Rh4JBG7EiPZKRCkcRgyyB
gLXh3Y/VAWNySZPMNmOl4rg06LB/ZgwG27fVQeJtq3JGDN/9XTmybW5FvNr3ctnA2lcB0G+9oEaV
VNiAaCcanZg9RY16jF23Gr5ovufXRbWN/C8aH/AzXK37OZulz1Gl33gFkmL0gpn8JfjEV23oV+EK
Em+5A6yJdB9wNrgWRILDkB7cPyejaKdab0TZWKmG/VtYZsM6wijE1YpiR9KsFhhM9h0h3XfFcm2V
hopkE9XwV/5kz/909cGNzXxX+fT/a44AOqM3T9jEulz4vO+HYF1P5Nw30dEZ31LdZIgfZWf6xrZE
KR901g0wwElEMbpA2FBgEy2PFhF9QofLCUpSEqBBCQ9pCvqX7PI7S0v+TIrC4PUGWTObIR2/WdQ+
eoWz9shhkMyto8ksMYMkufszDmJSSe0eTKWt+6rAWnT9IhTcM6L1S++blx3Da7KZrSZoGncNxBBK
HM7H+nu33Jd7eKTMn5sGbF/AIRFxej8J3DXXcD6huu62drf8Wu6F/sjMC58+/BLu9FGw4p6/W0sL
SJnoknhPJ+nQtwWyYf88N9A6MlxKntj82xWmLZ4CcZNbBBvAzJxqu7JFFzQwlWL8STQcuMDJmKfT
w680pqbEnS4X390v2s52ofcGLQjX+u3jBEKm0jk25mxXI1nnlbjkWRAUnWiOTOiu5rknMrGHr2/7
8ac++Z6AX92N45FnNqVHTUjNQqLXfmAvpssQ0vb6uqe8aZ0x9iVCq+8rR8ElZSJg2VKFCBsjvLBG
L85dS8m4SQggOR0eYNGQFh9KNxNaHZ46tsxg0dZP3fhYzQWSmz63lns/ooQwO7PnCm/3/mRckP77
vrV+MGZNVbNESXfiGVKqlAMh33wHqdIQflpborzf/U7ct1wCp56Wy5QhnU60wkL2iEjvugxJZ65p
lHgitN4F1vsggLqqs7Hx03RDYk+8ZKsD59V31ojIePpzv5GpJJ7Xk2vlI5c4rbRVKiZfuTFSh7uo
HJZJ4p1oBPBuSmXeE6j3IBOxSbblglqjKRMAD0qi+EIqbiH4uwSCGIsZfgi4P5Pp/8OaLgL1n6s2
2K2bCHxg7RVQjSr9PA4bNcvXsTyaPA9rVed9iIKaQ+wBU6AarQWKZsQH7Y4LoOtq4uQIfp0wiSYB
9YteHxfET7fIS+AmdnxHSUbubJJAjxhKUIau9o9wP683j+bo0UsX3XP4BYF13h2d1KuacWKZ1Tp/
6PVpwBcKJXXYr94ApiQJAlxhSL0umYX8llE7TiUKRjgI/G/nkoMmwL9Ss754PEKXSgBBWAqEPicC
QrQms3arG2MR29sfAjDoxs+W/MglBJhnXMbK00ErAg7JHC1Raru3pfPWbT4cQ/wsGs6tTnz4U6Co
etk49vGJ4n5cHubK0aT6RnHNefv2WmrmE1H7Uho9bsj4hMorns33PyiIG+sf6OUbRFh/r/rpBWNb
SQO7VeobU9YnjQN/tTnbUBImUSwHqu2GR7T/0tY9XrxfwgZ8iPikQKtP4ieU7TDiRBLBZR0bcmQ0
qsY8D677/rSIldgC3oQacj5jGD0lqjK/OCUSqJcIiegGOAisrdA2rur8HN5ZjUdR580JyQBmzkZe
s5QypjD99KO6eDJ/UAPksYMAau6mu6at5JtubmPtNYulVKYP3WSfmcMs1k1Z2+n84KoU7bhuFz37
byGj5199dG6IV0MkyGkn6vVFkdwp8lgAHEfaS1CfdQHLRDlQ48QpuglOvumnkWWQPEgD05hHqlfy
taVpIHk/WLgLgogLW3d8eLzLOQcnZ7jtsueCaOvjAGaTo1BEvRz+JaH20ihtv4DV08bngcHaICFX
uhKlIJtHMEqEqJRvjFdLjQqXmb+LT5o0xs2OpOwQNFaXxNUbT2FKNGTgZHKT45U2gC9CE4PB3w+7
GUxdFoKL9Yzxm1fp6TFJsppSDPAvccdbu8vULQnXFuSS6bb5WoWslmvnGPdwbhKpsjOSPtRO1UiD
d0uCW6RpjDrW+RJRtd4MUDjkMG3tIb0F4X2/ZxQF1BfL/O1+ukBysgLe40NB3YM4Ul+3k/WX62gn
qCNOQcW34Plk2AoudVQEZRHoe0NZLB9YJ75JGffVVuGDJhTnUl0pX96Xhjc94G7bnSmericc5xRj
BJ3kMET4B8r9P/+gQGRqlEqFkJ9RR7MW0OtNMMprsGNqU5HQqOMBqGngc4ggAKuXPUv0Ejq6k5P0
EBInt02GyKRdBqJOzgwFqG4OpOI6y5qRMze7JRX4fCqqIfOSQ5oYvUvFDV8Txk3+IDWm1srSYT9x
lnHuTqeKS7WowfdEK6GVq/JOFCPuRH5LWiVALlsYFeSS5NZ/uON3oSeqD5tnEUT0DeG995sHmcsY
z7GTlIrckddCJrn+RHJelgtU1iQ8u82h3LdzJ9YHqEzMZ1AVAy+PTh6EZExDRG5qjbgkh1kqAWT4
sCEf9w6EL06w11vwGLZZiSTT3vpPgh9loCYOb7a2WbD+d33vk9M82llGw5LmskwuGbTTsF5oZIgF
hvd/eeeHFRFUPJqHOIxSxzJCbYEpZWPqL1IvieAqWjK6NnpXwZ7Jm9NJyQmWtKUj7RNtTR2Nb2XX
3jFPJF0udeZDgCagE+f4GviymhpnzgD32oHD22c9PodJGR3b+Pn/dlP3EB+yOayagmR3m3l0DfMM
1EusBUp1yh/r4jhoa9F31uDq8Uta+jYoEIPYoN8g/Ea5fwiHxj1gmmDFGUJZW+v2+zUUDIwXR5Gr
66j0tA717kvYz8e6YNLWAZxfRXYGdn7k/eayoDwxcs/iy1rPxLSq0J4cAlsC34y1jALAI42CFXiz
AOKEkD1CSGVzBj9XQ4PQM5IozZMqu1yiV9JFkNI5gOL81UB1pupNKeKqfu8baueq4vqI+K2Fvh5n
yhlH05Cq9unMNqbnILc5CHl8kJPqK38LNSeaCwp8HntwnK5Fgd+JUzDqHRfdlI6bKARMmSkuZdIK
4Z8xf2oeAaaVFv/6ODhwsZML3A7G5i9CtvBz10BgL+E1rNKyru14KlEfSrOzSN6vx1Zem4LDsUPP
CEiliBfkpgE5awOzmtI43GzDeeCHS3OkHGh35Ue1OnFsVZzVRtCzLrdDyW9m2pyb8PU9V8kehcTD
DpK6ucUTs0Scb1RVpGJFoBX31r4MLTxJ8O1jpgwdnVDfUIVCP2pOjed3mdoWzYoMm+sSTxxqv2Qn
V4PXFXxFoq2EXcWKYZA09dYhVnsVlS7J9FylFsgVxC64OFyp5pLIV+VAKFuAeaTsRvVTqKkedsVS
79btF2LuWaJTRnVpFBB/54KCE+SLArUWip9PTNm7H96u56aidopPbHobZk5svvYLnHEBNv9FQIG/
2m5zgrxTCf4RPNOowl6ts5dBQKcCVmyi/8277wgKfwnjgVEJ3OQSGUW99k8e1hEj2pfCmf1HgNsT
h25GtA7oSs6X/PA5c8Os54fWqHzqIo03wTqI1gREQWoBgIo/MQodLHvMNNfCcSRyODWqc4O424H6
d942yFnsjQE5QrDVKXb7TtaJdnnZo4O/nCmbqLHyXBEUvhByx3w9PjgzzR/goJYBSzcqcHyQ+sdg
5rBshIChJ2i1jG5Mz+gzCR692AwAkAdqzBInvT0ZSMWGnZVCA4idihklfxvxiP7cE7zLjx+rsRsb
sQgWa7BNDk7OLIMRobrZ1kjJqCfXwmWfT6XQp5irIHFTwcFtXhs/yxz6LRB9M77zP2KR8RlfkfoI
f6aRVKiOOYqJDtVY+hAlOIG2Tx+TjGAcjP8Qs+OmQUwzaH9OZuVYZ1a/MsrIK8owjHXVFLWGrcep
fuwdiAIwg2c+GKkutEgnFrUoZ4/QBCOaIB4EFwa80KgRjtL7e727HHAYRXvhXHN1PpsEH7IFIEya
7qwGxUO99+2jnkw+4sfmRT2jitC71wph6GBJR/viYpS5sO1I4bMXMI5GGHbmD6xprA28KhMOLM8Z
zZuyROEhLyPPOjULR3I1Pizi/zGdaZWXFv1KR+0pjSFwXPy05aiMiwJ+wDfIBFwuhOb8FVyK0Nix
FS9B8tYfpqNe4jwFU47Pq8vQQ7vLCNKdyC2D6bDUYR1n5KRrUMAABJ8Jh19aXJMwhG/AinjPkEBp
pFRINXDsRRlagl6mWx2zC9I90zBFACthzZxG1vlhQSSo1fWS//qX0LOX2nLYPOCebg5IYDzy4Dtk
V8i/KlMjN6tT7gaCvaGlV/YtvBV7q9Xvg5tgdw6n/U8z56CJLON7YcWiNBRGRH9J0f/a2TYvdXV7
mWuKqQ9YPB8JXngRAV9ri9emIYlmx3ljwaPU6eNOnrh7M8fhCeC26aTZUaIts2Ei5Ry3FpYB/XwF
/sHrC9rtGkpgdXqrhxNTJ7/rOmu4B6oNv4UpMSpOtgXE0rjGdGCRN3e/o6wQFj55MibNCMtr8R6O
RaG7ntvVENtNsiYvyKL0q/9VAT2h21ObwRm3NLonbu13tDWzBkkqa4N8+9WUrzwlvA+tVAZWIrfN
kj9PnZAg1xYtugQrUZkSxFpH+eJse7k20f2FYrbTyZUVKchf3BjmcwAxRGTXEHAfHOXhrRds/2Kz
/965qmkaX5tuiJGbAeudbJQc1U/mTl0SAKrgsnE7E6DaOaMAInMNA4r7p7VZpFxmv8Ek+GjvBXzd
fwsjvGnqGh7P7KWVKRBep5CKWxKLpqggqgp18LSwtVNR0Z56H6O9dewI3bNYpELJQwM9n4F/TNXu
Won1ddOgGD8DAr3BXltWHsX3ZBAr9UA7gIKGcfZToP+xlL9ZHVZAEr6tur9N2T1sMt2iQm9vX0iW
Kixs6Tv3V+FSg+I9plqP5xAGgOH3QQ7cLl6QE8Ynp8vS+OCTAS7HBxVko2IDuEVa3fhS65F9k243
+LyWr8/sf5UXLzkz6U0RxDzJcVNNcFMGiJ/p6TPgF38ku5S+3Ko8r/cZ7+pBZQeQ3WfbcsZmTrkr
SoOIv6EzcmGDDlaV9ciumkRK98IClo+lS+ngTZvUks/XBlrNamfcriYpghLNuR1HIq1YQugQP0bg
C5a70qamq5quCtXTilCDRPXyQcEsB2QKtevKShHS5Qksg4Zg6T5pkfnZfPEBxy5rdUH1RGOrgJ2L
zDNil0YK2g15smuNgkuJWXAGoMl093HpCG0/9srlw5DGCYlM2I8D1qzew86nPmmJu2uYkOS9EEft
rE5Xe1RIqZLhOnSfhMbZuPEyH7lMPCu1ZmHj5yiyecZNMqDV+oT2f7UabXAhJ3PdXAK0jOC3PbLh
2SBnHJnLBxibl1qxDhVfU9MolFIIW3rmuIhYpRLTc2se7RK5CZ0I2/E+RJiAT31HPJwtn4js++LK
UJnkmtWmEu2WJ8SMaCvt+zok3MweR5p5XJYsX+U1qdFEA3i8s9jIMiyCzlquTBdNtUJFvSaiCPaE
9KaUnkYTaB0EKAxbJpbf02RxkROcI3zixgOI0292pksq3W61K/8Q7G0IXEF0J5NV7NB9uNoATlWg
YAxrgHN5SOChFN9Z36MJtta6WsnlvUMqMSZdmrUzNbQdwF5UjNUaMEUdkG+ngMlN4J34gJe7xfuK
I/mECNg57MBOiNV03sj1dZqfdMvSRDERmK4+NnDkjH5imCOw2e8sjBEK5HEjlTlHgAA13mz9EANS
cE2z2yJGvRyPqkaaFRlr0z3s5ZImnDrM82iQwTXXT15BGmCtXkvB8T9ei4r2YQziNnOuTT8EVJ0t
u82MCVjQnf7BguOgW38/kYFytnvanGcNHngvEPN239KGpggydD+sRT+nj5Wvto9cpfrP733Ga53Z
1o2ijZNPbrV0F3Oj4Jkq2UAMXmHBfL/JnvSiltJeJtsioZi0tko3Sq53CV1MqDgAq2uTZ0kUT8Hh
PWyEdvJDGGD/OE4AKB1ivAy+7Off7VwJixPpqKtwp8EpOZKlejTeYklo9wot2AcEScoFAJPHjX8Z
cAo5HSHW37X6M/T/bE/enJgDeMWc1LzRs2HzjIoGwc1yn4zfGvj1kiuTiUCrft34Ad83ThA597ii
pqM5+Gw6va5po+hpOUxrHt1FNskb908jbRAb24MeS6pqlpVx8BCIL5zBoJp5vtaiCTtAcCTr+4sU
kVVjaw+f9C5upAYvjnWCofd/DYvZh4CeqJrOU4hixLZN4ta+QRO92b1a/3fZqmJa3wRArHGDLZhC
uJCp972yErsQ9+Ob+zhQdV7PKS6ZnpPRWmhgrAbj5ISd3eUrzBob7d/HpJ6OdgzZYeiSUqAp9GIe
gokYoHc2IWC5swtSZ7b0Df/idp5CpTNjeVzP6HMEzvDoTV8UVpq5NIlZu2lCk0CSihEw/DvTaVtl
BVdK/Jx/HKrn8iV9KHfCWimOl0rX3RQrolaSS7h1PZYHTMxKt1djDZdH9O89e66H5HG69aixfMFP
j3PdEIm1BXdF3o1HRcdBIHmDelqamiqzJJwxBy8KKQmDfGr9xBE5l12glm7jibxjmW/3Sxa5tHPR
iZhafV3F6S5GZNqZRXmLBvvJRpF7DjGViucuNh2ZCfNaUM2CHQf8aFDCjMxIGM85I7CmQtL9Jss8
iRSxYUjW7umHKxkH35X3i0aCtXksmWL/HjIe19Uv/Tk2HG40rLnReDnl0tKk96uJeJhf8to+ZVEe
V2vfePUmHpcS0J6I1UjQqgfOpqg4RrYO8x+j96YWHDA2StOkLXLpcuAb6lvC8YvIZI/uAT/Bd+G5
xIEux1K3m4iTecPWFWMhEvDL9aiL2JMIa9NmP/XrNfBhGWRqlUuzmAlxuJZ+Gblhkfk3BDpvMQ9M
k2A65Vx44rOVB9Y9hu67QkpyMbsEiLNNwt1sUufmOR7wEI5+joMjPfruhsTJOnUiO+aXktb9T5yI
wuJONXiNoKnI3AXAda7qtsyIV6fqwa7N8JnUhBZGlmtQ/bc3nwJ63T0h/g5yGa42+3tL78UAQgpU
aA+4Gm9azfDMqs4W8IqTn3p+whkmzYp94K4zBBU5I/4fsAbQL0yqih36WEIOA+JcUBR5g8ya4f21
1955R7v0FHBD+MTWNGxDfnR2ubJCS0uM9Jj98sWb8TzRgBZfmxX8YxRRbMkPmpqyl6+dnHVi/gZa
5dOhtavTsCFvvHXJw/b04Mjppsnkp8dnaFLd2y33e4J76u++xH++6WuEWKdQWVud/6LW3oVkExwo
8A7JbSGS1Ur3DfEnasP/X5Ku7kFeW5D77hAKGJB8HG8vBH5OKHU/Qqh8JRZXaW4uKj2XK6jCcPSE
pOL7cqF9K42DyHSkIuGdG9BJPqzdGOB9hoBITk8OFQbi3Q7tOPHC0bsevXV/lNpZovu+kxEpKdT7
oxCvkfWuTF8oWpVWOQ+Jk/0zzhfYVOBjTMKCx9WBauXLOVTmrNGtaOcEl7AvjV5FKTmUPxMAVxTC
vqfKyYJKxxYzUwKoTAXfWKxOtBPQK+nsuMmGZM1VOnP/HacuburflieakdrlGpG/49VMvPva7E1X
KpUjFZyZlox0nQcnjbRH3dBSHekQYG45YUZOZhxNz7Q4AXFFGJ7MyeQNYhdMB+2EtE/EpqEAhGCn
sQm5j+PBBj6YhDc59AUU/G+K80TYBY1UkbIBZht7pzzZu8OtqPnTf8X8rX8l98EzP4YZRC25fu8W
0BXouhS4RgLBLHWtOm1CESiofqUCBwnx2rn2+AaXpzkWYswgkVFZNjskCtmN1djnySdUBuMRMn0o
NW643AV6BFKvf+RHUf/spzZe4YAHa/qI2/3xGt9WRcpglLKWjZAH5zbEM1MAUiaogUp9JJONEpiX
A74BIaepXCYi5qV3jRAcZvaibj4+KiIQbWuedQcZZSDpu2zbsDwITr6z0ToAuZTzP0q3Bm6sBLWC
3qLTHGFN/P06yNpK+4mFQ568sDlgA7nolPQOoamBQJMYNi4FNHJN3eVE2IU0rzpGNo6+yyUQ2GTg
OWpz4acLTOLhTiB5+3RgrXtjqOVHo29kMmRZltKN6wDSIp0nES0QuJH+N/+FI894W6kHWmgr9uqI
k3eBeJA4Rz6OrhT+pQNocqhiTSrU518GJu1loOAkFshZDoXcNQQDQeC385Qk6E7T9ZNtwkwCJcPb
k5p5JXNmC2omN37ayW2VoMX9kuMEy5OULQvLvPaU0L0Ykqi8rYOPUq0HEwt4eH0vuu7PLfipIdiA
33UQe5iHPBH3PVRpzbb4oBHf8VJGNOdA/+7rDg7MDz+ivMDMQGlI7oNqulxtvAROwXXnRTWeAOtK
hdWiQNd0Ca0s7lf3KMxQ6W0ghBMBZd1gNK/mb9sNrtOC3CdjqxojzQoYEBl7Hy/I2QwP6aS95Lqj
jexM0ahp7uxjs/IKJtk5Cm1lIjn+uXTwzfRJdmj8o4SMF3BbD0BkteacuXX2c7UouNOtLDF7ctoE
QqH0LfnUlsaO+66zq0UTL0i1qaungJU7yhRhnf06+VTKoqweqHOhMRIx+3skChHFrLiLlaxGL1Yi
mfJCGG+T/OoN6OZd7BgFlLuu4CZZEPXiN++9KHZNisl3ysdFkeW1tl9GPPrFoSdKfw0YIh9JfFdR
Me7FJxLr/TJeBkThqRo0lkAee+sIqhZa1FkmF5+rTrvGNJn0KX0+Om5rc/9DGpyxDgjqlzG8EFEh
MOMxHoqUyg/hAJcK30G0WFsALdjCxfUU1yWCXkeLe6Ijxw9ePYBZbQ1MqGhriqMRQ+C3QRR6wvbv
dvc4Y1VhcnF7e5PrzlMTZ8HaV77hXzNr2tEXtbB0xUUPAbMMHXwjDoe4ibSZlOdLTp5stWRYPJm/
f3ovT7hAllFZoxpD02MG8xBUo5BXxQnLaWc8Dg1Qg4avAVMT1KO3rUE2/AzQwbvQ0wmzDsLroqPC
5kcp9qaV+Erddqwwey+P/xlX11WUJbpqgH+0WgAREgSUhet6D7IxMAvgSoZ3dP8gPQOycT6GgsZY
K+midB9lufkoWJNlck+5I/tpXvUwEkazyERloi+Uo31n4xi2zQa900koPbsK91xEyub2Pu9mc+2v
wmLCdgfuJ/RzdP+T1ntEVhNVlv6+NvIj6gnnxuCQ1On+jtQlKpJ4iIsxCoKZ+nSF+qt19FSHLVAB
heliymMsyJhmiUy+8LVAvB/F4SxGmMWQWjGOiWfS9w7sGPU7b6IvfFk+nMJGJTPYoGaraGfIjLfr
C4GUqIFAEHUkg7lO53ToW9iiNbp32kzYLOYMLXJhowJbycdizWz6ILlIzkv+1p7LglZTz2rzpDbc
UnJxlTetSHnpURn4Bena2X6tSl5iZDcyXRxosqi7iFua2H3jXBQ/9SJbKwk9frRK4R9OsMBYO6bt
GPPKNjSyoSwkr1WDJd0W8Bu2IoKVOADIHagAMZsZgCelV0Y8Jt/JorbQ8LM8lpKFs22n8J8dNA80
MmVRCqC3N1X7A6hKFusCZDc7odsieiy1zFZrfUPHbZNpxNhMdWDKb+QxqBq2PeIln41Tmxw7sdMy
FqgtrNLgh2ttTMSUCrY4J5p2AQovLhlSCz/DZLj5JgXLGE7a6yHGx+ANuIypCFAdrsUZfnwi4fdF
NOo0FruBTHkNa2vjnVv3NaWnWrBcSIXwCPYFLKwrxsBZLc1JD5JvrwiXcA8Jy5HqR3jIPhGTT5AF
OWlLCOYUu7nLgOgkfpr5D2KvtOS1kawyY3pDPx3nJ5Xr9aEiJmKqNOzN7enzH0GpmXIDO/TTbCcH
6D5y6vBtix2fO7FBFrBQFL91DczQTD/DKvkS8rHFT62nG9PKWSfWdlwVjjPzgx9i9n/zKNzILuqp
lOoGBuT4dRZfmOBxjzAJKgnQ2ilYye21lANXPxHSSIV4j0kXlfsSMSvD2yLVnIjuJA2EeX7av1Yf
iliPaipONP5AicjIYNn5QsjH0hzkFKL5DsqOZbRQJXDmNJL79oO/3B3QYM4lb25yrLDuh1O2MksZ
sOKjf3alxMbmwvEXt7e56jIGPVO5FQ4p0Q+5TRzofW0AAWIbpx4eJ0kasTZGTIEZ/XMD7sczmJOE
un45ZihZ7yaw7IM5XEL2Pbmxbc3vq6EKE2Ee7ImTtQwQd0R8jCRIn/gZIbMJPqT1j9P9aIbwJYxq
FOLLmoZuNp+Bcc1j48x7PoJyvVp5cjAUnGPz+eUdM5LuijmY2/Ok8Xr2EDetjvvdf/kE7DKQgNpQ
52ocY0f/rI+HVoNrUsDRva1/U693WLK5DxLu0+kvt6yMiXI9DYJYATjgmv1+SAaFG5XC9inGSRCj
AMEA4vMWuL0rfpFoTS4H1NP2a24voQ/tw8HjtWZt/arPjt/GVe5xqZktrcFoiWcbdarHf/ZOLoWE
8p4JMVTL/mNyCXlkmmpTqeC34yF9OnQXpxLM/jnz3SXNtfoDiFl5fEZClyxc2wHZwvbRCs56yhKm
1UrgjDoBczJAPHgEqE0FPNTolukc/OwvuZ8Kd4iTsDlloSF8c/SENUbGc1Wtr84K+YfREO4YtVAW
15p3ih1kawIMdCDnCm9HnutfZDpbobx3O9HlU6DzdwNOSMqJv684eIU3+vs+EX7W+3l5+MG1bczp
p6DZkuaPix82NPB0mDcB8ORhGhklXtcotb60njitFMI6fCHkMkm1KgKac9gwN1STR7jY8Bd6eLHi
Rh5mMEC03GRk42bwMvshMi4pP2kOlgXSmX0fiJHsuimRdjD7BLKMB12W435lDouK4arXZ3ApJT4n
vV4iLqgDS3JWa1QmRkoc4muMbN+skOGvfW9DXTvgr6fJstEjYSV76Lpsg4y3IAtcDqZmHCc/Dfa6
VJUhvRNoZbWYSvmSroThZg9bK8DBniLYZdZv2R6o9dTqOyQPM/3TD0XKP+OiFc2G190Y8sZ3erXT
o4yJKyI3UXPprRmbD6ydcCdx8+DbRkk2w5tvXjfV+fsUsM2/wMjKuBFTMpKCI2aHw/b87CxqqmlP
WzUUBmhHTy/YVnW45qRp2Ci7CcCx7UPcCVQrMd4/qKRHc4uMcaQ0ZKieSeMKIecxxIdwYO0Z7yzL
FqwYOviQOocEqUQhcS5sI+KQW9pD2q8jg6d0ZJH6umWhDHhE3nY3NwZ9zDGLcWrbkGm4MW32AKnF
LZy9opy+4rajj5fd7gSz2ZgBgLMQjATgeEKtUxdhzwmVC33gkZDfA+jDeaWclieOpnQqXD3y6Rqx
LnD2XD9O1Begd1vHg2/nQq7EIg2eJvdnyyhvJdIbCoGAiG6D/AuVIZ/I1PWWm4Q0hQzviuRoBYhk
DN/NKGVM24gRM9e4s6jprZt+7yf094Uy8lnCm+AdjrOppncrPGqXe6ofl2NjnafkWNudUZIyVjQM
NuX9xtODENhEaD37G/0tiXU/r1YJqdMmdG3GlvDef83vnoQ4iFx5xhhuXKF22w83a5ZoNMh1sCd9
DLTtNdMGKgulHFGxmCwkTQktjzyV44oSqd4DEVps6Wr7FBTrGk/+ReyPLkkoWhpMc2I7FV/T41P8
Vjybg0u3BOSBufYBA7KIoS/W5OV1ky5qexV7bsaRTUncIrdGPdDqxc8fOMJ5A2JuXDIIWlFhnuXV
pelkTX8dlMr9BITrv0VCInmLqzXk/xil0nWjyII+kE6ts07OepJ9GWbSs3ehgkYDkphEc0ww5KQC
y8GX2mbPuT5HiDieyF1LHyGoy9nn5z3JbeQsEWF2h9nq2ZEkLXJRCdLgDPStrRk7Q0G8eiKsE/Nr
lYUWDzLrXnfq4kzjWMzIDFWRmT3t+AaH1bIM3uwbPM7lS2jY8mo1jjHrYcOC2jaCG9I7yqs9YMLZ
ohaoKH/12DUVdMQy6jvM0xBp+JtMByPHH1bjGeD7S9M+NbPfmTF+a+AMGbryuV4/JDkEJ4IY8fLm
rGHAJv5l3Pp3c1DDkc3Zz/yytsgp1qAjLrn8V6JA8N/cjQQwK/laOoMmbQcPMPANSh3K7CCf7Xws
9PvGednFfSCnZ6a3KrvqK8OcpNmzJSuHRChNhowo53VApodlzC2/uxm33jrUp37ccGBNlssVHNip
w5clVK08BnP2FLzRUuGrsASkUs6DgL4STa3+NwkvSpr2AmbyClw8xlM8IaCxjbimPXna+59JbzcS
XF31I2MPKosQd/u3ioVycMxuM7PVzqxciW69FG0sV6jzP1LSSZBZgSuZ7TSrMhvHZ7OpXu/V9cNu
bY75Tw78klCIWIMXmQAgb5uQr9Lb+HJc7pgrvIy0bORd4yijroJBooQrn1z6PUL3W3VYw8KzGIDV
5cs1H7VsXEcfOWOj2F/t6naH8RJ784v2etEH7FNBV2h1GjkSShKbIuCIWYTSZ9BVih7zlb337//i
FnQQzMZzFfEgIXsIP0FoolEJojwtyFg6lcTDpgl71lSNoZH5YEA0cSdbTYKQSBexz/qOQC6HeCvz
88HQWOwYvJYLBMwMhx5OVtwua7/rsCYQd00Ce8VOcAfGC/0WIreFKyZ8NSgb6jU4JHrtnXbNnUJ+
9Qa7UTpBvYWd44+muBgZBRrYOPP3KBNzIlPLZHHPhOENJk8Vw1nbwkA7WlN2zRNhwI+oi50sD5Gx
tQeSN9/nMOI8UYi9/TQuYyfTFOQ/5y99WoIHZr254c1rVWCXR7E9nqgPUoVGaxkdFuhAUwdR9nRL
31r02DjS3W4vMY4ckLYh6TlI0pSD7eSIqJuKpsiwLYP+5oWuMY6hqT8KVYU0noMs/Zlo/oWdIHqQ
W3Mo2bLCkrdFVi91EzfrgR9EGaelvZwA5TMSfAiQMV/W8w8oQ6DqUWHPlR0JpNy7E9OVF3qrLV1+
O1cWcz04hfkB0A89xxSJhK+VIt6gRtMHD7yOY1nY+1dJhvCae2ms9sHZaEs9WT0umD3rnC2dsJmF
U5J9pgSbwUNNYoFUw6F5P4TpZuoX4cQPvDZWP7Y6N+x9GZ8GWWWsqseWZdO7sQtHzuz7lXROESzD
cs9orXBkAVFCV1X0bxz/jkUNMLyIxFXG9FLyB4Kf+ivUQyGR1fr5dZXvRpR4hy+cBh8TKXJ83+xG
JUlqC9/X4s/lIjTowVLe/74EUQrFGP23SVfNaopCMmBxMzRN7eY7uFIWM00qQtOxU0HojMIerhdZ
+gicsLSVBqvBQvsHW7sLvWpaFP8HXCKyusl3hdbzF1rV13Yk8wcmhbHOZ4KdY2KZKCC8gSg7KhSt
QLc8CbxE7ToHIyYHbGjVoyE7YARhvF92zYVqSA6uYbkvPQJKAHNFXqbzwyD752O8ZYnnbHaHY013
s5/XRapROsXWwHiqOUEdTbAEqck0koyzD8MHDuZtKXf0G4r98A3q5RtXokOW4JjEUlO+bAC1Ft0z
ZGZ/2f+nLeK0pjhGN81eULSI+VezLcpsrUg9/wdmQoUMm/H81yhATXJiCi3qgazUy7Dtv8C7YWbh
XamZ3lJs2y7vc3+6Fo4OwB2pLnAxhTH9akpiIE8HJmHESxMJEBd9gKghVP7Ydp1AAN8z6ZusKIPd
MXANcW7uBSWziKvYnsI12A6B9Vam6jwU64vkhtuDXNnQMWZSeoif6NTh1E7j/p3Z/gqOFOgTYQLu
7ZT/73RaoVeQ2uTNW0SESyhhPM6sesRYxQHT18RnwmVrGsfIQycjE219Y8TUyGqn/Xo1Q64v52mz
DWau+HBrPEa7Zxizl3XLO1m7snrtB/IGSr7mLY2qSBHQbtvfjlPelyfu3YCNiPOy0vg1Xz8FPuD0
OJJG/fa8UjqPcGm8dKR/Kp9+MmSLA8haUB0+cgfxnjpOHXlAVr4RYIAIZKGcAUElgqkZXiKkd3vQ
HyiXgqkDFRivVl/83IVU5LKHNXtC94qq9ajmCpSAnoAiRomk+Vz2dnM8lfiOmYQa3Me+QzH3RkGy
N663WhvOezMdgt9s11iuRhVyiDbLbuiHz8lD1MMQQTh9dt7ocPn6Udm9OboMxJiMIbZjvCzlxwF1
FzKq5S/rjxJt6MORaPCgPANoFenw97Pl85NJ8yR9l1+/HfY24bN/rwEIOA94vKqrk7VzbblZ9vK/
9Vw3VMMiAd9xY4FuRYOgZ8YZ2l6lVs6HZEGMkl4ugvqz5hvy1VqhcnxTAf7jEG6pN6r2RbIJ5cbV
FezZmkoQKY8LJdOnmwX4bjPJusN/5PaXdC710vzGTh0puUdZ+veVwQH9zrRJCFCs0iJKbV0HU3oC
pcmfCOrDeTvmfSDH4UqAddETS9Ctwua9iOAnD4i/JD+XwEeWAyN0bCkpXdazZVEYHocFPqo2LhLu
AoxXG/Ja0TUQud99U1fcA/ZKOK6g+h+KMgJAUCFbRMruvrmo0r/66Z+HupMdMibzw+i/+5x+GQun
qKD03VPmZp//T4UaBTDOx7Df3+fMYMlUDXeQ5T9NT6fQmj21dEZD3lHO0muhiQA5M/Qzzhdp5OeC
mKE7mpva0PpnaGHg1gcGsY+NqzG23AvNlh3CTQ89Hp1iQWOytUbja9w4QYprpdVEMbJ9pAysTKZN
FId1idtSf5guEfNceTZxOQPsJEr/wj5uLjueeZqhqJo5Iqvbooxjw4BWe3/20+ly4JfIZ2h4TKDn
rtGxrPHPsxJylYrw00AEiZ+c3GVKOSTCuxVpxiMg9KXsj614fVW4/hZtBI7SO3fApu7TBonFv3dp
c+L6sHTRjhjfQd5Gf9gEoudbE5MU4rzjLQBcwJdrOu7R2Oi6QQWhlUm0Qwe2iwme/xP6MRTuF1HA
jB7ujkU7qa9Tbs3/SpgPKk6xg8qh44r/7lhvX/k/eThjvR9C8Xj8A3x3LRTeyoB6nx+KmNjMNJAv
uPuP8AbzkXTEdKOPbRoLA6Te4w3MX6lhNlpj202/FstpiMiauaEnfNr9nz3macDxht+0ffrZM9xh
accoD7VRHTNt4OLdYHRUfHKQWFmT7wG61CsOjaE/llJqeUifuRSANw/qU7aTilQISyCNwgf+yeWR
WxXrd9u0lK17aoYL/Z3fRF8wD3hhyGhICeGT77bVSpyxf4AS2FAa4NXoUtXzaX8fpvxQT8ISrOuz
my9BCJaTlRoxzJfRUnckW8oxtxmSCMFnL2gvfA3irjSR1UbM8X93x9yMEDXg8HU1pb0Bu1P9ICrD
l9lNFLgc86lk1pR3/VcFqqfiGL/oG997hiR5H1zso8Ca1uh7MGIurUf7JFcgBwD2L2BdKuJVvCT3
FTZyghziuE4J8/E/GPvCGe2aCsW3scXuBOXdbOA0ueKt3rhBKPOln1cbtH9hZBd+eZC36BitW41E
Gznat6FQrPE62W0JCpWYl1M0Yvvhv43+1eELYEpGfo6OqPgcZBImEisaTGKW33IsU2uzKjzayN5z
ytuiXNteSTENUr0wqW+oJqHjYaKYmecQ4dnfaeOSwPXBr8p0//DWJ6VOFyfotuiqV85DZUUjyi76
3yIcIJfV4SuUVHB39mMqfBmJQJ+a9B25KqHhO2DtCswvErBYUUy3BSYmM71W+tRCwv04n1vP0vTM
ggpvKXo3onXjWUDDLn1P2vZnqihZweqNILsryQ9xFwDwJLmNhHRv+4vIttzRmPXdZ0J0Josdrwaf
J+8qPcBqco6I7EZ45qLBxzc7vZDY2TDXgMTsjLnQReBoivu4PsMdjxofOpx3V0hUTy7CWchuYYyW
HaZEGUdrhtqLb6uoIf0pbZeqqrq1Nu/Z1K2J+pAiEslj1+QvE0Gz2LSMwnJfoSYe+sWj64kkCWN4
9g6gw3Zg1/OxS19k22VdJITyy3gHsFgbSDOlEwtbWcxCCLcotzbL/C6d9+d2sb1DR+eyMHUpuIvH
Fk25SxHvT5cO0q5jQWPAhqt5U1s5s9stG+1q7LSXANZmu4Ur6nPdi6sJ/unMADDulwhDh5Tmei1p
j3mz81lH7AL5gaam5frHuYuTuk9bb49+v5c4Dpi71kRMZGsXwT36LxW4QaKTxYVaEr+Txwk4ZRTt
Dojm+SAV8xAuSrZ4QZrd8vPYQg6N1UWy4laOdL9sH+06878g3ZLV0iUT8Myd8ieKAtjOqablLRpO
u9Px0Wuk/lT1mMDL3BRAYm+3HDMA1gSIcOzx3/rW77hmoIy0JTy3Fj6Vo+iYHYWnaWMpuTx5+Aih
0FXodTa0q1qqM+DXD1vdteBSqNIUYXy66Xjk/OABA1SLp4/Zq9OliL1DVpb5MmQv1N9VuO7MYa+p
ZOMWqud7111uSq7UTQCNesJbwgi/AU0lEl9p/9dXxgZMj1JPg/7sEpb6gswP2nRN9M0MBBnrRgCx
2Hh1lleTQSW8VY+9Bdr6yEJ6gWUOSS8ivC228g6WEYW2naofKYoFwzNz23t8Y0iZX8nn5zs7qedY
JZAQMKAMfa/hZTaTP4Ueh/rostX+nLDLJpYgg5U87A2dPlbVBtnbXJPqseFRoseq0rMYfW6UVF9F
j2QqMLZq6IQ/NfZ1iQVBMIXQeRGTfKdyuUC6os4H26e3uPuv42Hu+4Mp7wBnajKbNNZBlIHeevw3
id5Hh0Qi6jrmhNA1cym9piLjQ1FqBOVTlegWkMRH+/PpvBWty5Ouv3k7EyZ3H9niF0gbL/TwDOkX
gXqunr+0s++A+aoRwVhl8X6Yu/RowkVnovCMNSRj9vPWMe7txU//rPcV4MwR6BBPxHeZBwhu6att
mCJqY/CGc3+8ZmjDeoEvTa9RoHhj3xbvl5hz/gF430MS3PhFeH5IVQIyHxx2oOvbbsBS9+8EThQI
eP6ft8aQk3xojSWt8n7uITOeQgdv6e4zNqnsQpKFjJheQ8Ie7IKAO123T3/EoEZesJ8WF1ezW/pQ
5QB/U2mvHXSVDf4Rmh3E8o6DBKNaMznagrqpjOe33yXXH8YpdlmZqvYStkQlYT1dYfMo8bnHW3MM
Qmzbz93BfRWGgVp2YbzMjUarymaur1aspmxXdZFcBEpX8L3Z5ktuhcDLvwU2Fn8+it9GDgNplpbe
xr1tC2xj4Ghaoi5jpJY9WZlLrg0ovIF2r+/qTYiN9CTCc3iPreSV+6RJrJ6KI0kStZWkUOsFHWub
ALRicFTRm6nl0eLwdj/SudhEZg1RHUXdYE/MaTJhfuX6pzFilXZMgCNVqNK55p3wp5RDG/TViT/B
HD+6qOXuzEgEqj4AbETkhijtqTCC+uNeN0jnma0cV8Fevv1oB4+7u0jbVns99IUGDLmcXMO6C174
iquTB73KisEfcYLJA52glLZhTyhVoaFScd60Gc4SK/wT4sAhjXVCZiuD81XiJgFAmJNv/vT413Co
726hZjZJFGAnfFy6y+UZ5tN6by1yD67aGwxtFXtTULuMlWckiy+mHEHbt2CLBPX5lBFd4bH2ac1l
vcXQbD3xAcSb3V6hKP1ojheadW7cNiI2tuLbzdz6igmuQXrxpZ1wgvLmwTpkFVFSN+s74wf24L6i
tN6lxUyTSOU6AdOBQC1XsGfSIpQt2SjonE9iF8ABtM4eZ7Gvox0GWP0k8GCsAqpeXsMvhqCqyK7H
k8pJwgpNUp83ODUoxKA5vvG3S4qHdFqAFQtsOnmHKVp3jSA9P+U6Xa2WH2jcIb1pumKup3CaUUXo
Qf/PepFQrIk1IXtk8BwB4osXZ296f9wB7sv13t9WkAokmTFSee9Q6Q2SEORobhQMgR/THZoDqOkp
m5ogIpeCvwp+EGxzqtwbSkLbNHoQ2pzH3kX9I/kBq/ksRFQ+t0DVfEJ6wqpgiCM2m2gkR8SxXtya
60QT0e+mHXjs9AFAkw9epgGfUHPLC+yK7LjCMPbbVs+sivDfEqjFTR4FmRZ+Da4lwvCDmy/+fTt6
k00Z0LrkvKRNreSI4L85oNxAbsr7ZVSoQJ5l+4Pe+2KOI3Mcr/nl6E6Vbn1+XMfMaNIWSLT3Ta6H
VhQS++FT+J1qcUh9u7xNukWITNKEoybf/1dEdV+Bzw+aaaXnYN7JBWEimrhGWcvUP40SEQxfGXeS
AqThm2su/xq1TSWiZWlilPU2wr6PsMOwubvaFL+3x9hbHt/n3ZNgyPBGA6ukYRrheKG/3WiaaF26
WUX7Ojq/dvrbPcgCOzej1iCvfbAX3fqivUBPsbSgSEbTi3p5Pjov5WQADE2ce4ygePgVmprem7wX
3h9DgxGeDlh51oBRTw+H31HKIxWsQm/ru9LPLs5al66c1hDbLJgq2Pfz4ZkZi3aWMZ44IsMjzi/K
nvUdeSRNvs/pQ6oe3miCObjCkYsYgEsgPy9lSOg/AvMn/pVWEr9/W7MOaHYZ+/b8QrjvN1wOmYa8
g1SqV6V4iAHWqggTLWMLPRU/zXApOfNAiZwI9zLsoYb66sTAVLIED8Wo86JSAKygbOSHZDlOxl6e
TANGcylMjYyKiMsk0hdbtWop+aftUiUPfoxBs+O9i7whySXfxtG15ce7A/B/ZuSQTNxriIVt/AnD
p6DqUl4SDf1j5laY/FJlUkfwZ77cGp3WVi1OZEtINTmjLvxJp09+skpQ8wDGVwCBYy0ZU3m8Yd3X
7/g/r53wzUA2poHkVFajEf6/S1hmzkFQkBoMbpz8qm7IumjrjT3VPDk7VkL6NtdqvyJxgYxGlbHP
4r/W7Ao9GHJm0x9/vbiWtP/Z+iGepZ9Ntz/3SltByRnY5pVnbSGLOyC9v9IJZyKVVNIZl2nbM1WZ
IMcCijWo5h5Gds/g7LZPZUt2r2wPV2cPHP047aOK33NY44WHI+VKxVHu4cUYVl7ptK5ly5IBEa92
FNMGMmq35HPCctc+V0A3hltw2rJbruAtiThyY+zPFoCU90AiNFVYZEUuYHzohWC+IcGZSU1OD5SX
CH2W3sGXPDdXAPhrEOklpJ4AlmEaDKdS7RtYXrU+0n9FT4h7L52gZnbVFvHaQpbrBrpDdxqBJ+5z
wN1l53r6qRz2Metv2CdXV7YjHsNVGFdTvIlex54NneQjaGevFgVUId0UUt9IM6ZfIad5yjmI1JMO
EPhfDE7ajqeCL/BU2ZMRqsl2RLYnUoWrqIrUnE09r8XvKQVAGs1464HXI8wOUbBMgKvyu0GRCfRE
fNhxvobOShDkDsgZkw/YftFYpFaJWBKHti07WyBdq5x+FD9vomT8lhgEFQi8byv9ReMbURsAg3Bo
I9VDggh1yzosY/Iql8Fnow2HtqosrjEbHlPU8JAg5sifqJP+ohjyxRaN1q//sfMtiGTg7LIK92fI
PCocRXElexH56VY5dNGJwszUOWzfksrnjSnIGcVeW6+QeXKz78Dn9W2h2lDhdXniDb2+qqLf2ebD
Adi9EKvQdkoRtXXPQiOZOXgUYvwoyDW8mQhoRqOard06/VOHo2kjeE+9AQ5KK1WMYs60cipmfKG8
EML870N00VRn44nmNHk30h5ya3rr9MrQTNO+YRqEULV3lDyKNg4U1/BW0xMo0YZZdGTcH97rP1aY
F0HUKjzZL3w2WK0zcJOoQugF6RZt/uRMuLOitYreL3hd9WG7PU6Q7W8JdKdf5YyQUL6/TkY7MMHk
ZZm+EhDJMr25pvrmsszg3HA3oiqgJOXdtM6JOG8g9eQD3V5H3cW6YQbeGmZaVyLf80REEm3wda5s
ZuXUDV8KebYCo6/UbmPOQea8478ttgIT0mq0TBVbEGvryaJzn7SoNgTeFAvZ8f5qxVzjGYpb3Zli
whMncmg9gUmi/zAqlfSktbkwviVeaC5nREIF03mwROjT1dwRV/yQZi4YRJaPRJBhfwSORI1EfMVX
7y7vzHkTE2Qh0NBxMByAlp5FYwu7UY6qs9XKuhmbRauCVV8PbGwZYoYbbNSpO0sGzo0WSmYw933A
aHz03Q4aLg7ZAdMFnRXMnrO1sF31RHkKn0n8eu28GdUsr3tlGNhSPlMhnDHB6A9Ek5OGgRn0jPSd
O3QzhZNvME5sC7Ccs8jyGTgLFtlyVmovOM7YapEn7kdUhrz3JeeS2M7vBKwRNU2c4mztUU0eBbmu
8J0EeXq3Euh4Cd+ev2NRfYw3dV0+S/aMVxTIyPNqxYiFfPTclHtdvWzgpySOHzSUBwjDM6a0sOLl
L7hk0Awqf0N4r4UdqsZQKMcBFhnMAftiND+XATetMLofC2Yy+9M3SojtydFMBlgLWK8hV3rYRIvh
+us3AODLumI31Pna/C9mdaoIUAJEzNF+f7IHX+r5mjpoE0dEpswyG/jYf7CLZHBBiWDSICfldkFJ
vlK6blvw1HdmeFZPy50yecVzEh3bt2UOQ3ccXNpwLXgOxpVn9DDMXwFqcTe1VyVPRsoc29gEenBQ
JWjF283hoKus7XcQ2hQB4cKThTvsOpoli3XauXTOsqymr1sQ+kZgONyb+mwLDJJ5FZv/3H0874mA
bf/3aETs8dZeQGOGoCPpMg5JmCFmlvyJfDfHfVIzVlWDzWtUswGvzQx5nXF8JVTFoBo0TPgyjgkW
qUboECVFCOwFlWH+Ry8KYmZX4FzSjdrSYM+OPF8SRD6hKgOOXZ9meU86WNdEcl4cR9jqiwJlc0/I
EubRmfjiLTbWURMAEgdrtMaj0MsNlPzjdVhVVHpzTHD2/3D51YzmiOovjtk6HTSy2WgCxgz31xfV
9v4KkHgtMuPAEJpX6SUrrA9ORcPBA1KtdJHOZ/jm6s+UtQ8Cs6557J/tyuD7kFzgI7htF6Aht/2m
GI5MjEe+Mu3ir7/qvDk0z+eCFZAxmqXjQ8EQHFw0cnERXkuS2o3DYxXkkna/OjjIIwvs0h4DWsxP
MDol8OTxEBaqYefyUHtWlO62eyiVwhkcGWvfscmlFECqYGccsIAHLxvdCiragFF0gQ96h2zd7ZFp
Dcn80tK4YMnBHPp/xLjvtZh6dA7NI1y2LhUu3oR0HJL6AvZXnaovr1herr/fZZVppME+IXlbot2X
rm41epk5QWWORIt/JWD3DP/7AHb2h3zZlyb4yLlvASwPlQpPCJuvJcjp/lPtQWc04Yl1+XwGsV7+
CGZA0g/3kaWRbeUywtJcoFoz7W2qhjJBeb/DNHyxGcAB9RvzOKOxiZzKua/OMVwhqnvUJf08axAB
vQb2PlVQSAs+Ekev3V0GevYbRUUlcQ9j65+U/Vip/zjP7ZCsfSpCWiOC6RJNO2KtMBzw1ehWXb8B
YPJKP3njSWiqbEM0Leb3ghH/XgudYgNzDXWYAoTLN7vf9sp7rEstde9w2qn6KwlWJQDMswHn+lEt
Vonn8kDXWfjdCRS17P36AteJqPpgAanFP+DP1++McvcRfUiro2xxFsNPypeGq5UGUcTvL81Unzrw
W5pU+SSITcCtpkouLimAzyITEKKBZ/WPbJRvuvkSElSrOCJ4Ey9TsqAJ/TaAg6UFuieMYO/58zaM
6VbDnIa0P7qb3cSSyMD1zBbkZ5Q+F/kFxiMJcVaEU77OIE7gKtLdej1uKWU6XpD/Zo41ewAbUTdR
vvPhILDILCysB//Bx7NZCW7NQkoYBXGW0uJOG/oB+RlakB0zg6gc33ZWw/ztejgD2v1aJI8Oosqw
qnz7umWi27hcn+gKiMOs3SwLomt/AWO8knIkqQDroUVTjae+oLq3eiZNaMySt1L8LUh3ac3ithIR
lv+qpNjjW6/fLumnDRbP+zvp0J/48eTQPJLa9U7ClbHYmULfgNHM73437s5e9ih+PBYn+o+IbONC
j69haYr0uzIF3RiLcafiwPxeqzCCrdfVj1l7Hsx4RmOQLq+9aHDxSMjd9yryOKW0rrbW/V93ubyH
+PCkmu+Kz2hYIuh1VmChuOJbOQ86/T8qHkQGQsB9vHrZPtgmvcLP+EydPGKZ/SXYZ+jXP0vJF4Ol
Lr2iPnlN4IAZRcWNtUCUT9QQmuBeo8bzbofGx8rBUXtIQNJ7QaQLxm1H7+dVlM634vk/9uKeivQY
Ep90JrU+2erRZVAQ+Rl/iFgxMGB6pFJcST24xeL9XosfaWjhn9LWaANaWjVlnrDJqBcQW7vjlhpz
uXxHpB4WxJYEKYjBbLe8XoPe/wmAeQbbSP3jejhbc4uf4jHYQfj4KfI8kTSw/8lP464JMsKX4w0Z
Gl8UNhDWnsHK3MycdDz0dKi+qKbhTpt+thXyogPUpo68MnOVAsqeDLHMpzc9d+o92XcETj20nRoX
QAUGvfTkueFTp/MtZXVk8G4UTWTGmpaoCXIonI+6XL5ncnOKZV7RjWZapeVZkoBAesXR819COWGW
Pc564nrmkPNA/h9rqh0g/a8DalNnNn0OecSZx+DEAMh26a5oMDHCJAlwGcvutcpykJUc3XeEoYPj
AbbfHe9tVm+ive+UPqNAG4ZQxgb8uHYChABCZGTzJgQGmO6cdiqTp8pcJc7PryXWTrRMd9qtmHjf
hVPZg2c/muZ9XI0Y8CkuAzVRLSciealWq77Q2TWCTceyoy19iqT7S3CifbuHsInPwL8pYU0XP6Ju
TynOq/scgw/PuszIiFw3X2pBywBi8lL9BrQNe8WoLKwg5e9LQcOeobtbZyCmCcz4AL+ipsqbJoCZ
hAWfyE0g+oy7sRSwN8Q4nwAI5LHmnYcLQRa6JzQjaDSpVZHOS10uslMwy63cgFVhADb/rKEH+yDm
m0Mc2PUz5bHYoM/Kn+lmRATR4pkzEn+JR8rokjHmBKt/q9LT+Nx8gGYdgtaSCZACG8zFwTzNAKZj
TWc3E9urHQ5odiN129lqJ3Y4RMArAKkQHJLdNL5/ctMrPEr/sZAfEFXnvS8BNdT0WnfGmS24Gko0
16DclIlwu+zxu8rcpIse9Ao667Knu7gYIbGS147AptKUjYqG+nhz4UB+Kv2Y3xcYLi1joAqCg+t+
BC1w11LCASq8WdFmVcd1WsNpLv21KjJV/EZcItIZVI5Z0XjeO0XMqpi6SiZdKIG/V86Cx/s8mguZ
e8W6VCXliCp5p/eysj+8JCfd6SYmrrH5A/sEYurhBsvs//tMp2BxrgWCekkbxncJBqsqq0rEyvSf
a/a4eJR+qggViFPJYJ3G1pkb6pl8CQDkhoDI7j84cgZvJEr00g2fhBY4ojlm+ubrGaRfM2to+JsU
xjbEMIQczCQLtOQy3T6/RpW2vrcvL4qxi8zR3HdUOMHuHQrzS7QpDiMZfCvNfqkJo65Z7oGWnLKg
127XJpL1EzsH+ijxgihChO2nCwtFoDk/enahZVmoY0QorXXVxC/L4Ote8+inqGM8nfyiKHWurlfm
ShvhSdUMhQ5sqUKJwl7ZfLzSKaC3P7x0OwOoxe3rJ+9HtKIuf48lGb0eel4miEdMO9mwtNjQB3iH
0XyomLjsv9rdptwWswOUvrbSsTmHJA25AlgS14g5afPXULLP32fNJWt1zvpOfWjkifzgIb08i1h6
KD8aRrwL7L1jBrqDwtmU9lrHmzED/WOUGQb4Rw1NNGb5QGvci6HDvaS1ueTmX1ouaZoo7zF4M2eo
RxS79srt4VRmaRVVwiaBW64nt8gMlBCx2QNW7BqIbDSAqA4jHJWUNnqPHRgno+H5ZTDN2t08MSF4
gM+pJ/27koGdLTaVblCSU7rRaD+n2gPnkovwJP5OW2lH5+2bcYkL7x4HDj3gdGq3ilJqGTE7TfQZ
5tuOb8iyvfu4RcXRHf/hHXcCuGZz7lObeM2xWn6E82xYbwWOE98sJlRiPrb43ASG056yr/40jkB0
Qewh0A6ZgBh2iL2as/WRoUNUZIHfN53HkecK0xe/sKvl4S9j3j0JhDDLajPGKzoCgWEuVCD54SrU
wqyWqIszZ0Qr4rC2xwYneoEsw8T5VIcenlhCOjF9d1//4+7mP8XXvhLETtDdamLt04EibtAnlJ8O
kC3hr45wASfhjgbGDVokh1vOydlsAZLh4MfosZaqnn/Jso4fHwb0zKqMJadaLrjLAxXRERiYEICt
pjM1srv9Pn9+4qUOIpnNlVKc6HSMPUqzkP4ElpSDahKGzioJ5hxlZ4kJ/LdhKmz53fvhn+ai1e88
4PBd9chMJc4JNCgCa1Nx6zCWu/SdSVxwYJi6VTImGrP3JdmijIsy0hpDkJ1okNp0zvLwxHcP3r8V
rPBwnWnx4d7J86BA/KvFxNb8P1L6nvKE1wcDtOCYpmqls25+vvNXCz47SeVcLB+BTxmWrLitLb1E
vlD47ud1MbpUByjMoY5MuCtbws5Drc7PwI6TJV4KxMzTwn8KbNu2zUmGrmvaduRzz0zx2UkdSoyZ
edzlvJ/K3eQ6eqghBT5NhWgjCqfsDO2M5AH2XuXD/re02VfHc6Uqvslyo7VF32jPbIPTzgdd/Ncw
zvtfQelO0Qmd5+Rwj4TzjpAcBLfbDI2J2SAywQlBGV5SqzjsgLHunVp2De0fKpumnAOlTZfjyplv
BKH+W5/RlGlel5EeAHnk5Uz4K72+fVyDTm0F7ow7iSVwnfozILauThM+LEKKcpN0/Ctxr5jwrUs2
1JQZd2xtArSO72p81ix99JolcP8ICPkHtIa1YkYjL7cC11bcsFfU4vxTAc3f/gHqJyR83T2Id9SI
/9Jo86iojdLwnnpYI60piRtYdX0UdOrKhNImfebLooqT/y8IGfZ1jbKrVbYsZcAlr7CZBUMnZbRj
6lRaHljW2ybqderJ/vSQwiATgpIpGDj7bcLoveUbzkgogiRg7OV+zABSllkQRoxLAI04+JJjEy6Z
zzRgO+ltnVIzSpnE6YL8P2HogX+BaF15dyeQafEIN2TnaVljcBrGghpdUgDNWCbvV5COZCQxVKqE
lKosPxkM1R2FY+xDeImhKaUFqYd34TSBUuNz4s0j/lmVVnAHlysjoXdfQWqWW2AoQE9G1Nh8+W8z
+chIAiVTbFno/f5FwomWWDsC4ma4IXb+o39wr4LiPWWmUI0AttSUnKKV7tdLncHQnBDSYPJMvdCd
dhiKiQjZqGQR6FiXgmLNSOKlOzGRhO2omUcC0TzFmUvmWsD5ZJi9NAhBqWKDntqifP9euaMr3g8F
wsTwkO6Q3b+PHFg8BkgHcYfU2nPjcUTqBP5hH1pKdpfibXYn0plzpEBeAQehUiVqOXr114J6Zkl1
uMmSMNP8IrKbJpcnXsltVOUubmWqn3IYjcrYlYCCIu5E8Lk9yypIjASK8RDM9c5LgBWJ+eqKCrkG
QfXkrkMIf3b8G6TESr2OFod0x+rPjffZt1hN5Pv5kw330Hyq5Oz7v6ZyqtwGJ7LG+/JMV7EJwr1y
y2Zq1uecauQ4HkJS3xmKu+SJb6jhBB1aPfoWE0+pYLsRUuxPyk8EUzipMNP6PRoXUjndmpWcifni
fCimvfLWZAPxoZLUU+l71brUVE3eBBHWlW3/hL4oDwJeuipORBejTuO+cbE+/TujqGdwgv28blTz
0SsEQHj2NhvCrLoijGBIauVZPrGvksafPEUaXoHoB4BUUY96KlZShDQaS+bgooJ3C9KwFuA+FO4r
uMh8H093MEft+Cg/WNSJq5qs8EhumNSwFLvVNEtJAudwpgTHZtpSGu7ZQAXQW1jsShfBnX93kC3g
94JdqcKqg/Mj/CHVTtVGDtcWzouAUNlaeJNodjV2y4RHKf5840+x0Bl42q0fd9QHHN5vhBH+/cVK
waCtci9tNH6ZLMCH8bn5VAUN+pn1r5vIQedcUzSPcQW5rwVHq+HrWKHssnwOqUj4m+65c4t5DxpA
TTpzZ5/ceh/mkFbYFYue7uyBMtJhPikcSzmGGR43O3pO8CyU1+KVDtiXf4eB22whbDeI6HOyle4j
cZg7uCPiYhvmXEQU21d39owIryEQiuD2VIuJmMRaGWaGQegbizDC1SeByfx35OvrrpGxyF9kQw/z
FgDoZOyeXCt0FKphLie7ABU42wYyy4Z/7p5MY+WcsYNeNE4nj/lOqIM06FvDD1Br9FO3BOdoTYJs
9WSWhr17kczSOkxt89tTohdEHImsf7QJpTy1dyPVPBKZUYu5UyNqLmrllDuGclalTg8LuUOUMdKz
EyeF6rOOcXvoG3Sn3eyWVJvSlQJ7i4pBlz575vqJVdXzTqKfdaX+sAsYejWT4xIk4QYKaJDN8EHx
r5piI14G5gmyjsZotRStwYrbWbRoAhBZppUxPz0ttiwnOtBOyXADGcTDXeQgn8jwzGdCOXjtRZkD
ABAAcPvoOtfmZLpox5CBTDeSYOl8LXdCxndCDKAGj1zrQIEKZe/Tby6aR+rnJyNzUa90tNzrCBWx
xSMl2/oS2OXE+LH8IkwlhsmH5XYH4s9lOG+rC1JjNTOm+/5iQpaSSeh1mY65LZ+H6TvvLiYLBwaX
G7dhi5KTDD0OyFc/PczLzqHLsRggK/L8KWOaYfa16nEhOznY2Z6sVboRszMlvwA8vjGBnMGnj9BB
Kx7FIfpNoEuKhaKKHB/PSVUhxPcDtb7rrkgTzSXhjZrJFBRlZdUP6m2sCIvI57muo/mSYzdEbeWH
Qu+u3ZNEJ+XE6G1JQkBg40AQa8KMQGb69kRcW/SyuqV9ocnDkY8qRWWJYtl+iP79yRusECKEtCdS
pJH+eJJjAM5Gu0PlPKlYriysPy1/RKtlylq1ynC3sBbRbktXwYEVhnrk/WlN2DfuyN+IQcDK+lG0
1/QDWcuILU3V5B/sbYE4N2viNI9G9ORaY/Ac8rr7dq+QccKnRZAKSJYDC2osuPfb7qT7EmOPzH0f
LwHIJOQyDv57al6JE0/0z7GHpEMO4TFyHa3IPLuVCGfXH5Q08GUAYTFYO77eLCzOhBpC0Y25wX+T
1qKTEn8vNd8D24pqQ6llWPRWsmRN+FXc1z/gx5gxSL4hSDbacd5HPnf9ygXXZMr2zlBuoKDSYIvW
VpMPWNaONxrfx3Muv3wkLeDHTbheTz5u9EcH9qKDvlBBFUphibt62onl4KdidIGqXQQM19VUdatw
SW3QS5fdvflKx6B+AvQRmqHvdkM//8MzFPq4DXS6nAhOAFEe8ERMbGEyUHS8faogxEATrQ1LRTnd
uAzgciy2AaEn0xseEk5uQqjYGDLC75drQx1PSteexwBiWxtgVfQS3CWci42anw16RoQtvDkH7BRe
O2/TKGa9KMrEHDpcBUYHvbQ1F3NaTkWv7gvk8K4A9SiM7grtmx9mKbfyc/deeKTCAB2Anb6AndFj
kz3MuwVZftNDMjjemyC4fryQ8y71Do4f/sSeXKcyKLRL5ml0W6PWfctvJCMP2kjPuQZMHv1OZhNR
9R+u3TlfOtaki6EFGjQTjR3N/KtC4Oy8jAza/ZRHVjM2USgGjukF0qVE2bKicUdX7ej7S2TyARV4
obqErIglUpx0ZiYahYmtpOXboJYCQY4dFbsGzo0qmYVVYQyqGy64VRueT02gQ6CQik3EGfpxTfBl
6pRmdY369lvo2fVM6n7cJyR4cBRGwF73BGWDG5+EaiXeUeZQGrZlVQx5Q0nY2pafuU9TVw1fVO7E
BnN30S7ADBjq29OWjp5ZFTbDoHLnD0U2e/QLKOcbELAiIHQnLqeGdRiJInh8voChG8MATtiDnWau
yE4PnUD86OHtc5wGgWQVPJSIxkhB8mb513B1FDFFuP9GGeQHMkv9DyGZ2EiHRPKxU/P6RbsmG0K0
sCQbQbZtDmVM4hLaUqguU52Ezulobvf+gi5eygLwdQSRhRF60Qn0KhyPzXMzwQOqQCmaFA3X1/rA
gC75IGM0WOR2j+gxaS1tko7Xj/bm9QHlXlqdOrcv8ZuRumaGHM8um4aAZqQV5oQBHnpTd0Bm+fk2
GJHp4Q96IPjAkQuMy2VYMzEbU37c/GU2W25kQAnzNcXdd9atYEQjBzpTBDdEaUApLKDHKjBrJ4jC
VfA+MwjQejfV01u+XpmjmofV8CRSCKKQCHmw3bm38IzsZBZArw2ljqrS5heDlj+4DBnIM70200NQ
jV/VJZsFLwpShmF6jxMDWN8JeqmNfVaAsTOf7H0WqXFTK7VTczvrDbXyRUWcj6mcpIUhbJpbjTZO
cqZSY4BFdsKoqc6oTT7oziNsh9TLqCRADXUgZ7Ikk4D1lAjT/54kC+TxzoPzDYRWV2gmCAFSDCYm
/Iv8RswqiVcV2C+RQ2RSn3kENe14EYcp8uRB4eGqkvHOY5Pbbt5n2FHZoEGmKqvBhlsSe/k0y8Is
JU0EarOgT2ebaI0wEmoJP+8rG01LIg1sPxL3xJtG4w/n0YJ2gUMtYOAM9reEsJrHEoTiE2xtlD9f
hls46mY+cMcvNRKE7uYUkSu5Y4t3iToXkAXqKX2U1HlJpgYr01VxalEZvY+8BwM5la7JQLfH/5Ma
gMjmLc1IvA2msZCkBc8QuAFHQBKmpYvi5gyIV2r1OgEGb9SDgB0A0tjmVLN2LDGN/Uxp6qNPsD2U
N5xc3dkqVCQYvDr02ztkQO0UQE45mNB3unWQWTwoZUtBa4LpUAupi9+qOl6xy9J6ff8nYJatSGAw
7jf5Sr8CxjY+2MQfDO6CdZXCjiV287Kys5s6VCjEsfgRZSwrpH2c3vCh5Pla3wvWV4MdIe1DeKYr
UKg8MRQh3csdpB5MA+YwXMyJQlH8583tPhGvj+HOffgPOCtlt7Cv3kpGstLFh3HOyd+Nj/NdzNtl
IbGt9ys+rU/9nqfJSFDvGFesD1pRLBXGgFyFxmn4FE7qwh+Q/imzyODM1n/I+WHGbOkRwi/TPE67
V2ofyeLXfSB0yAIU6T6nxlFxJ4yYNaENnUkYCgILcW5i4lGYUiogr1t8nOJ31LtLLJ5ZcxI/64Yf
U4KtL/CiDqTEuG6gcly9+odNdLbOtM1BpBp8f3t19HmBD1S+gPs1g/OxYWtngkVJXIuiacfQzqSo
iD4bQAaY+eWkZgTE+SMf6OPMoMzjWVwwEL6S6DXvWLthotuQYvH+CC24q+wk67z7UhPCJ5ygGoQ2
3IWTQfiZT47pc4rFzwEwXipxQpsNirqI4+VWVO2bxnNDLk2oBTz9pCnHCNiQwK6T8yk76SMHwYCX
/HAHjaI4UNBtHrJ6ucZPKjbQ5WE26MwOGy50xxwhPWEabxQ4b+S2zvSmy/q7h7XG8iSbnWHAr1Bt
qaXMv14QtxWo/FEHwXAjEgvu14KYWa5tarNPZ8LVvZCWeF2R0taEkaNyIXAhACloup2Pl3h3dLZU
D+dv17U+gxoqK8pNibVy9xm/cwgr3cAYQo35fGXTTYbk8WFHcQPWXUDLN9XxCJYVB35knzCmeYKW
pq87XomNW5g5o8L0CL369ZoqDVM4zoxHEcDKxiSd13xqR53moqEK84bMENutppOqaIbgGQiNkhwC
ZXaS6eXOxZVr5CrY3ELyNRd077AGAKp3cLMn5+X3nWEgZSEqIvNUuP4IifscrinAcmtxTnd0SLWM
tvHcQnJUO5SHrEmIhHCPKy9Wk4tajl7PBvj5/rE0Qh4fOr+YUoAu+cYRc7Xik401t7ldkWgozVNa
JxE5E1f332Ai0uFODH7b6at9DZTAW6VhAFIYgS7A8Mi4JwGngIrDmgudIlmyJHMjP9I5As46oVF9
/fLazOlLb+AMEWeCOe3Rkjxf5A783Owttd86QYzJPAHks+d+c/MCqSitxGPcFSNtr1TjQbrsMOy/
Fn3t2Sa2VOswHhD2bhFPxrB04Mq/OAIFBKw+oV6kOmZ99hW6GPbO5atnvRm0hbSAbYC3BaTuJCBw
BdbATSKp1xMxPWswweanpubusPCt/YjzDMQjZxGJUUWT1HKAwfD2/SAbTcQsfV6TeLS6yOc2eW8V
OFXy0ufGppIRGmQaidN2Gn0OCoMiVLzpfdtsO8qUvnrHXTZY9SxtWA00PkfGZuuxis2IV9cfYg8w
idQkOedHrGGPtoBexGUVCx+AC5tloj1usoaLoqL5yy6xRa8MZv+6Gsd7OP8Ta33dYWBxjqTntHZN
UnswzNOV7fbeCD/YURshdLvfXJG0elVoYhFBTYG4IbL2PfuBZO9NL8Rz8QEkpvu8Se4aaHT+oCXI
9zaR6MDGXq1szAXZohVKoMD+lKB56MCTGCRW9zcEqntQu+8GqOEFO5HukwuRDUcxZ5jrU/K8PYW/
3Hyvkq3Ek2IjwCHJnn0LIikY4OFbyzX1mn+8QD9d3DincXfKulDorkmJk++MkwOnPJbkmKsrjfnX
svYDseMA2PGvmH2P2ie97mcLRDLKT7xqEQb6AILJP/FJEN84QUhq5OsWC0Kl2pBC4cxYMtMNlwz2
vVr+dsdiUtCdtw38ShpOePiQZSHF3NsYhHxXTCk7pnPQRXO/PRAWOx7AqFrPeLT8DZIENP1FW6Da
05TUcUq4PCp9j/wyI66jlbNflA7qEk2ZThPQsHEY0qjriYEMCDqFb7JSIgZEAQ1CElkqceQ56sd2
F0TrygwbQCM8u8eGIyqMApVde4RBo4McLMk9uk6dkBLoIVDL7PgoyJmQjLHgWE72e8m4TwPEIDMF
QEP8yq5HT3Y1/kzpSyhwfxsU/A3CLwa7/FLgh2BMnI2wtiN1CbN0JRGgUCLSocvVG6SxMOe6U+c5
6GdEaXNezTvB07n+hy1VXsFL/hf1DzfG4RyHMw8eegX9umlg5meCJlHhmOfzy5CYOZBNDOjdXspD
t1EMhL80AZ3vnTJDuYOWy3y5tLRF7nyRi0mXRSeAKvpNcBoMURxWZRmftw9QVGfFwoQKc9hbIb7j
BIUw8Fp/YTFGa3bucNaqsK3ymDLvZiv/2kNmeh6yZf629DUKmTwIuSLPZCCwSv+JwC43WxEMrDgv
6Y9MVe4A0X6nLwuFM7qPKrdmrPepi2ovMIBXpq1DxPeneRJvXsIxn8D6YtQA8Fv3TT6e/Z9RBqDM
AD7+jxT8cT3J5pZgwaPtPBDowu2ELEbbru5ZtLIqwxWUwHHCKJ7uU1Ms9FusxLKM48Y3bI++QQYN
A9L2t1bvLB3zvSZDPdKCIlsftMPioaNzVy2roOWoAF0mECzlfQ4UN3yZnpN4l/OagqXxPLTqkPHg
ddt0/l2dNluSTYnF4x8+nfSqQqQEyFIGC9wDWzXTYKXwTS8JUstofVfbvbEWFlEAA+1eHLQ/hnRR
2uJW7zx7MxbuzWF1PaOSSEAzFQNfclaUl1EhmdLRzPngHAWQwqSdojYMDpmazT1XOt6PLWZRnDEU
eEJbtE8C+isJqYJw3GOvT0Qmk3gtwPcpF5YCHzoET54Tqr0A3aX1S1+Kkiw+CHUVlf80SpO2cgJZ
1GOTUYlt4h+lyrYoIucfcQEqqgJwiPZNEIAcBqc8D3yRdLfun1m+vh0du4qGu/ADfpQe+wYHfOgf
Rw3x4Cg6cv++ow0jI3y4CBEZeC91d64R6slu+bieE6jCrTKlBgtqjU+lywFPGoVl/j4j+/pdDNnX
DtU0WL/OrpAgIplIl7Yd8CYcKid83h2/scY+SIcUAb+2X+pogNJhTPFC0smCKFV71UGmFpl4wjGF
KK9PkkJAmLDNdaL7O1BPj4Y76+SSM8BDUII/O2tIlUCqjA7LJwGlFWI2koZrZNnY00Pt1JbaJNLf
wwtQ+yD9wtQgIHYrdhZODzO9BtAaVAPB3yR3/mUrob/O4lG16d0Az0gkNfgIo6tnHnHoQ542Eoh6
V0gGvpMDTfF79isf4attWHaMwZJJCndMiDyB7BXxmZSKsrrFUTWp3l0j3DvXHcQGHV+GJRTQFNbA
m4/nvalT8wWt+GYd2+mHXJit1k/Wg3xr5fbv7P2ghh2FUJnaCncTG95YlipiMGuAXwbD8PneMejZ
juXb/0tqA0KBuBIzZSTgr37dfmrCKqEw2c4KXcnc2C3XeT5Z4vTvlmCfvw1p38ex+8n8OOu9T0y3
/L3ytz4wXjfnIWpTDhhB4IW8qeXcrNOTjJIOIJIyXEsNn/KHpL3DfqCEZ03WJ+Tvu82mFmMsAuOm
4+NcT9To7ZUZb50EvHw0bOGa2hu0uGvR+ge/9GtUnEbpu1yQldYyVUBxlf9dP2Cy5/NJ61WQ/NXG
9JtL/HhQ3W6Fk1bUJufD7wBP107JfrCY9wN7xmNiEaOkcmVp3MzYrl8G1bRnmsRzt8abPPOWE+I9
vlnega0mmF+llZ09aRcbzeOYojcUo4VCL1UEzFxv7ImE6Bn4KVoCDkNBnw1FjjWy/6vodz76KOGi
RiXVmF+N6FGjQY00COxALgPaV7GTiyX/bbZZdnhbHRyhRIL8o5oIX3V9Tdr8thrwR2yeYv5Otqlx
AQS4s+eeoSMwD7HxthowXVuVuvH6dU+bOPk1O4wyrCUvOTmEi4/C67KcMRmdMjRphiVxzKqlrQS3
dV3V2MTSSpnI971uZJWBea4tPS7vBmWwNrv4w9NmdE9xLHzxN5f5jBdViYsXkb7/ebB/cFLaBF1P
l+dQZDl00A15XCcemrb+pzC/5xx8PMOpgJXK9GH+z/ztHMqerfMF+vugsnIrRDeKNUrgRfak9KEo
EGBs7s72RVegEKUVU74quTwRjRHxBtl3lGcsRmLXRzF0Z2RBwJnQSFkxUMneO+WUOVvq/PdsTO/C
zZcevzUj0/VwQOZKSglVW2dDEAAhWqzBu8SO2I4/G//1NUR8AA7rq90/rjY9UFhjlYkof7fx4MTJ
cimCi+S4WW4AWe7VyfaX6qrAppE13x37z61tUOruqcxNla8sNRZb9rVIPov7qd7c4mruwtjNKRGL
OZwiKKFk34gTYZ6CsiwO+qMy+Ryy04a3SDHX6r4J2xS8YKY4/uCXRtcxWy7iQBz2//qn5fsidvsO
BHdk0T5/LQhaZrY6GPbJjrxIu/TJmv3RS1QIo+gCETIY2SbpNJagi+JSB4gCOGbCBpDZ6b9uA2JR
3CEKWfIbcXkLgnP7KMExWAWqaIoVboOr/OWEp3RCuZHrup3usNqnRWAD6YbY6Ip25McYLA6nzs/s
JexfRgICHapPhurYrDolqaRUR29jm6lPAk0gQNVZaVo2v3eWI4CONY1TsV0zMNUm5HTpGDmYOkK7
DENSsfQWW+agKNHzt9gjWCLmjOpfeez1P3D664OyLQYj+X8xqz2jGVOfrjm8tTmwq4FQWGvXtglk
IdJ3+cOp6eVyxNMOKH+V4ufZZoclNQ0KkCcBahg1Os7Hi0XCT5bWTqW4V4S58XCLPTuTUpaGB8tw
4dgAasqjcsnniVgRQ9IkQcWuIaqo1x74dvT3nNno2csiE1+3MholW0zYldu/vrExJHnWnZtBsmCB
5CBIpJ7G9g5B37D8cScQFJT6XFcRN2Dfsgnl19bueBfefTwTy/RnXWManwQxpJ5ifNOurgEaIgOR
4cTtW9mptThSQEoYKdVWPzjFA2zBdPwe52EEBiRUlbfzc96M8aaYXYHt/vqbQQdK6JOgCGzjumvO
0Jnr++mmtuGLlbzugjCuFEd0qWOqeoODZpsR9+++CdW9IWsnhYDpUdDn3fqEEWbZO3B4Wfss8lsV
gt4XwkcDTV6h37IdMPczHekHj5tJYuCX/h+jmzXnC1UutSoBm5Wvd2yTeR9gKl5NSTi4IkTlanXA
J0iO4GF6tz435ag8iHDxe8Wh88WI70NliQqsX/iygQt/vf1CZyUae9EKZDxICNQKprG/8SpswoK8
8B3AmrsG2lVHOsxofyAb31VcA2s3EqXpsaF3sxmG549LTuu5KvT1Nes8A5LnWThMUgacj4oYMgdX
5dT6kfarzQt5giHb9QXeTTLTcaqY/uIflPD4+UasmTpLBt3PWO6iGgoxLPhlHqP8nBU4w7B+553H
kYKgxVJ1l6xVm1JIYtqEvmOLDvn0sbtotwd1SHkMVKA2r1k2HmoBTnDAUjYoS4O9mQUnUAySApk6
YQSUrqc08cY3cbAOMYkaNMipGD24zgYiZlOPNZyUMiChqJxUwsmOU93ydKbfY2qNjXX9Q6gBVpPe
MaTNsHytvcYrN4ESnUKySGYTL1Mw1Zp1ta9X+8s0t507weDO6ENiDn3BDM85jcEyDWu7FO1bVMyk
61EHCrWC/HyygOvnVQ3DgJVOHXVIgFsHRBWLMQ665Z3OA25pHlFKLwGTCDb+YMD+o9Y7twAMN7Lj
qnX8LwiOwF9dJCnkXmedzlMM48gCEhCGPT82euMsbj4l90rrVDZali0T71K88/axwfM1p7/+Fktx
ao6KsH1v4gIcaY6axFbPOlMJzNwfACkP4kQ9XjXxjTPCNpOMGp+0FYS7wtAOOc2CjeC1x63J4n3J
2bLS9Xq5RHXeEyhUm8J/QCCdJn/vmOHIbh1T1fpGxKQw0+IAdYdjJTo2EGUDsemRqkYhQAk24GKS
pc1+HYHO1B+clf/eq0NwGQntT13n4t/3XT3Z4GxtIU7rSErNPQarNz20HdgIzii6Q9KM2XJhpTG+
FiWXNqAJc4k/oWWelsYv4c74cQukX5hkBIDlgbTgTSQ/u4BN2GHCbOETOlQCGdHClO+FES49nJ1k
tE4hAHQNDoKhwewC5PZUuRG3Bn94lpAPRVWgCBO5Y3ufuXs4T/SWPXJj1Mjrg/uWWS8BsDoV7fYN
kTK6MEOVAAiFXhBriFHGBy1U+jHEfj0eXx8gvBINdH7TvggZbHbT4HTRsusNneoN+D1ObQkHLRu/
gRic/PIac3JMGit4xlhpDP3FXQrkScPkhkBmQmftfArZsduFe9V/Zmnk/mGWGrdYL+LVwI/Rzupi
q01JXhm4dAf2t5liGgekDEXHMLJQS3WH1kh/yfsPaDMIJbqf7Zj8Bvba0M2JlFXm6ZVyPYtGdkIz
RLwmypPiq9Av2WZfwoYHDs/sGw4JShbwUA2J0X8rOnOLf4JMrWr6VGkt7X+vpe7/qcoFwuMBsKpz
aCPO/7NDHW1DPsoe/Ytvmh1jWtiZAJxgh6x2rSCABsEAigiqbAvmVccElWjw045sKnFdB52OmY0f
EPaQYpW8TwW+0ALKxor9FRjI6sdS/cPQnQAUSo4kSvkvaY7z4H9AzvceBZPwHZ7YNKcaL0Dv2aF4
7dEK007klMbOB/x68JYYMdkUhCaNXwpMaZZFJZLDSQwm6UuwzB99ISxRTTOFLYewxSnwXEi82r8s
D4wHBkgOadHRV1YGAQ4VxqtVFjXesVsTuzLIcgS8rKY12RSexlIih05hAA9UzixQbhlj8kmM/BN5
d1ljHThmpWXjuMlkLdmvzKBFk07jCFA9eiWhfAh5TBGAhpGJC4Y61OfbuWZxVm17ZbNnhVnVDwIl
RLaySzQ+xIUIHxwd2L6sB6SCHd7BXXuS4YptbVIwAHHe8w8JFTFzoPjR+Qv5KGNPmGqsyiGgAAvM
qCprxgwpvFucqSXtM3UWpqYmVECquCaHSxdnEyOM6I4QkB9f+Z732TYdC9saQ20tiI2dUCGnELnq
WJ8uApvHeSOCdK0p/Mr5/4Gx9Vk+uj5Mgm8WvHk6IEbC/TSQdG6TTlKtFUuoK7M7oXRwzrhrtyMT
XRChVzfyb6Po/u98aRBbrX4myj03gdqwqehEMxhvDrt16J9DL75bWXeOL2NBuCM1uzPioH04ZcR1
mdbiPHAmS2MyoQmsEeOurntc5cWCB9PNediEMqBI/DmF3Qt8KlZIe77UCANPLYZOudjdMq27KRhq
6TOxh6jAFljqulK0BSPpySy6DniUqrB32KJp7RYvo6qBl4IhwidtIdMXu7FU6Ap77FORCGS/klxw
hQ59HPwcl8Rg16dxkYEoKn3fTFV4/XKNWRyY7vByqNqtM+d+VFyvTRNfC/aFqQEM/Ks584gYReS1
nVfmc5Lf70SyLp+2LzezFw7Bfups5YVwq1uzl9L57Ojp01JFewAuhXZ3rmQv12vkMYrz5l5zMK1b
LcdSyH1LuW0bsl2Egp2KYL3HCajMsRR23u2hEkkhvPmTIFBnLCSeS9s4+2v4OaZrlqnq1ddGcwCP
wGtC0HxNNsGOEA1xhB1meuXpOeTP//F0hthXVBIwk6gy5aVz8lSsYtrtctBBnSd2BR693KsQ+zsZ
JNVGTkxBSTSl1bVfxZC9nCnQnjBhfTZRIQV5a+Oohpj+qLgQQhUaCnVj830qEt5LXFjNvlm+OGVO
wrVJRDBiJWr3zcgdfBCwkTUXgWso4l5A4B9Hk+1V2Haz7UjQ3gM3SWoNQYk7QqKyKn7bJKHUUNKY
qvvv/rmGx9hkPCwbGQnoFUwaMypY6UcokVrww30sJy6zWyHsYFO2M7sze4EGUsXAmK+7rqZqcgxK
dg5XkNloUwKqsTIRHAtSeSNchmxFjpIZeYjAP3lKnG4g30V3VDAfLUCyyDt58eYkGozrpgmbdx5z
nivHTCnXgh31oJolzUNFBuCe945sdoKqwKpU1keQd1GmvO2IvpvSgMU27dWWRiqnxYa6o8b1vzcb
HEWBsDhgVccPRL6yvWGZ977D7d6tfB6KJfsYr00+7s7mCkbyHpr++1k13CeiGKNdtdlhP2tybOVk
oVfkKkfGkg37/YFVw+YoJZ5XFBUR1RF5XPkEjbp0qcm3vtjneTm/DYefZmzp2osDyZ1pcZ90DZja
0cdHbcRgg+0Yk/8mtCc5v8IEhJAc4HIev7nS9sdjZP+ITk3L2JyTXQ6NewOR0Ek7Xdt9QbQi84lW
WV4tjjRRf3idXsT2vDUCbu9KyjK8/27rwIMCEVlTsqztsqwsjiIIAPNaYzhyIzcbnm1xUJmFKFOe
1vvCI8yXTHecQ8g02dmb8fxhAlrtDN6CVDnoEwbxVNM4mgtpvo9kHx8GNiZqQ/G7x4qLnRTHDYR1
vQIVDa79bVS7EYVpZbDuiMXRCOYiLvxdGrzozfGUR6BjwJ+/cEiwvPsp6EwjpJrFnt92Sqw0h16R
o5LA8xYBemtYabXypFcYkggpQMS2JqQvLHf0BEZl7L9tKMI4H5XP+hbA7vXc6gjB+qm+wmnYUmV2
8sE0BDCo/YSZTYY+sa6NmUbc3sZH8BiePogNeI7elupvjc34/A46FJ2+WFITIv+NNmV4zTKkB10U
yv2Jn2lhOtubzF4UP9BPyfJOMNfvy6hR7Eqc/y6Z/hU20maPZm04jtwYIh82aakSdeccDe9w6CmC
5qoFowgNOCIH72BNHezfUbGWmk5kcsVOwqcvW60y3kRhL3LCm9b156oMqvT+R/FM6iXfDOOfMniz
BUblcFA6A8Yhtm75MscORMS5ofFBhKJ07U5uw98euCf8rP3GqzWo1qEsOgtoXzmt17MajgLiKqQ/
NUOTIA0eW4b+DXSapR88eHzWwbexBI1v+Act/65Jn5lqc/BYfIfpmsqDSKTyPpeMbu9bztvmEBMq
ow3yeTbRGKUQZbfLn4MG2UeLynCKx7dwMxUxIBupTUASNpvzEQt0XQHFmch69xNkxtHcdKq2cXhY
aLthmEiSxzBUZ+dw7hJV5Pd0PKLBlb6cqVwb+55C3Ud8e4ijxSUBs5aNsPW1c3rKXWdNu3EjO+1F
UaeF5dv4qya0dOLP7FR3PM/81oTC/JAlElTF3m4/+ciIPpkzzY9ehOjK2Q9yUUXLdZDMAuGkq2Mb
zhXYfQkalgjlYBKMx0lRSZcd/FmfB5iEmpuJ8RhmqFPoYddtpMO3M6ki9X7MyDLpxfJUnf4aOgRR
HhmEaIWBcSJek8PRTnBVafWBJPMGRllq/szB9QAZabNObDsr03LfpSnREE3GdLh3OJ4Vr2TT9JgE
J2bjZrTZV4SflyvzTZ9coNawNuOubYJ34XaoLB5T1vPJcXUYCya7o7PfmxY/QQE5YqAo8PvCOQ5y
9/wf5T9NpZtN0pt2GjkspJYRrVYuYhFU6DNsjNTNrF89dFKfNsHXR/7yv1GuQ5jgVTe7PmdklDmu
ag3HoZHl/kFJZX4uUH8ABQ7OG9Kf4c3IkPZW9E/DU4RPd2nN6oyvaHX0JHv4AZxmspZ/vp0A0SYs
0EtvfAfyDw1IuSYxj0dfWX3jThdv5F30zaZUJ4Gpj+5FhMql/7X1wZffUbTiFQkg5wF65tbc1GSv
hPqLbxs4U8n843OCNNskLzX2V4i6+iFvs+jOvNjcg0VhyoKJ0kPNtEuKXwo/7w8LdqqsUA8wfAwq
Pk6t5Va6EYj5cyFZ6EsGPKFuS5Mxd/4in1lwwC6K7zJxRF0jxN8UpbvRDyhJQVSpYM5HvdzZF1H3
3qhf9jiYlxUxChmL9SAI7ntktcGean6Od9L0P84Wvk65qR9yy2yBosjapeGtZ1WKR73hOzB/2l7/
QyVXsJydl4OSPfYFpJ8mZnNUWdJCp4nLUgZ5E/aTQ5upXuBQBI7t5GGTThXxaCEqmIWYZBEr+SmQ
rQkLWT0lDvZZHIoUY1z5SmEhN1oRL1XymQ/pNZkkIUr0hd44qegdn6er9/+BXTxr4uksycPwR7hW
6y5ZNp1+TiPe1Cf9kIjcCmt7z3chGGI7H5wcpd5l0Dkqx5Jmoh5TeNU+FqyIfexH8AgVGtTLI/Qs
dTB01DuNQTe+zEJqfHLcybh74jo/eCoIwvnxXzv1CIWJfBeVb1RB+QB3KyQiq31v8JOCQsAT62XV
v+7W2OnGT3OOOX4+h5dueHV2QAKk3PyoBXygs2SnjvQtWNOK+EDIsMtI63K2IQ340RVo0NJ5N6/D
OfhYMRTFYt+yx1j3VwhC3Zbzeju4t/8Fg6qALH3qUEDHcn8P3NRCACWJpJPPpTO/bjPOYbuEGb1E
gES3+i4JRjirwyVEa33hosjAtggqSoAAmg1LcdBBdxo3bjOQ6oXPVs1p4d+GWEqIJsgW6DEARN5b
jiJgggraHXdD97YDFB8+wT4leZgxn1879E4xt2vWEfSBy+s+rlYFX5n/g1AYCI9NpIjl8v0j197+
nSAs73q0Y8JjR2Q/eg0/HYoLHbLdXf4mf90tynCgNCQszUJwYd8g/hx1VvhFidlNZ4I3R7G4bsWQ
HuOgXGqXTpItJvrf2vvXdaDrbM/Q7CLdVNm+T/dIIotkeFrwUOZeJX0RWPaTwOTiyu51+4Rb9AnO
JRYW4XUGV3Ul3/1o8hEH6anvNiCzxMi5QoN+QS8mLPbJrdHqUgSfAfoEPONPktxsIgjDXFn/Kh3o
WFGWyPX5hkAV41kQEnHqWkjo0FjBwGH7Gw64jr9YdAMSHRv2leBuWZUJ1Jl6PFXWs2iH2+ejU/63
kg+lhwzOsCCC3YWNQQum7Snf2Xu96rQrbCWCpnYaaHYooiwHCTGk6d3aCtezErbMlJPV0zDV4eHP
AOAC+Iny0y9/CmQY0fMaBdAUIDkvXGOQPevA8f6APAQElIemNtdqTWyVo8IpX6Xc3zLM4VI5ztWT
JD8kgg/Sr8X2Dau1l8nu8izAi3oDrhoUSEdDx+OssfcXHCIi6BfG/ViBl6nvLqdbb4FJPgVRvBKu
K4c75xh5e9im/eeeIwrxG2fjLRkNUfYvvDG8mixlr/2phL/xHhqBuKF03MIrs4L5Iqd7NjG9+D+L
UkZYHv9pfp+OgSYwNmnLkpijFVsh1TH+LCUAXEOjK5zwzdSqwxIR6EiEgQLNaIY97jcq5SUYP7LO
38s/EOqUxgNyHXR7rupgs/v1U12XJyXJZ/d+O4kogS5Xn9O/q1cxqJF1B1XjYsQrB+MVjEH3BSWL
nXmU8aRkjQb7aU21YrYFN9o4EgJDEVO65Lq5kjcBBDGIzL3sMXmw3udDSP9609x+l0vwHAzi8Lco
2jLlsYhboijMzlNhH5LMgsrNC5h8JFONhPsg/YgF8bIBziEDekPLG52pnqZiVZkMGtUVL3E5MAgs
LbyRriYNw5PFFaV3bkZByB/768+uIB5Ca60xJ2+8ZPkDk63UOxqJKdZURpxESGYG8EayJ6lLnKyy
m56jiJ8E7gnMAAl9h7cSJfQgP253CkEa3DYTcm0cVXmNsofTqymUqIUUk3vL0i5SpuX5Xd8dv8SA
zxq4OmyzQfPcdyt8Wtv4osYyFW9ZeY186a6IY6mraJ2OJqoKYYyZnltebvsvadg4qH3L2cxYulhp
SoEM9OxcMXIfZfsO4z2VLRCx6eABOTlNowPDbHdtyC8LFiovGc0ZFVHtH6sg3bbIZH6oesGXeYpK
Ne0kPdOPTLJTlmneGT97oCnt4hnRjrpcmKltMTeb/BV4PJrrhUgYzK5mEK17X0sWhKM20+aaybvf
Okk2u7Zb7NYUYEN02tD3Zi2ctVs9vYGVobUssQXeNHscRnBoyL9IxgUCfade0pUJ0WBzH6Tfp/uI
LfGR8q5o6Vdbl584mqzUTWbIGnAiYcRNs2YsMP4IZ8g88zKMVGMmqmrvN4x6Bq170VLwGarLmOAg
/HkWFKhpgh/6gtGugwydRC8Ql+6/uecA/IcCDhVybAzkrnF74J8RKExYUzPonRc59RMUgYSr+Ks/
Fup7ujfXMsQCGl0tZXJgvq4YOXdU/przxzhiz4OXX/VQypHNyuye3WARJoIcl4kZ25WF4ok+S3J0
rxdiVDrm9+7N+yBUVxaJOAXwuAg9kTbm/O7hqMaHrYdLtbxcHUHOrZck6kfK8EB6tjl6JkjjCbbE
cM7W0YWgLBzVjoRDVpdhowz8nbdeTdMJWhqv2MqqekspQNhs5cxJBzU1psmCCA7WZHDno878EBOJ
L6eQ+t2RpwUy+sQ4TWhQDEBr523IA6JCS7RR4aE8+/4N+ZX5JUzP6JZMyVF42X9IvXfoQNwUqHAd
+6A+Khg5btp5Deyp3zB/wFmKh72xtAgfpKJsHjDXSodqa2yrkx3A8VPZsBVWOuUo24/0Y4hHQHqF
vxm3Qw95POELWYNu2oOjmakPflPhD5F831cAAdPmybbFcnSppMd586V/k6FTivMYnSO4xytqiYEN
5Ev82qG531AJ1uObZk4B0MzAgu5CjVznbEpmOsSaCmhReF6MWtcop7bHlvGI4lcll5ruOoFsIdR+
GHfZYSlzl7zz38Re5X4Zi2omAxBGsEshSTPWA7Os8F/W9Ig7NRz29c/4EMt8xRN9fJCl7HNSOHvG
NQpqRAdh0tLhV6eGTQMqGieplgRF23h5zBQ4ZNrosTEbPWniQOUR3mGL63wO71Fo7CUTlxvkr/XC
zzwYuGaLVcNrG5iWzm60UpfGo5h4i06fhqTbl0HvvgKJ/sY/EkuTrn1/S6MWp1keF4blePZg2SfG
TIzmkiur71/9tV3QAUbOCNop3PXYDagkK3tlxXP1LBtEMdZ9EPSQBMJ1YIE4JTXSbU0jzRIB74EK
k/qiJJHXwEyGWtu+bDwCrMS3qVZSlf5GuLnXqgIWjG3ENbPcHrHMU7PRYXaJtPw46BOtU/R5LbBz
mjdz0jAbVpZs3qH9onpt2YyKI4jFtDSQS8MDtSG9ju8uO75bepyvjzfF32AYlg2+w09VJUxbjzFh
+AZIaNuNTYBuM+U67q1nMAEhllujYvofMIXssJrsyWvp5CTlUiJ6qQbyw/QkKV2gPQaQlcpUQrUG
dqpUP6XX6xRgRfEIXOjO0NcfOT5ecgtPUk6g6/bXqGQI3ft93NHMkw9zI1Tdm/IcUF5yUJJ+zLEE
azSHLVUpqloyqv8ot/CZTkcjAnL7k/Co9PoIn+CWnaBOLaoDNuWMoxJvoGURdN9kaPosrPYoWFuW
HWzJDTEYiM4R6mpe6Knhk/U2fh+byel/hxbEo6+bx3trS/fcOkNZY1BBe7BKrw5s1aTAewP0DUWf
xmRRgcx7Orsb38skU6ERVERj/pwIvvnnFNm29qWLP5c2fzdxEGhZ/BzXJpm/34iudPcWG3NmSvO1
64LRWBOFvorj0LARrkDjlQfJWHBuuMxFk8el3jNL8dZ1zSKSX9wEjtvmvOSoRpMbCUSDMpOlA7eu
8dLpmC2dm/lGHos/B8VxI3J/SKufTIAqyLJktL7jPnW+Za22cjmom0R+8ODs+ZnlJHpguxeMVmxb
QKH33Wqz+cmgpF+RsilaYIcQumAdoiwSQzE1kK1Xw/KWFJkEHWOj51HbxqPE3EX85NSLKcDcrApG
3vvCuj/OKciIlKJoxhmDvLxuGOcK4K9jHFWXOTEpphCmTs5fPKyhJXHyIya/0/Nmeh44vPPYQXXg
U812YODza4w7dizNajXcRLDzys0K7/uvxl6ysMEQi+yt3FW13wWvrpliamozzVxzgDNbxcObrPJA
Dc8DHr5kTx2E3dFwT1Xtbwo/48OqWs965I7TwpbEHhKDkYv/Ts3koaY8bNRCSnNZSjSE+eSaaenq
/TB2bzELdY8g27s10QX9aPaHd3KOZn3LGdjNYn4iLwmKhKJjYKuam4G2DFeCQf1qQ2qsnBUHV/OC
ibAO+66mFPqSxiJ6iuVupK9vbtUsffY1oRykCFVmNeQ564iDHULzbVTVLCAFwHLZdj5wY12+UqRN
IO6FvSHzYx9m/PExBarX8S//8irvPNoULAY8MtKHGMfqJq/pzKTKWXXhEtgrKqNjzmvXIcsI4iCM
wqgPg/YGc+Bx0Ty1E2M7pZKge2uUzaQnXXIKo4T4irkPN3sWHeMfG5tTAeOQOp+IzfIYN2Gcwv8n
DKQv2zCjweHPUnd4VBXaQRjOab6XZzaOmYGviXrNdTvbpGTI/YqTxmxJO1Qx852I13vqm0umFDhr
pPYFAbpo56YClSZ6n1r18Q0A+NyA6imUm9KJRo8Sya3yinNHrokH+L/aEY7ug+ULtoDok5cGL+ib
oeYLj1CbxJ3KeVUQYAbiEHGfg2Ut30dhZS5vJ7T3Rk77qV321ortmJMGk3/HcMKU/6Kk8t5NfxRl
KsOY76otYsuPFQG86bebn5FUwrJHEdhUEeIRU7HEW/n/tSU1eJI/FFjKX3azykY+y2/CV6dWbZER
XaHiQFEYvQ2IDDJgm7UMeQmUFjewdIKKdV4d3wiVLVSo3rF7z1SfTkxoegCC1ZaY/04emMFbQx6B
5Wazw73bhG+MHYhCDc15Qi4BqOA0OZ5tQO4HizkfNUGmSRbIS07E1opVdr1a0qkR3Vsw5R/HBw/s
hPVOc0IrwW6ECONvMWfypAudao6u3tMlaBpWWhm6U2ji/eS9dsfC9esjIZMREvqGirdGS2fINpqk
9okCNqYMSgZNTyhswlq7WaxqK/QdIYE0SqDgHgFZDVaIFJji180+rw16+Zc4DwIszkkWYSsqhIyW
d7cotIA0RPkC2Z7UDHA5/NMBjbh+aXwjCfCZJ53bPcMR5zUMbYyVBDZK5j2aFjHr2T5rLlwz+M5g
rb/GQkr63snHhBnpHPQ85+AATVcXgaZyPlzWNjB9/yMIvl5XbEpYkGx9ovg1vcsez/qSWEkWr6H8
9HnmkFSPRILcSZFJgknK47hVf3q4R3IWuq+IRQUULEdkPiYNlLxaqoLwh4sxrbydMTVDFTjVudDY
egpsApOSx4Kh2qRk7N8YeGhZorSAZUybFUcYdmee2iks97szWKm+S0GJgUb+on1rLyqKfQ1JlixC
pn2ictLcLC7pjLDNAmp9+VMAsyxNnG0ha7q+2X1RAGavjsUzGWaZhb+mJnoYiL16aTM9D3XgiarP
ZU/VPTrrm+p5q5VSifw2gE6sUc88xEfKC5mwy1+SFr1ygrqh5dbi1CaWsTnFXSRDAp137G+ovhew
LzpGGP+LgUZ6aKC7SMxCV9euFrhdVip+F/ieBsoFpmkMYFJUkXJRgfj1q87MmS8HQsoFXN/G1Yxb
6T0tQXXFTLqQqe9GlXV1I4TMQ9pe1qA5h2Y1JQwLw9gDJVDzS4lrqp8XNvINn8I/F5y0dPyO1Jy/
tfCxMxKXtmTtYoodlwC+8A4RHywUTUmJ+iLCjtXS+XYvam3ORVBYKnKfNXx1WsigTY1QTr0JIuL1
dVW2/ETiT/JG/9HmRJ3BN0JesstoNkO+dGa58JoYWX7TUaEqzwEhgOFVxxRuWeXcfUZkk68fA869
6R28uaHqWj8SQa34yksHn6n4bbpBxGZptMDyawZmKIizYPyUdRs16bsccCU2vI3C1YLcChTNuMnC
mnrCo+ChogLM3T1lpO24JPQyROH/VSzsJAKaqPlLpflrhX6iQ/gLmaRPr9ZyyoboFJ/skxY7Ackm
t3FHxYXaf1M74iggx6JcaeyidayFHr2Rtb921bviT8J3jvodSp1xOZVOtOvsxu7DekBT07Wrp84l
miavb1p8uJy+Sw4oatLwI4/Tsx9JQJeAhyCn66yQgJlSWQcfks9/WRvC8yYCXDm5j6wYK5yWqCtq
EwzpolsZmlzXwqofYkq29+AOJ1xJbTx5LSZ/0T285RPBlCSJLDdC/f1ivmv3JJ5v8AgZhZVkcstM
GdVp5WLUhYdeOmCEkIf5q5vWdDIFkthmJIyLt8i3sLAfgw0EfH1n8FVvOwrqYosazXyjpDd+fkrJ
zNL8KVEDiEIqI7rZk+p60VykwWaHUR/smWI9r/AKxaH5WO61J29fhIHJ/5UKivL2x1XOz2lwh7dH
8YFxmzD7LZi0Fr1sisv3mtd/AK8B4lxQ+zN2QFtVs8Ybwu6MZXCBS/UVrfqAbW/CcCpa5mi2smyO
uxc24TixRzg5T6mz0x2V6vuo20E1BgIFF6JrSQrUj6TJC0WRv2j7R8L8fL7xU5PRYU2DNTscjiju
6pbwSc8XO2Ge9T2VpKQKpDji4QA3wxJf2eSbDw/95M04Mdx9/bJLzrWkiuvwAyc+m+q9GKfXuixQ
QUl5jrF4AOzD2/2nHrlgSj2bVcPGW10F0I5+cxiSYTLoPxzLBUFFSgn9Bny/aws8XpSfzIXJ+ZNb
/TvEAp4ZeSkM6NWGzveKaYMhETL6RWdklU1+QbLBmhbiQWHmFOW5sgjQM2os1BE2LE7rH+mPxjxF
J3hPs+pwD7SFEwF1Lm0eVgW5eCGjovfLK7fsSDAaImilhWz0u9yW2BiVjd0KksaMhuOHQ8O/Ikn0
qS5fhg5guLV9EFOn23Moc9EfV6W84xRBIsnotw/uKvBySjVF281djh1RTcsxopxntsheP+5qJgwp
e8gn9q9RkjvN+jsPXM4lukpKJUxlnCCj8ne4SW2yXhXTK5y22YkfGFuKANKwWk3KcbuAfhkvfpbv
s8ZrlvJ7UfgDgdxE+VI+0jRNiUbuPEZoxklpexG2IlLA4EOMwv/EF9q0f+6LBgtCpjRpr9JoBUYt
WfD7/uLgLRHvJW9aYJ5yTThTmhiuBDytIMAg5r6UMquo3Bpr+u56gEnvYR0Ncf8zkUc9fJJIJ3xr
c2HqVdhIelv5r8oOMb5U3vsY3H7saGvwSyFqtvDBpONUPRn4LMJFMhCz1qEvRHI/rbM4m2tvpRIn
1qIMBJ3hOLC920rnKOjdRd/egaXR9nG3TNgzEBcnOmDOcFcD//eS7fwlgwj7SW/Tqtm2qvuLNbPd
Xjqv3VKjQOEEp7gdkV1ElmmGtMQL4o0NINqwCqbfLEpSuO7ToLd48q6YnjdMeh3bzicV4Gqx2JNz
8PDO1rjbu5s7ejd3cHwBS0WX4JvoROOKiesAN9aTF2SJnzgpwo+TIh1P7qLbIedRLxj/faLmXwKV
SkCPI9B/MAssDtnY0qOpwpIYOGfGRRtKd2vtVewZqHU4Skjnn9UDarpISFqCFZG8zGubfDu/i6cX
olADu3ShIfBI4MgsjBiryHAr4N+Q5sQduwSsOOVZ+1DdKxKkIpvHFLbW1E3BcGoCgksl23RfQK5P
5L0Ti+0lbdbgCa2UGHyKFqDAgzIADm76J45a5w8jzd/Bo56rU87e/a16F1OIiX/KN8UH/XE2uzk6
M7Y+CxqaFpd0kw1rxgcmtw5JzpFi8RM3/UodbsNSWedKCjCoI5Oy1A0NaoPSzcoswYjYJXkTp4Cx
6S2QPHU7ABAtPNLkLmdXv7fdF/xavLcxXQcGt5J6+YlA+lQac7QYS+zqm5oNfroPwcv/VThKDSnW
3YrLcjky/hNm4vvHEY9s/ig0yRZ4WLYUPTVxbi97BOt6mWNkZ6YeooSeIRoAeldI1s2AcKtFVgMa
q34SV92fxlQiuRVN/djr/g04byzEhhojZo2bh++mjtVs8hrus6whaFge59O7wm5bivb93KqAYUqP
+Af6zTAGmCfocEor5hmtLNq4lsmeZZX03jkqaNUlOoDMjw7oDnIrvVBG6FlstLmfyoDm+raD/TYj
IoDYBY6rxMOF01tmGSuXg4UIO2bZFyrBUGizBSFUP/NaAE/Gz/681jUPqh32TZEegYmK5KeCW5ku
I3v6uk65Vkw3B38h78X6y0v7ijvpgGgjXODGEnSzfha7z/Qsvu5Z7m+IexOlO/DdThIZxsrO+ZKe
6JEwacgbhpmCsrtoGxVVb4pX8yMinXn2HWzk6vXZzUIYLxVWWXb0vte8ozklJe/LdEY55gshTObT
wXd89n55SRW2KFge6yV/6PBU348E4WT0lu97JA1ROWNQ0/hKuZzV+wB94EGvwyWISK/HeB+d54RK
7WRHztOabHq/7XlvyPjZRIUtgAvjq/YAhhiExdxf63zEJ+v+tMwf/0cQw94G3tIo2s0zmVGs2AcC
di4LtJcZlVFTiDr+pCylBqaPcWl31Nf7E8ZsQT1Z4bGHnxs6Eg7NJ72GiR9JgrbcFvVIseHb58l9
g+gM1wigyep5cniC2Xg8+G9+xYT1wGaZUfFmHkm2ud8DSNtMdKJzyTNEFn0M9RgiysNPuugcZJKg
IITR2QFfohx6A082zKOBFJlSO5doSIVk3wygCH5AB3VJnZZnc/dwoN5Kce47QtoqsY7InleOCp4y
LwYaB7AIgEsg0pxuUIPGWZ3BF9t1/b0EupbF5b0WUD07qNVz3zDt3mEalz7QoBg8wkvAmtxX+rL+
xsrj5fC9pgvHHFLYmCBQB+xRuPK9+OUPag5a27N0J7P4PWoz+9JYiqLu5V1IvT32YhV9F5qunV7g
BFOo6fITS3GigubC7MOfQRT4e2SUdwEDnXh+006PcFL8L9TDhqsoE1+AnEdfBTFD8vae2AUD1s75
HduCPLntct8mePlNcCnW9CSuYwESPy6mCHDuhgBUdTWuY1izxhRvvNItpYzz2liilAqksgB8fJLH
hqpdZPIwtEfSzwhQ8XSODW2vl5LajPW0xfqoznfcOd2cH6x2AUmIJHn5WiSayD/c2qBoD/blvkrL
4D9abtATYcNuftbcWLj3jEstCp0phJIKbHTUB2baDosup0Z4U7wuQRmMug0ieSfjfdv4djt/YrqM
LoLECEeJpmdHaSfQ6516f6o8LjAcAV4kkkBj6O7TDmYBud4ZC2p4eYIjSs1kStt3wCioR2koJg4U
+ySdj2xOmRqKwGlfq1AJWrTq5O6EBMPHB/WYXyCMmW6eMyXI3ErqJCuPjj/JJltyhk2roqWX+WhJ
fxPDl1J22IoVWyWu/kCHikx5JoKf+VMoigN7ABchSXMIxtcirw3gQ8VoMLUbveZYHuO45C0DLM+O
iAG0SFWJZsZRKuuqE/cFRYgPjXm9nqoI0OY9ktcYImkGDuN+wD4j0VA7IJGAc5YuJ4M5zPzqvDod
pwqD+wBQgiBZEQNIzO0kb5CAOKkG2or5p2kBMGDgXUIC1lTK9uzxASKviyK3zKZwHHRuLAtpqF/r
3Srahio703/DonmXi4gzEn/dt/jmdzH3BAyCsT6FvQAv4DzzX4pl4zqWt+J91mWiA8mROM7fOcAb
FIP/5gvq30XzUDRzlIMFrxpzzy+22+sCwlo0BkMPA2fTkmDvM6n2nf9iZCpJVhzy/iB/ObFK04Tv
N2gPB7kALjuLxnwJTgDrJ5sZ5EzZtUnf2ouCERdG8v+dsliRG4c8X1sJ1C165hY6tHM2xjKLDj7I
TBoj6eZkXrkop8UUIVP8XEnwUOFiuVbp1aUweZaVNBPwFKti2kwnaUU3wTnzzue3k1NOJqrZb/No
xRhuYkivMg1ibITyzSz4JN1ka5/IiFKSGLNWDEEY+84fqdrgs4MoFzlzB++jEZtrbfuh3i08tCgB
V5f2DdDee+G0f/73M7tzkuwSEyQqc48/5fz1Llylic8jkvh8EpVPTqFAgIZMv4yvW847j4CxR5Il
PoZGBgNwD/upG6yvyyvrmvNYZ27FjdRT7moliUia/Fs/nJifldSN19kFMHdkxz+dmjHaO2r3piwU
YbZeOGEt7wLPTXJS3QIMcNgGR8691Y1v4K+4UExGXqW0taJyfwVyWfLaxn8bZ5I6kes9MnjryNlO
ThcwqyDQdVo8rj9ctod3BGfTPBjTgOE2mhiS61vNW3Kfo2AyYVRNSFFeBGRae/jqWeRLfvHnTqcP
RPRNkqUPhC+dil4y8pjQ9Nhh3lxN1vVB9rucedMcc2i+7OAgR2Zx3eQ7dwxSBrW3874SJ/62IE1j
JzUhF1AL80TU0LFrl99rQBAkOmkhsS1dtKkr01/CrN4bFQPXQa9ZJs4sMln706+QaBm5L7mLDUU8
k/zNlktDrIWPskJWV7lZZgDKZ6QKAUN3hGVTTSlsfZ6FPOZJL6Y2auOgD9iLurPrYCq8qG3lBULz
WOIn2u34Khcc8YNI9VX8j2OjPByvqXCuw/ufjq2ZEA6TZdn7PESuWXVNLVy+KKCEx5LZhTOhtF5N
Nvo3S+tRO/jwl7Q4YM4Ux1jPvuXA6gTiywc1h7/06cZb4e2OSJu+VO8ZJL0d9DrLOQ3uB2PZfRPd
FCw04i6MaG+N33n7NKMPSTJ8nWa/YOia+7Zsw72Z/JRZWohqVgzqbCsQ9MS/49WnJLdOQuvGdRES
DXnUk9CKcmnKsmPjkXjVfUF5Si85u1KCeIrNmPDOsBZ8obqlPPJ1qD73Qtt/Ysp04daUSUiyP0tE
5m/XrnUhHO/b0ZQTB0Pd/ErWd/UIz/bPjVERtyYI5f80yPBEjJ2QoHUUcfZjKRqUc79keG1KfFSn
dJkDy8ltPxqHZy+cd9SEN+IPoqlkQpaHwORJMr+DKfkhR93HyJ/dSc0sUyW4vOeQKRITMTnHaepF
FAFeLJkwtAweCF2ybH8a8+eg259r6mLy/cvRfnDmZn0pi6hy1lzpvEel+ziU4rrZawmugt0LUx1f
hSWDTrcyzyJqSYMx0xJot3urbswGeVNTM9ZpjkU9yExbULBQq/l95QlM7F4XZWgQhgAgC+BSOCvH
yod8kgJBEAMUPHwNVZzmz27nGt+ZWpcsdtB9H3kCFYIeolHf/CBwk0LKS+1mryzZN5Br8t+HKjaX
8ztcR9vUpuMcIblOKKv1RLsExmPPhdQNYyciEIiz83htizV3VYb1wsKdeW35NU0L9c7JqDVDMuie
FpjMrMLAJDUXOfbxWjIa/j67L86+hHImOD5cFb3jj/G0jp5nMLeRXtR9DjPhtj24NIInAkyUDUCo
MAbFghQOiPfKL4Mi4Y+bI0OqzYj6zCL6JCod5EX2UV6MI+0BEMWOQWp486YzZs5lOiP88cRgShky
7SDxzS5tYM+69u7CrMpdobaTwcm+o/Wc5vTD6+Bp6Gi7VUZuBRv5W0U5NvnjmCrCirAkq6AdQn1i
q8BCygeXLWiXMpwRWHLoFRcvffrK6pFmY+E82rF6GfYhTZr9qnUSIE4gxwjuWbHCzLGP49cLdKAD
iZkkf6B/+Z6Hae48x+aoafhwupesRbvdgTdtnwkrAWlbQMUMB46Z7OpMnxe85VoAsICZgnRJS+3J
EoSKerh6Nby4rcS6r7Eo7PodEevD5bBtP2/lQNglLWsbLI0B9ENbksd8z9UP7Z/XrWcqWbD1HiWq
HhuLkWhr7QPrD7xrme7ZFYEk4Orj6d+VlOdQXAEUql2FYWAv4CUuWsi1/f230Ix46VbzRdu3nqWZ
QrCMVH5m73D50Foy2SWzG0V6or1jpj9L3vIqI0BAQ/oQwKSljY4qPqMlYGVaJQy1YzGqwRtGOry/
AtHTebq6qmfNElNJiPInOhiu9mV+I8X5DjnSxOAFY12XaFRaDpABc4WRDRRZOWkKBkMXac4VCDb5
2OXnA71feYLRCpPR6QarP6KZDSjfgI/H9csvxUMA9RK0/bBb19OjUeCvry4Fw94gvO9HxgXHJP9A
wmpyv5n5Ce6k1ketfpECrjFvKMFjowZZKDFbEeTVDH1wFwPMUtyvEfo6Qr++dJT6V6L8ei6ULbMU
HIuJSq+87GDDoRLQ2EiWuMleub1WtBv6P+HuXSKIvI4Y33cy0GT1zBHrk7rBoBOIIrGM56uCcrQf
6+cj16ea7JcewIDgaFW5v7rCl3KM1V8/aMq9DV27PqmacxDVCeBolVArZaKJk/xP6AsyNRMtBDGq
I3yee19Ucla0Pn45vnaTz7JD9cCqwBIwpKI5yerIC/7sGvCxphacTPuRbnRMBufk8l7QLjojwd0U
FHbs1zRa0FEdADDLBbr+A3jwZQXKGlW0lpg+egvS2/xjaocHXcQGN5n5fBI/dobUCMzGnmXxgcko
mdzFKie+zu15iG+pQrrVVu1fTTDrsVx0nraEvrP2hpEUkVl8kU/RAgPAc8xxCuO6Z4iyqv0fIWlq
ZnutgXSBecyO3ycD4lhfd84K81eOwToJmP70U1rQ+wAmBhbZzNq9cE/r0HOxTiPBvJouSrWiXB68
56J88341wg1u0eJsKJPWV2D1RTurusqrjOKjnHWvhebcEIryoRwfzIvKqD5Kk3S9aFqV0CMZC/6H
lDcWOzL4lXrh0pEaaCKxyvUaPeGPN8u3FjcTAI282JuumtLVhhPwu0VFB2uzPxqScRxoYLOCWCtX
SHdN7mMQd932/5ExcFPDFNq8Sc+1p34SHMbdfgPgiCzQC/p3kFLBQoU/wVYBSdXCuOy/ahkTmVMr
49xj0ENsJM+nFWDMbYV+wxDWHemomwwHxdYtDSi+XYplemAb8zNttvJtqA/qTMKLn5l78Oq84XNL
VW0mL7ZpPVWmidTRdnin33w4XTL/uH3+XfwYutz7Dbi0weVHd5WoHZqeEZvJDPBoCd5uj0Zvlvrh
sSH5WfXgrHX0CTbUv5FplEmwW/Fz4zz0/TqQj2rUzAwxb2nMIujg0Odkx+4mAo3X9dFpqryC3Bv8
MQMKw3S5AY7tuOSE4FuCFxKMPVCc/FNy2F9zjdFz0REV9ymnh0uAGoiPtijQX+tUpprYSjOB1XBU
gO4aRAH2OAKwnXa2VWSlzBRJL7pQNoa7rfYLIj8n+LTTWtofRyBqJdRRjKiG3bgzLxHAUCidNKST
LZbAjSOjojr9bn7p1PmTAO9ex3qXCp2GAEsR7i7DlocDCgYXMtEIv73DJwmIq9U2LKaC4jQDOtaD
82cbAwpxzXVTrEgQZjeBkLoxMxMwT3FkJXLosxqnR9SLxxL15qmTUh/jh48yskdEli5VXMLwad9Q
KRyr0ybi7MqOK7pNbGJQ4BhZKOyq+DxqmFd8NQPJlir4Pi9rDGZqyw0KXeaWELTjxo0QDaZMQAMg
moWY87iOHA8oYCgwBYUvZKSO9q/I2UAAl5glpE8kxpxL6cj9oitpSkn28tGUapgT9XgAhC07URxh
m+r3RPeqrPIfFnvjweZow1k6DKW7Rnj6jDMviTsj9ImfZSmOzkZ+X8kmdAHK0jLwpuPgjaq6/TeY
UrWoVcgSsKeIG9ti6ev53fO66yy/SZ2e7fa3WroiXM/J7m3RtbweZA5PgaBeSdBgCOGyHRKX7OrO
IEnFPSdRUOfyL5zERmGRyEHaC0bicBT13Qa1GoNUb9x/00U/mpp8ggkYnIkvEhyQCDamxIG+SzoK
PFW46rG9y1GM+YszCUsu/BBiZwXA8KK/qEjhoKnOG61wB/5N5l5pzRKIfcHjZpgvLrnlXjrufkEc
+mP7Zs1FJ8tEmgkvPA7Vn3BvQBO6c/nTVtTjs+cmynzKNNXo4fqI+kEZJlNVHlsw7W2Q7pD29nfu
7WQptMeQ9vYyMIskhAnDS3MXR+ZBjaiDfvvIV4wAeuhv9JssOW1A26a1hlJyanVKmzGftfC1oJoz
9lhYXiagv7xeo4r3DimivsbaPjQP/dC5ZHym65OtWP5YwpIGBv5ZVfi0j1fd2bF8b3MwefxfKu6C
T924ukMqtoSOoxPinM8eLBxRNlytRB5tN5vkFaU1z7VCYBWbg6re1lSFzwhoB4iXEc3hPzFRS0+y
l1anap8Soo5BkojLE0i13qhYEWwfFOCDBbYBh2QLIAleGzlzllieCnbXi5CyCG8rrfUKP8eyhH/C
O5VxuaWbOOHHcdguBeDGa48ZfdPY/U5OCQ1P6BwSZOBFhr/ZBHhL6H/DxEgStbNY36HAjif5gSrP
/VPkUB5snQRHGLBWa8yHfou90TEVb5IzdXMvLuMaX05IKY4r0qK3cJYtX6S915M/pxpgxlAeXNf+
bB5ghuIlaZzfh392PC3hO6BjGMZ+YvU3W+GmmdhrmJF70i+58vLN77IUYt6PDw7Uu2tQq6JRcCQb
Hotfiq9FPEApNPKV4r4dVNRGegxfoiBCrhGBoXtZ9M6qDQcfR4fywS5ZJxeltNG8ag8Y35704EuU
nEXspM/40sj2d6RfwOfRAyVJZ9gqEU8THS5eFozmFUuCD2ExWjLdDGukwzstQyllQE4JqAoHd4XM
z9oEgdIwDpL58LV36OzNI0Os9Dbz1W/6l39u63J67hQl/VZD668otuYgmIzlH7gjNX6/0f3J3XDn
meNw3EJIFUyXB3s3ZM0o8WBWsqGQQkzcUhaWdYpLB5RtOi15QWJs5JtDcXJa0NDIw4FswAFJ07nZ
ofrcDK7P8m80GtdNrY5PYii+Q1KaGLlKkXwdVKPCZ3/8Sp79KV89by/sCCDMS4Oaxx1LL2FBumYW
pUwTQPfAcI25nYb9YYhFronAq8ZulBJ0+Buz3xgHi6IEaRqNFSvJ2RFqzQOZRYKL/N6LEpNns+gE
U4rPz5TQyOP1OYrKAp4GItxICNM/9Fu3SRf/pqipBowzXRfOeEdjIpM/SGiwx+2YFQOkHiDUwTXu
1mtdatQPmjBKKaQqf3kDNE5WhGF/X8/LdUh43tf+B0hNvRirSuNCXYA7L9Atq7IYslXRbuqjO7PW
XaRSO1+ayv3TBBve8nwtGXJNaactDba3JF4CLVOK5idtYaQ48Ci9EVwzem4R/YFWi//klId5uQ6V
GfOhYP3y0e8ak/GikU+zHxda3cSIFkya7rYRrNk2BmK1YfF8MEiDSMkDrMgarsGTSxx7gCtGW+st
x86rfG1mIw0BJ105A5+Zh8sZJTaPUKkuvcoGqUP+8d1Z8cxlRVzxoPOcgAAMxvdjgUOZ4cnca01u
UuyiUV7C/UtMelykauDzC+c90uu1bkRoUAipesyv5WgehOdJDzGnmuMOygefkFYv7yHEhibxZxlv
+dprHu981k7RYq2W45ai7T8xYyyKRSJ5OL63eenlpW1M4qjAhEH//ikHOTlOWqG7UXfE1A2PO52m
0FqyWfRi2xfY2SsSDgO71fgy6FdQED8Vp/7eM2+4C70H/UQmL5/oyGqpYQyqRMaFvqUS56karPHZ
AHPmK8TdLHai19nugft+wcInEMtxJWINYcBVbPic4AtAd+Ka9OZKAvx/aLMAupxFALvtHME5rMc3
LgZ2KLpTuE2txApRQ7dNn2bqR/xOoS2FPhLlDKY9KHyuvuFxTEAC/WFlZ18YzQ8DzQBCNisvHL4U
9yA4WMYnfTF28K3mzUkr/zd8z7vPABQNHUEK0qb+0x3pDI8Hz7rDNBdyeTEzVxe9NT10AAQXk51R
2QhXrLR/XrXRpiRBk2LdJIOMNIlq9lKMA/bitH8aqqkCGV32lw7q7CCtGlsRV18Bt5tYIH2EunFn
osR1eyfk3sOC6+/5rp+1o76D7kwzgCCjjRhwNxui+Zm8YioMIFs8j3R4I2/40mmY8rpkp199xoE2
Qs7tCJi7TLPkHVF5tk+OMngxLaJeRmuBETxNmIADP37yZ46Ga9Gm+AvyhhAUsPBZwHTIG5OjuSEC
OLCtzhMtN3BRqDov7sDfkVnqp2DRD3+gD/quCrnTQDsqevjOu01wFP0wCT88GKoouqSfRUOLCj8y
GMp9K/rUq5lFTMvOGQMZNwZaDsh79tVP8D/5SSZcI+RO/zIAbzKxTW43DdFLuB69NoacfpFBspZ+
hyjPZmXMNe9iuUNYSNlg68Gv8sOPbkpCKGb3sfNsx7ejbGU7h2aCXkTpPnyEsSwevck1dO8rcFdl
HrYNPmHmCGekYQ353BPOVV9PNpf0Ba8GpoxOTE9xe+rsJQXiAmEJHQC5jhRAfbkcr+ylKVeWgW0S
lx0umcA0n6r3a8g0/8ZRavfqgPy8E1tR24pCSgCM4EbAHwRIZDQAicxTsabFc5seyVGms2f6LKMu
pBFPFbpaHD+ssB/dLWPoADpDXonhB/ILgh0US9OhWMtQmPOSUR+O2hXzYvMQ1njLTGtmo10WD7wb
d9w9L4jHxFdoOnIIzWEOjxbCnG91lTyME28dzaYCM5IavnO0YK+sEyOKE5RQvSBwJBwpnJGu/3Z+
Ttdl0+38N8vPIMIfd+ZK0AsAFBpdLJWw/Bo9De6oofnDpB7uzo886YlWfLXbTJe5/CbxR2HA5get
62vwnggslAMFLGO4FHFWOx5A4XpuRqA2lFHukJwWqBd+lOQ0YVQXeegoX5U+hkxkXn4BhXhCqRcd
pjJpB3Mf2Ivi7XLuspnEMesZ6t5srFmZPhqMMYAe7RtKNeFcFWpxG4tT1HQLBFkguAD8qs9TJ6at
EGpduxsldm/dkaHIilE4hPjG42IOrHCqAUg+QIiaTEtg+Z43MgB9gqnJdlwbuvEUYU5LpsKMPYOE
df/FqoVy+1JvPvxTDNr+r/1QhVRx+l2bKM1Hval2HsUEKc1rynpo9VOyzEapCjegByjz2CjBKlJl
7ooy9Haj0WF8wDEsB7dd3ukWrpJ2g0RKnD522XV9y6naguqXBzNyUoEuTRTll3gYTUaDotVBZvEa
3Cn86asg99wrGFVD+5HOrHLPA8vyfRKXiA6IrjgD//przx1hRPQg1fkd+1rSRkpsg1qO5kVWKEVs
HyrbOpn2aukL0O62tOUs12gUggKb3ymMM5whGaFwEwDitUUBBEU6bcJ02h5/AUWV/LBTHnW849ED
0fbTV+2GkQIgXJ53yH1xCuVAY4ZQpSpkASDLk5OmDj7lif/UXlRD/jfj5v27qApysIFSdy1/AShf
lfEK7qhnuHWM2U+vzZrPUuS1mZkfRcS/RFPP3XOzB8L1Ah5cU1GKkOyWRwpPFlzy71Eq8QhsaeVv
qxy6KExpLTT/dwtp8CYb/WzLTmO+EPqJ21kHgxKrhLuuoEYOdtgKyJKGydZ6+xRMp6QTbM/G827W
qEHMi8Y7fGFtpJks2DN5SxRMGt2OgZFIDt9HXRvNt+4IzGpI5NZt+Oh2EXO3zh/Wo1YxQbfudweN
+OXNWl4ANHXgBj70DFE2CsKLkTnX6Iiab2m6mHeZQNw7AZAQyVnHwsK3jbBgyTEs8dJ7v6OBswV8
W13HOUT+0ogQlzjHVikQruTtUm/Mai/mfnxMQ/9CQMLVvEiw6emyzEeSItHMOA7xUGtVWUADbo/x
jHDURL5CUHDdCJRgWeKyht//vUwtfETQHa9YSEKDbpDFKbbL2HQa05BOwH6/1keD0iJliGsAmQy3
syU4vZMn4jQufIMGZ0wa0uVEcO3WJMqkYxlq/y+qkns7MFgf5YRmoRhe+ph7n4slIZtrH5MkF7y5
M/xJ10coYoMpi37VdLy4imOdJSe1Arct3hCBVkc3jHU/tOpXjdtJtXWL16Ca6QoHEpZ/2KmLxU+w
FOdNfgS65zHC9K9RoYIoEsTGhUvbb8SA9goE3c/+iuvxCfAApSBRqWZ6AA4MRtdGpOlQGRY9fjR0
I5COA0u/TkkyXrC5yO54uGX/6whFFW0vEy4mmNlUkI5XkrcEPvAGkRYpw8VmD98msTd2pfwFRnFD
HjuNRhRYtp9ElCCZJAMttBLKldtv1X59G7zk5fAePSXePofbv53fAky8B6ARZ26nAzn+POLx0asn
lu69MfJkuJNBlWNTwICJt45N9iCpKVGyQOtQnJxgWW/DNPLaRsFF3V2rHMw+puNyJdAxEObHsOjD
OmcW6q9gAaH8zzJRtOCTklNErM91jCl8WfJiD9Njwp5N5a1EetsX+51iVFiKUHTxdxKeUwzdZpsW
Up8uL0QgKgamo1foXLg9pkdfcXXm9vgBg4ELzHUhvNvWp9WsqwnAkwNWYuX9+oDpHx2epLA8xAOh
B5GmJM6MpU9tdIut/GWVlq5a3wEwP+xNsgRkQkPJuRAiQaQT25u4N051PyUedw9eo5WLZJQ4kF4m
5FQ+fHBAq3vr0B85j7qTX8xuUn/6bZNJ+cS7qYCSrNsEMtGYm57ORLB6OFMN6wsFRKP8IdRY/WzD
Q7CJSW/DseP5pgpIUSAXHdqNiYDB9GNFDY/g5UA7IOfykZIt8aUr5dxtitasUNUbogIdDA8NtVDk
c4i6Zh+YycbhomwDaGZrxaNYVT4UtprZXNnXE4D6TxLi7ciJlqwyFRXH4anlWUnA/WQWFUu5B770
YPUiZzgnEyHyHJKKkfn+jsQrG0/wTOLXR7yg2/1knayY3oY4bfYOqa/pAdFiDRWTy5gGku1j17TZ
SH7qgPtO05kpuR8ob5dHQX/e12PSdoxi5BX/SCXhDse5TMj1fzWmxtv5NLISYic4a9HK4pd/B+2F
PMM+QKK7MVGtxhySfL563LDXOH/dUmlsHEoLkEB9V3ILwYiY+MXkIBeODueTd77UZbQVAOcDuf9h
UvX78P76cU9+i3t+IDZK0r5j8m8LTr3AvQtea/m1UmErfCe0j5hfBCGh7qFY0XdPL1W6XCZBOvu6
nDBfYcGHCYwV+dYKvWgcI+wXfOaURn5srDwoliWuD+DNmY974S2+5gAH4sZp21N87vOBbOxDbrAk
5C7OIZ3f47rkeBBqxTYaWCWbYdSQVAb6lLhLwr2fzv6YDCuYyvtkK7m+nkt82fTGMOeInF0QyG1c
uPrQsxqRdmPhqO8Oc52A5hoPPgb7FjKB455HpC64P0OC6jlG51eKFq1qZDT9nK4msbB4Dr79oPPf
0HUdZlemJ0q40ycFKYxSb10BgzmB2bl2NWeFtGQFEHY16mRSyg/VZY0McnZIZzHcivLAZWRwamGP
X9XUfsl2NLRmP5LDA3Rr+UwIy9pwvRNvAI0Jz735GqUXSUK14q2vUcSCJBb8jBKRLR63o/PWRB1w
PDUsly1hAbhZI9+J265dLsPxYYL9mz2IwtYXnqIdN+STR3D1dfoQUm/OQo85q/UGQzsm3+WniQOw
RhL7jsFmqg4CnKfyT48Zin1bj9/zhCqoNwB1v8UrjJF4GprSjWYk5nI11k+qH4JfytKfUVl4UtlP
nwSAXpj7kETyFh+9WaZT/ofDwQmqKeqZ5tw8idDc4VdDr8XRK1/rj8hGH0Ns5+ZzdDGTzFpOepu0
spCCSKMDScLld2rlZYtf7Y0Zf9LKs9vJ3MZH7K0hqsD2In73iHkbk3EYeQJTjNh3fwON5qD7zniI
z0v8iuhR0HoFkzWfYb6VfcBeMFOhDmBXiGYvKnQH31muCkkmnD+WBy+I18kvRR4mKOqc1AZxpTiX
a00OBdrdI+sJIqSOAr+JWz+G8tp3wE0cYUnIPX+WerscdqCSI64sD66BeN4Ev6nRTfegVN8FFUKy
CAc24uzjdMlUv5uIzAdXYWJdnL6plHH8sEsJ6aZP0z1BeUgkSzq3mH+IHZ2wkjEQe6Eg6j5Q/2er
7dOSwudgRHnSofGNAKuQXgQoUXZU+0CDaFCUpEVmjX0miVruOkOD0l1HenWuCG4Bqx1BcdFtg9B5
YcGmLYVi4YoMeeytJIuPHPLfIwbzaG2/nrWuxEUMxODgls1TL+AxTuHDvxoPbvi3IqJP0fV8+lAp
xdxGdiiLhSfJnptrYrz8QQmp4H2fgSUB1fnEg09Z7+m299r8eAfkwp8U4MpomTBMErIci7ZmLr32
BQQll7Yb8gzYwdf4hId1j6tFVAzdyiQtp5XJGwmcnLobBiWd91Oa1VGnf2X6IibXxxkJ3M9UYqcM
r5Io2YGuTzQKx0kevUKpg34j4gLrXntRmvTmhQp1/xK57W/h3tBwaz95aXzpvY8wjYwvxAchjIKn
U9wEd5mA2BaBkAdnzTFxdgtkZrR9bIZXyzpv98bliYqlAQz+8OADDT5unqZzoZWKqxB1B01n+F4I
fW9cE26taXo/H1pIWUHZq57SzErOZi/zg/Jo7mAOE9YKKpprPoKbV4GiuiB5H2CYDstN1PkM1fRK
ZiFy1VVW1OXI6tu3n7XrmJh/pG4rTrw+NsPQR/h2NEMB48vHb6qGXssNAOIme/u43FesigqO3/Ry
oFyT+wAUKevmIyTPQ+NEXrzLQ2KPWp8HBVUer558ps+nMXNwu9Nk+P91pQe2OO+rk3eN8EicWLtN
4mkscDTdSrTHuv/xMD5fU/7GdeRey+BpZv5VfXfkq0x6oPZEnIfYPk6WqO6eEwaULt8yD11pprsl
IZ+m5XoF/v5v/+joUC4KM5Sn/oGjofhisJg1m3PUvJcSQa4WDgRGDRNMN+Q1qjza1VxpCc1olitM
kkAQlVH8fcWIQbnuxom2KocrKkjEULjbfXDGAsUJIPmjqqbXHOlVewD5zZupWjnOuVzztGJyly6w
0QrpfTNN0F862Vr6aHsQVh983zpRB/x5oCJSC+KbnNXijWDTcl/N3JahEUzzZduPR8PupWRMX34A
mgn2wC+Wv0g8F2jOLXsDCbcwr+HEI2TR1LCf9gJ+0JAk0xG/mVOtiHyz/heq6oFdgh2FM9zGJYoK
jwV7qwpBtCVwmpvB/R6nBHyrnRLpeMQZpgzslyejXLptyK5YZ4WOWdBe+ThCMAuwGRFEfk7Rizd7
KJ92hqSz6LUdxmPcd+PSPWtpGc2G4492FM6mnMmiELxS816bakn5YDDOYWntkWQih6DBKdRESZi3
++RvM/dHUvLYxLVwBXNoPnU/N+MJX3qgR8nmME5guh+YYh2AD/gvNK9KUrRhcxdQAEwpkMpce0K9
SJZVzj1omRPnJsscVckwgaLv54CW06aYFILUFgYrMp+u2c1IUVw7tdUmb3c2MXj/Cm8Ml+UP6D0q
6aj6eTL/h7a1zVOqB5Vh8NeHd6xp0Rp5TW2zF4s7AtWU/sesgkHhCtrtWF5gYnKLjSCm88SynNL2
JE0KVWtIy/w28nDIvLy4QiOxn1lQ2qsHNnAG4YMhedu+MfBG77L9nZt9uKIVfp+/r4YXsvuQ3pZ9
Obs9vLlW+oCcIZNCm10+BtG4Xtk9ez6hz0248QsDbq+6qax8nOTgGqPVUEKyjLFyXyvdHy2iKQB+
mZpwy/EPLkkABvbnikBsX62sMeRg+xkKQQmiGnQBDETBbWWRkOGL3yYgSUkxhk0X9q1GHXeDdkD8
LUV3Pd/o2XbiKRwvID09/VskECMGnghIxz5ZllnmCzi7n3e7gV6A29JjXd6oU6r+C/shSRY0B6NR
VZQVt2uqjXxLOIyiH/m3OVcC1sWAQH59WgHOZm89Gcp1CH0NNzLr2oLCBkmW5LUcq4y6AvgE8f22
vzn31wlP6ntJCCSD02odBaop4FuOPztrZ9oV1leqPzdFxt8lUkQ41oosuWdqGTpv9+UswaX6EE36
WVkQ28Dj6RDM/XosrK+4MwgsaISMHVkbrxgNUm2LqPcZpBkq9zYfSe+uGVNetTfaC+5gj1Dv2AHc
klqc5aM0+d4EQopy8VD3wtIl0EvcR/UMznfkGQJh+bJCmDenvUNvzVTE1IJk7+jvWNCeuC/uhlIV
jQOUecRzrHxXKsNrLsrFHuPN1Ai1VyNjsB+LisRkvwvlNZyUr53KJpFPANnYg6G5WrBELDXNii5v
UABVcLIk66pp1SwOUxyHzyAkwStLybJVV6QMM72uwhwTjTi19oqE0VQs+XozwGgTUqaF4JoZg/Lr
TSPhBsUOSQHPjgYXDLVwMOrwin3IW15kCvcA8dVV7UlktIwsUA3MKoaKVzyoMUKvRu8rokZj1+kP
PfmhBIF4BOl/znW/Ukz8bn4vyatA8cegV9ChoIlkeJIU+jcQcciXLFDGig38nnsX9Kig86NWoBUh
n4H5thyVBDkQnA0kEiyypPSSnbtYEV6DXKhFhdD2qBR4h3uR+WVOs0000jEmg3r5vsvIcUsMXnyI
WHLoRHYJAVTpmnpmKi1oLOnjdVa3YJDR9rLrKzyT1YKyNzwjAUrh5lLa4iRaGMit1EbTT2ERkJFy
A8POOB5C3iArG5KRLjm8MWfmp8iW2f6hbakyhtyo/dD3iLyjkFMxQzGUvJmA208Q6B/4o1TUBXmz
tgNG9EReMwG/5iJhIsXIvx/d6J6Wrv5kmdf8Y7s336s/O/8PFsKowTKpF9eW7qzpEdhO/aglqsV7
z7p6j0AOYm7VCbM25LtxLXqzgcOzVPlS0Q+kvK2pN1qvrJICyxAIlUPdg907eR1LN5Z+VJXjWOb5
dWwZh8eTQwgDIA3vHb2MwLlEi09wPj+K2Qlx51SOGBdjRLe2aCRUR9O6Fuqs8uTK8xh2Yal6OZPH
h2ClajnRTNh1UkaeXaAkINVXi0Rn2X35eXcwEkpURblGRUP12okao8BSFl2uluC3zZ/spI62pbxZ
kvIt0sHwL5R29pbFU2DqLPnsayHSOZFpYA4PztrYEp6mgn/q9wC2Iv7MOptWUo9YlytUP1YVTDA8
70JmlK8fFkYuXUse27NyuIJzP2b25aw6lrSD4qq6zP1Y6GU8UD6lwwtx9fM63yqKUcA7ZHJWVIbZ
FA1BaBosFyE5BI1lOo9LB6/Eb7o+QdK9lyj2LBKfKxbEb1eWtyR8u9z1ibLG96x2LTxhNOQ06SK4
E4O6+oKEusCBCmLPWyIzaETvsPm1qoQyWSQ5Fur/UyuZQNCd/DRyimYPgGVaMF4EIb1hZ78stxnw
j5vpT7/oTcXxK89n0WAuvSMMAKCwsBbKma3Ce/SuOd94nZLf8yetKCvfiXLDjNkqG619+wZ0AUV2
/uGb1HT4bLp1EWKLObq69z71BUPmJmbBMA4Wouw2k0IE/WS20FZQY3AvzJGjzOQ3gVpYkuXij0Ps
UkzFLVezVlsl8OlFGytmjrUYzTN54en2hum64Yxl0Vl/cbvzB/UoOUqk1dJAK+ypBTyA9grqGoki
1IJzAVlrA1Gf5/BP40Cp2yD5So62tMk1efMCC460oGQYClFtbkEqAgObTojHaW0NexMTc4XjZ4zW
NtiPI/TqLP/O+99QDR0U44Gq3BC9ZAq9XdOvm0qgoPVBuxXY+NvD00fe6X1MOygn30EpQ/NSXmWI
h+34XPX6KKtF+ZTnnj1r8af/zuFL0QKzDDJuN4KL7ww+VVFUBIUGXSAU6ptbosqL47VPx6YTMGZV
e+WXFt3tSX+Kg+lFpxBZcnx3T6pa9JFzHdj1lPAibtO4czCnCtKZeNSXWZClBZg2toXuLehoSHe1
87FwIf3c3fRXsr3lZWw9zWcYqOu8QqOhDWpxtqCVHXgie1y4o2n75o7G7QqoajIttBFGOK6NNfCf
kJTD+ast9jzYFI8+osxbX98qtZdDAjILkNWay6wamMAT9ulY8kCdG2CP6Sgxx8DDFhmrXTxbpz5x
T4yO1AjADonwMGzqJ3xa1larv1OwrDLEkgqLGPls+HUmmtgEAHxhEmDObuGGritA24HcQ0/38vUW
2cLu4NP9d1UHScuQIFoSSN9Eyuwj51HmoY482H9KV2IEZKaDx+s6iGfknm8y0jkLjgB5fWo8ZKxH
rJHUu8Xg5zmL58QnHF6uXWU9OoT/UbZzygejyci3Hboq5H7hLhPL6F8ogzUMhQ3i+r1e7Bh7kQeg
8EJob7FHRdMu8WpBb8n0H6YX7eFIcelMB8KqTIOHsitc7g+hwc4DviklpGjSaizoOvEPkoUqAYWf
xmnqF/tg1/u5lOj3zM5jEZyjw210jGgZkHVYm4vUO8GMGlYKIG6K9kmYR6e8YJ53cHw1Fr/HkdiX
iocJGV9b/ZFXyO3mOc9UPdk19BKVJTgjxNrRC3TLI+GvwlEALhpoCUWDQ5i05d5KyIfcTL9LqGuC
tkXxhdAIWo3IVcB/S/GW5FIf/MSpWImujpkAoYAG0f4p7mmY4iOWKRIXc2LPEpRdxzUy+auJ3Bfc
OWPyAJS4V9hOQ7AoCYAx58Oa00YMAlOZJXO0FDjMeLKxj/GRVAVvrxCvs0YaQQMORe3Ad9CXMoJa
QdnH6KNlIrpMbWJXmIsD5lWKczy2W1zfh6B6KfTrOuicYBa8l0lr9a/C79cU5O2RLYoBqGGqu9K9
zGPk+3nnRwFhL8wHpToVlxvxPRjz1Q4Qy840/0YxjgCo7v1URhOmseiP9oHPvOr++RYR+faMoJTd
dxbdhIyZsFgD1ZqLeF/2DjLU9Me8mFLIrU0BttB59ewJ3vAp5hFWdqmJ+dYAE82OPEk3maLwh4la
YvVNQXwxWheafYVhbiNHBdMOln9ohSkz42ARrDePLUeD5ZvfgGYMR8WTWXINP0YEUPuTxclaoCru
vSjws3drqFTvmAWh/ppEcGUQ04c3OIbJ+QtTmybcroNy4qK+KGtx7s9Gktn3BzsD/Ozi460NP20F
OHy2GsnRnRov/K7dq9sG0vHoQ3dlNnUli9k3irzLEcsonAwqP6MA2MRUmTdVu3uIRpMjxdxV4v/C
/VtFhTgKvtrZoo/7OaWeY52ue2SVU+/bK2spLapNdzxylVXX7Q5EzYr29NVKFHphd1YE1s0eWX79
teslY10rfieAN54oYU/2vqgOwQe9TGl1Ixdv060PGxV2NyPD3lU9NZIDBTDGBokq/ziR+Y3WODMx
xugppYstz7oq5tZWafSwn9+YVYH9Z1qdnnm7sZOMSSLjr2zp2Vv8T+yd0va0c4pvKrIEOHATk145
gC5xVCRNhuPkDWP7RJjlLG4KK53uakh9LxyxaoEedJ+j7vRg5GyAhp4YE3PRtOIjvCrSuN7XE08g
jUOSTKmc9bBgUdA3j5fJQGpD/tJZDqlRTKKtXlsGyqLEg5mqTOTQVx2JDyPU3do6Zx+iahT5oiuI
x1cm3uesjXo6kj6WDfTM67YTPtUJcQ9pZ4XHPupSpF54IKYU1ztmcEOR0DSfaT7OQt/UxY25a9cD
8EEfZ8Pyb2FPIgCgPoX6HE9dQF2t87Wmf9bBtCYIt4BUQBwKvz+2iKXTYto4RxczTmAsJ8GhlmCa
YRkFTRfbSlZNhEjESjmJgKMGAIlsV6YQWyPify8URlesfgnPOXJKVNbuhKhStOVNnCZ7LmhPxXyS
n26CoNMx7fVjmvxoJ9wiVCVkFSJJRd8OkHxZnBXe1kbCBgSikcmvOR+RCRR5+pMvLcOX87/hW5+3
+YzRyF+UgfUkQHtlSxTHJvffYfvaZO2VCrLXQdk/vwYsGKHKjJ+K5dPp7jkWnRWV0K3HIIckHUMQ
uk4aoCvhOczFy5+CH7VnVa0A/lqFn+6E+Uzlhdc+EmPLEe9mTJcJfHwEMnPvVsuUnAsqFjf/i789
dqC7QOKYCV2jPerjVLOZr5NLJZ44loxH8ogh7DzweJzyY1E9MJzb9KRc4P0x3AGHRORLJOmQZjpN
v9cnM0Dou8MW3KNcWra2FaFoX3Bwc5D18fL1eWWPrdQAWbAAqYhyjvxzZ8qxw2wsw0ZA/Liodsfa
07T3Tb3htLhg3ZgF6jV4L/uEbsY6XyUOjh+goLwdELz3NoYkpMrlaCjM3gnbcxtTOvqW3x5eZip3
L0ahH6Z6ymXoF2Fsj5ZVS4cA5my9/DwtFNXB+kvPtcsRoi+FeMnRC/Vhb2PSHcZfFtL1LvS+Hp/L
OzEBS6h66ApEMW/X+FJahjRnwX6LuvvGV5ci1tAkMLRG7KHo1mlbKm5rsQ9B0vAT9aCwxsZAXHCA
liMDWL2JxekL6Os31+5XZUgTJfnmvIT0iOie/nV9bTLbSXVUaFU6Wt+3Bg5fkX13q3e4Dyb/9l24
6qGjEOGoDt+d7U84YR0U5V+hiPshQpuOD2rIeCFAJiBfS6LtZY/RYOThIAbc4oG3gGUVgpAVZ4ed
poNQ42T1/JBCoPmQWwTi7f5IZOid1k7vnF7hjcVFqN1DYqv8hYyzVsV5UKj1yyAVZSRHlEwUhVOo
z5AdCgA06w/JudbwW3iuaO2J9xqvtU2COrpfcKHOGokfqCWmGzhWoZd1E/45wGkMBwUqjUZarQWb
Mt5O3GK5vHVx1GtJl/ZIE5VytddwXw2RIuKbs4VzGvnMqUti/7/FV3ztCCAMcAfZpOkcdR6eNRJP
7aS4q3UZCqZ/7xgLM6SPanFVuRpMDaqn8GnCvlL9932lbRs6aWrbSCwQpPbasJmAyxIsn28sap7k
0R9RtrnhfWLqUGuoUEJPpcE3Wx8EUhAB81ZpN2tKws+VNKaMO9VRdY+dyy6JVoG5JPQXwAD/OwAJ
mluKyk4cXH2quYjmVT/XPHswOtbnuTBt0uX1y3aiZ0rQ4Yjc+rp+RUFhemIfGfMqLLvK3aT1qbts
gOOoCMH5srZNwflIsVPBo84f9/Ahjb5TWroKheRo8thkOW5p9jhxswl9XUb0m+ZpoXn9LK/KHRNO
yrIOpTo3SBC6bG/xaJUvCgdauy0+UY51nUHwDC97or1iyaYWz4d8qesG1ocwanhr4kK5ADWtxuKF
i8w1sdHtuR+m1f4Sv2fxi+bim2+IR4/UumjDi+pvxrcqkhK6l5Llo4ievPscAU7E3w3V0qREQmgc
7ysXr8LL5A5wDXjHZ5Zthe5j81ErE3SrSgKJHFuIGeVNqU1nM/Zf1eJVOwC6hDxqnFxry8jPWMKV
nLdBpxGaJrB2rPJYk2hPz6yko4bZV6RonOEFeR4MBeGcjzdg7ip7mVUh3U976T0Q8zWs9jGndlrH
tB9toDZMByKWEKTfcYAYcery2x2dWPRA6fQsjCz0oCjjH12vJFGF3q8tLabJlvDzl1Yda7lvI6w/
NppoA+ElD+X5OJUQ8W8XDyP2QKT1PwqeRWV6proAQIuUwdxHg1N1cpxxvt+ZUWGlXXHKD7qReAVn
UdEWfRC4eyp8nCqN1QN94ixeYO8gtMszGb/jLeXH6CH6Y15vWYqf1nSg50gDKcXEudadvrkgXQvF
G6VaU+GODsfurXsRv7JhiezjJThdI5EIodGIwFOuT3JC9pD0bqpUTywsh5UCN+YgkAjRX/pJCEV+
S2dBmjlRplF3XDX/TDfZFBvaS00502MiEm8rbDfzgdxk4cKbxeu36KvQrkZdGxouR27+FKnCuAUc
RirBUecrpw4l6Wh0CuorL//1W4aC9irnsbOMox1jAr4SSMdZlW1FIJc2LyfCRX1NKyndYi2X5Riv
M4ZnB0HzQrFp2rofYG0oleptF1OLi1752yOl890U1TotMbnWIZU4ExEEdGqhkEwzFkEStCmVt/1h
pC7LVDW6Lfalo/JU714h+7C9qDpP1hQkCq4cFstU0d9xUw0WaxUmwR27BAMZ3oC836mptfj1vxxN
M8zGLiW9X22aQWVx95Vk5sgKNVBIz2hSv5Qo1lpWg01LQ/ZlOw+CIK5gsIVOS6YxO5duTJjR4IU/
ttiXlZophJ+rSKrEwiCKRWAiCQqNDK9qDktdY3wLQewRWYzg5yIExC8YhL0E3FnfQywEY+FBx+GB
9AI+XGAMw3DBuHRdQkChjU4fPnCgj7Juo4TH7yNP2Ect996r1RXgyORp848ce1IWPKMxtzxvJ6Aj
INb7VUEOm9VY6Fb8G/IdgAPpi1ONvFM9ZvjznXEOENRPLMXC372tWR3sRNWsbjqDGQOW9qUvzLv2
HOF9XXzNV9IdqRD4gRLWlmkaNCfEuSNZ5u8D2SQQwZRM/4AFD7p+r1WOA9ypduYY28RJ2aR/vgzg
v9xFO3/qwPJzQgaGF/yXS14OGgB6LkZ/Sn5L+8/gkC3eSqrttPKc+1vR3/uXpRvB5aShSHh+8gx6
3l0JC3eB5hOixMveC2g8B/ShIx5SS+IQ+40bCOLX93odjXZdoejb5tiD+x6dWwu+gMlY5OUcBx52
g/SBYRRd62BNZzOThyOL9swvfwmDlJuEk/I7kod9vuiPwKEcedzl8YuW9Sk5XVcr7KKUXvwfaELm
bzeWWa+Q98qHZU4s/X0qX+2fjaFIJzNWRNI7IyUa8L3+EC89Imhu/KVR2ABeNTi94ENmNz6T7Cn2
zu/70qa4TKYmpcfgy+5MIO5M5H3zAufBAGpnbjwOllI4vVHXg1ryh/ZOj/FAIk8s589UuE5NE1Xj
BS4F2CieZTZUUX9PdYaNJioJqRaKdBdjQPJWcbvpSWgz59FGP3mSzvbiMO8zyWcRWqplqpP09cHk
H/TkdoqH2SIflevkFxfl0s3lZYZ9xjXhlw3lfebfWxOARRUrERODAjvgtD3oDlLwkxPOO2EdyOtN
Ste9cvCmmxYLXUyN5a4V1ufLGelJboNF04JT2pXaeHPNcImYT/JYxycjZKufiFDQXTlWF7SKdxlF
bEi72mgm17VO0Jgn3H6h0RKu0xSnUnBPob731yLx/yeVKOa7G/38joN307GTMvuKKpQEHkS1j7SF
L3/OyJyGm7Y9YzQ1fWmW/h7KitIXs7upXvfF8rv1ZpdlyaS34sa9/vKBP1rbFXAP61lQsDjsLgTs
jx0kQEgqBx79U1f4HnGQ1k51Jn3JPCMW1E+Q4YZa30bncHcWgRQcHHNS0WpoZLMTM9qt2S/nNcEd
Lm+WZXlDLvPb3LX0iJmE1ZuLr8bUUjHX8+VNi47eZbl+v41QmtLBVwvMt3ECn9a08IwIMf84pCbS
SEIm7HnR2ReP/IFhRzf3GwGkEnGtJBCADqbtEPC3zCIJXUlhSgoxGQuMUpNzBBEnTvZDB4MTSmj5
qFtYFRBQhTIheO5+x2bmiVrTSChI+w8zbhZdt20VBd04hSxzu6TIX2nnSaP5DES22Ox8ogrLPlxI
fUPwOJ/BcZyDYFc30l0QTHqRy6eVshvZOI3RyypXA0kAYr/N1Jarwz6x5JasH1ioWRfuATgmX3JR
Fx0ypMz+nRJDlHqnVDtaIl5gioZDnXbgcP1gwyhFmwR78lNaQMu4sl0CIg4fB/+mrLkH2lWzfkDf
/8CR8qvykYndsWOh82uTqOxvIFUwAEhivKMl3DmZVEd/WMeeU+PiZYG942vsgNlF2uhDo365AIMp
QgfrqnAh25GaWvpPZryihmKs2jmuw5asb+8WWMBcIo0D1KeMHDmmlNDFaYCsAHcjTv1b/qsfOUMO
EcqpvpCRtCkzXgr6OkDIOYx8Mj021HwGIB8N/BTWmew2kOi+Tp7VEA/Xh7Ox2F7Lh9r8kIEEE3+C
Xe4HDs/MaAq/528UIqi2YmTyEzR0gHSo3YEizQ6rrXLX8foT+roK9Z0+C2aLq1JrTYjDrD1kTHZt
HtyHCjE54bHFfzVCpS9lqg4uTzixWu/l3x8TvDeFkgj4fKJ4mHpvpIMyjAOG5jyjgPdPJ1B1oOjF
Wek2OQpJdT5j+XTVZEp4OTH+5NyQWRJcj9bs3HyQdOcnVU56XWVeY0BZRd6GuIEBYEvkY/KWgvFQ
MazPud8V+MpwR73KKFgDQCIT5tQfhbtKhyGYAFq1BUabwxkcRPWfzuP+PDN5Hb1EXumFCh7E9zrK
a0Dq7HMnHXvIkQHtpk1lLW8bivCoJBQgm1WKBb7FGTk/4iq0XKW0Y8NYD2+8ILWdOjfWj83wiLuD
ln8XyjR2jej3LVKtjeF7qs5yeU/YZ0Lal76DjWAkPFtvXiPgNoxoYS8PWF0YDGF9rA8BPYQVj2wr
0IR80b04Q0AOPxBFJbmzXPzRs1bav+Ft9IvkKf/NdwXGMGaPk5oNPmJBtJwm2pzseTA2q/9wXgMV
QGzakvJ6DwHwHo8ohttVIBDEFDYY12Rv2uv5HokC80yPWF+IGm+6JXwE8dto1mKt3s1q4zcvqbsx
+/DP5xULp1RNzL6vOAYxUZiu4Ry88+3NWojPa6cAYpfjXmnZfXRseKtfSZSvgN+b4wHXNwWIBAO4
nR6eSrkRuRLEwg0Tgbdd9H4N7cK93cRr2frDQKinIlvEcdofFvSBROCNOenKCP4VKd/vKSXUDg91
mpWHRWrjtSYt0x1lgeyvksJrmp6Qm/klypt6FYEK1HfvMkH4RhzSo6CTxUMtQxRPJ9Z57Ni8Lq3t
eYX70FkNVm+PCBLiJYajMv+8CYjJ1lT54lOz4oN0rdOJpySxeWoexUHZw+PH4YlpqsgcsGpAW7Q0
BdkQvCXO40GFW4VKhOvB8CmU1UbCp9g3I1UszDYffq6BVt15g+31BoxQQJk7z5WAxvUVABzdWvRc
Q/aoDOLPRYhHm1FXnmkthuvXfZDossVRV33JEIrCwH078zmxPYUDCx4cE0kCf1zlABeOcY1A8avN
PdXYhZp4adgoTd0F13DMn2T4P//0Dh7Pmbwne7Q9/nolOXz7OnnUExVwVoBIaqglHmg7gd/5AiRQ
dy5F4E1NVDGRqTFaTo89A3nOqXTJb7mZ70zNHBi8q+xo3dCFImamv/EdWSsbtlhEsaQrW5FSLvJo
SssCghyXf43Z3Eacq/GoWKCh4duU4+/oYyDmp1Fa2kTmbpLk1hnc5gcf49h8HS7c/reowY9XgW6N
/YKKmAv1U+kHM3NG5uKEPwShRQSK9E5RkWs9DnrB9yp310LXpkpe8/zBm7DBx1FfJYIhGx3xjZom
KTMOUkmgOgFAZk0p+Ej7XwZ3fUpHepeXkx4mOHquTaC0q1x5P248TPxjELtZMooEMEY9e9b7DXIH
8R8ZPLd3riAvHKC8K/koWHw0Xk5UvLorbP4EsrufbkjUqwwE8qKmH0Po4mHl4FIh1kGVqhHgoOhC
bkbuAnC39nF3Iq2HoC7GMpst+tk65S9tMZ5PwWXgOKtxB4W8HrnUvYVeDKIl3LnLsYcXv2rjWVnl
q3ZjRNG59toEJYdYM3QUNyuzIYvY5Rw5Q7bWO/rQ1l9nFoRT61dohu1KDpoAUy2ekAkoqJZj/+pB
NS8OypRrR+32KZ+9Ghfc9rQS8zVtKnblIYWZG0Cj2aoxmxg2VlHuwxtAbE1PlxOzoPfBfIWT9K97
LXSznsff9yRSRK9QWrJo//E8NsdxwX0F6oyVzSmBcdMmGuSjjLXAkAxtnaESbksN6ewSxDF1KfkU
qBFh5N4Hbt1t6M6OwBkNd3sZFK040e+AtWNORTAgzopf/4/dsYVBMiSjPOQcOmS3ZStQWsH27Pby
AbndB9CiTSSubqXSgzke1VDO2gkcOcgs2oiG8wTxKdvuR16Hexs9U0jp5rL+pKoV41naRwTz12DO
pYCpBS7pOm4eQ+ATqOEcuosXbU07kbm1wrPQNQ7Tvuz0mdPAlQbmIWaxg3Dafez2kZ50gXNGMKhH
iW8xM4sAFC6GgnP4SAk48uuAHDLIBmMDgN0R//YOH9QiJGGvL1msuwdBsWSYqjBqMfyXK9tm6AJw
+d36nJpJeMC7aRXSSpvu/llrf/u75NMRsAoU306WFZ69WZfPS6TmPGBivok89ewwjuTRbWmsX4d2
f/18Tk5NPeF/rmuzvIYuEfFNaxSZHL3fC/6b5ZnZcqgW2VsFlejswWDj7qBwqyUfk9BrMRkOpylT
inHDiwlJGl5VWy7VcWuadW1izTFxwIGuvn3Bd0mQ86CSVnUe9NoTgrrWxoRaHyPbiVg8dadMMrva
bydavUyC65IStZvIiZdZG0qr6ApNKWyLEYr/ACRd3ge84yCuju4mcTZkOtTs8r816NBia8xnvDBd
Mikf/Pzll+G5rH8WFCEzXPu4FsmNe8jaIF+YgPgNYkzIguZNKAwk9bbpKzGsN5sLLRsa5PHf7zjy
BV3NbsmZspE1mdCqlBqOGN8JiK6Pys8SPhYmPlRwy7wl8COMWgKmupovpgdaZDD9KmzxvBmsjo/F
Y6QDojok33B4/SbyhL2oSfPT+EzbBhu6r5KxxITj+Th+b6XnttTRxjwEkO1rIvRsxjW5wAoIFwY3
lC7IHhujwQ6aqP098rtlgutkGWYSf9Dv+zT88A0o1muBiZjqqys/eZWewY/SjV4oUa8nUcEvaG3f
MIf44CouMPBNdfTwpLEOPMSqHrOt8s6Gew/nIM7ZNxlvKtbChoz36i2rVl/RBA8cddLtXwsh326e
AOt50CrQx14B5vr9Jpwq5PCAsE3Xmm4hNY+QROe2DoXgYQ4U5nYqBTlr+6tzTgCD0ZVDP+HsrzhO
GbwYnglj3wiY5SfeSsETZ6DJdQj2DcyjSV1QBTUNKVb0l6pIebNY7VnvghVNDfjggRBvftveDufF
WMV7+qL+Em0Lnjy8u6h4OLH/9cwFJKEuQf5r/vtIwuxj3iB/Uxa4nndOdhxOeHlZX7XJa1NfQBq8
Xm3+Vg7d56huki+cCc3PBYbeG74nglqpE1fM4Zxd9luH4Tzagq5Qsbbr7YMRhOaXhT4WLGve8DHC
UZVk4FjBGQKrz5zuUUmM674FUEzEiLCRt/HN+YuA5QLctClAQlf3WHOuTv0DPc7EvUVxitgTpL8C
iAcJkoJcwVr+gmmEv2aQSXhf6IA/Bzm2ZgBQgnh2Qeyihfm/5CsEN3kLGWtKhVO3l7tDCRiYIHNz
l6SNH4uvFGbdmZdIHKIY86GPX3sDMNYuo9aqouVBOFd1IsZ+BYtM7uMZSc+wfS51+2ibqeSSCJh2
iIYSokGjFv4jamiQxzlMthskwrqWKVRtlMdRAFz+aGgUO6ywOw7WeKZS99CVMWcP8nm8qskCqA6y
jI3LMITt7pHOY47FVw6LtqWKpyN5zoM24Bnsm4lwNd8C9dqU+6VArH0QGAf1C0ea5HuJx6YZuYPP
f2UE3+IYLi/ikmOprD/0TOTffaKg5DxlGKa2JtPXnQIMeaBX+YghtIf34zEU+AgAsohIxD1FGY7v
lIdMPjSn2u1n4riY/xRlF/EwikIS+odHtqIwiQQNGn0w4VNO0FyXgDtDqSKfNILPtDrrxCt9wzYY
Rn/9vOeFoxd6dbKLQsaWy+sithliqXFT7JDaLT5Kg5snzEqmuGBZUlfn1b8+V3g8FxO92xSLk2Qh
bxOOJl2VbydFdBBSyxrcFvhz9RThxYrzV8qsOMi8O0+HvaZ1SP6NWJ9fLzu3t+lZEPjgW9UZ/mz/
zGkk1FW8/Y1UNUwjLz0wFSkD0XxH/fLegkhjfyoL1nWkkPNuwSTZnytsc2P7LUPWlIzE77JoXpyl
wsBPibv8X55U8JPsoq4oRC2CBmiKJWyKkV+LD7KIOBhXS+v/EWPyV1JYiZ/BtjHt8TUNw6M1U3AZ
0ogHfdAG48e2D9D+1kHuffp35TqlCNGmwi0Jd2ChAGnMxgtcxLli07IZovIcOUwwlY+DOdGi42YE
lH7g1SCLtCtETbJNtwCtpxgtnqrPoQhdxiusWrua5YyEk211z3rOuhBnRxUxRjZ0T2zQaj32tPVd
J0FRsxCwkPSn9WdwNMgm4tvu1tUV+OMeLiOfoCuJAoLJbWVb8Lq2GmI6UH7tN1RuON3arjn5dUu+
gxvJb1f+pYgDajtSpH+P6kh8n328CUNJWLufHH6G+5jbMLRnvOiRelLZC6Yg13IpjuQnMCiB4dFS
MbBxq7q6vGle5x+RFsjSefKMOABj/haISQYnpr3VOrqH4KuE/EcovV3hYnjmrffSndA5UZTOIPsc
vyZopTMYU3tvqMqoZmtV8k6hSXt3f6zQy1eJra1AB256e1nZbe+Wr6Osb8ko6xnf2+swcYMSu7/q
nvHP3PUy+uo52Y8hA+P8XkG4ib19Nq/L1d9Lmt2p3hG/Zq03McZJUVNtb0J4vTHcH3lYGPLRJORG
lNw77E2EU3LjmYJ1YNFzjWiVXKBrxh2+NIIJ6EoVPYnFecXeBjQ/W0ONqeD9Gm+02sMdB7b+hqAN
H01PB5AU1oVD7XYNITizD8EzqmuRVKlUKYsXmjGl07PULexJhBv7O0XQ/E0BVllqJIvwaFhDqLLA
Wu+Jvv1eWJxgPTrRcpsGHybsufRiAUtM9LWX9T7h/D8vF409k8+CTDBtQxEHiw7cD8UBJOc7kH4t
AUyTorc8G3jFzwto8PIU95qgmN4Mhj6YqxjiyO4uQmWuOjrlxfcnkpgafwoPh+6TyydC93vldEON
xJhAqgWFYMzeSPsgmN5sj7ngIviNyKfZ4EZcJX3wPiW0Zlsz3Vgobmz0bj+m6hHm/qIrX+LtrWLZ
A9oVrmXrNxEykBkX9c5jZXNOPs2Ch5mLAgtOjcLh4cFpAjZBXWh5jaBPuR58dFFlyztry3Hb1Drd
irU2SkmsrPmlT6DUaHsrdl6wubdupfRAcQUik2MWzXTu/9spsDPqUm3Wsyv+JvtLbgSt2zYtG3Mw
jnkmJ1MKSJM7nV3I98Z6CY3I+JGbgzVrI795+IWXlN6bvLJ8ce5trtyD7BsLmecC9sKkyfd5MmG7
EWV5G5FOpn9PEvkqhB/TCoPhfghw/szz/v9ehphbspPpHybWiEqZk1JPb65tSCZU0+r98wpMBs2u
GWL5s8cxu9e6VNQKZFGj+2ERBOnkELlPJqf1XN8UTJv+Sh0+trEqdzxSzImtTDn363Z1sAU3PrLj
ISWbYhTMSdjPjB3He5dsQzkJ/BkpKm0W/LB4JBNAYFeeSk4renKDKu6LHtyEdZtwkiMDM6G7dVR8
U3gxQTmhY7fVh+j3xyGs97bixgucrTcCfUEvbz67E/nwWO1ssNlEcTG6ReOB0JZmTjVZ/XsJwzF8
STqlavA53oGOjWOlHrLNNzAt1kxIzoa6MMwIPV7FezRpgHlTdSVdAq/U+LlpNgwYpJMg3q59DWpl
D448dbCHRcUxoGvqnGdA9TS8t5tEY2/CwrqFqvRq7GV9GZRk8i/F5BCiDAbXPu2Y3x1VEIJGi+xq
IfzDTd5k0oQ8l8NcyKP3c7YHZ0taAXt72+64KQGz4Ki/znL7rvUyzQjei3+dA4iMW34xap8oMP1A
T1hcLVytk9ixyzvgKtfVxlcjF6xB+5DXXbmf12ay07KmupSJ1lgwqEHd5Qa7/UMPMDfkwVpiRo94
7u/YWDc/SDEmnP4SMMFdBoH5Lz1utk7Xni1qNcpWC85gn8IS8LIww2lXVWxMGaG8cjHe/m7lHekp
tjlio486cMjN93YgdL6hSPeWjAcRsd+O+t0bbMfgKPBf1WSHEP+Kx6aDbzgOiPMvqFlrFJe3jeUC
+wkWTrRXXMZujLZ1SzGakeysZLK1AnX5WMtsn3VS9MlSgW/8M0nX7379AfQitg2DIXmoo2rHfeil
q9a28h944f1I/m4oYUE/iIS0gTve8eSl3Qy59AzXLx5Yz9fZUQ01gw1ZDvlJxqTzxCN6kElQv0CH
aqLj72XF6o7RxeVtdoUjrwuyOTSoNSJpxmdrvA0vneFh+53G9Y56Cgw8a9Ntli26qp4oiLyfjm4C
zWLK36oT9yndtpnn11fe4cpFlczm2vciGx3KkVDllgyPWtgowFBjQCozfVLTY8SzrwOeFKhxiiMj
3DLC9iea9sZdWZ61idNMPFiT8FbX+A1076+7lW9GEFqPpWzeIX9yu6Q6BeeiFbRvCdMBnZ6aKP9A
G9ELOluD6EYaq/jXXizWbnYYEPgFaPz+JmbHald6Zn0WtDjgqNg6gZ4RZht/NJh18WQ3D+SueSZ3
ynROo9VoREixPg4/szoiW9OnExX0xNsWMKavGbJcQVh/yCgWX+HE/N3ITHLKuxVfT4Yq6FFLNoXB
3BcMoiW7GZ3Vb4ADGeO4NkqN+5IaR4DV8Jt6RJ2HMwcxJo4WvgwJvMZOpi+eWtyuz4v6e5B3xjNN
I6Dd1+pOTdBmeaGB4DjXzdMkl2JHU4n3qW+Vw5B3XNbGx6zrQ44sRNDexM/T/EctMDxJCsnCpTjs
M3RHmRKeImG+wTNN+f7kgvzz/oDwyg4tQRWCjixFQgCdPfnx/6N6SAaMxOFPRrZJ04SYDjB8HXxe
cAwhlLuYc84z56Wh1dZGJ8sWcA9hW9VE9wGmU7QJqQSMjBvZWlXd4kJWZghD1nUN96dt/xRW2sR+
6pNQupPq/ZkMTdG7MYTw3MCIucQteSwm3QQvVm1ROCgrXlCQUgiJO3HFtsy1dqflU59+rCajgv14
CHhIqnWX8xhmH+O4lazeYGaAei7P2M8J3gK8XTQ2DFmLvh9AMUTgPwEKsrDMekQ2Z3/xYi4XqVAH
1HptB8T/SLTo22Cj8/tDQZaB7MFCgCYO3KkNcdorC4MV/lO9OhvJLiGIPcERoNmxvma9IUqEdApV
mpkOH9paT8Q9+raBsOa03szPo5UHyRYtt0o8S+yIHuT47xbnTn25m+PtFRbe7yk6Gd/rxuBqPXF/
iWTYe5kPT0oAXAISiB2ph/U2nMZLUAH9KBuE5g6gr52xLSny63sNSUbm8u9tCQqCK9j8uzs6oHc/
x1s6d2jHwdMu9cvnpwJI+i1Bfn1+5IhArg8ZB5Xvcyb4zSqZGW0KE7DBrxEsZeYJF+rRBdZR7gWt
1MaFHQmeMwWfIRKFqzRQ6pBckWV0vi3yxn/xrUnGz/mWPGXzFK8TK6vV/+jOSpkvOzqiJVnu21jj
IlMo6mKCWKxwbyexu2SUOgodXDbIBefguiq/TifuosPAj92l4EBhRL3CDIOI+7dMIzQ19uSXLttW
7IL8Jc6yJo3X4KCw62A8Y+KZG8B0oh7yK5nP0D1a8ZkDSgrh14HacUBgXl6OfXa2Td24LftVuK51
kq3zcakLKpB38H/SjiYqlgJgP2X3qVBCA4Wxav5Zr71wd5Mueh7ENgUheBtZLmAMvUyy92dkEIZI
5gfRT5wk/mXW7gf8OzhdQynKvhdJc5My0YSXC/VwZlNex0XN1DTyEXBVS2+Lfe+ozc3q6eGFZmjR
63N6d0smhBgFw5j75KCacn6xuRlhvzkM+3J4yDHBKv1QH+SW7ipcMFcHmvwh/xV/H6dr1fwBKtYq
KOUpBgPNlLg5+5XoOLT2/YBbEdnnvBjCuem6QIitRXLtziNDQPRds5Y+gmTXvGGFlRQhVbFaY/Wm
4qeVxbmRJAKdV/gMp1Qk4uEKC7Y5apHZXCk2+B2N635fZ2nBqcVi4fsW4yAsjbj6+cpRoJRHN3/5
OozH3UyF/Nfm40KWNGSrnaykNzsfDXSygffI3mRXxzG0VxlJ4HeUUvrPtSh36sluRd/XC1BZYJik
DqNmpGiOU4ksVJ0Gh2z2QyjBSb75yIrGrwu+dQ5SA2AvEegwixGLVlvlfqW3INQAfQEz+pXGjnl/
DRG8zO3O+RzrDMsqaD67QxdLXC9fVstS5eEJeX/kBJo9itCRIEvmwSKT8Ie10y7k9N/rc0eNfKaZ
UhUEYoJpPz/n7/N3jrZC75wZB89KZKLmLnTJRzxzdEZLszkx6KgSSXoMsF0AAxD23locNdyfNfIE
51SeN752PlX2krtK3Wzjfz36ZNXiSS6BLvwTnyOOpI3FEldc/Xq2aprVhQ7cF8Tv+iWgBVj1Cpw7
FQVkrtczbnGSEgQ6dRqvNNUlrBXmeSbuew05bNVHEKf6rlwicIQJ8v3eL4JKiqKLlGHCOGmLKKP4
n5yhNmCRaGXrLJGvlcSVqEcVakxf2ZkkqIxc1d6Zk7u4OKESsnONZT6zhH0sOxPWUx8GTMqM/aWn
jz1pS/R3WPEP98dvYsyzqvqMSC5nFiW/BeUAOn2huv5hfI0cDBxnqNdxtwdvp9uSbvkIJc79z7s1
iSIKJYWMNKoam89w4muCDvNMgpArA9NruoktGdJW+RAp35dIgOTey15WxqUevIwDiEsxR+nKtFEN
eEmtJZcLfx6npy78M0m0zEK3STltY7Ev4sB/ik5TRdAxzcGhayYDHy2fmRyp+FN6JXFyIRrIxTms
YkpkIQYasRPFTuSm6fra684gMMu9CkApk8t90G5WHNRyxE8xH/wxYnxijs+Nufqpw/t/x63LGK8+
jM+EIONrQRABJU1S7nJVWOpUJ91NFA2senybN7fUrFComSqZHTjEbeO9x+Xbl23x6W5LGa6V5guB
0Y7fRvTDOSOZSn9MFuKMxF27EAHEA1y+iKhLxF9ZD55qKHBCAjiRznUbDHFOnv6abHKqFFZMsaTz
o5vO3GckYrAB7sSIo+e1M43SjGdKFOdxq5mZ92xMraOaOtUkpVqGCBkpdjkZYMjKg6B401DFsf5m
f+Im1e5xxRjC175Ch4hgZDcP5yiYRyOQT19lOZDiQv4jUFqhvavVlYPjHHTbgfBzxIDDhlVbcTwj
4e74h9wIhBFpOcgmnj2RpdOEenc0vioiE9nTn+cDnSCxPyAqCpCpwYa3JD/6Rrcr+EqNBzLQM05c
/0gwZuBmfXNOSE0kkqIY0tIt7oM3hpbC5H6BdHNwzevJcIn4ieoibjEpfSNu/H44nCMHw6jAhyLv
eRM939sIYkAQzUHn82MBvgOuEgxBcUVlCwxez9XS8mCtMmnn0fNYqWjLCc9I32ZbV9IRSUtFmFtv
UVPZBpcuCbtP506rhMv4IjPadqROKVZ0VG2cMVE2NsOncUbYgcVUI7wy/6NQ5ntvsphskXLA6zyy
GDDdRyUYZl3XOL7LnZLLF5PPnLi2g9FDqfnre94pYEI/xBmFJcsx1LBOBls6riwwlspF4oLFERrj
TYHbPdFARBUurHn8FthreoMTNO9Evqcmb0GQRgCkb4gBQHwj6+EOAoIplHXYK7DDavrr1jOzkzWC
A3sCWwk55Sa8tBZg7yAW/EjKkFZEZMhf6LKXUhpfmWnAoAM37SytByIdOq1wetBNB90vh6bvpAoc
aHZvqeNPHFYa4cJNhAw2mLoIHmlXPGDS1XKEeaYZeiLn/rKlPYGvkG4JOzmHv5z8QcYls9qw0zP9
drt255yUcQXFWD2wPQ2NAn5fLnChu0knDUnJ+xegwKtlQkQHSW1xbLhHBtoWqa+JvXbdGoS36WvZ
Eieq8PbJD1q2mMb5RGiua0F8+geSoCp/y7X1sr7tHkHVpgev347SxFEAyqTnGLsUMFo70RNx4HR8
zwTM73qydwTGPWEzdHtvL5tKq1BRZyQmjMTNccd2btOInL9bouBXwo+recR8m2hqTOzYAxj+PRVP
AkgK+2A3z0CazOeB68+mb7KatcBmGPB+OXbZ92NGQJXIMlo3kLpYYBcah8VGVrTD1q32FWnTalUH
VDnaZp37c3XbVL3XAMRBz4ZoXVJ7K/BUodlu/26W8+Bn8XeaeoVSc82UhxQExeXT7TMuvy8MF4S1
F3xMLsHxS+TC1xnG0K5UOE+h6vuR59Z4ho8FVs+gqH9S88hXAxtjo0qaqcNTAZsWP2HcsmWnpI9b
T0HGTXYyyaUpCi9coqKRERwxCqNlDVYtA1UBNxSS6SlrCvJ6sy5oR45O2tW7fYUxf26wlWYAuNPL
vGR6EbgaPoITrecqWVlcofWPzDFlMAa//tAUeKWHNN7oM+uPrY3GM5790vAKWiMSIAWT+4U/OI6W
UjOMEOlSZv5mb43Cmewe5FAqF5EafKDX6oDil2+bG3z8NEK93/aGLakJMGS1VU60pLu0qsoWZN7r
BEgIXkiAOpKwo166rE17jgr0XyIdyMo0eoijFjcPK4FqOsl8t49yCGzarD5C7T6z1vHLQB7+6qGs
Si+KLjW0jalRm27KnM8nOqhjZEk0wiQdKkrUob+XVWb6uTzTBx7un6Y44hmxwHe6gKvnZJiIYV0F
Ogol/iKUqZc9SLKPjCjn/abIwZzwfzSjrlyOfpEyg8mnFDxkj3x57BGSu4p/6AwDdYJA3eFKmi9X
G10ckX3bYRTc8BKYpP8x5Ki6hvhsbaRl26iDxnxwBkfLRCztCx+uOwm2STAzut3wlI+ATiRnnXtk
nkK6Zme2RoCuzWO/ZO9G3zRbg6de/EB0ds3rlvS0S/5CjbI9lccjxs7qcHIabFDbMH8KCJ2whMfg
OjawKhkiYafmjiYFIw22u9ic7HRkpVAMVZG6CvHSlSnvys6okjN9UM91meJtUvoG4aIKljW22mwo
b2KSgZvveuRjd5lsMgQstPHN1lbICPgGRI0kAvvH9Uuh1pQKmUztixIUi1xx5jyXJme6NqA7lvAt
bnerKH+m0dscf/o1x65K6QFe2geD2ggPQzcLZQAwRjSvdfHoMPEN7tjBUZCjA1b3ysCR+85NGOti
QYexUXCiAo0mIuP5K9WhGTZHwrGvwf2epGNicAQth03jQHERD2kSk7ct0531vripyx2pt4nu7/jz
j3VM7Fws8aMHgzRTIKxGVX5+cx9SEhqq3STz5NXWSnG80eVYzbzjH74aH9FoxuyZtAu90AWy3174
kFpnqihJqXEt8WtWQ8nURVNQOfK4Mf3rUrqJUfzd1BJMdIAvSIOmPyfnoMcs9q5oNl6h+ezAzPsW
CFST5qT2yKkjD3QIvQhlzVhVsX9GKaX9m3N00Nf41Y2CuU8yowqh61iHShWWvaGK1JoU39d+CkXC
BNUB6B2r+1yejTS+2K8YPcwI/vKUMif+WRLWmljrnwNyk2OZDLK2i64LGAYuU/t+HEO90+6jGXG1
E+MLW+aDk9bjSRmQcGBlmiaW0XjhfoCVBQSjgxNISgzw1FZB87GO+a16lK/npHRlHnri6088lVVP
aB1kavygyCIFGn0hcUQBxYXUE0pqGBBsS50ZLR059OZrPjS5DsYsnljxmia/t9f20tE+eRI+zaOK
g07QFtJBaaisocMHiBw1tBgEF3HMgK+njfn5F48i+RojT8jMAQcnSwDvR5O0CEhCwr5xm6l/ZmYI
wwQ/Wzztx8ErQZdaygFAPCGXfeO74G8burL4zmFr/qbBrxb6tnPzjnhT8OAYoJiGITm3kO2bVJ0J
sQnv/mk1KD1qapYreo7oJpICKcd1UZxb8B4uLM/Nwu55EuHseohm7Df9cmrONb4cbRWzJmKKGS84
Fd/uhrsjVnBE82Z4w/EJTCsz1LgxRCj7HavkRyJbOum4IQcLXebWYlx6f8Sc5Nq2CU5vIHMZXRW/
vCv7EiTx7JSTTWghaJAWdxJT/A2aQY1tA3b1F0kFrZRl2cG9QpZi4JQraDnZh6IHe0UjHWZEhwgQ
/Ox2ozNFaGiXgpZCiduQJBpNFRqVbk8wU2+LdBp3oxNlK5JkRARa+ediJ0No6cbyiiU5g0X+O1ty
DBZeCmzW9ZPo9NA7jRbXkKTiFoYqTrdzjGq/NiQJYPMwY8bxn/ErjlLDPrb/BPs1OrqdmTTzS7e1
bgnjAYJR5Aw7YloIPiyvBlqVKZePqncrB7QRyXn7Ys2BrF6YybDvvKOss5MPHAWt8LQNaSdXbmV3
g8eypzE8Kzv5wwq/AC7Ct9Fo6nXnpeNujoW3efemdTazjC+p05ehh0YOqXkGb1LSQ0A97PfJCGzw
a0RMCxZ4n2iZBb0K84y5s7CUU/aGGPovdS1xWi4+DL6grttVp8FusvBuOG59FM+T1OYJdhjIpSmy
tDMUaOv/rTCjdj13aEaMOzyMTy9PA7Drh+lUI6sSX/GhBod9vGbjNDzSQZ5weyxuJUw3YF4QE6UD
xyqsm+fLb0SMoM3Q11cWBJlazVj+SpyPCvqXTZ56sViOmy/057j6SUCMjVi2/bpkwpm9yajjh93B
ZcuHJWojG3an2+HC7Ak4kPFJq1C1wcS5EY0teRGc8L2+obE5GVyrm6P8RX0vyATyd1ueQckk/RD9
vNv/eicGC4ygKrGtkErfBZZeq0BycGOCriOf2B/RkAL01Trhqh1lKpUt9wHCWTtL2aVkwg4vp6gd
kZilStCdV1/2tISNVx2qiO39TTBRKfJ5yE4b/eXIs4BzvWhZSkoyQIgzXTuJnLYxnr1Y5PVpOW/S
fKzrQja5yjUZmco2pkei4YheGjCTytIr/a5FmaeKkJ+cQ66jCwvPfQ3mB79GSMGhmRWOZzJM1Xyc
/KTRCQ89TvQUTKnOhTvERqzl/3unqK9zKo5tGYDZTyDciUszg/sWey9J3Ui8ksTFGJdwAwgOJdJK
IdEYEIR0SIQC+x65W9fdkrkm70JaSLhxxVSkXd4x5ZpStz1kGIMQD7QOWiXKKHh3CGXQ1u83NJuc
xNMGH+DJiJJhglNeX4ElTYz0rtX3sCI3FYB2Lagug/Dsq6ZVyN1egdZSFz33Zl3SIf7dAs3Nk3eV
F7mRjpHyIrD5R90f8OywNrG9HhjdSlvTLfkJViDCcno3pO452O/Qmej5IggA088h97aj0L9ghl7k
iGhFgm0nVtuTLgSuhuk0KEUVxQJ3mFrg0AY49tHgWXegXRYw7DFncMEn0c3a2qpc7ehpVJ5UKALg
jJhWgGRQgK8OprMiNA2mSUjQW3Cq4+MIxixuWu+Vm+obzan1Uy1zIdUWYcMgkyEI+ApAxOBfvuRf
mlYz+RRn7wFRDYV6mo8TAU2lTOXa9BeCXEcl4d0xlCVAvWn/i9vioLxjEJPvUlImzSO0DwYeqyf/
oF0w+ob1yDZjXvyukPWB8NTuG8/TyHD/C2jTRsXt7NRdceudUekkAUfkd83iOfcNUSzWxubd6az2
jphgfOpJhtN269+retGR2DicaLRdFa1lqe7kGsu5ICrnH6T55LAR14zi66uUfe7ISsiwbQQcPUXu
aB8Mt6CRiOJdyMUpDzIotE6jHtOk7NBaEJ9oPHrqaJvtrA5GVBgg9DWcLIhyo2xwSpFDHvuLHjuX
nBZZLTQthjID226acSmTXIVvN8oOn0WVlTJ+ylp5eBANpVjMr6O0+okUlSMAv83LFw0AebeDtbeJ
zKb/QCWc7tS1sP86AwgBesrcd7wRzRN9h+SrX9vacdkFFqNivC7ilt3xAmpZnWsI+ynP3NknXxEf
3FK6xf2tNyBnIfiX3ot2rvtVu5c0g40NYFPK/me6mW7YjTrJoYmYVLDyyKxmfFnTslG1L1F7PlVY
2P1ljWBB7xVRlq740nF4CqrFtFIkE+28N0skeAB/wqiwURkRXNiQ19JN7/Cd+B3Oy8x4z+JB/nCL
XfjM3C8TrPr4Uz/fqILl320FmXTYvkOwpZge1z289UD0DtyhX9hqDYNmGnjtTzfbs6NBB92lYmEJ
Zr0KPjPJPbijYIiF9Dy96Vfgf298H1GPcPlYu1HLo2xwjTiRPYsyO1ZlRBKeyI1f4J3AaRiftRal
xDPreFLT2GAmz7LwPCDxYaFRKA+lW3x+7ipkflPb4vQm1GOCOzINFKW71Qbt26sPxdSzwchBvgsN
1woOItfDbPZZtF52o5PX3DT/okSSPSqtEau164VwO+GJRRUGS//T/OBz8oIJ7XvV7q6ZyY6EwST2
AHS7pBVnw4S6p89F5ZHlM2q0o+heIWsA2UYor4JjzUwZyNCzS9p/jIlnm3VchxbJ87bwIrRCEjiR
48DDTwcmJm0BWzhg9y6cbnfXJ9NzfwHfv93dJWafsiCVfKchGp5taZ5U/GpEacO7uPzLeRR0oHP2
K1ORRvrfxy1XpxyhmIq0Y4jOFobYUvkvTkxEr0rnkYtlONv67ilKz5CelLuQoNhkS2H9vnTkUNMH
LOHPHuGwZv7vW9AdSa5rYJ43ORVrrFwpdKY4ZklNUFWA80d41+gVjyjoggRJJ5aijDea/lLIXsLb
qqLTcG2spIB99l62q79Hva8gXtjG+WHDFWwTCc8I3h6uNL7BLad+eMXu9k6AcRD2OoRF0gbLIRyq
AZ/uXPuYDRQpl6krj0r/n4trZOAVqMMKgy0Ovz+6pk+oD9E4Nl+pEbIvJFuac79ZMqZTlSbAYT2K
IEq6405t3j+eQfadOZ6+kadRPselTRPIjmXeSMNIZm3bgtqKGodSXWXC90Mp2VtBg1YQFGy6bvID
kGA14zsBILeZIOx6xcbEmWag5uCdoAJoLP38OMh3DwIERKZzNTcX0ImA3K1FtN9bVYHXaHnaIVAk
n0LV/fe4Ro0/qvfag/znqUccwBxocNU2n+2PYHBr8pnNxNa41+NNlgKQqE7ke5GfZ6zbqZShcW/0
64JzMAqunVGe+B0jc6o9qfetkrxjSuCwxQGL2Ae81VisOaLUaqMlyj3YtIfjHPSANtgePKdShaul
j8FPZG4Xn39P9Jc6VcF5Zy5y3s4x1D9pHXH8KdGzGDMjh7J/euTU1X0RY7eTVci5JwRoxQr6s2AU
Fb+EtZ/vof7KKSgKL+eLDxhYLPU0JCNm6xOWetP8rR6g9nnBRo8YHe2/r39qRumqt3wb17Y6oM/W
LLB4/9gP3m9SMam2VluELo6ql0dfKGcX68EQEGAjMYL5xUziSRLgJxy5cOKoeAnmhk+RFUab5Mi4
hE0gG24CETrFZFIWoQf3FcGusYR466z+KSC45B2U16zdHe0fTDojsbAbZ5YVkDeRSfNCMuznIjmB
vaa8x5vnGxL2RAvv5gS0ig4ujRvE5Nmi0juq/ktbu5BER723/pDBN/59sw7xVObuVThOJFZ4cw+b
Cj1hJ+cP2X54O0DZPjffo0uHZOZctdKhUaIfqFfSrqNMcq72YhpHn1luRb7AYtr6JROt58RDC/3L
X1ilewew78si8BL72Qf+AnDsocu6BJF9Z/yh/NhQfSPlZ8/9V0YsxG3SrbZJxvd132c0pV6ySMda
9YzsnuRy5yMmczKtJFRHpOS+oJ2cfZ3pGnpnYH+lyX7WqZ03v5p6InvBAcc9rM0Vjftq48nDlszQ
OnABZZekjzT24+V6HrPjOfo3KGcHliwHtt9iVfE7F2torPrmEF2D4IrRmjmXPUgCTasmGm1oqh5+
UB8wQB9OHuAWpNBfdp28nLq3rssm8MHE5JqXfuDu3iedzhtltPr9rAfRGz/kzOvnHOfLoBU212mA
riuJ7QLG4C60MHG4JMZn/Vj3XEdNHNh0lb61yKavYYG+QKrpSFHPeX/usRVTD7oPv2qDeDMPHZ3t
o0Pat2Cd5T2YC+M5RNFCyj7JcyGaaorf0ycezWlWL9OLMJGRsglqN0Jli9mWBc7cb6YIkNafV2JO
Y0tKiowdRnuujtbu0i1GEXHRAqj3RELiQQjnWYT9N6Cf8upmjpgrf33Wu2DMDZZGTz/cU2c65pFo
q2SrKkNf7QLN5OF/xyKLt4hpObzAU4N54sF6HMTcHEsqI1zReowVUv4hUOo4/Rc6MHGSOiPMYZrf
5pqVE+BGWpLjkDkqHhYDq9Y9JzSeiqUQv6tzKQ9vDSLLIDaTIVBjWEBksWpZ3iQmfLrtBUzs4CLa
iUskBcE4D6Mr3+MWx2TDq4ySQkIBGW7yBA0SH2kwPT9Hwysj7RDgklHGOKYnwQtiD2HORIYGupUB
XRaDYCLdoNR9dkN6xyDjnd2FpDAO9vGwBRjgNl2u8ojEIE5DoKvm2gEPi70+nkAL0dBTPUhRy3UL
LsVx6x1MOdPHwmmjSu1ME0GCAnVheA7Ih2ENoFlXiUNYQosQKXWo9mBLAMCOifquDLudwbxrQoCe
5rdyMTtrGNkMyh9I8v/WEqgLRfCq6JZU1oUk7uqS98K/o7xi+AjNMs+GXxytSyuGe0LPjYNMCUAN
E/pAGyCoAFHlfW22YJYIxY58F5ZGTSaULxjItZLCofflBrmF0+HLgL9COvx36pmBefmSPBBgnbn0
asiZhkcv2pkVyKSvOpuNJRQUC6Zg8AQM0wLzo3LtEwSo4DeTE/1tu507RycRJOhqVyl+xDiKaGgc
q6MvjZCSITUPbXtv4jq76S0JW3cFUqJnbfPCnz3LOdHafRcdYwgBXSeL3fgF052Kw8x8uaCo3fd+
lUy3a3YToy761lI3KeABMn093ZLNdYF0poocqhpB1emb3l3dc+/iXUQ1Aa1TuZW8rOVri0yj+lF1
Tc6x9PoLSMzyQA/Tjt72T60mED+8SLRiuV6641VC9LwAw/1UxcAg8/3azIpjzwIeJD4A96OcQRNj
8wZFhjgVPAh7zLYBNENZyAyBz/0u2edg4gpVmvSNpl+y/ilhuxIMScrnk3eIq74een1lxjDKhT9S
rnvYQhhWd03+XiFq4y4KFi4OqudFyYDHFd10Y8dD6kbq2g/P3dkJx/xPZBG4RcA9dupHfFKhsW8E
yAbORmLUYgeS0t6hGfqWY7cCdVDXjoo/7/pMoSDKH3Y0p/fKga+3ivw2Z3B+ZEKAryNwPB2GqnBw
rJ5XOYhvW4QQ4mAl9JHH3mWTsLqmARTW6u1wrUzD15TDZWpyro7pTH4hi67IOQhkeB9yKUSV9ALa
ptnt6Sxelr6ndoTL4MqN91NjGDrKr5g//b6EnGGq67vlKIVtHpI6EudF4V9oxwzWmA3PG0Ss2mhS
kb8FB6aGToEBTzQVSA0lV8hNVgSw3hpSrH1AUKZx4ew5XwoJ3lh8RN1q5G5pt4WGCOJ+9to1/Wcg
/lsYuH6fNKfgjAAmjKHRaWPhqNPNKWcK15bD9+IZ+wmMrw9dx8QWLnIeLkbVxvPKIt8Xl6wd2eOd
XPzHXO1TMwLKkLsrhel24i/AdlmU0LiCXrhmmhL5j0j+2z4K7J0MZ/rWegkF0UyDdaNzeJpdj2w8
VcS0H10t+OLykFDM1e16iOCSxjPNoOltM17tKeacVw0oXLg13CIeMrS9VHffEMNdgwR5Bzpz4Zzd
63C8XcIcASApvIjmJxCgQd5W6rybT47ZE9sofAGnznEcUrEIzoT505fJQzERL5r3IMD9dTbqhCmQ
ieEeyXcpvv+gLFFfTxDBubIIZGfMW8WAd/5LyUfHZ6HuCfCLrZstnLctA/1Vjaaeg+x+5I0O3kt/
nltparKCTf0fmNRgj3Mnn7r780ajvRmIHjvI9QAa3Xi2V1xIEkTkg6H/6UVl+h5G+Rcj08GsKUDR
76wc4NBbjYKydPHAqjO8UcsRAlaBrnyO871Fgq3jrErley+s1goQ9TtjkdhYvaq7GPXX28U5Z5CQ
lBxl4w0RbDbbxoV0W7Pgg3ewFWME2OpLuTMBRUrAq90uI9JDSiHlx6fIh2GQaspjKUDSXmmu/Wqb
TuHclnOIhDEOKTCF3VWiloa2ywvdhzSTu/XjYXb5GJEede2Cs0G8IYF4d8Yfn5eOQXkwT9TSZblQ
EbwmXDLTGDyQ0JHre36vcZ3vwqqFoDIpEArcU5xVPIn23OL1vRXcLD7YggRTKps/S2pOENp7egZB
QwQ2gwIHzV4JyvEDxlmssKCzpJwsD19qUWabjYwgHW7to2JOQ9htz7dWLd09dGrgMq5eHNO58a7L
3/V8Bqp6ayfp9QcFbQAwx4+dFNabqAAaqd97NT0w5pwx6nwjtxumEf8IPAP37TMHHkfi6Yi/mlsU
IMglrm0eMiUGY4Ya8YbJDL4bgPJFB5JxxCMFMmGBRy3EhC/alH3h7MK5PKlYCyrPn2x/rFiGRaJL
UpGWDstDXGuUr6NAoZa7SjQfhqAL01QNsC/nSqV7eKwrapAZMiHuMAQxlPCUD/pJk+QSYbeq6Ihf
lBKNsbOc1OPt1WVSeCn/FZWI8giFde30TqJug18cYI9Rm3JajRy7LFwFlKuKHxvI48WSh93qxXKI
U8BS8MkmLDQd6b9WlE2/WhI87mOzctmYhR7uKNn5i4JLFhE1mhcm2Y1cR5VGNi+rqjtE/j5rXi6S
rJrD0xcvt1RuouuSGHVRT4W8loMD5Aekg/8dTx4uI4NdKrbV0rDco8V1mwoq9OzHX9i2XKG6zkUh
Ib7+UB6upNJo9a493+eP5znnmLaF13mThaH0ondk52w8aZqrmS7JuoES8y9SsDuyO8DesxSVi8gI
fLTnbTQ+QgmFMHI44f3XNUNqg7Wt4AJqcxQFOJGFZn7p2xxTpPrfqeHu51AXB2jLo2TSdaea7I4V
BQzaFFgD0xXoEBlbzK4aM2A+N1G0gfEQ2yWdKGrhYhSHcHkkKXrA1WYdM2FZwCpNlvf+WzQNojCr
hZRSA2I0qnqGtWxePnSzoERP+HsyTY8r8yBYjI21MB0xOraL6RlYmB4hP38cROqfMLC+CRhW4E0Z
cZK82TWIfuwUnIZPMn0VUw2fYJrL0GwjNooDKqH8nkwVrrH2Bi3F348tMLWokhsIuUcdSeYJyheN
A472D/q++juGLv8sR2o9kvrR/HqJR0qTwhJW9kQHxsT2ULZQXlhLMYgD+nXbvPthyyBKiiKbMCH+
LLdQJBifmbn8eUi9N9MmJSDWhy8yoju2sybzGIGS1KJkk0zqHFOc/0htDBXFuGoCBaM1x8bKk1XV
WiRhVv4NCIL2inCZHU2mHzqg4Cu7rKBjsnJF/8Sgj5Fu+W87ov/m1ukKC4/5OHkiOANeK3i4Wdw6
b6YaVLxWnw+9P0uUsy2h9lefd8VEAKwmSz/4NnfM/goc5v1Hds322CVRakylk2cTuj7qZiQ5pa4Z
AzWxgACuLmddE4pfrH61O2oDiXXitHz5ljhTOzPrGUGCikabfrd/mn5IsQoZY/KtJwTeN/VqLrRz
UDBRK2zON6J20tttpC4iBesupdX6eoVk0++vJrMv8PMD+uVhhll9+pl9DE7AS/pf6s+y0O9SGfbz
jFVXicb+0qoi/8T/ihNXV9XkEIwqndxRJ7L9MuwljF54RHoegNFJVy7dVMOr9dALFNCSy6SlRjLS
RbmYRsOX4BkSLK2HX9rQ+YPiqy6J1mB8Kqhi6lYbtQCOL8m1yOWRLqHsSGgakptWqeqlyHy/jZqP
yc37RwVOr22x7Rj4KFiyG4q8VF+fmayv1fuBOJuXUVa6Zet/WMW2B9JJyx7viOwVFKzE+hhhCetW
zTNtpTPzw73sNWRoT5rXYhaVunOz6rdITGUF098y6tNryHFynxYgbja7pZBN3REZn5jX2S2caA0I
erYgjGqL064TgP2sbxyeUrNYi+5dOSF6+aPatu3itpQhMrKPfWxj96V7ASuL5ZRx+KS8D9NfzM5s
wKps92SFPODCMfM1NtVsJ5cWapT4NZZUk70A7N+hILAl+y3J+GAZXo9sWbUTfDLN4Kyw+KdyHwbO
HDq/piGQmu3Hx0eNhn1CCUmthisUVQbGoafFUcJQoSqOkz9QLAPyi6RFuIe17wue+wZc95DlJMhL
wIS0vEV6rdB6eWHESM3lYOg2D07070mp9+cpJXVmnrpovz4grSYxKztlDZTm4w1oj2Gc6CVMzNvd
Lp69p0kMGuuk1ey4AmfMR8YHPv2TFDMSxZyUJR+/3oxVQ7PKL3Un1wzse738CPqaPmvSQ0zTka4P
rB398ZW326xD+yfJN3aIAPjPGiaN/hAkbC0HVPm/ivR0CzZb1q93DEvBZUb6D3IcMfYpC/dX4x8S
Xe3qvuVIfHHKWVTDwnbINgOV1DGSqtepHZ3L7+6pcwpwNAfk1CsNOckXPZkyBnUmK7sQbLN4xEEd
Fz/PfzCO2GzcydqcvzXHDRcSx48cYVPsfvU5zPDphtqvuyBSxxajhLzjglVgkwU6ejiZPV0Rx5+g
9Qn66BcXogNz9BbTbEB9s3ngB/RYEd+FIQHtDcSLLrhjI612iGxCMY5lnw2FS5U+fBbqH3WmeXUp
IxiumFXo7Vk3eeAhOXdyyoViD6QsaOxI+HcHe7zFGAGl11dPinvIXKJ7YsGi2iZ1ABYuTDu/n+EE
IlSYbAzDBaUBy8XSHalsYAb9clE3xe0slFvwOVTHDAMQ95BAEax4yVb8JqKErYfZWD/Y1pNKOqBk
WXQgUe4bEYWwCtESSc8d2RjJe3+Iq9g+y1YkAFKZ1ok4wbXaHCgtvlIl+eDOxFl0QtvRbi0D7ZsC
80HYUAkeRnUZD3s7eBJpSuH3eA/YPAgmTcRRYV5h1waNBRGomsaxA59j8hGEM5rfLKBKLfBrr4xc
PdYfDT637S+qOjr6rxTlBJUi2LKQZTeoX04mplZasaxLDYU8GVZHHXeuOilwZLeQO2Q5k2dy9re+
uf46D11cdE672Br195GlFIGk4VhBPOl7sjAZg3tAGO2jDTFAHLBAzYLXQ0C6FY8dwKnQ8JQfePir
yoqXr67sZeWD/r+k+aF4lkystNmcJ3K6y+Toc+bsNdzWQjzS3FmO+/YleeVJEOA/TTv24bk7+UUr
lqmEVMBM65JCcsN4AmelW+jpEtrtybtKSPXjuR51QyFj9Oln02qGss/a+vr2oh7+m4eWyWMmTHHd
0Y1CNDTkjnZGZ1fyFZKO1Z1Iy9Mf8949JnRlUrpH1u+BVEOFVoDxe8E7sj6zNVz1QEIVbINIFkJi
eodvj0YKQNHS48aCQb4JuEY/YDuk+/nce96Ft4k7uWwItN73ICjmMCtdNmJ13mooEmM1ZzQ1mAAL
nMz021exHaholYMZ1yFz18QGupYGMOjuMTaY2jTHFF1stenhg/oxY0AlnzeKVptv0BJFx6Ug4kpy
hBjQ6lnif1crYuG56AiTHYkig8yB67nXRcTcGYSBL/kkzw0zPtVTO0q1/S8ix0x4tSziI+oh8yFG
NDkYN58A/ngiVqbjv6+C7o1MEpWA5NEHXjNSbmNX+imW9lJOdhCbNsYeFGK+7ksnrdUQL+BoJvJI
gHBUxYYmBxbEDlTf7Sp5T/kJFKjIkjI4jdYiwPARLruXZ83OArXcOHP6Wwz2xP5rubpFser6sgDa
Ge6QM4vD9haMoaBXVZhVdjo6OqUKLKyE2gmOAIihGKcl6SD70TExSO8KCQe8xdqU+xb7NYjXqIZL
+PunjKPINPV28G6tMizsTclx2d9/d0p0MYMEOe7qz7PHzDwdt9G/U/QrpimG5+kk3H/hsR0eQYq/
T2A5wYqtR6W8+v00BTWQ/oPiFlaHPANdHO/0gtb2fSWmx8VCh+6ofHmcibGM+GEpM+rgRXVRNw3x
Zfv0Swk2MCsReNTrMcenNOQwR1ODoRfDM5e9f0fy6M1lj2XSRLlycCwkUL28NEI8pEBp6vvclpMF
kb68ZBSwNqd3pvxrT8/7mDb5fjHZx+eDSLvnSnr+K/T1saxuSSP5Ieh9VNRvR4i+aKJzGJmXNlIc
da4X1fKBPfs5WaxCw05PKNGjbeDWo/UKDHnOvuRrR09VjI/r1Wx5hMSfQg6iI7MMNFSiTZgUof4b
seZGMoTlKpuD3ipAo3xhtBvm/tKspxpR2ozeCajvYS1AbFjufEt0npslKiRy2RLIAbN1d7WBVcth
QCdebSLqfnHZNFPCEcbroeEza/r0paElWFrKabpUQ0i5AiAxMp2I18U08D3ub1CJoyNe+vHAm2k2
ei1sx4ZT1KPJyXAcR5PkgeRzGvTtz/2dAZXv6wqhjRcnYBknJxXJvVVRFg0u6kQ+rXEFcvRsIXA+
f2tkG79Jl0PY0DPCzOvRNGamt3wdHVjNFxr7T9L2dREWl+11nJsc+scokMQW7chAATEsCTo05l3f
p9RKKSAGt1Nov7MHbV+tKHVj5xYcJIAkrusiyybUvRTBf0dFW32UxQIoA2ooMKB+gJigOWMbOTEv
JmM3a69mJCUj89ShOPYrxI+8wWQqLryY4SKCMdzW0zeqUpzs4caxscTcvpS90T10n1RA/qV1D0nN
IJ5/Qx06tXMuLntoih4zz92kgpF8YkyIhU4FHTgApGVeN+QRXG6bWpRCxJIXV4KVBPC0+2I8DlQO
01QuaUBTqPxVPfoDq6B0aXlN/SY2QFxvpb0LtcsRy0Sni8rP5za+as+BulEU/FbGWyYXVW26oa+W
HIAMRRKtjQK1lmiVpH33jugtwHjj4VUSErs/kCJg90YFJo9j9T2XTzWdgNNByvxCFZ3ayiG/DzoK
HOGx5D5RrzzgUeAr8DpJKfU2wPP1boxAVTvalRNcs2kj6ldMKQhAVS1EjdUPq8f2WicrHcHgoo2V
JXA2I3HECzvAiyYlX1lMgduIBk2J6tlYlxYxqmwBo7IHAsuIkNB/Jzc7+PqkOJFkrJjnj2RKuvII
djd5OrbVlH6Hzx0eLEra9FVlzlSqZ4aB9SY77xJHCkknyHCmlnmcnaxPiBN9qHLgt8DKQAtVxZIx
jqR8UFYJD4MkHsAaLgS07nMXKxFbxbsxaFcntIGYZiRciZOJ96c8O/Hzx2f35lC1WXf9+t1Nv8oJ
6OgAZgeU3Z+ffw1J2JQvVd4AqvVc8YP6ywxrl6BPvySVB7hc8tF63Ps6paPxeVjBA56SJ/gMuJqr
tlsMC6QNpekGcIiWb6oNMM/5/CVLhqSEim83OHjmaA5Y2zx5+rhYjDNFU19gnr1NX7iBYSgMm6rA
ATZZPradLxHCoCTrE8Otpzrb/s3R1Szzc8UvAK+XTJGbmeQwuCrwseIiyHqPK43ruaZ0sGfT1BsH
v4d/DI3JFOqfDKqzD8csuGyjYdYYRgEmkZZUqKz77kDxVguRG1WnM2ajzyOk+DhAyunMRcjPIBgO
8+so/yddXziyR0XpuOG3s+o+Skkl1sB8PGyRhzazpI041BlMsOHHCbTpgF/nw0QC61N29nx+DYZQ
shZogRuBlGbefLifU05Bztg7keYX8cISexx6IzaG5I4MAl8LnGShAgIhXNDRHvo97jWAfQ6wJ4Zc
J7GLmGyjs9mgyi4pjsWNzN5uDcqyoXiyDw5vCUo8gqJy+6Ww2eKykGk+AuscST4P3j2hO1FIl/Wr
+rVh2NSHUDA3v8cJmEb1oSlOcOs+8abBpKb4+zoBdWN22T6+PVlDW+FbnY2xlB3Af/rwWHkMgwyu
Ls7sG21TWBCQJroUGI5QUcQRXjLoNAwwW3a1jmCutFP4GULhaxR13Wbxlnd7bZ6Tb4Wd46lFveYQ
i/2DMVnF+h4jfrsL1pFXXVPX0bizZWsCAFjlHm+7lah2xFCN5LKMRpFp9gEJaCbBcNCS0WKHL3eL
VHNwZ5d0AokGC32NTms7bn9Vd5sLSH/JiycTfMAoKhuw8xZbvQbBcjXTSNDdTM/8kHiAtkeAiE3h
wid+ZxwMTntaLuq0oDnxRc0HBZH4zMH6ITkGegOFh7pS9onI+QobOUDI9tBUKDJrSC31yycsdD1K
aeiwVDPG4WibAmbATb1lIp0Rszopq4KBgop6m1q0ZTpnsa+tJ1NuSpeWSF96q973LYw58wEUQx7j
mKU42SlzAPepoTCrfyFR8JdTpO9KC7GY9Lx9225tSwe59cEk/Tk38M8clJQmK/f84lQ+8s5BmkwP
eYUw+tgDmgS4RwEV19Wq4HMTiyT34MI9LU6sf3pdV7dt43bUPm6QhDXxyViLxLUPcqd6G2UPtHBC
Rip0Vl4r7DGKFJYmbte8rAvLh4Fcenj2d/gfqD0TS3pzmzC+malYMWB3xmZmI2HjirVglct3sCiU
utowYrgK4ChyuBI1uuKuR0czwt2O8Kyzx5zdp7itPcFAGdQEnqxDIsPQOUPKUQsvMEtUfQeAfp5x
HKFlReLFcfxEGFisv8U50Ih6+fzXfsajR7/vQNJyp7Bh6iQh7ZYPun/z+D6FeUUa5j7AIRWy6y7z
Vu5DM2CfSgKGrXTLJGmUbK6toYfUzFSVbRdLXJNPjZl99HaXA+ez4+g6t4hTXIOBtcFRlLoJAyuQ
VXEqtupnhpITU87xkhcEUlsYhwETyFiW5mS3IkLUBxUvBMlfszUOGEC4veRWyTOcR2i89yWxkfpG
2A5W+JbsYz4ISfsUP7H+kyarFSwUgk93/o9gHO9zYn1eJcdEiMdkOtQIAJhLX5z3nJe8PSF28tad
5gmTC8DoX7IsjkmiE85xAu5PW+qIAv84c8Ofn+R6Bo4PBXiYzSnWzQJ7VSkgv0raPCnmTZZb3E8/
ksYPfOOXKshzhC82xmq43kgZBDIdbHC4YEdm/HpAXGtgQ8GkNeGrgxeyH7qeE04LFrghsIHP/1H7
vwI5vNCqBqndC8P91AzZNocNr48/odjCROllnVlAExSOJY/k6ce/cHNA0LovXtXnPBxyfkVVqs1t
Z2jgIyQ8SDx7R+Sxe8sFaY5WE4Thd2x+DofUilZoz0BKfovlOg4GOreJMY0bcVBWfFd5Th0syEAv
aTS/wX+MPRgGf3e239C0SZwU6FXbOKcOV7SkP6tnkJS7LIC8rOzIGvxD1UkR58wsElxG3q9m8/18
4PKL/6BdXAYInQ+cHfl1/rESy0PgGIUa269/dsu2ILJyokXPIzSLNUnaaVZ22ArtEAXIZ/+mszwu
V8g0Ddo2JYnyiW0I7igHXlzCg3wqa+WhoqKh2BZdXP3KaoXxzqhabzGqfQCFhg2V5aRBykydLlmE
eh5B947JimulcfzExzLJZSXgfdoQ8bkDOlKxnc5EbamPNr/0Ho2PkkyJLN0x+/6f20hU8VqEc+Rw
C7HwA/w50KRD1wKuM5+64IaKiLPvbzRvr/tHnY5yNZJ1O2AKB4nCR9zVA77Pbuf/PZWqWCri+ex8
WPPDRSRX1qhD64fUkYu91sddi8nmAmKk2jgkXOQIb7UbL1uVgaUGT8qzDTHhUQSb3FLL+Ni0wfGc
rd+ZxP1O6B4qbNDY8iJMy09ylOvJhjkQWumJQWeIjQDFpke4ROSPyc32uunY19yiFiFgWg9YqEH+
PASIQ3sFP9Lo+Qko4MfH2C9Vr7pf6D4sR5xxX9VB+cxizLlCJRrhrCNp1IYgj+Z66L87NZtG3TNN
ex5XJqGp15t49iKM8IldIvNeSLq2piLuqqw00IRCnBbc1bCH6M+1VaLwKZJqe+6f+B08Szd0C1J1
CBLyH1xafDMwdjMC2Oknt3G13eO8uYuNq+VHBwEUE4Z19p5MNEY1XZWzNnSQnSR9CKjv3Vc+cSjH
g3ZJwBco6h/vPGp7y8So+i820ZHw9ogqKZbB5qbbivK2s2izuDfBKz0uFfo1TFVVMkXhJBmwLd7J
zXXooleBSkBX9f5meESqeUm3Yas2nb2IplKFndbNNTSFwIVSgxLBkdjlBtgoIwzOBjOte6tSDMtQ
calgvmVlsumJAZLHdA91lE9OgXe+am/QkqeSNCTW7DTJaG8+uEnBzKoZo4elnnBjmuVPm7mv6Gl3
FNDg9yrAWrLg2modWlNIkl/YSsdbbM8jn24IwajzpYKzsgFQDo8DgYifL0LohgA+RdIk5L6frQoM
UQGf4LZq7RZkuhDXjYKsrq41PjODF2F4ru8ZbKWjAGf1k5hpaZrEE3GLcqZHZTK9+Vzsd+1EzHqo
5PRgg8MbcfYdk2Lk8vZlzKhDzRyu/AAsFBdAD5CsfvOVMDCV6CFEyNQrRw3SUuZxoS1cUz1ytWPb
5Ip2b/U9L1sy3oWvCYVhGRXW59HgBtZCQgLrHLwquDZtnSBYb0NYckQ22q9xwB+dE8lNlVFtpFnT
uGy+EusSTHNqSIs/YUncy8ekIB+uQOIkrXXx0V7EmWpPUFdQ+xxyYIzLZ+4gEuw10TbeITqoaBXY
uUdXnKLRObndA3fZLo49IginaJDrbQByI8HR6s//rfTdEsw7lcP4uLcYwbeQ5eGRJToTwxIdOYi3
ALzC/5EemKSeJ2ztM4Y+qhHWFx1WwmiVCGYFv7YtQGIdx8QYj1/QhnKJ5MhRyL2FeVuMRIDVMl2L
ODhAuouGw89VYJBVABa7gZtEVozrMjCvSY3oPsTkqL0QSUwDDoTVDAnoaUWcDJVuRzpGADA6mtNB
Yc857NyP3JeH/PJFxA21AKd5s84j/qkm7oYa21l1tb1FG0oaAlAm42tWroQOrEDyH4VZOx37mo7X
JTejNeSgxodO5yULB31D3nRQ/ko2Io4I69wSfB/I4dAN0G4eVeiugPm/do8gKVLUuwZkQFHqR3AI
V54h8UWlZV/ekWusjrzT001uGwKVAFvZcfQou/m2RPQzlkgsLtxrIXQAY5CwYaNQzbNHVONqgZ6N
tPv2axryvlGA8VQFbguhOe3KPfa9Ciu50mp8QbHoB7ZwYE99fLfuBCFLw3zNp32oa3NFfjx93tu2
ZXMK/PWI2wdN2dbXtwRjFutgheSXw1XWMvG/VCn73FlAPjwIJMGa4LSke9Q9dp9FQdXASsct09WI
/5qBT6fYzz9+rq40P7RJWzmy9Q2pXnLuwKrvwxfblVsjPjFChDbkcPgEY4JPoHLatY5QIok/xdnD
2vyHlFR9NETqBiwOHTTR//7hx3uhDFn8auV80vxPD/waPVF43YMbndAqHd2YKoHZxOxsF0iORQ2F
XGPKLj6h24g/9DU08llNwifNt50w1Hhj9mk2aIyT6v9VIRyp5/CC8M6qkO96FJLW83Sqe+9yGgzM
bZgx4NLxNQgnHQ8ywGJLhncT7ES1ytIQUtVLHT32F1iCMpx8bs3nBYVREIsL+QK5brVKMvv9HVIv
c1dr5QlV6WeIvZ6FN0mqL7cwdzTvLWU6Jgp/Fxu2hEALzhGMMFWmklt/Lk96rqmOIY/gpj+mdBfj
f/4eE5h9Pi/6R4uRZvLWPIB/x+VOnzZPfKDkrNNCU7OY5/57EFFkHoPdTphsJhK/kPDbaLSyktrV
gtJ/TodXeg9c2BeTMb2BjywNNNtHCUYXSTvh8AUmQ13TARluGk+cHiYJ4GqBwzatkP1zwMUTVy+Y
ouYncwDqzMPK0FU8ZLPOlNBOSUlH0v6UxIK2di8gL8XnwTEpImWP4s4Z3WgbTTb6oliSpmgmjtBo
3anhMSRrPeeIsUpM2E891f+w5/bcJW8HXcLo1WSIpLtT6pogfRq7LqIhMWO6c/wduB34jai9HnGO
3NbOzD9+H0+vKOc4rj2WXhcB06LetlySY+Al9VW9NKfWZYHzPnl0cUvnLpZsMzLW00fAUMlIXuv0
WYD1G0tXlTDHo7WWrMeb7joECG1ToDsEhzGatEf3ZY65Bdeez/EyC1I7cxB9K0deNkOyE4jmnlfT
5ZbAXD5FkuICVFiVWSAFDcZDy7ohnR5Gj9oOzbQnbH37pLpU30rLpeqhsVZwFVT3p6NfAfLzwEhb
S0Q/L8JkoDHjys0tWhRGcMBwjYpkbfJlTNPIwdICIV4yPAdKYu1lhdPoxN+oO0iPYnTCuao/yan2
n64sVceS9sUM186GgvTBecAwfthQhh9/Eem7h7S5pw1u/MRNm4bzuMpguZcOO1ElV+kCz7vbcvbP
XqEcx0DAa94tRvXQvsLNp+MB2ksSUQuCO6H699fRQiUY0zqvS5Zz6W0EG84zcKPpAL7uJnvQYRA+
Eg8+Of4z20ZUtzkvraGYWdkS5vjEkRcgAUV7Kdj1kdria6hOP7P7fDFnu/QeSLX+i0MYS9Sl+lne
yTLxdQ34Dx/kje7XKi0Gm54Pz3wom3zVZFOBOpkYlGzTParvQDuuKRxFpoBQ348nuoxPqetghwqI
9TQRZKr7851vCEun0g0iAUBpXqL9vi0/hJYO0u8owJK4+gIXcqrYklfirs35Uh+wNp5vtZNpmmC1
meSb4LDawV3ZwuN6d74iDk6WS+jq5uceOz8SaNlqmgJ495LIr86t6S8OE45uragu8H94NJXtCfFJ
0Gfgsn0M012/LgjC7JzKhyeLCOqIqOs3NdmeeKt4jHaMGwK/pjw/MWWHJYV8lbnf9nRHM4I0/Yyr
W/2vsS5kTTuYV05x+2ZRblawnxuqaeICksGvMu6Z2URs/TrI6gXIGv9lSNeUwm8R2qQlgKxFLi3g
ZW5bMN4UJ8ZLK+/H1T5+yw/LacOAUsgqTUm/cU51uXFQp0LphPmkMfZmFQCvraHhVKz4fX+pkEfL
Tsp/9+mcKxHArn/FfoLBN+BwrxSglMuYn0m6zjiW/4wKvjts9lZHOboJhppcDCFWP8WbTH5dOqfI
0bxeqAOk2OhHAUsGD2zGQE/N6h+hm7NwmcxiRGdDvAwQk35JedHdzo5S+XaPkVuv7nXDuIgN8Wnr
3U/X0pVsD4BK29eQI+yjZUPqYI3/7RiIw+I2x5edhtSn1HrTWeGOykpJbuoux6wU7tAEEOP/ZWTz
mg69HlgtVlIGvuvNFsKCSdPq0mssXfnkN4MXLiQ5+eo91VD5r930BFQRlpk19tB3kvQpS1hnSpCp
N0RetGu4eXgP6O16tLo10k7hXw7jbUBvUGgwURvfjHjAZmem1Z8DM7b1cPRXEezXVZ8EGiIeKcdi
x/F17NnVqSJ3tA05LvQHxi5cE55IL1AEvKeR3DNnhdNdrMu+SjC6lA/W3kwIFCT5gcdi1fsQl69X
q1RNcdIPBt4lNMQHcB76kUEkPl2GzZLq5Kbz3Nl1XzkhzBP89Pf7S10QoKAnBvWbsOFfaAc07Pb5
AVdNOcOhJnHLR+JqxrVBnve6sNs3H4UuYTCNXGUJ9p8NcC/Ynaa8r8v9xrGaBddd/uVcx+EwJJiX
MNHiXXaKtMT//pkHRBFRjXDTFSCzp8sh/1wpwIua7mebKH0FRDB7TzRrrDIjoTH8Kph17LsVCBZw
JiqJZwmFAqwC/rN0iepcPNU+IGyXGnf/1f3/5Bq75q14SYnPhRnRqg3D8QsrpUwHqu1Ys6Xk6Cfr
IHCH25EFie2eIEltOBd5CV8Im8CSY/oMHmUUt4lMiFaqkGekb2jg3hZawEAkblnCjKnYbFm01YWP
+w7KxGNkD8ng5eibKp2BRA3VolwMeHVEPLMLpDcNwfcfszV/pd6DOrM2oFIn+2u2qI+XxVQC5uQr
PuXsU8+B01yTgHJ3vgGOWEjJaxgqA6YRkUXPvPO+kAyczwJGquPCEF2/b5wW/PJ+DTBr6aUmLtby
LCdnp5VF5T3vqu/ayUk2BoaGlbQJSgBUenEXv7q95KUUjMKp+Jrsf55Cwnnbbg+jAMLy7QBfsPKm
fKlMsd1QcCDUmrucrLeNeoDxpWFV0Az8B6oHuttUhZ8DKcg8qvvROft6FngkSXKG7OAevY8y/UVu
B/pMCuI32rL2gI/1HG1m39tGj1TA/io3FbT4skl7o/4DD/clSfc3MMUKhOrR303iTeNxuQycvTff
qUYEc+8lQVEepG7L+P8RAR/NNBFHWNLdkIgdOnryj2s5CuqPXdMZBu4dx0DyCI8LS2f4bmOdZbLD
adUY9Ax6Ffk+oZvIMheM83SzETonOAgFC7zsQwfSjje9hmV4EoXqFQNYaRbC1z1QcMn8+Y0trBxs
OL/0FgzckwcKFGBwdE0KEOCj11f148nbyFwkJp4qtK05PG3uqE/meuUj4NuH2dFHzZfaD6WrUdOI
vRRZv4EjB4V1AHS87TL1z+KnbgNqdUcNMbxaN/vpy4+A3tk7Vzrd7N1p+kZO21EpF3Eh/hYMctyt
sPwqUh1WJOsz3eJdI/e7A4YAX99giDGH/RLgP3L9/5fMU83q7FNRqGthVzGv8ZmSdfBTUbpG6JJ6
pSljWmvPbzBwhKA4VUOq2JR+25is1PRlnLAnDItuVVz2pi6btaqxol3NdsTceF3WU8w+mMD6WgIg
SidZY2YqwSGsctHev7mWO8nO8vjaec2FbwGyeIemC/evbPWG5s2UnK/iOMZcqoDcno/l0bSpZsVo
9tFmmWvcWMKeFa92LBnm0KiuvP+L+f1g+KB8T7E51Ph9BI/pAG1berIGsvJQAV3AWePnoNf7+i3G
zpI/fpeOGkCOU+2TteURlPOv03LHxpjQ+m+SRcRLmVA2WBvE0gwyuXHwBWNjJIlQmN31G8dOzWoq
47LFCB6Cd9hJi1FEsaQ5pSeGOsUyTQ3wowNqSQTGyMtA03pp3gq9lETjoYdu0zZi8cs+o+EDKvF8
bg9/SYplmiU+8X4DvBTH/cZFCPgm6C/6DliH4IEqyw4jCS3qwXIvv94hyA4y8JPPXshtsWaw2qbl
aXIed1QFcucW5MY3OGFcd3kQUq6fMleCLf6tatlcpzZtk9uiOQfBVOiG3aHoEQAhTPfUhJxBvCbb
PYUkKVE+Fml6SN8NspEip8S+Fi5rjKWb8m7I/PNUqhlL31xsrrrI+kkjuK5458Z4A9/5eNRmhple
IPr+GlqkE1RoDjra3p7hz5M/R7paNmBS/cylODAq1pfQravOWWyqh2OXgqCw5bXFoRFT96y9ZXFY
Rw/qnS4S2I/Znm7pX9uCruFDMwCAoFRFmBbiKRIUoWJsjXd/WWIsra4MurlFHOOfKERlLdMWysiJ
kLREjEJColIY4sMLHVA+Ic/uiGy2gCMcnLjZmDvPALmomynSOJLOvmXHDDppWG8oAouXWBDgFaRd
Q9yxk9N6UD9LpXLKr8axUTrS6r/40gZDTGn6k84njfIMt/U0iXRahJgkzrW3MaXJYtt0WgYxr3aQ
0w/7GI/VHqWW8YXmIaaowzLEpqyOW5ZlcXDSaTssNW1DO9Qq0vVEYRg8dmh+yUy7IE3N50UFDdIk
ZuTIxmy5A9EHb/bv24Jr0bTYduCZ/l4W3TYNxdwYelps5ri/n67btsX9fqpPA/Fo8Yh5rFRc14Xk
y7q9S/HEdeLP3zvjf3aUdMu3mAXr34H3blo02miUpfQaAcZvTLUjnnhkJtXViDGNwsAxgVlUO1ld
UIyy4MSHb7bI9rnqCw7e0q5F9DUXuNDI+0U6/qDHgtDXN9x7vIvjCtIBdBL8pfZZ3anUN1UvH2jY
/O5YV9qWvD1QalU/Y0xqLrcbr44ftONaQOga/JMmNgBjHf5e9HlOpokVP5awtCa1VBd795QfCd+h
aOPNxSuUy5xiApibYBXqsxteNAdRw7JE9O8r3eTURTd7tMNSpkBgHnkEntqNe9FRcc5vwygVQOL+
Fvwzolh01sGMfhxAPO0y/qN1E0WaYtuMqN6rxkKgB5EhtC8Glw8kRaf7tUkgoCGwCIYnkuV9ZBwt
3i1jf5vYO4Fo63Qc4rnIvEjHGlQvpk+8JkIRRq+jOW2N2tEwE5ucJh29ICR6/8QvOCCybofmcF4K
SKJUeZ4K7ZddS+OToZnZbecsrn/uPh7c0m05agRa7/QNkGAgS7KoCwUYlDWzNQ5IOEbCObTQbfmv
qbqxAr/4UWQCftFObf4p8Rn+xhLD9k8h9HREHvu3R/XSj51tTIODIhloZxUu6T3FqUvC9s7oG7tH
O2rFm/98SJ5sK1WPkNv+L+SMhsEO/EHJrRWXZAy2OV8u2O3dXCLJ00GMn3BJu3WiPLUmx3czQ8Rs
/9EYMs7VLkluavl31BX/RjnmSOg3aKjmbEirjU6YGeC9zhD5WYU3lZS1ZQxIw2ThbMFxuZ6bvl3U
OdtH3DRuYBLHNhsa+oe7g7j8STOzYC+FFOKWYgiy6U0cl4yNWT2ulpmWFLT61BeP5H7LsGFynfr4
rxh/50n2Q8XpBsv8R0KKJaMXWw/j3CRor+EAXtaRiXVOrk50sCkKCKAMQudAr3Chabhbvu/OzUnu
I+wGsMF36Gn8Ucy/Z4ve3PHJTIoO2UemOQakYkfPAQIJu2+n9pYC83MHEmc3H/E77dKhynKPRm5T
fHngAOBB7j+j8RCKWzNCTyreVPxv7oQatt2BQ6kzyEQOxtwfTgezqzJY4ao3ZiVNDqiKGfgtU4r6
5MOAVkPzNNZeSB/5w6BRiK9a+bAPNj71BldlHw6nyukHYrroNgcdP1/kqThITMh4opE1A80YjXVN
CxzovO9mgOOrZz6AORFGOjZsCo0FIn7qgD05SJTQJIXBcelEyUbfJnQelGhe0EFnFdot3VU8AGTm
fY7/XCax48vZiutG0HONrzAjfxfBC1F6UXK10NsT4lqR9zGbB3UAuObcxC3/d86srecpaxrNJ8Zg
soiAWcRD6R5+Ju2yrGWkdiwRDE4Yw6rSOhsYHcDH4zTp/AWCYur0xZJ4P4kKJ7odKYHRKpSlEvZe
6P4ulfo0a3iQiZK2qVdLimk1lg90uwrgvEtUQqV8wuKuQBUsXQUHNpR3bmohqZBoIg1Rj9hFs+fY
eIlLombnqpMQZOBddEfF4W/Bkhn/KAFTyZfV8rZ2hiXAS2gniMJteMpHuMLECZNGuM2GPUAaqy7v
0ItIcA5wYPEt5TcFeDMTStKgdZ55tAEvuirioQJhwNrnXuNMp+SATXtf6f4lQxdDS3HA8v8Uu57n
rT20Y+/B6HnBpCVNNPe6Fwlj8d0JmpyI5jV59bmCqk7n4cwDy9QKV/n1eVbG2NqBTXbmt4DTAeRC
1rsgQcde7Hkh0bbT9hlmq2vPPCuv4fkjSBXkAHWuIyMOurQ63kvm1ZxJxPkflBItNWlJTWi9Pnna
sjpfWrgo1wPbTP4ktsor2NS/TT/CqAQiJA8jiqB3vpEBMse2mahPB1yh36LSUmk3Tbhy/EtyQQ6z
Ak3fxnK3P+fbzzhW/EOCK/SMYEUVhaj9+tSfusDido5YaAdqLP0Myq2AKq7mANeiPQZjxRKXejfS
cAFDSYg3KmFfB9767rIChVjZgU2RmCmakz+ILuV7F0tfmhpFy2SveWWpEPbToOJFaQDqWYTRQBlE
zP9aC5GcI51Yxeqtsab6yxF195fTWeVUWK/jIOvB4t+Lm2mnvL+CfLP1hqeDxf3AhvjOyRVSj3oq
F9kPoTnr83Pkz2y6czHWZrFOoQWqBvpwkdGj7YRaHM5romtOxB7Ha52BtMxO3qcuSuVQfxjCPjB6
Qq81z+z307qHBB7uhZ+3Ul678O3JsZGIhrlHS0Mz4CdQ/yPLckAFQhGI44KAOWuJvElKkiTZwA3J
whFJgDVWWdE+rYKpV8DF1Jy2wsYgPf6iKUUcpBtnDkR2Pg/SPyFb5L2Hbzz1nasysC6JpCQ1Wx4o
srLmhHR75VA093RZ4sjgQPakwen/BiGFCi5FvTmwebv70Ch06Rq7pu9pnKvtcUkkkU/lrXqdPhAe
L/t7XSSM92QudiveeF5bc8NpobDp73Q6p3CQe8KW3hkuNWn+0QydaXfLVk3sqkiqzJtWhCoIXiLi
5j8CTIqQI5r2El6xb0jWiy3Bd6SUNYmqtyLXyOYReiv9p21/QDP7IZ4IYpOq35xMcjqbQfXGypNC
3Xu/CiX3v6bV1YSCjoolISAJrjpg81xuV5spVn2i0yw1bSwJ9YcJEqv9cYN3QGpcOb/85w6RpPEv
bI/r/bx45jkPueISMl00lBu0Jeohr3kTnhdVT3kCTwh/5iD09HX+WTE70hyD8K153tpo87Y/10ZS
oX0K2TZC0FUl79xruzTmvHuCOVj0cZT8NQWZGNi+CezykslYkVj7OA8ecgcphEbn6oTgjpLhKf89
MWSP1vqDE1k5DwbB5ULGlflT12lZtR+7oWaYQrynEQicAKn9iFiVdey0SNjbjHOkl35RndhhI5ZZ
RZV4ku/G8K7PmmzZubiZSITRyJcq4SaLvY+bxWyNa6u0zLMYWc4R5ZZhxOJua3OB3a1OwuQ4AUIK
sc27Qarxdivg5Gf8Cw4m6k7r3mmYi+IsjKrnfBQ4+6R3GfO3MFhzmAVG5IvzCDRrZgVvU/yNbRrD
B6bnaguv2KZjpTWCpyfUvRcVaTsNgaPJt8IhxG0HOiGVbG7uQIjpQ1xwaDsbTw3PjIdaCw9YO5+g
GvfEvjMvAwuMf/7HuJ0xpDAKH+EKS+n2i5KpuGJjUoreT5LYK0HaV2+EWTrQM7jTFV9cREoXKWKg
MBSiIkbqq38gYm1mZGbDblePKsuZSWy331y5dhD+GKOT8X7/ZmaGIvMPChqIuIlnLjwqWTDkuRJL
3Gr38SPfb7lHsbcSxBRTXMDAcLlSoZQp91hbuZhNn4wXB1YMhA9eaorwilsAlicfjG0VhrD9Pm9S
jIb56FepnQ/f3QYd7Wksclj7/cf+XGwqG+EcsWcBfwPMQoVoKywfLheAdRtUTpvHdiGPybxXXkdN
0qdUEqGdW33dq8tI9nG6Z3JXtbFFQnE8QuqNMk0znlPuW602I7bY5GbipyZBmi/09KywyXnr77XL
N4Qm5W16esDjFFuuLal+3lFN1J0zj+FFNbst4tNCalVI7Jq44dX4I0zKyGVD50q4VfnJNyM6U+z1
oMmRCOjq3NjpSSkGrhcMGsEQ6TbuvdXzARwE8pCgF+FuzQrUfBtB+jXPyGnKE01XTxbPkfTipbBU
FAwiRCDF/4Yvyn+zcddQGhsDEySBasmmcu1cp/7TuarqMRg/Ch9PfoM0xq5Iu3AScVW6m9Uf/H54
UR24DjnfCNgQUjp8m5jeEGXiW4lz2jizdhkgaWkwO88AxSXKXsheahV4LMUalpk1WTjWsNMvUbit
3f6FTVOW0BPxiOaUqGOEqyOLYlk86T7vchI13LN8mLk39MAwwgUEjqiBR9Hv/XKeVN4JNCO7w/TX
yB1NQPrnwqMywV/tsyX14ITbsVu0ZgFG0HjFhnd2ZEHGzDooSmuNCmOQru4tW8gbkYBZBBqe//MI
jaiBG+1lV2E6JF/y1on5WWn3bp1GZOEUeIRCCDvzERLfnMF7iVLXlYYNC9xSaqhoWYLTRxgD68Qw
9IqjMIeXdt2H79CNEJ7+13zd3bX8FqKBW9pNt+ZhoZSawAccHn5BfkaO1xfgtA72qeRiYevjm5s/
9ZIbn6SuB4KrYQWfVQzWmzXDPsR1aq5X4FPhdKgWey5wVjX3spw+BS1TSmgWElvVUefyk3G222L9
VjcLaa/ZSl2W5K+Ug8HI/XkhtBdFcKelj369RQaWXiTSHaiR86RFpz5bssXFysZPpfZhJu/bqQ6C
PZARhgWEK0OSLlFcyopKg51lmApHfn5XlzieYZbGj2pCn3aJ8KevQMVo9LNnkyJId0qXDywk93D0
u9srfZKIFnEI6FAO+dKJzccbamVv2F4lL0EdXWiS37s6px2fu26HUqvEStKNfL5Lt2w4jVBsft3a
UdksUndf2GHD0x9IyErvmhDFeGFr0z1R5gVMXAsqmqX0NHowfZ+lci2Y1mTK5JOpDjFkls4P+Jn7
0XTg7/oNSuM+afV8MghXpGYhNcMYykbnnaF2ZKshRSCiZW0wxHVhTFS8Zmyvh28amQ0rAuQtJCie
Fl2I4dW5rrqLVYXKarR1BJQjlaw/1xUZOh3jcJ42TVRnKIBfp4DSa9IuNevbL0J5HqOtaeueD/2p
ib1Mwwp5n0OZcFWoSBJbClQAV3HI0K1a5ra+G3HgsjqXDkZXuy1LFOY+lcFcMao/OZo144aUPqFp
hlGdxStvO4h71KQV3hyi4E3cIXyGypYfMNlxz36Dj7DCGxGan83oOKGF9SVx4kz3hpZznNsBMg62
t/OIXy6loO1MeJuE6TXqeeXRAqKOK+c7Jpuf2/T7OWUTQgszlWsts+6bTtDcsd9Kp7uwEgE2El7T
K8A6sWRkuTqKhlLbmAC3GDrRilzZ10Lzp2zFAqo21FOiY+tgSr2IY1Lw1+2yfMuymH8yH/5Vvc7k
cjx5Nd9w8jhikiqepPLES5hrrqu/zRRewcRvmCM9Bpc1aLqQZjkKfMBr2P05lCC8MHn4oLKCH0V4
L4+aHW/tuE1jdw6JvuglKnAMOK+oeMEP8kQ4P9zAGZe/2eCsW/sC3nnvgKINHXRbmmD8CfNhcRhV
5MLwtQq3RpCpgZOYPoUEwXlZdh3u3602ONXPpjIJ/ANkdFm/siDEd/270mo3CHqWjf4v82rpNqXl
qWlLrljsPv21W4LgC9z6NRHqH0LxVJhUIdk5v6vGU7kkHYJ85diRf5ytcM186g5Va+SHopf4Qm29
u4Olc38NMOfl/nFvRFDXfiLZUZmyOomySMXgJdZbydaVHL0WPaIarvaUzeEt/A45oZ4yPW2IRuQ3
EgaIVuYPgziqLaylXl7mQUPXwLLo8TMbiu9d+hDyusQ8eaywELtvJ9pLAjmFzvUyjkuL5Wq1m99t
BYn60KTTGYPHXlkDkhk05AT5X/lgQxuOcBJ+c30m20ZxjI9VGpxKRg7USNcnY1skVpgj9c6+f5dA
XSip7sd31g8FRXPBhwo8BclQyIpvNILPSbqLqEu6l8RraAFiWqa0eFo+PsFjOqi38PNtExmVuiEJ
RDstCL29u/rXnC18puttyAjHyQibOlxeTd5v0wRMlJ4frgNT/y2rKfRzrBto2rMkzd1cHnQ71oCT
LIC6fi6V1mQkrYGXtuNyPIpysbLCvX+4DDP/PATBVkTEdD+YrK6rNx9E0tz/SUvwx5+AwiXz0ZUA
j8qzI23eyNoCP8bWRkYm57uV4aZYUtXfA391of5udhsFXsK0ZmINpkN0v7a1PYQkdHGhqdiYAmUA
9Au/M0RC2kOcl1+0TcXcN9nlGL+QIOUVeQYNdx9E3yV1N9311PauCHXd7VqfHcAFX27gzwj3nDia
rqZR2AOws/zSbNMlXRgFG2lYjl6IVx5rf05viToDKkr9aGXaSoCTDi+nUg9jtEUZWVlwsEbS42Pm
LXZe/fMAv57CnNmWZjwAuu6D5uKjDpi5U+AnwrDrxMjTABXTApgQhSjNhmblOHussrsQP+H8Dk4c
sprxEnt2X6Piif1OEIZGiBDiuBaWr5Tl5Lh1fzlbvgXmbjZI/wMGNtpA2rSdwFcele2LQzio/U6j
8MLeci6E5IcqpcSWAxnNpxlXPyJTyZZ2/Z8J0GPz/iupgnyuds6NUMmMVnBAzNU22ajMfYRKUZHt
XuJz5lRL3hnN5r7zLAw+83J01brHMh+IfP7h6PVkosI/t7Q8dW+QXOKksIwaKuMrkVr11Hc5LxpW
bTSIFkX2CeTsw9M7F3B4cGAbQf/UULGj+YM4oX2jkm1sSWqCl8lcAoCgyFvtFsKiexcpnX8cHp2U
XFVJFFC/3/oAPkOZFdhuJ0Z131CtoY3rPYnYyk0PaAChv2OBOwfwXC1tfj1LOSftP3/4nYrwu66j
gQ7Yie/FQxe1sMEi1OMzoZvEpr9xzNeTuZn132gtbpA+FO8YLm763nMZeQqr1h/TVdn2lPd44D93
BvZQm1DUmgcRJCjtfbcPZUz/CHLqEIZvV37RchuC5wKEQW/71/cUACiIDo8cTGZOgH0icpnuo+WF
tG2lqYwG9ltYHCR4Yu1TGULYckk2ywVi67kOI+GinTKhGvUs45t0uAjnaT4Z1DdPXOeGqk+xkbXP
QGjE9CRgoQciAdNH/p3P1I1WqZb8vLqT+RJSHGy6f4HEtKEMIvUO1+xoWakhnSEvLmaTEg66qyF3
8wwe8xklk4vmEhaNcxp8N8WeJujeyipHzLc1xjdjz3l0RO8iRs2qNLRQkPJC+MCfXRb6bwTVcO1W
HI08WvoUsTXfWdu7UtLgdpzePujAcU+7PSP4vg19GlJC6DyfmXqNNkfX2O3RvLEh6UQcszHVR0b9
syBSZjueIVMm9OKinsYibpBZQeg2iUzCxBTcm667VfsVPajHMKDdR5QBAEx2pV3TVT0RCjRUv2xx
q9ua7sRhLQwL/xhYS1E6hg2Mhdlev7/84pVbjnwAO5X16ngx9u0PRsE6X1svCki+WwS5jo02Sdhb
raV89OVRoYEkLTFuUPnSziMd7DZ6R2DFVENDOugCSJnIooCQPMnZvNHiGpokyGvlq1qDoGiRAe6r
HNo+TWnXAH2Aomhm7jJLUzjtMylmMZf36VkaPgu0eqru3tVjp2pexfSEngqDfRn8iLPsyPHSWCfx
z2PlR6xTmzYy0nJg22d0mTTkbk8gaJ73oXJxrbkB2h2TT80UPjpCGmlFaI7bg9b3zxMPCniL/dSg
GXKulWkjp7dCEpQno12leNi9S7ouxbf+cXdJvtsIYNghGAmXqwNhD3SUp+N0XZPmPS0E0SHmwiF8
4IrZo8EO/UrynN+MYzH3Od7GrjGBn2Ayi4AOuSFbVOtT6jdLczKJ60QNNfFWwix+VSyW3PTzokbn
vjsrWDfgY8x1eP7f2AmzmYkkysiXBlvaap78PsZ348e1Zoya4qTnvAOvmfXAdfgOHUmcCKNkgG3A
a8SfDkdl2yer8z8JPi3hUf6CIXalYIHSWZt+CiVITPSY7pcPwILXgQJ/NPlnxYYe7etGeOZqR2RM
Zl2RixnvzxJnaHi7J66fEwnqBNdGOgFis/f8VULrjGbYZJvF0ApXnzS/1L7H4T3rERMBa63Gz9Yf
xSzqo2hkPnOmFp1eZxIGmLCr5rU5Rwum7+ExCmGQvPgJlAUu3GwTtiKhZtRr4VkvknKcZTE278rZ
xn1snLh5TygzcQzJsEd8mospEslvNR1IdGf5LO53Lo82IwNqnz4mECafWePpYbzyFTpms6TPSru8
NH8dR8WSMxC3803etLujdJ6ESns6vHwAOtfZpBrPok64d/saSBxSOgU1NsnsXwrGq/o3k02nOpk7
PInZ/2Do544y0xzxjr9ASBsDdSD9MhVCnxo+8jyBTS+s/+piqqCbqub/nn+PYWh0BPd5Maqqwjfx
5IaUh83oxi0KEPAQ/31pvz7uW/AF9woqFAZRyH9vi4u2uY5g4llm+vdY2PKKOtlB4WogEo5+V5CO
dUg+62/lnmMdIjBA9KvAxbERnaffDQ/2FDtKLQSpp2BhfRhgXZVFz/9ZJvgym99huRFbz+sli/ZV
fDhcP6AwgB0Vs5JCDkIoQlEALNT/BU7Nzlrq0RVPy/cN6EPW3i5MDbPGfCt/WfwGa6MduBFI9IQf
sbzoWCvTAuNWvHZK7R+Ia65EJs/SvBrEYh1X67Qm1Wl6lRCqIF/fpj8i+sdE7743EzvfgZpkO4Zd
9tYF0g9lA9CH+m5ZL2qNolMKLnMwoL/JPJs7LhBU8FvBTpsUPLQQUHwEMDljBbl6t7Iy4/e9kJ9P
owUVGIDxQtdOOeqgdsuheyLrDYbbNbDgfhbpItHb2O90Iff9id2Z36lMi/WaX3Uw8IzZlEkm/zdV
9BqUfhsMLlYL75ZcyySozPa3Zx0bdXi6KnTOhm+LFt8T0TsjdVhMh3RNfHgCoCwKdgLA2K0ZEUHb
YbmX9fr8J3tem8ShEHmoIJVieNdPVLV07YVLbZjPETHhm+QvexTRotiSGB4PSPXhRZrNqO9fIc/9
91FYK7BqLLqHZzBv8fkRsdIYN+9exrtVK3delZxgLM0ih25c/lb06KICF8mv+zkVXt3czG4j6gQH
CoZyxKggoEB9Xxllcxe1wgtX9IexCIOFl4o93LX+49IvhVRMRIID60PGyV6csA/VXO5XmxxNcQOm
ipr5xPRqkGSJQIOs7+sh/q3dGRFPpFEo4xW8CDKHO37yutDvPnV/1iY4xNz52tIVcmXTuTR9V2kK
XGSaWO34MaMQ9E6T5mHz4MhKy2/LR0PsV9J8PgrwmGcsWy0pzPS8ajbCAlb6MnI1vnzFwvWRHtiv
wu93DQZbnrFwjNXgAu9PBJAezQQBco7D8U9ynna5yMZ6Rv5NQ+DNCurGSFdFib6X2PRp7kgS73fI
2ES7TUpC1/RJJnRgc/I6/xdrWZI2hHhJ3yUwev46nNc/qz+J7dzCN1efI/NjhsiZgDr302xlcPyq
30bDMuWKO+LRktvcMa/DaIv+FeMR6JThmwD4mZEAfdmiN7Nqyw/XKltWnQZqpoxuz+nZQp+xyjeG
P8xQM5Es0jXHJQWVEwxhgLhmsqy8j2ReBBFgbvqm2UCSTiF8GN/ItB2WaL/c6p3k/qtbVBTyyut8
TK5UTo6XhnaiZRSa+8b7UKRQU24MQX6gTRRBEiFTMEQa/MP902lz1TSdv/rezybSu8gfriK55qzh
F1sSLZ8YP0kGxH0FwU+RHOd0z6sJMNeOAcN2yHQONoRPAvgWAs6BnGgi2Gb5ygyN03lZvkrlvYGY
Isr4J/X3eP1f6fj5RXFlJkqQSIHL5NY0DVCWaFdjvzYYcLyk0TgGMbPv+Aqll3D4OIfg8/ZlQNkZ
wni2fE5mLLLzCBcx6S2o/kWiJjg2kpWo/Doy8ZczpG0rBdFysONVHqCuEK8cO/0wCxi+b0a22jmw
dPKMthc6HiSL/H/rUEcQ5BvaX2GUsCuY5TFKngCMGR4y2pBHb+J0HY83hCaACsjiITDnmsDsMwKt
m9ml/KPpTOLR5JRQgAwVab3Xma8e3bdYjqO91Q9/KDNAcbw6qa2FkLGGdv0GKYCNEdkPhTVg/xD9
1ajgPO/Q5iw/kdqxcNwPhwBGwI0epDmToPMJN85YpBw6OdIWUJxKZJU8jHoXEGrKAqpS7Sw7iKvI
BuFSvAsVTZiA7nq1MLkU/aoGN1yPdCNKgvRItvaSeOszPJBJleGbHx4xQpUxbfCXhb8mnw1dr5KN
R7eO46w0depDpezQOAwXsYUR4ms3jdBXQhxBGPS3AnPxZDm20TYOn+m0kQu1k8XNoIHT3RXaWs06
vy9KtHfvvNZXTGRKBwMvY/vNHObpIW7pHF6Oo/3ILkxDRrOhGj1Y7wV3aB41gAMSAiLysQeoUsxb
IAjdenrZ5FmtGWMMCIfFeNxaCJAUXrpKjIRWubSGoOpN6CE0Ecy15B4j2I+jVvk30Zwozh9FNtKK
2Ia0zOJ7LkW81osjNvp8niOJ0hcfdPbLwmAFwz+r4fWo+brM8Dkn3vyWtPt/jmhSYoL+im8wNbcr
5dSZ6tCg1XdwmaA3wawnVsCnlxMr6QEWxOJ/5/IpETfu/365Hy+FHAVx47uuahYHnhDvUkEbWkLV
Pa25BeVnQOtd7l4JkAJbtbg5tuOQ6WLXKecgO4tg1SneHkYHMEBnowAQw7r8gr7NflrJSS4IKpPv
E1A0HTB7ZsQT+sHo7q5RaTNQ42GdUAg6OkVgK0+u0yT1KI8ijK7uoKFWq8lq4G0ChupPDq0NYKb5
mujotiYCilQE6a4Nhjc7LMN6YPZvPsvTWK1PswJV1QJBK7yBpliNy3JXzYA+bYap5OrVwURH91bA
ASoI2c6O4JB74XnzhxcS87EpPq+n+kVCGGHaDPZFanlpHqXVRmMfcDB84Uab1QogiAUUzQ9QBety
dZdXkEf4jMefDAQDcvMzwIHynWbzflVsKtx6DsNJwEhqqBf8rv88z9Ac+0jYEbYGiB5QAWJ56aan
iA1V3mjioDGeEBHKWuUv1JXlWFrN9qatIv19+kd7DBF2+LqJPTKX3EhjO39Z/2EtR5VljvMp0/DX
hQCJ043eg47SwoEwo5Wi/IHgB++XvO20xVsLn91WhTfUSJs54QhOPT64wXX/feFGmhp6r0lXJnxz
DjBaihedNb5/QY0uthGaSsEzXnx1v4MlIhDim/On370XqNjtsSXSveZ2mwQIRsOBGrwid45ziW2b
aVjq1WND4USJVr27u6HTnPPp30om98x5jnWtEPTRzxS/NMxTvYveo/WIOExwv+Gb2Dh2kOmLO4h9
YXjO4DN7eWFFS31S9yBrc+SF7t7G5f4FV7mOwBfgWyoxMcUZrrl/YzJp0+bkMiMWACjIc/t5N1ra
sKZ8aPFUBK7XcTX0+HLrapNwPVrSejzYCjijpzVHycAGUSfQrhIcVeseUiUc7ANe/t7wWmF94YGa
pXFNTHP6czj8SRPFd2uUVeDIRhhFz9ALQbsaEcN0Ih64yOqQb63c12odMF/dGu2ZE175WkHVNv8K
vnSe98Zk5IK/uK4TVowy0HDlrpKPjNOpmDezajcF2y6/VHB9vt644XoCChVh8u1ZgU+errCudNCf
SI0DKSu7zBVUt5ipVZz2sMQ46IlaCkG5o8tzsStdEHLf9fL+5dVoaRA5Hyo1bI0+EBVCiHR9xmeR
eZDdryeoGrJ4TpodEggGxhMf8sF+7Od/xxNnDV6NwUuMzXsKKEoHEDAqioHC3csj8zcZzUcEk/ME
jrJUOnC+Nkl7u9Qb/8bpLARz5Ic9jQvntU0YZ8I5m0WQ4jq9Q+96wMW4SsM+cDReXqz8RGOcFDZ/
T7rynuEEIytIPtUqJjq5Z1veUV8xcsjxqY05o+H70UEeeIeOqGKA3yM7IZM2wsewEGTCZ6jLHfbK
x61Cb+UIvStqW45LB0VYF5eXTZs6M8oRDTwunMt48iqc9XZTwJZlL8ESoybQRCbn46bkOAFznmvK
l1ehn3d/has9TPGQ7Y1SaBh/p/ot4tGYb23BLkkalGUILa/aTvXkiJRMJO4iCvP+Gu2VvzO7tZx+
dfyhIQXwzzi99JOYVLcKubT2TjiOjPXbOu50SdmBs3lPZqxDlXvAqHl4B4QqBKwbg8SBA3cLE6aS
WESJmCIPw0DQIcavlstT4nkP/QrvR3gg1X7wej1RY6th2TCs27gNxTnlDpvFEb+dTe+CVJEtzDH2
EjzTbNxV+5B+3YmfYWRi++JAoXgwz22+tmbjDDA2Oo+mpDcGz4G9mV13BpINHav35r1K0mbNadFK
IjM+xASL35WaIoMuJS75C7wllY/6OOzSSgzLhS4NQFICo41VMTyVWI2wBcowM3cFIeA8sTDrCM3i
7y8RFvunC4Uk67AhLjKHOyeiSc58COoodLPO7mnjBRuFT7GdKFGjUw1fIsK6vt12jpE+INmgkhU+
s/TiOzw4JK9ByvTYsSFpXyGyyVLe0inmtUz+J+Xi6E8pMjZqYgww1dPl8xB8YVmYeeKJWH3XrnNA
K/zMWn+d9lkPPOu8C+ojuadV8KreaHiicpVWYBhtGB2t7Dfs4lrcADQOyVZaWXw3j8Bum5DEPs4D
hG4+cjgcC6hp29Fhqre1K6rKxBFMiPtseyZHw4K9cNWxW0yveBDr7vorq8MfWU6M8Nt1CzA3Yfbx
ZB3OcUTTZoKZ/LgcgQnP6CoNJj0r52FMhjyWBYn8Vd8wGg0/F+vnDIjf2osniXo81EULdvZGU+mw
dmhR4NiuFZ+zcOZMc4vau07HuoplMAoV08Xh1FCIkyEWNfn447Tb2xLvLLcYtna3xm59Byvp5jFo
04UBGVaSGnxYEz4zCqXb9+X12YH+bsRsPJL1hXbMYY+EZpCyZt8maTjBsugOwDjsyzgKhqQ1uSPe
rEi39rCQ7NFWANNp+aSwCBDlP0j0bJHdUwCfJd/8S1qPtOlfF5/i/akQ1cNdXNa9QWUqXpfkD9sP
7UCP+ouGujbyn8mUMmiwz4jI6NXFT3FI0gcKj9pwC51BfFalg6rpph81XFw6oF8pLFPAcEzTlT6N
ZvWeCQSVMsSG34B/glehxMPn4Q2Zpl+ixgS1M9/aHAZ1+4o7AJmJjjojCOUbTvK9UCMLGF0GConE
0dX03uoRNAnEOGPGKb23B9tbwhsSAHxbrGLOvGckuDLGzQyJ6Bsue7G9ep/8QlLesFCV/TqYjjvJ
JB1kLoj4OzGIGtZUYf13DQIrZD9b0XoI7BIgu23VcHTOXLiEEVzOYN7VmxDtPtkx31wxwphdS9Xw
+rxGjIZcjaWn6/x1Sx6Y8BjWuW0A4qr5tMZtgR5L9IJ6iq24G9x4xh1laVXPr6iDOLzOFAKDuyFa
XlP8KHE1pBIaZqXA86jL1ujhx2Y2Y22Df7287M1x2bfmE2f2EUIsUJFr5JKJ2sXc37MwmAC4nG5y
9OT6L0Xn/ATc2wqmqCipvtYVEuVt8mEffac0F+/whKOEeiRudBGKKaT2SoUCSdrCR96aeRDu1Rki
SeubkovkW/wZ0WyHMgIFpabE177eXRJPSGOHBnJS1wbgmdJLwfwhY2tAwvEuz23XyRsddalkfrSi
HdJAwLxhr6HcN8hU8pIhEloXuStkDMuME2yY2siIu7hK/toBsPWLwjwJ8mYz7eTRy5yUdezUByVw
JIgP+mW2AD6L5LasMoRf/TZiWvI5uHG/4gWslDf6wGM/tmy1U99wHPhu2T6zSZtWsN6in8YNJ5A0
vSCnc4FsWulVsE36jZ2KZNjV2mCMzVQhQsMeWP+MgRLrQ+Sw92KSL58hmgU1vNZyWmFGLH9574vU
kg77bQWdaZoCpwMLxKuNGQf180Wv80dcWHHKXuGXWInvOGi036y4G438T+t0dxEeG3m58NDOMKao
UwX04OQXfVeBNKhaMG4iAI1gp+snT95/YDHKP6VF0+OB1yebpLKuK2clGGvBANYRmmEpSVwiF0Xa
U0R6sLT1f+DSouvTTnWW50F6RCAs9MlsY3hZNeYRcEjDrjCW1nMyeab+NliPrcbWR3TWhVgLjbj9
vopG0dyx09QNxbI3Db6ihLlkJ7TqtHg0XdTTM8IQcOjLl4rU0VVOh8VYt9OTKaPSBCXJWMV6jFgA
w5gAq5h6RP1YzDGbhd1swZq5/ehCX5ZSJ7nHdOu3uptBjt1Wny7MkqZguD72egoJUF1UBdLGUCJ+
E0LRa2GInP3UIOH7x2wb+EsrwwhAVYP8f6aTfKuMRj8OiSJbDn54CitwNfUDgfuim5SAwLHg60Ps
XFXcjRBUctZfjJp4I29av0XYFEPsVoBbDSxR1zpR2rhVdakSYtT4y7Y146WDbNy53FZHL7XrC9wG
ImSywjJFuUCirS6n4hf+57sWPcnRBd188F2E/QSCNtlkt1pjfDf2XCLraPwOXUcRUbPmpbYh2fRg
FCOa3HR3qhTDRSR+t5pJs69xnJ4DRFpkOdxbPwBMjZOCD1WQ7UBOHDsTomCflMLXWOn0eNLbwRNS
NUmEyJ23Pw2Iobr56qvyHW4FPgNe70cwJLVNaZtN+O6Pz/k/5EKHV4vZXC5LqNix/Bdsn8u4lLxX
DWM9rEXmBbvuYn6/1c2Fmi9BWNzBWLoLJ4vz6AbfSOsBDaieji0W3SIWKQwvUdGbFcCG01E646YP
CkYthRn8yrQacRPEV7L8ZkN9orssJA6b8vl+CCzP0QGG6fFuGqfodYR9QekGH/AwU8+k0vBMrt1h
GHchPg4iFr/zmOETAV/gRl52usSnvXtmdUeC7ZsSCRNyaTb8wRnXC3+nVj3h9w595/wAjQY/asa4
+whwHtTNGyvelSWICHBYpShMHT2i8fxN4L5GjWUN+ozxhBVTxJytxXtg2X9yFHwZPxguxrD+jfxm
l9ksda3t0kWwJjQCZB+SZbiERodYPFKqqcGuBnyBFubrViXxeIBqfAbyJuxuw1El8UAQH5wc2xyD
XmJTqQW47tQEcj4SkTKep60KfT481fBitcoF/wDNZT1G7h2rlNx1SzsurFOJZ3VDMy8rhISor7uR
FVWBy2SG7OX7jnX5a7F17DIFskRbyjMIFHVW8ZjagoP6yduyWE3qzHPdOACo5N9RNjv0olS/oZxq
0llyLmvLyiJoL12pcFJfofeFGrtqa0rPLZvXiPOzTeFCMm1r7OFBR6OyWnz0VUckq9N8kUtjI38I
BFqG5hM5/0Ko//K/VEeLHPwnAk5nFVELIEjqV0yfauKK8ptJsGcjvY6zdWgcCIKbdFVVIRpwJiyO
FRTIJQ4YGOfwLdA/uXqkTNsKyHY01N0eahU4HEdmmjUBsNtC7AtMVmwUdoWIRV3WZed8m/A4p0e/
jT/jZlEE/sDhdgFHYjbSD8s9vhGjFsrt+4xNay8bMEYQIKsq6+MR+bwDQoc1K+9QbAtaI7Kr7gCV
KXckRQv10Yjd/Ot2iR4F+q8oM8mHZtIBhZfld6kmQJ4GI0RTGoZaJI1gHxYsotvCshbTG4iyGBHj
UFr8jLrBEqSPyutuWpuYxJ1WZePhUSRsRBfGXDVz7TeplxztM9zSs5GXTrp2s9k0o7eT+FSu3H+F
FbIc6DWNPIHsngoTig8zgl/QKbaOu5P5r8KuwpYTj6M3yfGp+ZZEEuevc9mBStoKMIsiQ8QkKVlZ
i5hewxJ5ah950ghrxUHUV4ZKMqqzoqvgQXvtM50vAfGLaxtX8JcUMzvEB2VIw6XO7vaNf0FV2XJP
2jPnL6+dOTZ68KqimzDp22thWmQEWBfWoY16BnbP7zEn1eN8EW8Na72avmzSffy7tqwJ3DmQWorA
LdqrRhjImoEnvAjU53yfIlahEEQT6IHGW9lKIirixU9P3YuY6dMB57B0Igj6ZG7KnmZbs2UhEMpP
rBk4acbAwp4jWMqc2hmqkTAa3e567A9BHoazTmHrOS6WfppSrVZykJ5a/R3LvFTm7xHdCqqH5Q7N
3F/4WYipCccejuhBypGLlsZgzCXsP6BF6PCcQTAJmV6e7vEVHd6V6ltwbg8mQWjZVn2ZkEEcsLli
vBFbeUhgBbGixNepUNP7YGJGgs7+mfws2Yj78v2hFD/IjKtIf7F+GMOjCDlBPsn+dXMv1AYJzw0B
thzInKJe0odBfl6XYLo7T2S2t7mQdARtx3J1Pfe/1KA9C8MJsnRWO84uHjYUtEpuhh3kSz/6qDte
Yeyxz5A8wcxgK3GVirXVdAFqfZ3MvXc/AjswIYumGlbDlLYOrIADXKoktzsOOU8P8oTLi3urBWLg
/C79TID1j6X2eV7/zDPVZLE+FXsjS0e3sm+d9S3umlFdksi8nXDuNf0g9KQWQd6048QNvqABaqjE
1JT+J5qnA3h84qu6L2rUA+EdMCe3VFGZwOtcHhOFmftlO7eMwEYN5VFRGN8+eV5PRm71afFTLSr0
lZRgVWFGnaJLmXQ8TJd3Jy0xIvrRdL/NKRP+EzXGlueKIFiTmPJdtQbkqwIzulE9uo6i8lnn0ftX
kWRsC7ztLEeO8g6G6CKJOt8PY2AwoKdLe4mYigc2jGcXfwPpKJy5mNsVcW8agH4Tl7IasbY38sFS
NzoIAtFIn08rGBQGU77ddwpoFyKEsETn/8vnL3gW1VA98uF29y0wioeTizmiSXyb37NL4C2+CJni
0d50c9JENTDXT8VSt3/Tz+q5VCqqCyM228xr19OO7Op3srM4f+FYmQXOKszIgoCzm/n/OM7NyRBs
wcWQF8tXrnFPkC8zXb0ccgS1tdBXs6ifjWzqNsBVpI3psHThkSn6yNu4/3IcUS8JXCQZ6BwnuPEU
9+owFEtoHPK7eFdy5rBgzqd7dHiN9RZCKwDnJXFzmCr9bU9yo+jWwXYF2HdyvHzkjL9YPSFp1Gw2
CkXuZEOqaJlVtFY1Uq8TYf4pRq4O2zYE9ZFvTFw64x7Ilmqmnm+Za6z5sqyN0GUNygxTxDzYqSnW
a1g3RFDsNjzdRAxY3dT0c4ZN8kMZ8OKcjMvAXiWgNJy6u8E0ibgsSzrDe04336OpgjmAWHfpJm/C
7kYAjAib/qoWmXP6MlGS1P/C3xuJW1R4sFETjMU06dK4Q6SdMrVZwAK88KE374/gB9FKBVDy1FE8
nGQjW9rKgtSvvobrZvMgoIQGBbxaaMn1XgtEWwGrZGK/XKyRM8SdJiGJRc1P7ithfSXKAeOcNEfQ
sXog5UXrupWOvLyNeDOWB2zfdAH/8gT33/8ni716FX2naH2fUKcYBrObF5tKE7a1LgCUg26HJVn6
WKWueKJlt01yVJZIUNkRkwXuFkJH/u8PMp7UcLnYyqa+CXZBhauYJGZWkuVLXu0nfJwNxtKVSGQu
VzxVN2+bimMkL8xFb1HC9AEU20KNQAjcxapCrZz88flS1sOscpVnSItQrBz2A/0MLq2FQFUs23aY
+oFHly5P4M5sJaDDFtL1cZzbsVj5VzzWPu4FNQVvEK21bMGwUDz/wfiyVExAcornRn59ELreN04i
cD/sXRmkUg3GKJXtddDihOI90ELAHUhtmhQAh+NUeu98RjVZyMCdiMvb5tCXtrsWqHaGis1lrHiD
7dI228AaYyU+dfwZiDY1uKTkluJtxACNEydys/DTUfdl1/I7TVSRZnt5UUzD0h++5BS9lIY5rZjW
VgAGX55GO2vQxJU41uJ70iIs+qwTk9WT5WY2xkw/EzYnCVMeoYUdg/QXOdycFMu4NpN8Sl85wrpS
FJtqYcdRQQvUiDBOCMndQ9Pu9EKpDH82b5LAT8oCY5OxCCSHZSp/PG7HInZn2ua3Y/Cdf8ttTpfY
VRXQ66HA7/tjvmjtAfdIjA2gpu0/5f/DLr6+v4OXWvi0nE1QZBjH7yCeZUDoO1cnEXyjyZYXVuiH
VM9LwiZgRbqc/v2JIKkAR184YS7CasOB4ZMPCoDD/2cvYYSWFo5bO+lw6RmF/h1aqC5DZqCYd6z6
cYTk0HeHxNO/6cYZiEwJqZnXOUg0gbd5fVx5QA4QxX3xPno7Hc3wHU4bWZUdGEG0VG6231xWKhcz
l14aCVI9H1oAkWF3xfM4K3pIYcbBHBgwD5dt+BqrVb6pkTnxPni4kGpiN72lMzkyW6japJSPknjU
oiYG2MzFuMT8LtXkB3qRq8wyImZCFcfHRDjrd1s08HcYcqv2rFb0HfsjxStYaj4j91AQLxm80VL7
41BarctDSTD8CzHbjFor9dcatATUz8hegOGCYCWPQR0rINYlm6sCglwCEdOFDsdahT+r74DeuFxU
o7IHaenqGyarh1Aypu+Hnuvy+j/aTlCZRvvIVDEQ067wcTBUeI6LtSzoyVX50jUhDYZzmIlo6mmC
o5SvKkGSrKePmi2nNjjv8oZA2Fwiz7zPBYOH8u/t+MYA6SuVbUoYfKHY4o/qhzgrtWbdyJOYb0GT
FYatAcVcCwkwRrIDjDk+V2En3oOGFIoDqwgGBb3NaVPyVRZwawF+KxJvqVAAhgJfnTlsBKooHIID
xxBP33ZjYJOCQE3xswkqnQkHB8gGT36eYFhzO2/bDViJsxwHeZccDJ0o/X75ztWPTuVp/mvaFNV4
tgXOr9ebMWiTHw0aoFWtTiYyw2PLEDmV2YltmGDQAnmoOFjtwJr8/gaYpKIACJCqDHVmNHuP4nn/
yRNEJitM44sW9mHpu55syhjfF5trNb7ynlPc8eDGne/kTWTZTpA4minpQQCAwTnzFHdsCHzjSxEp
LMy0KHHT7ocLXfbL8foH+2owEyf52Vy+8ZARUFrxCAS9UGce2E9t1m+7HeKcVDhmvJ5YnBubw+ER
YZLScjNgs4aLx3YbWESUQy2Htl1qcRswwK7QK0fgmuFGtvfHmeQ0CyN85EAmSqxSsJCerHXpnA6k
MUecAtkI2MlMCLjmhUcIrXUKL0DAIZ76Ddfwomm3e+xlXd0unGkJHwACH25zs0mQ385p6YdP5zDP
KEdBrBTRdO5C/efCF8POnfAFibODrQ2dAebmMNCEm0yHqmmg/dX8UOzgxJBDlV5mR9Fci8BCd3Qz
yW1p3n6WR+tWaekjGYHt+PR+w7WLVnhe46ZVjwuE6DopvlTCVQilF+AEMOHCAgI2tg4Mui92XUZW
JvSLMHxrwE7uFgRq5GFJQj7yWO5ryOLwesPeztpijzxIob/3VjXU0GoHvZo7MMlmcvrhS2QoKqp8
kKuvJXuoau4P0q3IQ+/mFHBev98mfI9p0lHaj85LXx8da3w9DrYzh7IOCbfQBmjTkHvpk/Xq7BiN
hO9SoInooX/wFZNQiTizHo8qNX8kC1ofP1giUzvxTfDWp/aU+OQ3Rsr4JOZNmRmVTElgQjB7mVjL
bWXSv6VqK2HY/6D3sEJ6n2XgxPNc1oNrAXEw3S5vg0XsY+AWy6kvVVD6T30jk8fXJ6QNA+tqVB8h
b0oANbdWJGyW5YP0BMJx3bBHGKp8K6vvNbIvUX2y5K81z6TQUk0jCvC4HNVYqPLmWlv/2woKn8T2
17yvsPc/5aV+lCYQ5pxSq4D1WlitHmETPid5u9fFpazGjwIRWfjPcEQhuDTDIMJa2C0iQX/5vprS
tx1zvVYmnxZLSBIrtFkNI+esqV3PYS4Hjr7XE87gp7OgsgeA7uejMl99YE/1MlsBlmuXVEatgdv8
J/dfd1Tx/XMmlWR6gEcSpmiq52O/8D8NkzZsrpILlu+hBYDFf0nvkFVSgDPr3TPcWM/QI3RXGp35
aFZTyn63oa/ClZcgr48Y34SNFcWRToVJRisX5Fi+dConVRv67bLx5vPOHRXNtsesd6MHo9oFxijF
l91gN3V7C2FEV+6lbCrOEUZUxjy6fgffyd+6iS+OHbLgPK74DLixfumIVft66DbXavL8x3uaQJ2D
la0Dk8dAL7jQI0eRtqnkh9VDNGXM8CQ2jPwiMFNZCXi+ujwmC40PfqoPv6pFKLF8dYSycSlrubOK
TqIOT8IQh7Ycdj5TuCB4k7tlPcYbFRLFTpJhRtXGMsSJkcpw50AbCVbNf9KZqTGIxi0GEnAu2rIs
rpd80qLsYhMSqRVED5vEkXWeClLj99Qp8AglEPPeAUvN+VbfxYFJp+/Mt5DmIz535Q8WC4iQQD1Q
PFLmLXNl/waH4D+yJ3LipvEfBR9jazbEGSK1I8y6QO+FjsW+1Bt59rxMhIfRJvHyMU9oJzMshcqT
KxLSSgyM4MTTRS+ju1CMUOhc1CIKqaDdkVR861J9rNpG55kDLyejSlF8yvu/8Wdhy1re/QltGGsw
bqn/IbX7a0Ls/bxf0VIYU6JHpxuXzwzMpQHywbPCNC3GNP7ULA9Sn4S4L8h43CmHSQ61FUWL/u2/
MTE2xGO3Jz06hhzlch0gukifLNkctFs4BiT3kSWuRZ7q3qzM19j1/ZlGs3KYBFccsqNoIpeRwDWJ
YQi8eEwyun5evKM2u28FyJFGagK/VKVN0IOAWslXXyjgEbl+kg0PKNItbP2eRB3O9nF9+hxBGOB2
QB6SyTOTO7/qz+kMZ27V5FxE/LGhhiCV75fwu9EOWClh6w550Wlhm5RK5pyqNZakVEUMLE2DxTOf
MFdhJDvpx2U9zbbJ9O0dTY+DgiVh9dwVFmWemkV7bCXtSEZstUIV5KNgLFYiovnkWyeci+dVnchi
7XDULODuFvbzsrykux6iTm+tpXprCYclwgY2oL9+4ygJthT1f+0aPH+J9p5jXDwZoITj/deiGXhA
sev2w23GtSIu2bMJjQw/jfAg6EwxeKeUoyhu2EgDEYMTOnOpGYyc6YVLS6z6oYyEfMMxtY0Wrl/1
+pH7zJOQ5FFKB2TPxYqlos1tRReMTCUAKYAyXV0tMTmMdK1nZqAnMMLhidUELeyIkb4ztI/QA7M/
JwUgyomBaDzKxvmzMiV8AJfaauSkdJoixmE8z9DhjOo9G1/GKswSLZGPSe2Sr9CR0P0ea/kEvHEE
NI7s9owgV5U46jtMC3EAA/6FI8AYog5q10bc11wE6cau+mGnaki6J1CESgF9izhpp3xxVbP8FYSp
i1R6XKGW559F9oUGRePRi5pShQmzjEvog6jDnVFqgC10i7yrzI5IQsYgWdUVI3tkA2QjGKEWXj5E
bdyKSgAmaJ/D0qCB94je9+DGwYBysuNBw9qCweQ6emqJkfT0BNs4DyXKkQuy9OQNHOKOjyCI/Z/U
t3curOuh+YH4TVFxRbO5fR6sp0soFnkmCMTQzdmEoi+7+/jm3eoqeg7gj1uLG9NE0WFt11kLu3CX
4yKIePLY9MV6+xgECaaQP0r/oKN03ukPUjTX/j/1ixfiYNbEP19HYEDHTnSXouevgaRjsRrcLHJR
wcDe+uE83EHK8fOb2H070m7ThCEh3BRdGYUvEDTnIpBaYiVEJ2ndeV2YHP0H1AFv64ZfnLyiNedJ
PXbe3DTLTTGYtQ/dsg3CrThVIw4q8KerMylr0dO4g7/33TCM+XiLagIxQxcVipPYtzFR3UCp5e4R
0wdkm1Ffk5i0hhUB5A/srMv2dDVzMO1/h1e2dl3pXn1wknub/64HSxI264lzOyZ5EvgZFeQfxT6c
AlQxmWJcAfa1XqgjTA+LQ+0B/Sx1Kxmam5JvL/zHM9OIty+Qp32BcHwa3laKO9abW+LaYqEU6ftv
RqJJWauboHDTXS68YkegZNt8S6+4+hUIWuQeJQ42VjlKYRi9QT/lekktm3H9zG8s6WQwvAJmEIyp
vXGGaIyvotnHxlu0WZkQ2hf1fGF/PBE+zPQX+0ekhPAbBxg0R97xep1BB6A1xbTc2LJvq6tZTkTl
rBjxvMO1nD73sIthH9N4KeeAyWhhhWjhggGF63n0GUVbzy50bTgbRddjvaam43hualNZxqAlGrXE
SCnwxqPlJgkuIV9l9LBcTkdXb1p5VAS7K0P0FBWNRRopecawTiLTpn2z71/FshyJlPTThXrQyXgW
E6mhJns7KyX/hEi/MRgXI7SqM/8kpg/iM/9knB3MXpLpPvIC/w3V59DYGDUSeEsv7rOF3qI6+apC
Fm0CD7ElzL2Tmre6HwFFWoO74E9UiAJwwvfbRYrYlRxM2I4nEQSPtN3rhwdGwdxEh2zuXy7yUWU+
f7JgboV2IE9pBaZ1gcZP5GAd3rxFBxbTJ22NVi4ED7Fo8rdBCp0tVxD7Pxvsrw0xKrHV8EhiWIKX
CF3/MlAhTPsnbSjiVYQLrRC/BmE+IpzE++ca3KGbimFAJLT8xXWurPzOnN2WPRRC6Yo59veQpoPa
SAe7mW5DxnWft8KF/2i312xS/qCMwcD1tm48F4AmGeJbfxTNKOJhSgXKeV49vy7+GR3HBgS2DAPb
VeZofsBZLr8p98CP9lj0BSdeZ8gi6B6QwrMTltUlxvfypSc/n6ro3UXHC1U8M8tDGzYoa44ccvxi
ni0u695slYwB/q+g89nOIGy+zhqFndDvhj3M/DpF9Wgvrl3GpQEx3aQnfHpX331uz3hU27u3U21P
LPduyua38Hw1Cy6NoeH2FCwQEkIQ12rqhWteTh5d/UNFksWmVeZ8og2e9Yco9sM7xK1rk4JPzRZe
7zEBgrccAdnUU+n1TAOA9WA8+ttQx3EFjZHb477FSq25A1wrtxb+HB6ChJYohBBBajV8gaUPztgP
S0cD40m259Ml/etIM5f+J7CIiCJhtshqe58z2RAASY4zXM2THdczbiiSI8oeX0bvPgPXj07+ZunX
9GHcZLwMxLxQGTnT4PskAct4XNhuvRHjxzImVh8xHiT3J92zwsZa43pxlVetbuo8QcNTrTyQ+7ee
Q3WDa6NZqAn8rv9T2bvBCM051wq8IWnXNXOXEnMR6UY/sr/D9Jbnh2KngvHw+DD4P9RdehLEtX3T
IL3xykXNGO2MqSmUlbbhZZ6Go1PfHCJTyRl9xKs3yCVDno975UCcgkP66n1LhvBR1v3mnbf215t9
atTyr/4Ws5gXheGmIAijtAEykJqLh3GaLV5gkwdpECYrdTu18K9vEpwHQVAIqXlPhcr9GOwJLQeD
NVYsmDe6BoeNand9IyXxcE8zroMvUu3UzXzkbBL1U5yIZ1LVaGLxBM3/W3lSOrHcA0gFm2l+PB3q
j+3GJw0WdLHrOQoSne8mEwgTs2D12wUN2ED5huDHbVwSKjj2NgnZslvYaUq2d74BK20VFKirOpSH
9CPr1V2GDyBIalwgAUGDRKC3EiCQOSjOVqR698yfBjaXJ+aEx2y8thSAv0/HiRsdJLg0tf93M1GM
ht8sp64vhhYJ1s1bDhZCWwIZVTIYfdAqVVqdPmxF6zeUG7gNM/f2Eg25l0LJx2TbdWKMibyCjOMQ
MFbJU7v2do49mHBzog5FobUskG4bHelPb9Kq1gkd4vZrJsfxRbeFAD1qQ+ZuN7FN5m+vEcAvxues
EF1ed8F0Lih1MVvizO0fmeTAMqXonP965BZKCGUQS+Q5WbdZGnppndQiWohuVV1wZjFj6tY1e2zk
L6u6f4HfB4kcGBFkIu9arlzwYBU+vEuaC23zXPwYETNyULT63fbR3deyyRF4IooyQJRwNOYzVMci
q45/HgCYT1Mjlbqv77JtslZdQ5fkb0RgrEuV0ygFxE8qVHLOBD0Z8VohkU9xxsuUSM3BfrlLSFGz
dz2HMAGTnErWf72ppDi296WoJUOHUB6L7HtF6F9mfYl+/XJUSs9AurSBBla9NLpFlG+BsOiW3ZL+
W6Wa4pnqmcboMZkIf2fhRjJrXKcjNMjP+nd9fJlrFHJW1SEZ7xPUGTLTJXSjx1Kr2GhtxRZL5doq
FdrbdxTi0zNSJ/SdbbHpHTsauzr1J6Jy+BfaPNiOpLzCbOtuJ6RY/DXElYQkG0vFNobDDiN4kwEf
SA4MJkMlSSBbuS2fa2SgXrqp3GwI6LvOTozA88UP272KMkctFd0MtC83eBbIMylB/VhzdwWtWdTA
5f9Ro6P33PpZLSoJKD2EGbtKkhVa5Is2XUyBTIeRE1anA9gPEWGnc3C5NQoGwBe+eQ0WPno+3gfi
sJ6aulagRKiOs7yeBoRz646/LR3XY8Gfn+uYWCVSHQGaZyYhy23Ntd2jEmOoDkh0iHKmM+fHLfIc
LIItzee6Llx0h54ZV1a4+pd9g492GB8o4IDWNKnkXIOrQvn78qutJYknxr6jD9eS7Ogk4GEg04iQ
Efv9cRNdjB2fW/3Kwf4ZeT2nx2JDJJtQidpLtk7VK7vD6B9fiLqzeBaRadQsBrAf37JjvOJ7kbcA
gU5u3H094z6mkk6PU8+7xcc4xgdUZhmbu5G1sUjazZ3DbHS+b1oRDsu/59voWH0RhFo+crAC07aa
XJAefypHff4AhL3vF7+6ZynEZbED7Rxin7u5BiR059zMSwc0zGoCl7IsTiu6ozJMJQpD8VQtnuAW
k9sVxuWMzlSqaMSui3TN7u3VjyDtW/4uyYzr5uOCKAvY8PqTTGT1V4j4Bb4+y98J4egrO5yYLqPm
48AruBauwgfD04sI80WLTkIjTXa9/TPMvQWrDWDIVioNKCSvdjr9dLRvbpAE8ewWpXNGaWiOLzxP
9qWYrqZABs/ca93sxnSZhBu4zJNaX3/hi1TgcU5XUrBGk3o/L0IJW3RkXHmhVSM/57QUsS4xTpvq
GdpyD1qe25Qd56NrADs5xZJ8M1Zja1V4TPQDQh4w6vN2Hf2laGIk+DOlwZeeMqb7q8QhT+h6aAwV
W6TvuTNM8c7CXqqqTJO3G8OJxrN81NewvFjJa/VoYOtjdJq9IMRry1sgMykx0IXJ2C4JUvFGZiUM
s9Y2M3zlb5flbT5DMo8tkH78YZnC4Ax2r94Q/9aVmu4ZqCYjyq86OeMIjOmqdPjtkkpLmfaB1i2N
+SArJ2Mo1RktOD3uDJdhbuM+mpnw4ta44uQIWK3njVl7RKYjuxOjaGpFgJ7mXRR8frmzEoIdl8Q9
IdGqkYLUb2k3nQFaB3HekFIXYb/8sH33Qf5o9d3v5BtHboundpN/19XFvLfmlRhH/qVhydPbX8Zz
s45mzseAdxTk8bTP4HVDYlLtP1gnEYIndNdKkX3NHkxrDLK8kP1sRRnvKc66t/G6deZ0JXRHyzWt
NnEdqS0TsXpjPzJX4BvuxTQltZYuCoNPj1cDgx0xDKq3Ki+9E1LXtZhlKIhn36gOGBSkfhBfPqcg
OvodQxNivzAbyuNfYtB9ZNE90U/spVLU+01oozbiZm8r+kcNeDSiuoY5jBFj0Yny85ng8kf1NQa1
xsEII9b+BNqT80LvudPjarRDhHGYABXSQcM5SvyH3Kc+ayZRvsIIsZAxFhOyVPz36f9x+Xa0Z5AD
lVCr/69wlwqr5UGS1TSpweGPmW6Zh2B0vhXArhpbzjXTXql6P+j65couuFM9prApTpq2uuzgerLf
m9FYvsaoik4zPbtAbb8eRw5rKgQNswfmUjwU01yWhZLasV6rqRG80bBdk5bHmzZEE0ciJ84Bn1gp
miT06yHqq9WBaKLt2aEUBHuHswywkj//siNj+fZY4zon743OFgLBoINHWcALxhVrICyoMvN+WsbP
Ue0JvI9TGCE5igI9OVqGrQ7F7KPLfasZwppo7EPCZOU92YuDl3nWlUexHjUzb6Xkz/a25/K9VKwH
OKABV/NsIj/zyP6lB+Edo5eWaAyd/P/QmYUP89Ocq9tfSO5XjBZYYw7H0d/fRXBxwc4jTtLd1+cK
iPJEcQXSbKv57Aksyd6CXq43XPcQ5O5/HtbjTQbF71BCD/DISU5HMttahNWPysYWJJ0LTL58Qy2+
RC6r8Ah+VhOT6aJsCq6hFt9f+NnJLGggbg0wn5R4oiY3ItNoZkoAt2zgTfD/Rv/3iMk4wDgmWNOg
Nr/t2XiUpC0pGSa9w9FH9PS0Hj5T3RU0JSAVrmGHODjm1cb3dqo8QEMkMyb1zjlxx10Sshxt3VcE
xx/ItUbk1RbKLdP2+626FDqGAFl1ALnS0C7ErbXW2K/njHLO0F5RpmOVi3Ad3IzXd618+sYtCwiY
89kZ2uXIWhoXNI32uAhAspP986BjPt7bbi2Ynt/1GDsyJJCKySr7sIhbrhv59A/IhsTu21AVJRef
11/1CayRW+82/Aqbq7V8QunDBrCdwYpHKq/SaCjRCgMEyVr8vvtP4QzFhSPT+P89Od8M+Zrhyzz5
5vMUKdJaZQR6Vahxduf/cPn6SyvEkCNMRhkaA5Q+Ch+U/zX4t1wlRJeGj3emGxgampIVX8v85Tpq
wwa1yq7vW0jctCPdy3SD5q/o18r4SOWt7POjEZ1Lgw3hm7q550poli1kvOX0h1vLR1YsNhuLXuhl
Qx8JFfU10eiz+WKPD9xJv0RYU2kK2l1lcEv+buy+tiTscQGm5GaCr/HMyG3IidYvPWmXuXKKVLEv
491F+B+fRFaG/0Gy/nIZsq0HU40TGhDKiaqD9NLFrolf48tW237rJY9WlBmjaTY5Dt/BbKpDkPa6
RqIUwq4XrAwb+3o2yMHpo4KnJTlko5JTL7sCGLdRyxK+82qFZlcExXKfVHJynSg0SHV+IvK4fHAr
rC87KFuHV22U9KjasHGQLWA5X8ugtjSr3DDiAFnJLl36DjKMyHjJI3JXBUT+Xtf5RPqAWpOHOe5W
NowOLQJcTfq+vuw3TzGzsywmvFVclBMHbLnRZZL8p3YJMmpxAJ/tfOOfvmejxt7O+L/GOtnPktng
DjMXJGjHJ1CDUnOM92C1PmBickEk62jc2DM8UYRBE4dND+czS12JbxCcbXWofAG5FQWwyhhz+/RB
09tlJ23URwMWDJm3HoPn0EU86UC78jJFrWAxU7ZXLEbnwjECP+hwqHwVVUPmWVeFQe37TA+ZRxc0
Dy4G+vVY5XSE9UJ5hd0qT+WJSDSuSGXhoqtToltELfix0rvfBsLc5lDNmtLcxkDtF45R/XhMy33m
kkhK4FC+0DN2BY5DF6se0/k1wdhRDmX7IL9TNugoWUz+kMoE9gZDZACORdyofrceydZyTAEAC8A1
Flj5cUfJZyGuzvqMOzXjiAiD6rb9DNGE+tjJXVxTy8/FMDpfWDNVj8kj6hLiDdeUqxqrIaY5iL5A
lMoKW3HegAIQ4HnTHOVBkP66UDokVQfFQgqfQyAZXRiVFVAXMmWl0zvgZzuYGDUHDrcI4z+lsD9k
zhvwg7qTp0kj+m9FKtr26bDu4KaGWM4C7STDH1oMWD82myO9Mt6llwzHwR7D/2GpclKkuxruWZAz
3dyU0q1bKDVT5gSaQE2oMxqMx6WHmnHSQ9CPDfH35tbUZNArL9Tj3eDrlb9iQ2NTLHLYBePO19ts
iF+l1kxX13LuzjSCe9J+SrDXsWy+dp4TVCXtSa5eE6L4+8lXXEPyI5VcuIG61+oXQc3ALZGbl9Zc
IALhrwLYSxAFlZ+hkihUdBorso4S7O3pXYcsLpAQB47K7gHonLR0CUj/V6weh2u6XB2WkJiZAsxj
tz8k4dw0YjP1UMtnPAAXZAXQIrmA5PZa7MyRy57a2s9mtr9+ut+jIPhqapfMikTKqyzLDmYrR3OU
m3AxT1kNtjgxSd0uz3AiVtRlpYqEzogFntXi+8u5U/S1kzIAU0Z2YfxfDIiBnPX4d6H3TzUckugm
87Joz4z+vR0vwvDUC3l+Oe1shIEvwYFV3WtZGW1zweWu6SdDrlWoimvqH/BoH859UOXA5yrAs6qm
TDYNJlv3M5dMH+xx+y9GMm95ORE21cKVq4j0tChR2E6ZOniz1No6gmh6zc4duU7K5U4Y1H853Nen
ra59j75kbnYhavnxAhEPrKejVI52jnpn2ZQ39GeKVk/ZxA0Utx8pmzPyf753fz9lBIK1bu6YGeyz
dAtVhUXmoUCN+oCcryw8sqzbbPuKu6EACSntWZW/wVJujJ98TfS3bQgfqLc9v3MxHxPya6tfPzsZ
RigfieB6dqiNS3h6IlV4sno9jcB+CYDi8NLGmRe5BXaXZDwi6vxITec6E129CshCrxWXwutqW6w3
16MJUdtJ6ptui3xR48Rq1HAy2BTgdZN5hEMIsfZ2W3OCY2VbsLgVEjki3D6fvhU6ggnC2GtMId8B
/5keheFKxJzEgOd55Uajva1kwjDNMjLpOqUYAPLydq77tB1ivq4fF/nhH3m7xRbieIn8yxcOAuCW
AKticEhw9EK6xFtHAMLCeX5EhsvkCrb7uUdi0fRTtlJfNj9Bn2Hq5a/OQJ5xL9hENaIUctvIcQN5
ZlDKOCJTIW+NqLByVlpcQkstB/B4F9BQAyLaqjg8Ix9W0onUQYWvDGgjiq7/q9jjDXJcMlsT8znT
83HHGuHWhjd4cVGbUb5fhL4HzNfbCDRlCtfnx/rx02Lm6kzStoG0D4kyR620Xo1tzsCTPYnfTXNA
hWTCmum4jsig1suHvZjJO8KCkuIxnaV5pzau9f3K6b7v4EkcLYGkmvIqGsWvq5UGsvr3ITS84fj+
B+sOYNvE0x05UOIfsG26HFag964Ec3EA93gK4C8K10M826ds5PFxmorESn7v8iaYy96FY3eumh6W
e9XmoHqz+Mu+R27vLVn3gyDJkbIazOrvBVK48UEOc+V7cKrE/b3ht7ZhHMRkDECJ4/6SEIjDrCrs
nsupsPrB8s/EHJy47KI1NSTLfl0OjaJ9xhdWX0AjxALkSq/BtX+19sKnd5lcvt6zfbIOICGPam40
a5GDAy6G58ob9Ypr/tVJr3M2BmqyF8qlZLjhULaeyEM+ubs9kOS8eznaTiqrZSK3XC7B3IEUHp/d
j01yp9mztX7DMkPyGRcV1gMKyGSr5HDf1XmmNSajIWw0N41n3wHMELSEsRrWzkTBYphECXAMcuNn
tOhKqnSDWEObPE1ElG0LtVPBG0bVjldHvQJ3eoxmGVLnK1L94DEfX/ZiXslw3QaGMJfRy/+jmsZb
ex6tEubequB71AHHJeTUQjCoF800+p0pvbsxiU8tQvViVlWpvOf0mWWfIs+cjOqsEw55Zsiz6nlu
QRGJwSn77M/BeP4h+bbLI+KdyxRCEVU6BjrRNbBr5YmEZoDiGFCE0S2kBFg80RGdM887gghJIBqt
bq8Tyt3NyLrXNgs2gIbJmUyG150BmVeKJQywtdKPEgR0kRYSbylQZntnn20NH/SHjfaI+hz5pSft
PP1lQze91JKtGQ26W/5yM/7HXhkDG4uPpBHSkWI4YiD9e9FFhDSv+k3cdS+eR8E62BNIqDV+Me4G
eqsZGfGx1PDHA+TSeuNqRSJK7SRv+7kmSqkps/5FlkQbCnaaQ9t/wFbUAP9QgEAylbypSeUyr45d
ADJHvC+9VNgYNWghO4rmBh17cwmT1uZu1M79qEHNoG5EXxuan+Lk/p7fXBHnrdMBDVQKSzeGKB3c
uZg84Edz6M3gRfaLTzIDFGliaUvpqWPxcsGBHqFbcM6/MLUBmP3xolYho7sIXJS8EhW2mwRPYA/8
ZBbKWdQ76rGzvcORu0Cl4+LnSPeov4QXT5osejNUfJ7CT/5PN0pzOM4yk/d6RgNw+WhrxPbQdVO9
qHNpMuvKaYDJDdgQ7IGSY6EEndBOvlqeE353Qt8wni5xtbjs+oA9LA7qMawkEd9zUBdcP4ZNndXo
Peht66oraeG1uJM73tNA5p8q37axXrTc5bmCAeaiFePcKcca9p9M+N3vb2L1MEC87DsuL9ZB2/vo
vAcTeDLBQUC2T3Q6WHeo1D+Rb5xmWOUBDi99pG80jt2W2bYJGorGjNL0Gm1h39qWJ/SWpgHa6J0J
24VntBW6ijgO3pkVhcj9liwnXEy6DfP+7pXch+K8XUWI++KqTqlVQj5rJt9U+FqOokAUN7YH7XHM
FMerAImsdMGzqntAnBdw41xg5WLcJfQPTvlhX/oW8t6QNKL5+4C0ovQGHrGTYlYfJxLC8jgfilxP
hxKikONy5PD+BcoLlej+q6OvFKknV+0/rP0eEoOJFMCUjQMVc3f/G+JBPglWJXvVbIDTDhJltLS5
jgbHFWfpFmvOqxN/V99G3obYoHsrc5arcuCwJnpRY4XSRSGkjivLC/AxzLdqwvuF7lzAtutoJAWC
O8zKMJq+vI53koyOHSFFwURBtHtTLJ660W9IrpVeEZzSORGLl3aHvV+V0QQV1r5trOguiznKj1WV
Mw5cTSpi45hXZ/nKcKSxata4gFmGSmuSLL9iz6joe3hoEFSK34ksTFHOrecV1KfACavRnlgy+yTe
e86GfoWFH7cqnJ46LVmg9f0iD/Y8IaNxeZq7HTOet8DlHMJ5m+DDG9/eJHF045vIfk2kHszqBZJg
/KXyBy+ndMkyrLH45a4ADf2Raw0qiauts8xsBx+lySj9pQy7sdaLqUxO+t8hgkBAz7g4OQ5ViGwR
JmxJPrtliCXPWuQpXbXDecxU1F6z02Us1Gccqd2uBQNCCLErLBCtw3dLpPWCXgaFZKDR5uv6MZPY
P1ATH1wNbSFVNtOXx9pwLWl+vJvvadH1f94Lgbk8e8bqeLcq4Ws40bD42zG2qhdf/EIAE9encQ57
HZ/c9jSH9g6OCCgaNE+834zPSeNdmC0lXFIEHrkyGxvhokNaS9Jv26c7l6Xa6a/Hx5GLUc0y0Ubm
qM12YY8el51iErbXrzTsUp6kz06rUb4hJS9jF9NhtQRbgje+jNQvTpueeqMSrdmrrjpCGX0fLEVC
YKI+9zo2XkRuEjw6PwrQBy3Ev1ZWbennjGvejMd8EM/In1h2Wcdgk57JAEVLzsDd3AsoDPI4hEwt
yMORfBUVPm/x3ZsVSj2436PbqX90hnR6wu5bHV7ABxyOoJOaTMMgkIbPAEftnvMHdXHrDGfUfc6K
KwrJcJ0+PsaETqBxuhHVB2k8GUJ/0wjrX4nUdTx+r1+vkCbs5PJ2kVoELJ3vLhT4xcbrHI5g1Lip
dz3+IDCdivk/gh2CEghTEONaAs8XOLpjN+3Tt4trjVcWkexGW8hT9doZgTP7+sVcxhHPjlXBXirE
K3ALXMTplzHd8KxG660urU7hJbBwUBWzgJTlyf/SHbWsGC8dqVYsyqjOwJQHdYePv001vZO73+YQ
UyPm2oHtCd+VhuwhAmzMqIflhTexwU9eij6o4C/KWiSXi/BcFeXJge7sbhkC+uVMBrRmUA/iptYE
DfOcsrp2Cw+PPndAH4Urj9HmmZxgkYfuw+3YEtr+WGSAN/5L0zgMdkwVLrf/7BZuMPIo2VFiwsXt
0kwkAdCVpnIKL0QY93vFiNMNsynMP1FQB4extuOA6q44MdmgJn1vBoRLUbb8JHm0CFA6ju9XMU/E
1uwG+jWkVqe6AiLMo55aY3pVKp0epQdjv6gVhcWOJ+Npf/L+tEGz8y/6sn7bnDd32yQSjmh8jXTU
+KPM9zMKDX5yrjtZVdE5s2D6M30bRfoElvk/i0NKc24YxfmxcTsoYyrsXe6Yf+nW6gYAfRAtb9XH
KQUAshGPyvJzfc3hYzaNolBz1uJTzyse728AIcu/SMH41NI9izZkwjnfxMkh9m9BJMJtsJvw+nca
kBZMdv8YEvdxV2ngJWtSOWQdqAPtSIOVO07lPT2vJQXPe3+wdpqXA7QNrJDu+S0LGg/A3bp7egqo
DcxgoLv5W2D75PVFHsHq2xNCEFWqdUDK10/VROO7ITzQzPAonL4uDBy0E0Wj5L+LPAu8A6ES7jTp
IDhvQcumQaes4SCmKQwOLw9fc4RHhAibI5bQBNskYM1pbP8EH9NE1lroZXQdvFTvPWF2hVRLSxox
ycwKBc5cQiQiaPrzfyvt8WM5VrILgnSy0jatqB/bf8AX7CAKRNv+8FxLzDA2h4pdgyMrP5ErXQpz
jBTsrYws+nV8aaO+aaXr8o9aHoqRjT58jOKKGmjVPISJVdaIdU/sxm7Po0ki1UaUJayAzlCbwrQ4
U/n1koS4sE2mduvwwm5yTfLbb5GaR6ZNosCCZzq/yl82jQRy0rO+VqHT54fHntw/lJU3tYat478u
YXVhv3D7PXzY5pcw7X+3kQDUXbhyDmYJBKVOvCBs4prE46jT+RYCts+rvm818DHqV4FLDQX0ws4f
kf5Frrjtb93/5cWLlvkH34UCAxoyJu+TGg6LfzaCPCAeV+9TTrTLn4we6978HQTdc9aHUqKzPzUv
ZTxOszEEKpSzq7Oxh7ZzUb4JANAG2dlidd7jc7N18zQt9pI4NA6Cb+mdnTW3I9qcSG4F404hDRPr
xVCDIMJbnPbuqU8SXw9p9hmVI0g3kB/ECSe8nGB2DBawBnOvtSvDJXg4AKYC2J60jVnWNDNDUmBq
AFeicYUfnqTOftApeSkiGoLG9d6YhLp4L5g447o/AQad3KawXXozcRPvwK+KaYuQ22w35BrCCWFM
L3Cv8L6c5VGq/vUg09KSSanDeY1oLX+C+ODvrCNBhvN7+YAaFg0J5zmSs4Qjo+TYvv7nIlSOur+5
Upw+mJuet+uPcZnkByRhvzWNrSYthwShCWzBPwaX79wyesOKwFRQQGYBtJgrkocD8oSZpGlCeXiM
Ld5EenVMOGb49ue0feSahd19J4CeeCnRq5Q3oZw8pFSspCYLP97XCpCKCDfCE3vpIUoDfJrftNwV
05GkR7xp9Sw/jv8GBVF0iBxK243DiJxTvCz6c81qyQ7KkRPRsYJ7xi/4B13+Q2MG1084DVMvqKn1
aIv1TtWonlSpHOn5ykTfzx1gHCopO5QKLYlO81gZjeo0AYHGiDFs94m618g0VaDwCdBSjnGx4hBg
x8O00pKtRcFW/RkYuGUMUYNC5kJ19KgQUsEcUlfzDRv4s8ZizUHzdE4Du6F5etfZ+WcMRBStjj83
piDoK88l/9a14L4e9/8riNWyTdw0DqLVhXYFePdCdD3RlNHcJ4IDxDljnZ1huRqTdW2Z4kZjdnKA
zMFmJiE/kmQfATxSiSmbK3l8xstZxwfDIGyWK7KEAbpsLjNf9+e3sYkrqRNakx+93PIwcxQ32G0c
flS6udyPleNrGpwcFA5wYswGajaGnJBrWeSDHs3s0tKu5mu4mLiGC6/h51LVFHNr6bO9M7IBUji9
9z7aAmH/YPEuBEhch+3sQ0x41nFLMw8VwIhNSIkGnJ3O6mv7V9ryy99dDeZg83VdwAWWIypZ1bk5
Tzic3f8jRRUAGDQXTpEs6iAOTV/V4hdgmEYSullp02CmdKbfLj28EtDUlxdvSsLGZRnUh3Wbb6QK
JuFBlDajqX4nKAdi5uuder51QiFCIEkXURaNp1OeWJBu/fmY1XuzFHn/8jcvzFqmreqjSPRNaJ5+
WhbNQIdfTe1mmrmg1T6BYce3P8PfryrpKk40IuU14qfqkZfGpCpjQXN6Q2dvoVwkZEfGpofPWM4A
2gB8nCuNN1ADI6gn426SQIXR5kckISuYRx98CXJDVN50N3Svhx1sBrp7ZFUYTPsi1VFmPv40Qj92
7HAHFCS/aFYtb7K9iLslbR6wJE/T/SJ8FU9iESa2uPV6XqIF3n24p6Au/IzfRpWtW+NubshcrZTI
XnuHJTBPB8m+pTREaDrc7xxksiGzxrv2V+Lb+r4LU2FMwP6NgAMF9St23N+cxQY1/aMObCttGlCl
jWAt6onbIpBMv7NCJALY958mkm+/xT4IuSeT01kK5dh3PFzqk/hHfgRJ0/2SSsImwvAKrrhP+6aA
+8plEZWD/HUsDZTnER9eyczjvOetasm4RxgQ4nxRWZoJgzWj38mvTP3U3PzDCsxcHWA92k55d2Fq
LR3ZLga3s/OFHnDk3YkxQgZRh6a/zQxsvfCXjs2//vHqNNtWLlVoLF7etxS2wJAI6FdSfmKW1JRO
I7WI0WYLcEhfpjkTSgWhPg2oFTwQTXVLHlhity2uHqZZHci4IO1bazGhTHpCwz5ebW0VdmnH1Po3
u3NuAWFiLGpbnpc8Y+UWghiP1WcW1y7mBJuBpUbW2m3KfxKyIRUTjLynhDw5pIhE5lpu+P7Wy75F
strJD/VKI9Kxcw6nNp5rReOdcX3sButE7w4ov3+niq35N/JbuDcTvY8q4f9O+LLJFLcvg683SOMx
OkFgxTdptEqPdGpPzebr/GdapE6xwrbpthpVXP+lnzGsMwGsJEhskpHbo+Tm/dGJSIYSeLvlLP0G
/bSD4Jh5W/EaLYdvr5a5GJVHunjEKRtmNr7YzSWIHdLAS0sc9VL8PUSobQffJgY1LMYVG+3U1wAq
14rhuWgFK489uF0MYvVmosNRIEX5EVPL6a1+Br0Y4nKy9Zu3Qt3q2GmK41Tb0gAAD97HYsFueXRM
magI4ujicWlsVqYzZz3SxjSXKw0LqMye9Z1g4Wwph6s0mvBpZSLrjbsu6+IK/7Qbk1Qw09qRJ9kj
m+gFgGAVa5S1tqOecpD1bnWuciFnsv2nmj8fMPmrCQMu97S8pZ/hnTnj2P+QRJU5lQqSq12MFRKD
8OpXgWg+z0IPteW/mE+lZF3WhfKpSarqraGBmHmKtQ8Mg6PCEv9npaW+ngJ1J1cMTPk+e7+WY1rm
nfvafn7gVaxgy0yuTOxfNuDWa9UFEuGEOc5KYt3/kWqcUXPts1IxTGaz5XFvkPzPg6aSqJBJu1gp
dvueFKz6i1hygvUQcxJgXQGugrTfl/63e8AAdUnlvfD/ysKSwTTxbNmjdolr8aETB5EZ2fkMqAex
2siimhKos+OOC4nKHl0+C0/UsQKrlb5IXErunJLPkmbUSxpaQgYE4i9Evb5M+08Gcyk5NVKYY5Z0
2JOqhfuNlk441/ar/pHtkR642RJdn0ZrR0jH1ArdPnabhCZYpjvEOJlfPPcEUEHCm3Vh/wLtCQbC
PefJKhLSxfKCt+3viG1aumpFy3wg23BVJZt4tesifC8O1FeHx7YlIRpJJwd2WkDHkRYAv2Ujqlpm
Qq9bP+AbtS46G9uCVdFgWSr0Ko3TQjJnnt6uPOLQWmZe/xAmLAn6rUzdPOqk5w1m9+GkBts6kO6I
ZhXQVrUTTcTib1yXcvHTFhskl5MDZlQJO1iBNWWTQMS7pVh4lv92D0sPYmEoCbwa9HkFyV2l+9k7
TB9gYseUh4/AZagg9IA9C0+8gRVUqI+Ik0VBoongfoTqixUzGYt6S5EYbEbyFMrQipOYb+giwVS8
x9xUq5D36zNSgRScbOtl1FGOTNCzf5ybnVIrgcPL2jeyloKcHHSZr7BuzVVHeahajkKSzBpdLPOa
fEOXa3RRjGaxD9zhwhGi/2JTnl2WtQ6/6OTFZb9ZjwZnSYEWcP4thK+Ni9UypCpoMutzIAZwZMSE
LZUgo4h/QIv6sEZ4tdcwmnsV3hTfWZPbcOqfey20p/83QgQDcaw/Wqxv3+ueaodOrbvPYCqJ3Beb
0yL2cNvxHyQdgZgrKrJo+3kpmvhVtlavp8Fa+ONbiuFSxudS8KvI+Rlhhy/wzlN0huXR46/raV/L
Wz3Riir9ZcZF+3thUWlXC8dRBkLbE6dpOhRSvbljI9nSExxF4fdkRTLrfZOZLVyiW6hpgUghlUYf
gmZzbwr0giMbemIezRSKG+4PJmdgbWn6l4SiLVLo3EXnCwmuvwwK26ob5Fo+SLh+jNcTp38T9W9i
2U4LbytfiEU7mll6I9hmsWJ5dTlXUVBwMHwSVxJ6ofjOFpAf9VIRe6BzRhU620bcSU50WINQQrI1
j07JmLM9vU4qs4NlbBqecGu5MwhozwksQFQG2s7GribV5p7B2LLhVbnCMwJ2f4wroz/EvMyHW7I7
xO198h8/K1/6GD09WC7AL8KIWb7mk5HRvKQ3DdltaDvQUKU5a8MsMtUzjLaMJBnqulzMlrAXDNyB
73NcPJKF375z5HPlC1G/8XAkf5WE2lE9nngGUY/djZ+y6rWuoAgmHGtyhmpYe7WTKJ0/og6MzACJ
Rg0fQJ/cVWnuzeGANLgvHGg2685snyGftBgrOVds+O4l/YFktEno2GAISlJehx07MaAObslJp5VA
rR/oRmXEvadKmn7x3ieH4BiUcRv1X+EJSiW86NhtLx2x0tb6sR9Ue2TpBsKyLc4HleM9y3kFoG2B
nSpLn4FwkdvUQAhmtFiNVYXHuf7CYipAvakPxWT1VojdjMNSAhuG28Mey1NvFB1eLtEQsYSznHwx
Xxg9uWi5QnrcvkKsVZExfgnpkzlMdwcNKrEUoo9OOz/R/XMSr+0OLkudDOoe9FIhn6fgTX0fVHPT
Wr9EuIyLz4DXjj36jPKob2N01FEF8XkiQG+6fxzhRYrBkpf28Pz/Nlia5Do/rCeU0ZAungTU0zcY
PECuuLeJhL7qrxUmI5gd9VXK8f6Vn+pA3bNqH2qSeYvIqHJ2pX/oySFtE3oWaEzeaqbYAYCWu6DD
OK7CJrPICgobwB/bVz+7J1+Klf1PD0Q/1rJ1Di+TTXirEBO8m79fELlgqSIaOmHYn3twqHlTXs/c
BHcjIjl7Awa8kNDEkHWHgfF1wouAkqS4ICQv6SwZH2ZrnEGTwhbQq3tPAbi8GBqvCCovb3BfJp5j
vpBA7KUV0x9Wea0mAyjT7ETSgX0j+lG/jS0I4y5FG8CFcBcCdvmAr4ykhMAXFrE8a/ef/M5SDBDi
lL4eYd+HIpNknfSTy8YnMVreEDMuUp5MHh18wEW3Gl4BcVcS4VVExEIr4j7dcbZYp/hsx56IRzbj
DQn6Pv2zg4kykLbL6Pajm6OJJdi1SbAjGjJZ57J9KGxscnuvZFGtXfBQT89rE2f7y0eydIAO9JQz
7PeUahR6NJ4pmsupkJImFXKQ2tzZVagxddeacAhIhmqFfqW4QhTiPFNrG9VWkNHiKdM/qRz9ME8X
PhWtTaEkfoWrQPE5TvTSgFeQtARoMYf4hn8wrL1hZ1FgA4wsRecL79uTbOB4SSevBmDgioD6R04J
IbL+rAgP0/08SEotmR4xPXdOEPQYdOii/6i1gFaD4f6u684AMCR6GBI1ZAucAYtGV+u+SfN3R2AY
3OSArDDz1AdzQNVElwmdU8JZL68wQF2Nyn4XbbGt65LcQBCY+QhRjnunzbPvy5SD9UCDdpwK/Viz
j8aYyh8nYsHERtz/QLwQhBgf+BL+vOjyomA+eZG9irWJyWOUIQilPfUUkas43ncWqK+vPx8xRDjp
Tos1jHIOiFRB6P/CHHqz3z9cDEtsGsJd7NxF5ZTV84sM11d803wglBxYvpLh707nARxKAqNhD4xt
Hu+zc5I5rBhjGoB+QhzUnYrdMFy7mPqlyfZjuM011bUmvLOPCu3akM8AG6Btf39CZGeWS+fyCEqX
E/sCbYlikCoDUxqq4F5QwT9XOWNfRJNBAnaUzmISwQtpoLV8tqcgjoOe+YkeyNRlrFuNarZ3E1hW
mVDWAzCd6TGSOUCnY7MmbPiM6GVOb4J1Qt8U7Bbn2q+WyWTaT5u+joJToImrtKl/Ggpj4Dc6BRoS
aaKZy32qDMKDfR7VDuua11qbVd14QY0HIWFFC0M3/FmivqlUP/c65bTsXcH5ebp6UHJvDoYQvUDQ
VT+DQ174jeM3lP0L7+G0U2v1LLnx3jSXW4KpOelNBwHJXLGK6mkP/aof/tNDkfY5GKA0f1l23Yeq
4ojyqPXdpQf3X2nX6i+LSssDWpzwiEbeqJLJz0oG9pGaYO8rlJXog5iR8dxTFyxglSrCUNQL3ayw
YeTITBGhryEtD74WPYYGQ0Ll4Ywa/1zPY8hAETC6ocqmkjYiuicfhUNBr9HEageqeOZ5MTADer48
AKDVMbqR025VVVJOdtEc5ktTHb1urV+1zJJVYCCihsyQAIqtTLFpTTZ2+OGniOT495zZVreuj7+M
OiS4TunBvt1w6bCXvJHguHTIAC2VYn9BZ+FFyPFI81bgvGH3HPBPZiwSzQi6ScW+T1PvUjqu3ryk
z75wXnBTEpzJqPabp3+dg758t9d0Qnu+CR86Icb6JCvxBUztRabENFlfG9Sea/tpakZVSh1ow7B2
ePRvrISLeRoEfPlpPOqaNi6aU/7Vd5HexrIvm4crYy17ei4T51z/bDDMpng/9c0nNYE+GiZlMps/
2cJ3I1WrqGhGqgZghQIGaQxwxCb+JIriatkh14A8tJfLiRLTu5RQg+OnJFU8NSFUE38RWcnRyQpq
X39HjNfcxpKrc7qQbkyfxlPE37tWCaN4iV9src7WCa1JaUDdqtTEhuocHxaATJHocPtlzoQZOldr
9NCI5rj5vGiPptlXtGL9/3QIcbKXmFSbB9xdxN890nAJIAwwMT2xkQtBxKSLAIlHrMqBpOLaYgKm
Wq1i/lH2JqIa7EyR7ztakCKCXaF728UYnQO0hmSvJ3vDjMROheXT5MR4wtFnrksUlD13cvpBzO6N
lcvqJObJiG7/6lq3P381SLqVtyqS7v6d/Ti441ul0zwzAYGCOBPAzoFiIA3ZGdmFENVpVPOU7GdP
9zzxPiC9D4b/sNC0Di0JoKouy5Kvg+PT12/LlmA95ey/y4hPCzL74QBiguQfzfr30HFDKHHXGYLV
loo93ZDtVfZfX0BD7zglHpxLKPDpeMUQzT2H806xausfD4wblr2RytzbLBAe/mCuUQstxFlrOJ+E
R2D8BW2oo6pQejbAfb+qEjdoh5stuUiKnm6+xG24SOj4QZfqvPV7W20Sf/eIXf811Lr1jlTVWZg6
V3Sm9YhhcJpO/kU7h3Yc5kXCVgdr/DCMu1Wb/cHl5NG2uhFRxdkeY0QXPID3J5y5zPQnrNaD8jVW
x3WKOfrJZe6DdnH4f6O891F+dYIIeKciZipXL4Qa6sDn8Zt5ZjuUbTKQOeG0WYCTDw3PeKbtL3/v
NBzlIHbdpKm4BrLA0ECjjlYpugNqJKipo1n66CI8NnnK7sBcAA4JtlVBdKdUUDvXQDUo5fQB0Mf4
TVEi0nPFofGAEJh4k2xbrzRwXpLnVkK/3oBXzqpoKg45tv7T1qEhsABkTJ49e4T2YrjZYClTUW1N
JVA7NQdjbiX+UYGJ1HuhVdBMmiqUSGKxLuqTrUYqXnoznQy2xKZ4Y6rZsn7xOcTBzCiL/vXsZn2k
vekZ4Le47aMuxXlXs1+3n1mxVl5FTLHPphGxqIGTxzUHlC+ARzBtZJcudSyqR5nNpoSISzMG6Jqt
wJoUGUFSjoAicK6DfN7nxrrvyPhSemYEa8Xo1DG4mlP3QyJW0aXAEJ3Mg6jl3vVhGozYZlAKUVSL
FGxQzm51sp32Y26Prg6LlztMDu7B95Gf8LlDsDZtc32V8IJt426zGodu5oNsOqzMbrmZMXVXstBi
BtTXyxNwfu3i8det53ad/JxP9UO/NKzr1mEZQVwEiTIICXY9iWq64A10ynk0MOve6EfUit5Ur9iS
uR5b91q1s+vq8aOraWx8wVNOkP8E1CFu+5rXhZX6JU58rjswTy/YP3irrkKasIE8xm2fHAyY6hZy
HLM/Ad7LWTcRd6yC+RicqjD38VRY3rod2yF6cG6O9Blm6ZGMK07EXsyR0naIGLGEJmw0+S64Hd6n
Lvu9RFhOtyFZ0Vk25TfYi0NgIq52vNvgYyOAp9epG9sgbg8rql1vTN0xvRquMAHx0S+dis0nAmmc
cs7Oo+ENzmNizVmhoupal/3fDv/PZkKDJc3KQuxePt3A5/DDP20l5270RZFsXI9dgcCGLUooQcKm
FJyoHuwCzrm1pN6/9DsZv/54pFrM9NrVrloUuT74zO5MeMCBk6kCBTVcz9dtmHEbE+vUOtIcar29
y+81pfZXC3JKQbEEi5yDp7zzduAsSbTE+YMdFTriXWMExzSHIKbKkVtLaVor/7IrjWWJqdvXiW9r
TGThRgvUB75Sd6VruqPAxkTJakDao2T7JPZlwFCqTRlcCsC9mF0pIEVpw43UBMB1BSqpA68DjKou
nCRP3W2Nce+tKyCbvipMhIE8q45atoD89slhQJPefuOqpfQ3FM7eE1/TG3q2pdyxZ9OqEWaVfEFl
Eg2m7Cd9gn3kfM3jY9mp5bfZ/ndotAJ4x9s0WdxTfMfK4G/oL5cN5SsMR7R/OR/UC37omBNoV+qa
sPOkOqfXippSc3DLpPXnpPT8+KhQOI/CzfkA8nLRmyoAlutpXLsyFFKMH1vNim4PV7jF0T309RMl
BvrymUSBRf7DOFafNylFkPRWBdDToBczhBsk00DLHTpQqsg2uforOI/gcT498E6zSuCNkB8HmTTY
DahBGZclRo7gJIh9NsBFNz2OHROUxFiV9Vx0ArZwTMB5R1jvy2lrmB4mTawjWig06SyjpOKD2hje
pINR5JxEboQ7urUmH6l82nICM3SVIPptTsl1PWZVbjoHd6xsHQ5yBQTEJ0P5EQ0Wxr39muvSRDIc
tSJdZS5fvPxfV0lRco82XwQlM25ux+2YZbFeW94P143X5f46LCKzMm2YerbQ6a5CA9ji1rIPFjKT
2RzQru9zrnAKOV9LBuG3/ylMaO7D/DNGhO4VAOYPbX+3QAmUyyosePHu26b2bJ4+xP13r1zWLYYW
aMljck8xKYvH4mYcc3f9i/N3t5g9gDayWB26id8UOArMBxYIB4AiqUEtCec6RR0m2naIU0cOYV2w
EKX1//7THgva3hcBkHbzZOZH13QlMXKuN0iweg9Mj82+Mxa4wUXewRSJV+viVblrqKzaVnQeInAJ
Ee+7fgQ/LksUnmqgU4QfvlIn+O3W0SZNV4EEswmfwz/L7jrQtxcZmcIFjtE8fsIJB5XKoRxjb4WY
5gwy6DrauRMk02ZeygyzToTcZ1BeN5naSTavHl4he1XLOVwR1DP+on9xgRF4pKXrzXTp6B5jyCZn
F6UuQWr/Fhk/V7dxTcPg84kbL6vdMjoeM2qaw+DzflgXsPBtOEGSHysam+k65vEdT+HQr9KRWAF6
nuF/NH00XeJRoubiOGlbnjx9pvyZhqmdqMiv9QIZ9M1vNlgn8TBjfgczReajDXWVcU+Oqc5ihDPB
8YpVEsrkExIDWHxDc1CwaMojQ4cgN59iq1jVPHHRZWoJNuQnJY3rG4j2DfqpFR42mia7Osx2rKUS
slKwCpG8Ok4KyrsJpw1MNyiJcBlis1D8D23jNNIzVrunVjc5EW1m5XVeymJRin9hJYQ9cnICpops
u1ocQVTHbV6xE21SbiQbrQk0bgjH3vpFWjGiMTiCGOTFpEbEOu23or8SPsgPcYXm0it7x5FpTHDD
5tXaa5H8gx99irgPoL00oaySRmA3sFXBk+xCSMD50FwEKedFPFbKsrlILoh7LDUQK/A2JqPCefR+
XIZw4gR/PUFYwCU/9x9nRsl/MPGRC2l1whDChWFNg6EJQ/06egWe9cNaNa8iv4Ar44XG3/yg4Ovk
/6UIr38fFftamjIZKrhssR9QN2M+TdFO9Mf6lY/sQ0/+Hu3KloaZze2Jsa4+NdHLhivWjMOtCEQg
jjkRldS6pMbBJqHdw33nyFqkW9YJHqTF29ojjnnw8TW3uBKps2pMVECm/SJcdXRw3b6UW7QS96YV
l7O9IzecgOdO1v/dDNY0pgJSDM/e6HrnJvkVs7dKip0XdsADEuz7sc14vMrPCxTr7PwKu6h9Xmr4
j5jfxNbw6F6PZkSAP9H17UTvfgTzYTJnY3SFavEsOV6bLzW1IogO1bvBNkj3gTApWKwufpyDLY2Y
K6WhY2/3NVfrcWltc8e+c0ST+oeB7sxQMGloTCkvUM+vdQJdH2tvrJHRxVrIhSyWPM1ZfRSJFjx7
pFTkYpC+jcFMp0B+lYAY6+i2gJpWEymltsvCK8pDAeO+Pz8omp9XuWGoLakZrEberSPqXQJYJ/50
qAzZJcn/YSQgmWwLL/1ZQowdCKRSbqFOJGGbvHPbKazzy114ygtMbCqFs5mZNCQiAvXVRtNspbO8
r8GZFzMsveLaCTtfDvQeRuRwLjn7af5oWCCGRS+iMxVnu7aEvemjH7r7ySqKZ7IF+nIcp5z9CMEA
lOCQbyIBXwxGJOvaVaDGrcU1C+rsG1oGpY0xepZn0QvGfXdTHZMLx1JYBHNQ0ma6UMDzry9VelNY
xbkdSrtX+EqQVA+Mt60eLXpJ25gCyK1cIN1Yd6QzftPGL+CqfZKUNwsApqG8Jfy3n4ku8aQfCy5j
3LyALxpVbUh0s1mwu7LznCPhN52dHkeWBDK36ZRzdUPStwII0xWI5X5vj+eU73XvnhMLbivOllPE
rBWzqf8HL9+DopkF6hBVrWsslOw94fbnWgm1CWvIoJaVz+lOzGBawAE/7EqMFXifRjzgl/FbGHRH
B1ldxG2nghrGXzyb81BoIlFS6BG0NGud/2xTFHv5hrV6Y2MKHUZtpCbmtrdBGFpV+szK6TpFz8Ib
b58+MrhER9RXE0PmRvnv/QsF8YD9Mfquo/qf0FSgWDZ3aEYP41bA+LsgLxgP6kKDpJ131/tRop5s
9Llh3XwhXDlRLSM0Aw3ZD78Hw797mKMARD9ahpvaIajmTuTqLnK6eZBiAGAU4eCFHqZGHFkFaOhE
J7571iIy+psiAbWhezBIDUiu0eYMsF6PKaY6hWa2x01H3mO4lb4l3riJSLsDwz52r/crfTFtFqpX
wRT0z/SGe73HFDmWEsiDJ9Afc73//iRAijD8BsnvNI6R+/NmFykn611UANYdR7wHCcBSatqvPe77
2FOsPDE1+6M+MXf2A7lKHefYCmkN0TRiG1bFCkFfniQ6X5zILvg14UGGjLEgqDS3d1Yg2LQ9cTlV
tG+kEqDFpDip6pvgiBw1w7vRl7OiKbKtxN6X58qrTkwDFtMxtds3S7xbv37YwPaoSeaJnfndCcR3
DMgM/LW5nUGx6bM3JxZPdi28OztxIvCCXV+F5cBKw4ijtrAfpJZHtRqZw4prGRjno0BC5HNbsL1V
KDU1EqmBI9bF4ThQiKE4HoblgSpN690Kgo9SedOntIvYfVaPeDkLRlAjkI70bOEjIsw1zB71sRB8
Q2LQuWLjse465QxLbcDVJ90h8Fyn7C6GrcZZsW5fzZj92pvTmgE0mMnWHSW4sIaNov1aIU6INUMR
2w7UNyLcwlSSIhi2e5iYLFpH5xH3qy2aF3M8rGTmKxaD5vrUIM2GbifaTOjP6Ra8p1f3lH97n9Kw
svgJgtM+nENTWJwStZDU/jCjAf++jKeBftYqcCreuZMyTyxc9vcYSU2Jg9t5I4//yjnZJTZS7Yu8
6r3AGoxl8qCCFQM8MPKlVtgHao/II/OlinUr740rfjQiQQAcV5N16m6UnWeEKPuH27jhWaSsOJBu
qToOMrASiQRMUghRBy6tcwA6FK0tZR3mb/yrTuoX/aeu7r/CvjvO6Iy2s3QXMvnUMzsVz9eRfo0B
p368uROe4EQ93S8X7OY35rTC6pG06cUAOMaiLWnUjPvuWYEpG7SpZe/lO7tVxldUTG0yi9w8fi5k
0ok2pi4wVu/0LjcemP0Tow4QZlq8gdYVzbRCZxUp98OaJDtO9TO9esGXKgIbL/ig2M+1A0IxYkYK
PLUcachLDjJOLbnqiWZ42xcbZ3oiPmNEcOfICVRxIBQPyeykYPVvO3lF+b4D20TJ6xEn28Ogph8/
TnmQucJlcfENWJArPdDVk/VF95/RkjHPyccOD7J5Iu2UtVrlJx6eUQpZdjiuHK2GVIcRTFa382Hr
GWYngGFvbF/SGtsblSrv3Pm/Iz2FALRp3u7OGGacppjid/2dL4078+hqIJ85KavIWpbOALIJ1XNx
iBcm9ZYB/FKCDmtvsatN/DYzsWYiYMmSesRp8N9MwaDFy9SuPpK4p0N9fMhCErULfV0obrYgK4C6
tBt4lYuz3BYASWY+O/r2nii8gVBfdN6yyiGrGcI47Q8RisI7imXC9omsveryAuch7RpXHWGMzgYt
8Iu/Z5RG9LuiaSYrxZptFekS94NMfBBytp/wllojmTWId7aiBPp5eafcuG0iKifll9wrjpN9cGGk
OCkv1eGfXZ9rYwXDCgPIW8PQVcPAl0BvHqwisrWz4EjHVwS4V9gyKCqFk4gwVqlwJmlw8yrytv/h
751j1bZ+fT4n2IU5waOaue6Yh+Cj43B11WG6yU9DhnIriGRo4lUYIPslmCRCjLDuYUJmQIq2vH40
/flLkgLmPcukuthPQ4VGOVRNW1UH2wi1Arf4wOc8evOA2C43Vabx9mziEpMNkpfp6Z5j8+3DcIwW
g3uyw253C/43hDc4wyFrbqppwBKwWYbvY+lwXxKwYwIp2RWpGnmho/Yyk7dwlwewx9v/DhhaLgjJ
/8xjNDW47gSjGVTEOvbM5IVJhlli7CVKzb9YEBfuTsItZV8G92oEfYs6TEElJKNJcnSO6xe67JVe
qmc7KRWz7fNKQjgldjJ5WoVJrJ3bThrLWs/k3I1F4Bw8fB0EsmugZ/yHyvjsW5Coc2YihzHm9M4c
3wFFdyHa52KoU4m8XoaOtafydqq/I707A3aVeYD/xGZ2s9dYMeG3DMljjWSOnZkM1UTnZCQ5JePL
fPVK2gE50dZmBpMNpbpjkdnxgUIl3uDBoFPtiO/3SCAYtVu2xECGqbBG651Z5IEY+aAYVlllkryI
LagTQBSIS6hTjfA98UqdrsXSchM9CxJ/dWcD7MJgf0KVjgDphlz/McfVA0U454cMLOZ/CqycNv3x
nDDsankyfB50xUpzf2XJGuDusEIRV+g9F75RIcztghUaOfGQLmLTa4VuxrAv7YAL/BEgaxrSaMxf
lIlnliHcCLFlMtpzRkuA+wv1M9mQjv/ZUdTyh7Bog8XirYV9aut1MWhQts/MFmILccKjyLUv+REn
ZTNRYVIOVUw6umkDFKkQ0nIdu24ZrpNLzNW7VoD6tEcuYdp9OvNspfT6uwNsto/wgUW1WE5WDwgh
8nxGT2RjTOtrAT8Cjti06VmRpmtTJsc7oYn/cXr7s9vC7dBxT4sMdzWFIyE8EeZxO+0L/pPr9piY
F/+xMCsdX9gOGWNsZoxjQiJPkB3+FCKUmkXniDrfdfnCnI2zqYrvmUh1zJoYVJX5qLsiYTfKbb22
HWbvOxDQYiRAt+AdBBlGssZZPT4KPr68nM00Eosk0T9CQDSWQn5MFhpc1nN+Y7EojdG9Scsc33K3
nY7rm7o14AXnfpJ/g7iS1P+EwVPdz71Y4lbI59XHnbKycQ2UGffhwm7N8lXxlMllWK4lcJuv6IJF
tD5Jj15oOEQ/hLg89GhthuLBV15Ox2MX2ng+Cl35hoAxnBrrgxtgseHsreG4oYnVYkqQKUgrS8XQ
OUEPJV7CgkpOFXmqDmclfIZVDKnbycufzsowK5g1Ip9VfgDyUrKbfw2PfAzvD8sjI+z2amZeNFeN
FSoI6att7+Tr2l222AfJp0WFmC6AetaTFeAU0S8DhJoY9XwTPb0mHjfIH8ZkYfrt8/tDzFhFh2OT
nAIVWK7mx8pMvuHv9NSpJd4AkehGJOpoZvnH+q2tDDPdmCryye2w7PyqC2alJnBsa7TNtHUA4nk3
YHCrD35BBaNE5Odvia5i/d4zSPnUYlBK9bo8f7y/zf3sxOCHUW+pVZD2dnncSGPyyb40jPfnbkfb
hdPeD9AfnbrpQoKstO/w3zZ82bN9sY+UZH4ookGn5BLIAoBMQQGfBJFT9yalkyPc9TmCedoEu0lw
fbgUVaQgdgxeLLRqX4n9rJYJhfywcBKHtYFxYQdAjPurjt28vm+drMCOy7Mv6b33uILQine0Haah
83TbwrazsjYZHER3IxhDOtBsF+2BKz0szRJRWWOolWp8px35ADw4Zfu34rPHlO7Ravp3dBamKKsp
y0bbYelW13m7VFXKQDB5M5nrgoBTXjx7Jm7RrA5yjV6Xf4z0Q8UZHERN66nLpTujYxXqFYZnrK0Q
jJ/hsci0HpcG/xIfJcinnQEU1OtMk5oJQQbzMRWCKiAG+EpHzHO5NQtFd4UdQfUgesy3UXszEtiQ
XtqJy7vCPPZ5osVvSSHyGZyZow+HD4CZMgiyNPO+g0cro6d5Oav/3y/qJTqiwZiOZ7yWUo/ELOfs
kDQ3DKJvBBlLJAgBDfAUFUFw81XQXFeJqzinejWqQtudnLsy2oxTXerpPiVHKQI5K3QgzIlFRaG+
qIwOaOlRvm0JPgGupiC5ufDWHN5zB1AhZRFXhkbVlnSqAEpW8G5+cvRoJejIoYdk+g6qoptXVBTK
9cuwSgIbYWUgHaQJv0iUToSTeh5/UUhfqJksyxQi9Sai9Ii45UGdC55ESi/RE7h3gkysl4Z8SUxS
J6UBe6AWfN0oN/yDwtMbMw13OEEqk7VgQZMLqmetxSsXADyLHgRC3bsaBNQQ5U4mjnCNNMU23JTl
IkoZhCXbXn9kSL02OnK9UC/vgsHGdMft40tHuDJk9fKC0CdLfOgJuK3JPNDmR1rJ2BOGGU337KsW
bSuJr4x0otQtF3kcieytsSIMyPDrOXvxGSaWXACvXGFs3X/VV1JhPzforvoaNqtZ5z//F4k7qYIa
RySikxQEsWmoPGUv05ofBC7NhujrXlQ0nFSzhQP5Fjhd2vDALhDRatv9oUMa04cdruXeGdIaUSVe
v4BJBhhvKfCjjKfdjyD6KEdWHojLnuKCiZ94THWGvAY0QPi3FxILcbVW/Kq39BnpeAq2cBis4Xij
d8JVNequi4ahgrwuGVe/g4QpKeOV3nWgaDMsK6kw2o5iZCWlmDF9X26AhVuuYK5cv8MQBmSCh971
boLpdFdUj5Ow5tS/4tr75uxp6MXiFZtz1hRM0gHyS3rNCw92JV7zaOyPjKeo4R1zPOSOtTtnYi4a
aLT/rZ/E/5OwlNbvzWalKT0kqwWM1FpA87+fqSDSpPAw+UAH6LIjEVjEpgLszwxqNGBtC5qS7h5W
RyoaZvBEiOmHoJJk9JhLTvl0tBmQcwOGRmCbdR0A1rRHjpX4DGoOu7qgjWw0KnC8XjkmT96s8Nj2
mBCLhApsWjcJZzkx/d/KXxuC/VWuN7yG/mThEoVGKRkVCGEd7DfhJ9bn4o452YDLawTtVdBpWDnG
jsiyeykiC7p+tb4Hs20Ualz2l44hByUgDe7oTu2eIqQuvU3Lq55K3XLquQfflYCGPnCUaI7S5N5D
Qn08tosSp0cgNbPmaUv+ZOru3xcUNPWJz1riR6sOCGFZEPDD64mLEFeSNUEGwl4MDqKSXE1vyqB6
2+IlRl4mEv0OswgXYjjOUhc9d1x1m8gXLRjZSatUlxVRSIq9f/DgCCew5Ks8YRJOOnxI8nCcUWAH
SKT/Zyc2kUoZ1jIyIvg6iEF3cXrNjdn1PAJUupeoVahQD6aBvn/r3glFR//VwNBw3HrHSc4vaytY
gd8T4EZqlwzS+aZkRQPFqREINSIjdxVybioWvf3OBXqSA5zA8yBm9aWh36/QLlnnufXisqYIk9Pa
w6KjyUiV3uuMP/43xVE4C7yqn91ZDzN+I8rEAZQfb3BgSTJ4IWkpZqzq8qxei4KgB9j7I89g7tco
98sg38TXJ2JRscgNBQjLBj8ou7qTXQXtZUA2hxQRg9swgNkvllIIkGZ1JbMP3TVMD0zypbftiBt6
d16d4VyUB+7x1YAE2tcwRXdTlUa6RQpRc2r5x+g1W/wmSZsa/9dmn01S+muhBAS1ZhS96kgpFCJD
tRPCtBvbUASJ+p8f3C/TtvpHCA7k77Um5ZkPgGNptRtagqjfxFGfyDURqYsdkegwsWsDyZ7KZVvv
Sp5mR1cqO0hIBzMwcFK66BvS8UUSzdpN12oC4L5D+pTnMfqvndwuvVBXa0OSMGoYIUzAgqKx/M/d
4H//CT/jpL5dyjjLflR3spVnJuRWN51vZEFBBPCKw9cvAkYNcpP5EH1k0COnuHIT9VuRs/nsf7b8
p/jrqWOHy5uIOX1qDQ+KxdFAYhinAA6uzMc3vu/G+ML8bby4Veb6rL8XKzUB4j87qkhV4/SMBoeG
NcMX7oondSWRGCzjbozOiE1IAleB4S2ylrax7RI/72yYpxeYUE81VvTOlVwTqKwDiUJxJrWWAVJB
7TMlZO6D1D0zLtZ3jV9TDd/7m0I6a2ZSuRQ3po8kgjBLLKLEDGTgCP9NyDUazbltmmm2H+JnkcB5
xyCWdf0jmFOBjfszWedWRK92LqhnleBdbAEpBD0F+7xoo/5d6Y5cJSKPIIlNPjpuaXgGUV1VdAaJ
xX5XOGAz1o5tN/jbclXnFtvC3zMlFsTHLiLEAnapcWxcTRJL/kFOH9BuPXJKzeTi+dr/lsIoOZho
LrHoIZYqFfM5uZFtetIZbQzIBri6W5uamFtElAiUaZI8E9CGSgggbeyRdORXtTCP8wSmN2626BAM
vWo60y5rJ02WzoivWa04PEJjH1xK/+eYLe0Qj/Lrx4ELEDJl7q6DT4SfyQt9a0U8wK8vr0jPmoai
NPnC5xWGUWfIyWfIdrqW162t1KEE9q8HZKa3ElG1sqPlmiw6SKNxL5dZsoxkzkTP+RWLabY3IC/t
dkwTWplQJQFntvOuz62i4rPZtU6tTmwxEUtovorAltORpepKckEJyBh0BV84572H4EB51TyMwyZo
H795KSSd1LTccOFNgClHhroUFtM6wFmy862uLtx3E1IF5aIT8cnitt1EzLInHduiPqch/F6kwA5B
7+cb9OotXQ69ZBJOjFX4WnWJCErixCGt7zDb8V6C7YRjmAMy+eUuBYS8NV7D+Lws2c9/5B5nu2R2
7hAX8EEA0U7ELPEm7Z5Pa3KPmrAsv+8lhPHjWjgSYdIaue6P7HK9eGLLhOMQCZGBXjXyH+mq8f8c
2Lyr6eBiUXdlsPW1npRtnysxD7C9tzuq0dSGysiux1dY6t9Sa80wuR6kKLgjOyFRgJb4ki2IpVnE
q5DRHH47oyKA9gmAyc/dU8eilzSLw9DAMHCOIuSK7infxhWgb5mLadYVlJmkDRFLWm11jVSNPtsQ
oeSCJ+TliNPAwdEe5LYprDcH2zxkxU08wrS5nefaExO13AQcTsyArWfdoCE+plC47xKI0iKOfWEj
E1ib3TsMSlWYl7HSIZzzx2ifOnuUK5OIP0cj0r16rdE8f0jvO8pqPmyQGBzuPQmxIFgORHXc++YA
dG7LJ32JydAWtyuPiwsSSNi0Gwynkt+VJVeB7zs0zChquMEATtvhafn+SD9kBsPnTbzMDMZPYMoU
LyylifkFCPik/bvq7S3qOIPQ3ci2MrypIm86rj8zrNTCmx/Wb+HIDgoGfE/tKtuQskGhaJM1RSvf
52g5hZ2rkhd0goZPbJnqzYi+SP82YkuECoat9jY/OH62atOMnk0tBPC5As7mxmUMlLwTfHVA5UBb
s0w/7g53ZbkQ+sURFHvYUnvL+pKeKfbtzZXM0JdHn4j9uzyl4rd1d6l+wl3IPNb4Ne3zn2sBKtUs
HCN+y/ZiVUdm5AKOdQI5eM7qPrLIMnRdbyGu1TMmFTqzd+4bwXnsWjdqz6g2iZUD9Vp+WfTVw7f1
2xC+J89Y57+wGpfvrkUH3k+3iavKnWY433HbN/K+5Esu6FlLaI7HU70MG2yNAJ9flwV7ezPb2f7S
KRZzU8WSkvK1mRyRRC4k+m6tiGqMYeroCK1+SLFh9zkQoutYXkHfbai81CBpmwQsd2IxNhiVNncZ
f+B96Mda+wTb+ypRXgdvqqE+Cj7simedow9Zmw8/taMBOss8kFxjHBr6BDA2rwXLKv/SB71PvjA6
XXRVk/vfbzKt+MAhyYZCbGkXSBYKryhO7WV6WFAykXvaCW04lMe8JmQ+BZ+cWMBqNmBXHuQK9gqT
Z97LzPuLrScZHGot3JdCTX8mJFnUe5dTN8KQZjffNxFBLZNM6hcnp8SFLlgGFejBI1BIi362yj3E
uJaOul9B1Ehavxk/1ZRW4eQ8+MYyIj8TiN2SlI5tj5Hs3I1l7czNvHB4Z+G90KeBR9Olux1DeuE6
S3HQqPVwcB7d8zGVKFBTFnFCare5J45sB/jUpOaHExGShxP3aaehuK/YVTmgraVY6vrXrgC87Muy
T+bs/Nen9nYW+5UtjdWCFHDx/KBgR/l8JMXkaiNsdrrTbGWR3KilkylniELkZdslkk6vMwhkyt/C
Ux9sv4mfDdUs//c14SVsRenvRSRK0vtQR91gHxRJy+Q3rbFpioL1ld9B1/eP5+fJfSBKX+K64Jr1
WdqFEwUnZpjGeUmtnpsyRTp6SSE6Wbnc9QCiq96ahSgmcXnAzd6KAi/VJpJFgaHhBmqIk6uYiqmQ
fv9nQFf6XgsauJu0JyIch5wEIzJYCY97ZKr9b4aQwaoxwj5Gz/GmlnuCXjMIHV1U5f2iLTeKguZ5
Wt95UjMoBslJH3g1XAgH8dZT62g93PFgE+Oxh4deUszjdUON/8Fl0oV8v0nsYVbj26PuhIvtEYbw
XnZc9NginIg0BRcSCDorPuEjZl2yLMjY+Ck8XFAf4O9xmOWtSCmEXwWhFYt8dokqwd8tGJiDZNGf
fmXDxLblPhXzyH5uPwrbfaINyJZuDhEI24nAN09V0GckC8xggwa5HbTrmb42P95sn6zvP/4ZwzLe
691M1C11pG+ZsHvyuDt3D6+FNkJjnQ8Fjb1rZ8CoslgoMzTMOtlI1Y1b98rz5fawBJreLc9L+fJn
AOogvO9Nmyycdq9hAmnzwyWio4CjT6VjAJ/bKU80uEE/1r+LfWLtpq0zTMRjZurOMs0MQh/gi6YE
zgrg5rDza7E3wRTcA731qTpJVGT1g79+Y0wAHzawp6laD+90IZjQ3a0ZgnYbXGaKz8Fbmaju83qS
ydP23YZ1KyflOGE28UoBpDJ8uAF/oSoIUaVt5hZAEPLU8SEh6YuPbnJQs5Sr/cmBh+Tl2iqSZ8PJ
3ceRaCixs5vaD50bNjwEAs8lasruFRKnTozjxVq2CEC8rKLiMueYK43BcociDPiZCifjx2FUqK0z
dPlvoHFlGD8NDNYbt1QJGZt6zIRrAt7yiiPPH0myOLanXQVmsKukrM3uzzpcnzxXx5k9PACGhLng
Sce8O3Ys8ITVqssTpOZ7qrcK7K2mmtznAMmdns2wPsx9+GITrRbZChNiWiU9nuKxnDB+cdFKUFWx
/vlo37arKefOMlYizGVMzaYMBtbT8uoDhbhQ8BBCJF48qLd2pojdG8hhqL1sfNzs4AMtI+yQmm9p
3ZFIgKjOtHa4KVKbDauZOM0sBdhiWe5r6PqRa7g3btmmwrgajh2Pn4+BAnZr8E35U9qp4jphR56X
vVeOlEI50epJ9QgMeQNxaYBncReB6a1eixor+3mam6yVKzk6G7NNAL8b1q2X0XIEebUx924Avt2V
pX9VnzeIoP4At398QC6Z4gWebKYUQisvrHQUJrhAji9iI+JptUNt0gbiWYJTCp9sZVxGhQ1bUImT
pCraDjJHqvU01TLlMx9PGHb73GEh/R0b42Lpr6xPIyjjUIqFI3TpIDjRZoD8pH5QShziy0l30T6N
QVw1Z3gowm7Mcj4r1RzU3rnFZfS59Cn3XcqlcQtM5GovUFtNXmZxbKs860IxXgDITVV4T27dH2Cs
haSe+9DGsO15C7XZWVseqixOGv8BxR0+AQ8WDy+dXPcwVXqPfRDH4M63zPfz9aV9bwiME7M45l1J
bhzCn7l/DDtl2BV+1uY3yWuagXNqG50J6GzvBBrLMoZTtgM7jXP3Ym22/Rk+5GjaYvJZonccLQbB
2V1gMYqKg90dcmiNGF5REAn+gXIp5tBm1aidUD372W1h+/KsryDl1Pq7MkE62OBwf0xiIHzdAhJ4
YK1NhWoXgOH2rM4wlGLJlmiZv1Kx6MjdDN1bYp+ZbHkrMitZlHfylComa5jafLtc5M8WoxGxk+wJ
mE9P50etNKaDyXy8yQMkilnrug4lxb5BpnC9K4mdPRApeoIurYxKcyGB+D36gnaAfH2TWELkzl/d
WeZeOxF0gZOzs+KbzA8KlnB2tKYJgPgumxiz0DiWz6nXa3DyTOzP4vQjHiHh9RZXJZ58+wToDO8o
PnxwDfqKFsUCkBzKegDHO2OCzZu84CcmhWc1bGCbv0ilYz9QTjuUCZ0ikNhZnHiJ3RsTWtiPbIrL
QueqmDiCNB2la6YCSvgv5Xpv1+Qywc7FppXNOTPptSbNsg7pCzssf1vJBltjqIsPj0lzDq3Px8vo
Mt7apqo+GqKswZ8hdPT2DDLzyZAlSBhTa7mPJQ3UJE7Lo/l8VWCBnuqTaeIZ0ZLRBbTtwU8F4AYi
NbeuvWRyITaFDvKP2tDWZhYIHkd28H+4oEot4HMET0VvrbNvQmqDJoNz/upSsvHbEShppK7okyb4
evoLzGH+MfvvXHAoSYnrTjsxHfy2xqhdHeIIBGWEnAPRhi+cgSssEmqW1xXDqkXpovpX0lC2kpgE
CNJhorZ6IfB/CYYJcChPZPTz6BnE0LW4xW9/7VelQQpMAROQUvx6SmzwVYQOJjKwrEr81raxte9r
slWaNrRO3wwx/m/eaLNq75ofB90wbRtXKAjiJMuTyLjM+hZvmF6on8vFUC2UufdgiE4mk8r8Q7ap
na4s75KnWzHs+3lMFsC7BqDmo1nWO8k+MCQzaMGa6u694P1gcVUqIgbjfQvEOFAHNU50/L/Mb2Oa
Uq5uG+u3w8qECYP254EG3x3+ACBB6rm/WRd9PZ6PWm4nVjHBHysfryPVbc8N+EtcVB62eGIrQN/y
MHC31+eFwJSwx+o80qiY6R2uK0CBCL+FbevsTeR+Saw7aUgrfSSe4n04ECqCUfkMGXjufnSvQ8h8
haxQ2BIZ4JIZMVsXiIY0DpdaQv6fiPtvxMY7etUkpdy6zntHZJonZKiRZ0pjrHEXQAzOHEOhZjHU
SXgDXS/sWbZWQ8vK7zCDIfbyP6OKQ39gk0jmPbnBjTRWu591FLhBd3w6206lChTqz9Kub0HubKUI
HN95C84WYZojzJtMxu5wQn6jx+XCsMFLjyk6EREs+3LD4GPEmor0CvWL+12HOglLHKBWCiwZ0P6G
QCM2HPGfyWjvRMFUdSpA85GBk7DIorY67nVeOMeJrG/15R3b4Xicm4S/8v5KmP+AHrtvmZpAz6Sr
ryqWpimkV76cMxs8b/o9dVBUF1iaJ2JX9kOCOxbiFMrAM7UjqYaPW6E/NbGQSBGP/RKXCcK/zKAw
T4c95MyEbwNaHMCpSTI4/Kzp9FffgE1BCUxEEEfsPXtfCjHzWUSehvjXfEQn22b/tgRCDdJocBOP
0/41im+7GzTqTnhNzZv6HLRopELh6FtQS0H/mhSexoZl5hNezUepUBFcT9TdAf2UU2JHsqykEGGs
11Cx+0FlqgnW6zP6YBt7WOOguuaj3PYxWLmf/dz7aK2KwVGiCTlTTC0CDZ5SktNASC7QOmuqaXp3
atqzat0Z/EqNHLbcgEhxa8JI0wYI5aLoXuNaa5INknk8fXmcim7dJeMwiMCGihKlE/HMeEkiX7Ij
BgKFz6+nic6UgtC7U7ey724VkXOJi6cAIPleq+QGymOuBb/CfVGy4sUuntncTHcfoasZ4MG0b78Z
8LHwokkN0FLfGBnQm6Ivsk8Z1OBEdRZmpSzEntITfia8d22c9NPADcYeUlBi2mYKsNYA83wurbKm
VAQHrpFu7r50sGoAN45bX6mgmXB48N0NexgRLWFERKx1Klc+jg8NNLmyecE9m/hdvuDD8/ezZSXG
Xqzbz55guqtgGQTvdXUL9gK/NgfIXiF6CiibbCjTpyOS9m2WYRQZ4faoPPy4zIIU6Te4RGO9uFEu
h/P/vPTAAP8YRGtWoKJou60xVSdyhZx/5FF0FVb9BhHCGHJVONg0RY1q38vwrs+nqoGoaWHa18Ng
M6tF8PCS2wcTQ7fcJfTc4nueQhhpKtKwhbuc5AUaLSysyxZrOm3WP+UIx6y7jZBmxjpcsRvTW3ym
FFFkRN2hVh4ZUuXNQNIJL+XK78nDkv7zBRr3DCHmChhMQIXNCnLdZv+Hu1T7fzVy+hfwDSm2dSCT
5h2HBlr7GsX4TO7tvXo9H3b8NMOUsJ1LX6/TPGG0VNQ0SwgHezxEuSyehfSpSu7Zf9/xdKz+ttF0
pVi82rtMYc2Xbz5Y099LoQY3EMkKPdnfG/mc/FGQajFY2/OilVkhOl7/tSHlu1VMkMfq2OTkXNXG
SApTB8a6c9+do+CXMtvVmx0RercnlVpwtiq+phuG8P4aOf/whYpd67UARG1ZemE3GsFht2OyRFD4
FKRZ20DNbfDY/m4YYRiWqBq7FN50XXnQR3AiP2uwOw4oYHoK+egGkDdhkf+MWeTIgXqLggHC3Lee
Xjq4ZtswLYNMQaEV4i3w65Pws/kvLD0btfg0lKb0L3j179naa1X/Tr2BJbukfnM+v0WrYO3IhInG
zmoEfoObr6Y6TlGJasNUVOo0EXi8KrvK0XdG+s23othiwCAWQv6Jjqnkl2QEsr0cyZe/DXf6+0FD
qQJfIX5QBC3VwLNFdECakluGm8pFMVyyGKtmFVqAcFku0dGmRPrqUnnUqGx6rQN2egqbi15Vzzb9
uoIlDVU/u9MWzxT63NV5Ol65dW7QPwh/ghNgCHnYCcrF7Ra5ThHl76ZdFoXmXtAzdT9bpQHn1S8U
CiFCaW+OfzNBlccluBQ5WHr/Mg5N/37U781IuZz6fb61FDWxT+f9KgANEWSdEu4tbo7s2Q1xOrp7
0YaG/diMIYZEAij4T+tM8fz5b/c++m2B6tlMa5xOjWLHhiSksFcbhjqbwS8fv7yKzQihF2llc8ON
R4FfoMurM8Wv6/ldyALrahvP52Qw94sjUlVD3g84syKg+sSrbEdAIJcN6pWb8Fy8SyL+SaasI6+G
Xb0AdDb4WT79NVM7F9x1qk9wn3FG4Y+fke38Pvgwuc9zmMQsXGL/57nAQ1bp02JwThBjgxfA+ctp
+kwfiag6aUzRfucTKcdAV746XssxD6v1ZlW+s896SBa0ekJKHk4fGP5+UcIjnj6lUtpDzhBf6wzX
LQhvsezt7TiY/H2I6n2Ndyq1iN0NbT/Uf5seXDb23Ixp8LXepgbn9nnH2oYJn/d283tUwXoO7cdV
G/ao3ByAGYm+A7AAAdG3/TDsCIS8nzQ7Pv1dxS8CPPxnFvxdQAAeHhepRiPJcgeg31Oy2GTAnFkP
CIt0bwCkqOAvbWQoz//cLlLFxW5+m0/0AUP/H7cDiBI2cTatrKps9ffRleuYYE3mJLcSbDoJD338
nCj6pnQ4X9vZh5lWsSSwJbDYekp03iEhXNkRLDhlFtj+ziVF9tgl6jUF3JsIQrq/gxeFLkI9+MY5
Zp7NBrQ/vVOHov17vUOj+4SxzbQJAwrgNe/UdpjcqHj+ZaloIrMCqlhJt9tg5hWflb2MIAC5gsAf
hK2sMwnGNK99giysAb9qD4Q7Gfjq/6NhsPDPUQG+p8rwE0ZofpLucXr2aDGjWPWARsCcEgddR2XW
52wEKTGmeXGAjCeT/GZaS644UjaKAljiuSzfHA+PNkDIcdEcGb0nBNRXWqxbgEitBkd6wXgFGS1e
0R/PH5m0QR6hRbSSZeJbysQsUOBSSPeCidiQSgB6vcOA7W/IvNDQiyZCz6Edt9n9nTc0lrn4RWfh
ww5QNskSehsLBdEkUuRc1sZvR+uIqTZ6l2XMbzkZV9tMp7bO7hn+s+c748BL94hIaqnwMkqAy5Ee
kSmRCESud9olmDLszGXrsT3zuf78nfKrUeXmFgmcZqJlA1W+GK6UDqN+5wxsnB6y6aKR0kyWP7Ud
6e5M90CYMVja1nowndNKnmaa+xJ5nu9XBKYxMLBoyDyIDRjZB6FL7KjJCH7fnT8grRo2QHFlKXF7
paSQdWXZUnxTz35y31TWeHzipuL9r2/YKBpO6Fu8Kdskq/5uKLw98wOUE8p0U1nLesaiC816uf0Y
Rj+dqrX0tdir26kMpUMTN5CIZnhQE2RRwc8iPyp7ocqvGWUPSKGWD7IxZMJ5sa8zucopAvzNb/1S
YRFyei89DMovVf4OO03Xnb7qa+5P0juMIs40VPU1hgm5bLM2iX0FJZvhKRFPppk6LV6/vbjsyQPv
G50uRHgKRwijTJ3sPTA+C1yBeahsfpuoBftUcH0RtK6OFGiUCTPIgZ6M+AStLyUqqoVntOsvVs3x
Ya051Ts4z3Swoqgao7d18Tw+BjGYPf3zikocihgw3zgV/kJNrQRdsrOA48yHAySlsrv+ku74V9Wt
H7OsuChBAdYhEkhAsoXxfPV0/ABXbS7/8HJIlDOacKOPCi8QKQYLJXdx3Q7NBI8xavWfwBUogY/i
P48Voic5l5B7WViXit3UXG31QoXVvaw11b4LV0X9ua4F9cGclbEV2rRLu1e6Hy2qFdJextkMeQ7O
drdtLqWTTQmbLr7pEfMCtWMoYFCbiH0LO2yR5nbFT7Jh+DRkmQ7uUzvAS66kK3I4uxJdVUiXyyTJ
/o9DrNDE8LIuXqf/NkY0OFrpfARq7ogZG9qD1J/E0exkzFmF0/syRDeC7JGQ3wsoQovi2JCtCy3R
tD7XFJCXyJACZhKL1ry0Y/K6Pqh9AJneMVbeZ7d3o4gzHq2BCSTxZW4i28Pjn/iF9vogj2U4oRi+
eppnkJW0HoOVVOzvw3SFZK5j36tINO04ig0vBucW6Ip4Tp+vE+KnEJJO8TkwMRc8X0M6dH6Tw6mu
TbI543Kw50kU2pSz++Ln32cAvvS7T4MPr3oJITkjeV9lOhRWsEkPmg2Jy9ipe3nvyzI04lIIBp0v
ri5+J/2ZphG0efDtUcOSvWhFlQPXpMqaVJNEOdZJs2jHEp8W7juKAfHlIehR63CK96VMkLVGFcT3
jMF+g+jpeG7jMWGUJGhtDPwi7IE9oKdmrA1tc3fGblk9qvPpZvYgbeIOXJJAqfTTlc0s9lEmwVl9
UV/MYOXQB5Pnwq30hJjBLk1yujHtmNVZKQQgDN5xFhQZDr5XXnRCtAyOfI8q2s2mjpBSyEHTWfw5
Kmie0Px6NCOxrllJ3W0gp/aFgyERVYXpe3Mpk449r8dXDCZFcgCCQL/w41dbtCJpTWlbr3itDKFf
a9/SF0gwKFD+SZkOo6FS5UhlQPSt8Bq+1NI+HBSRQKphcXF5xBP+QuO5Y/9k+jKIbGtor+h2dMCZ
cNgDOfc0dYJhrn/IYMHfvNpBBgHXgC4muB7nZZUmPv95KOTb1xubDF0MwsG+kyx0QEcxkb5Ku5vI
Mgf1pnPP6RsGBEB0jWnfL3BDQchUWtyWdd/sReXbIagZJada1F7XEiaiiosPNlgyaVwbsxQRngjQ
Hddck7tstLTnOw6/7vl/+glALmyiFdBiEXXiZt0Cl/RqYFD/mTDfpiuwrarGtrraodR2gPG0Z963
90Ngvi3wDweS6dmd33CXlGdTnqPf/iV0cs2MlH2SXFsZPP2rOo7qOmQAc3Of7lQfXzAlv3Zo8+JB
/DOPdAtxYOYdekRWCFsgm6okfW3HzkTp0m7b3XiH7Xs5MIiA2JFNzrlwoRctWE/zZF2H8g6uM+r6
W7xGKMWnLy4Bk4tuABq1iRxhXOGF4cgbjrFg5P0v6Y46iAqg82LmpofKxGCWgIak8F9RDxkjKb/b
KP7sjsupoGOAGRBYilYOZTBZM/sZm0q3dHSyGy0jSpvCt0O1nt0xnsJNe+zd/EhahuMlcrJfltOL
qI6EiJ7IGqTQC6S2K/jryZTa21I29OFPk9cbXjv3wivvshVnm5yGgAjHmgvhWT42ZRGU6bO8mHlA
x51KRJtaH9aVKKStf2ivDKls0NmvEZc7LNQX4Qq4JlGxfVnesLU9HTUoCP+OyPUXhD6QpBaw+SVe
N6MMYd7dTdw3tZXV0kz4SGiFCP2JC9CjFS2n6/y9MnqWqeJANSHEHrzG3PsSX2sR19df1zQ48r1F
DFh2RWJ6LSbanRAvLSd1tUJCnCYHEh/dznSrgh22mQ1EqHEPV3dv1NoNkFNPH1KB6t0TDR9RJlqn
lyuDxdiYCZUND8324o+YoyJmoAPJc2s47hgjGjZcCF1lse+w+iGIXCssN32IX6wsPgHiITjcgkw6
+dJzlldIptM3mBLf0mT2kRzfkSgXkewDoHXXxUUtBtsnz9JjjFf/N6oFss8iak9k1IXmsTm3B9Jd
qznu3Wa6ROStmHIlW0FjQO6O0d6f3my0tL3UCVQvDVtK2nG/Hxw5B2PBBmDKlKVgHiVrTlStIEMw
/9DTPUGAH/S49U829wQsS6ZDmR3isA1+QdzlivRAmbAvOWIO0rXRwg8/7hiIF14j6LRXyiFBrsG7
nzRI1U+kWvEwDTAsFTZRweObeXkDBwastZ9bTQbc+V9UonDxjwQWdtz6UJNOiLHuKWgzIFU4eIuP
SBcGhNxFr0MpJUnwUzyeAVTOw3xAxce8b2hLbmQgoE0TlTxY5+677Jn89nUNH5uJTw4dhL2zb47I
DWIfuN7A5QpfsgNLs1SPsjS2HuCwC16J3R8DnnFMNkHDASYs2upX8WS0oeV/bVX0wOzr0rPWI7Cs
CWl6yXJmi9twSAbFm7qA1ezC/G+kazVqx8vV+Wc1A5eLoid8OB+sVfogqgl6jum29yA2T4CHJkbD
Y+TusEqMRbZqH74PLTfPCpeYqeyJBuKTEPsM9SJytT5wdipF3HnPLHtUlYU+9on0yTWB5FsOaHhB
1FPKgTSabvpnfggyTGwt5lXnf1vUKuVKOZbbS3NahDif66B2ydbhRi4m78NiaUwd/y8V/WqJR/lw
sM07ViO+Hib5dAyjOCMIFIy6cRDc3NEMfvscXaF2SaYFt3OKs0TaznP79hVYX8Z4+YCXPYJI6hxf
FpLcwOe6RmP4nDb9rVRx2Ow0Y4gQiuDA1Q5Jhw0/BJA1nvenQlxiaxR2InhhIN3K0va/dUi8ducn
y0M/5hPJnXEV6dnyi/o65KDilJWthXlPCsBBxU6Njt2rZ8jHP8wxZMEqhBa47NVgRnyPa7VQMfvk
s0gaIUIKylK8Zy2X2gEgdVWdg5E46Pab5b6wkMl8B8asxgSO19P+APG+STyFmMfm3WpQF82BPmOJ
d7mitgRuxpBeFHWl8a69mSe/oE373Y69scxqTaVEHvH07TP+b6FUIg1hTicgEFcdF+I6ZBhHJM3W
tLbMaL5Be5+R3FgyvOTr7atkYp6dWn5vIYsxV9mfVHAr5pkFgpKm8oPsmEvSx9jQg9OSnvSFvmp9
vyefB4MAXaMLwbuly21wmL/WppIQ6+x2Q5kJKciaxREYpwR+CNglnOSBk0Ogntsmmkrs6EA/3vJa
ZJXIaVYFxJdXChIRvkEHQYFFYj0BqFBrMcsz0mrDRFcrlzBW8wIjncj4mDT1uZPxX6Uw/75yOSQq
Pi973AqfXbw6MBW+0TOtzN2mzjt/qTDWp5qFfpl5eRwwqnIQKCBCbx1U6atv8SjDCjI5sNnWfds5
Qj7h17XvHlPNEUQaFQ+KJmBVCiF+CZCrhcElKD6rCyG1IuRs/rCyx4mLBrJPZu8otHxrAUMZ9wxC
JqGvlCnRmFG0eMXWSVDDx82J0bBkzZTmWk18MzonPQgzCruHN0l4cO0RzvPId9ZT94lwsC47jzUn
KSfcdOeblPslJTQNmxqPSqCU5fzwVW0kqcEo263OLjDc20RHvMj6iO8uNS5y48/KKZSQPTFpLSZS
CSkE3lAfSFjm16ZgooZARZ8jA62HQxvWSkPujrNWC2cLlA9AeMk1nsy3BvmJRZsIfq9dv7P67eeW
o8E11ZESDM5rIBGBhVPboPvoI2tbGje/kKakMkOf6o4ht3IujLtut9gzLdIEDzpHV/BLt26qNpAg
FH49ubezN4NwvZrk3xOLUMSFpqUkS9qNST4n44XQ0rW0dvIkewq0v1WDvId9TP+eeJYqoZQd34eR
YgcwPDuX5KBxx+U2LDSRrlBhUfVfswXNu05HQ/+LO/ued3/hmptso242274sRGBXk9PvXqTe8Jtw
B3udgL4/J/IiR6xx9PD+iDsQ6y0voJHe1z2Lz3tSO3a/z9ebeNiLnCgelesfmXp50fDwvEn9Hsyb
GDT8ZnIj9CMPyTcfKdfMMGtCFcSnPACGQ6bgJILxaxbQgGOS63qz9+8w/qp9sYkSd2b/9EBnTygr
mFge0xmxpoucIwVJFV/BuGaZjLOmKJ/GD9+SJzByeDKhgmEI2tsrYD3AOFflN+F0zGAbA3JS2TfT
BTYT7+Dy5WmpitCnmTix1zXXVQx1E2PFZRm/+iyBB6lB0oqLCQi2hRSTVa5ba6yxxIrKksUskTGZ
WNEyr9Sf4otm/o+MpAUIbRSQ8yRnLWSTVgcFLvvCkHwlwgn8c+YTux3hMODns1+Qt1wiEv1vnwvA
YEjgIuvpSEVfR8LM+6Gcj6W2QUdYeeTRcuQnS5KriUDYVB1TrVZ+Q/ajP/dD+bTYZwHVnUs+6l5d
fy2WNKTz0x/mADf4lJouh3bVgska7ooV7tactWnsNcOXixtA7WzqXcVWmIEO9Qkrnmz3bzldoSKu
avmJ49T5eTXe/o0DfjQ9Ib3jZJJYuKuOuoNz/j951xvLIg26KGP7SLXkYYVVcmT1vmaPFTwTPr77
EoliI7pabBBoI0lz+75ydN4q/PQyjNjMBRRGFSFWddjbwcJVJFQZryAuWv7M8MWV0BMPg0qiMIUa
AKXTmjWeV49fd3OcGSZRmAPp/oRcHVqcNAYOg/hf5F8CFxDhv5EMEB8FOM2z1HwzuxuYbaw1Af9u
ZnhT9kgiFkNBLZnV8pYcIC+QwcqSuwFiUNCH2BQgh2PWaL2WNwbgi4eInm2wEsLmh4QmlWMHuRqE
+CRhHsA/5+BI9asE73rbaGbCZ3+dMTjKPV0BajsYaIJV2kr+finmjR9dEQsJhjJMebn7bTRjXQp9
jGpaYj0AuQ/1kgRSZx1OgD7yxGZGP5eqU/MnMqd5QzBIEeCRfOsE3KaD1rgCRw5EGrS3Oa9odkvZ
hwoWb1bfqJ57GvxmzXrexJ1kPbVo2ju5tc2MYyiQ6XFNOKsQqrwUs3iB3tomIuijy5ybGXzU9pX+
7KDxCs+I42BVv91J15HUJq6aL26RR7ZlslbklyZu2r3AIzRN1KrMbLHDoNpw+l5sdfxVnKtGMvYt
mvjqBEA7kQ+CViwcJg7zLHsoZSCYPKVUfQwej2fzvwgXs/e/puWiA4o/l9JcDWMkP+tngDIN/bay
Fac3gBxomjzetsq2vyWfTC+f5rkHN79qK1bcYJJavJ72uOIogXkujGnaam77Sy5QeHfd0B/Wv5w6
d66a0Me7BK8Wu20/KAvR2ADtxh+A3IlHJGhfHOCZS+TDstpyQ0u5r4yt5Xyzxa7wSndbFYzGwUU/
B3Q5C5nnDZH88ycUwFCu4AFEVwBFLrmZ5GGlUNtvnNA8js67sNdYpBJTev61Fd8jgNY8cMHJMuTi
4YtuzNdo+tD4ianHqoEG80UvRXR0tsRexeLn3CBTZ58Op2KMQ6iWqDUMMQf/rf16ovI7AAlW3jvm
mECO3iQUVCoESC00HUjBeD9uxDogQc/Q8ttyS2raZHs6SYVCKt4VcNmbe4ye04LoR1cnlhb60qNU
jrUmS0YJPSImFCVqRvtWhhOmWEAZpOiwGaMXJNvAspXbMbyhsgWsWjahstPllM9aHq1mP1gy2nwi
Hnu7SIiXjGnsWN4+vWEMsBudfkuD90/WY0V4SSAT1Sy1P7ReFzcqYZSLakw77B1WA2nutbT4eFSb
M2KkP7n0fbGAyDFL22Cob0VDciGpqSZpdFfLqpOkw/iVeNd+Jblz/0w83DPVcorIQ2ZYoC7YZayB
L0wYb+4H0N6Wk/AMdoXsvXz2olLBD2Fc+QL13P9j7LD5h706YCcddPsRk3KPLPdjwYG9vBCMXg7C
My6Gyc3BDFmHU0oolRF7fMtZZdDTU9lDqOuL8EmMk/Xs/sk4QJbpjky5+sklkHlAJW9SJcb6ghmE
kUmEEti0SksKlAZDB3lomMVbcawD2BvRMZ2/ghCQkMKmpKPDiKckBKyGfrkCBKJv5TUbZ7z9rW5N
nMmMDZFMmSo2lT5iv1JQJJnfGbIkXHFotqOLxSZFU3f/1So5ADX93OX+qCTob1PHDqps/OXfZ3Rd
/C2W7Dov538FKRQ2k2qb5QneQpun26rjnxu28Si4uEOeC4T53xhYSwMEdxOgu23bciPoDfGdb/m1
9zan4caSUSZYYRok8k8GphjejgsdbyEFWVM1C0GahFjFF2GNUAQYmlTat/sBBen7BOB44ujxq1Xa
jEPRWFnLIyQtWaRr+qogSk+tCuCv02Y8mJAnrbtZbhjUk5xvHLM/1QRyCCT+OU224BsA3yzbx6L3
zZ527lNiwpHID9gtJMbiablXscUqJR5ufJKZa/geF34y+clkXoA0T3wqahkGAFgr0544wTtn/XQC
NUByix8MeUh+liKGoEBkbqOEf3kkJ/zZztV+2/mOQrwNyGdZFuPxkBrZ68BiA2nAWKcU7uBAMmcv
y/GICtspO9AIm80v/dHnH59u42S5WieTlw6bzPnymOQ3QjW15jCzIihEdU+YZY8bPgA3x0viCkLe
H6RZwIEaRy7BWvcIZCrqPGKDjg4CXVQlM7zST1sYE2blhCGrirGXrg7WBkUfC1G0ZxoTySACF8+4
rn0uX5icXdy1cfygsX5tHjKYo3TqT5CakcJbtdSEkSjkCoqICz3nWcnZ2XY2DmT4zRa8//8OTq9U
BQN310oBWFd/bTuPzzHBzQGGJwb2GBJYVa5jUa1atGctf/qLO3OiOMf0Ryeci9fYSc+Q0511IPNT
mXwSFbVt3OvyhpZSYuQ8gtdZ4juuXhoSQLw54/cPUYE6l/NdB816xEqpC+MBEIrv2WLFbjHVNlxW
QWiEe+BnWO5kYcrA6q5qaKdD3eCdfF92pB8Yy13s9F7gCSsdUaIEm2rucfk9y4GI9IEJ2lV5fWj1
bxGnNLEBPUSQ6hEm9MUifOVebiwXasQClfYAwR2y2JluKDaOhbZbJ7qFGn1KcJG6oSIdR/M8ayii
WpcSByw7vR9NR56f7/noQC1zcA5TB3owOE+MPpzPRtMvhaArfPL4ZWq6ifUGiY8E9CCvuh3Uwnd5
/TJXu1aUZ7Rq8wyQnMPrIY5l8RXm5n+VDzJ8UiYHyxVRVkPHJLaJHY2GCnVMb8TqmiOPRMYliQE7
egG5qUxohMLRxQWjlr3tZKDfbzght1g0cvXezf7u7UjMuk5qrmsYLAm4Tb7wZix/utS0VTNIi6ep
K9rqdcdB1+sMt15YnyrNBFG18OMAZxNXx9v2cydvWHAta5/Br0jTTHQi1YR9p2swtYxubPeg59b4
G8HYPNxJIkUVnFIbAf19RqyRGOBf4lWW/FZFY9FA0oJ8BsC+N6NDUnswEZ9RzQ+8mH0XIA2vblfT
om+qzsLaIl6C5i5QAgB/18GM3SILCM2QvVjK5GKm+4y1i8zqUSZGaPc2NRHhSR4OwnN72fGWLXOW
fGPEZvG4I6CjvmLsaT1kAi+kGESsZ3dmK2pLpms1AoVDKL5uZ+epjhQgai6qOSWFubcCtPTST699
0SXxPKOHTVKeaISOdedVc8URe+Fjxr6/lPvuCBgWhv01mFKMOrSqOTpie+R2A6NhHKcKs4L7iHA2
fbOtcht6ipWX81PJJuLWd3ZAefZ+nsIXuYD8wTiFst+3+KNsxUpRx9Fg/8LMkVkHPuf/mcaDL0Qx
Jw7UbPGsSjQ4rkM1kGSem9+YbcJev4O/cmu29Dz72tMsjYufs+PGdUKeLXdzio1A29MvfUpsFcJS
M9vHba8/oe2SnIQgwGWLXwzWydsH8XhiLr4kw4YBZKcalPmDeVozOS4Aii5lFlo5c2xBOJWItC5K
w7Cc/OWr1SL84+2vYt7TEnDIbZcJV48Mc+18o1hP+k/+8BbrO34ZHbOSuQy6B3V0oxOmRBKdP0TQ
TSBzlWNcv6GLU1CK2LPSSOAf3fhN18bZhDKcsfmghLVd+AVUi22HnGiv/8xkipz2XpjZWQ2CqkUw
dP+MQE8/OVdgLjXEIukSTyElwn6a8k3ApsDfVLGnmeLkDmeI325J+K3zXkoA9AWXbwGbAdFerLjA
CWxhYcwQ144BtVhm0m43Y1pu2D4vP/plKlDOQaRlQ1iNsBNCN2TxfAsHGjT9w8BKdMebp5rBHZmk
41ayJ0udjZZRgWvaTu782GR+l7h6CSQjVl+hOQbyV8Yg9c/cFH0qYhIg3e8O8gj0teGRX9UjIs9L
GEoR6T0AGKdPkLvpX28zuB3hggutuBQOLxNS7QU68e6wH7TI0Kz3Omm/uMFSk0GfS/0FM4OFVezK
S8zTSCLI/pQW67DTMReOMuRXYsxYiXHBAoV+JkVgQj/jbXwVG10iwfb/oaerA3ySsOQ+F1eU80EH
mvlyLIKnRdwNCH27a4G2oJin9IoOpY+yt4KSKbKUJWfFTlMH38LT4nyzXrVPtZwVMIvrmwf1SRMY
ENaeG1vtcONyUCNrd6tAw7jeqrMZrCWMFuAzePNseiqoqkV6K2gs/TMDdOzn7Q5SG8pgkwt5fNrl
FOEKJG8Gkq+Eb73UQTv36b7m1dbNVEmRUVcV8m4A65PZ8aMcTufD7iiT6GlDVL6HW3TEeovjJB0U
Yz/6k3Ebp2IUICLodwN1y4lK5HZswI60meOW+0T3T0qK3xwSMaQJdVjGuWQWxdwKQBj078cp8Gpf
7hG+Om/dtZsvFAmUnZsZPfF+8FKPmsAc+Pzf/BS4HrGafk0eiY1DpF1NtBGIb/Yl2Yy7Ni4ss7Sq
xtZcTE8XWDby6MpoAl/qAWjpetd0QLETCYHVwKfs6PEgmHrrg1g86+VNo3Wr7nt/+Z5/sppIAoDN
Pviin+gfAqigDx/DaTnoRysRFoJQXjO5iV/DEz2GrlKa8qHIt2deiqFa6ULIAeXA3z8JnkCjUXQ1
q5vXBUDoX+6sF/DvPIPboGGseZFJ4DcmIAjQJdxtXCShxKvoOgR9haHGtkJkmHyQtMO7NlhTRY3q
ejmEhJhOZk40vw8Mq9gA35Ypvrw+zNrZCkBmiAhNo1oXhHqY10hslnuxHGLva6LfBNF25zrAYdjs
OE2/K7y6im6rQU9rk77QNpnzqaj1C0WwKE+QYAuRKlRxXu/OKQ1N/jcGS+9U3PMupfVplRPbz0cB
CahiAw781BCNgG9KjiDTkJLX4KVOANfBKbquO58a5ziBWpNakLs0egon/4f4HJk6xloKbzls9/bV
KmUpq6jNkRrxNdRG2jON3EGHQjaSmWMPsAx3SQVxIVL3DfD0GdvHW1mjDQLaIOe3j/6e2b0cQDtg
TTuDWgdnN7q1TsqTs50WylGCLj7IKoKzW48/fIwZ7VhnFQmD2zSM1/oiFAw4+VTIuhD1MVSekqkz
udSBcEvvKTvTVH4vgKWZjkLHQ+AolxXXbXI2nl++WvhKDas5yY8/AWNs2+TOL747pt7+fL5N6GsN
6P2fTW0NX8uO2FYcj/bBDGGFLUt/FQgsjEIKsy2e4VqMStwBIELIhHPJNbcBS67FNkerngRP5LVU
6fAT9wq677QbirQvupRL/iUnItMClzP1XVSYhsQJ0DqhMXW8hl2NWlPbZb7srXwjmENzrHvdbJAr
RWLu2cMtGko+BM7b9maiTRGKmvJkjXtnJftQSuuYdVt1+vQeXxrJm5UD0s8sEABvpJJK+TxAMPwq
ORd3U+8Coewr52y9IKmEXKPoFAJktHTUbPHONkALelcJbWZwR5Ns1AyodoKboZe9TS+fv8Sf+wpa
LXnk4WUGaiEvLbqhhkGcnhATTcVx+TfSiQENUWquhDanyiiitwmPi6fssi03egjbshvgBQRVi0p4
0aihVSHRFFYagn3+pGdMXLHufDdEdOEql8cReFDz8yO+9RPfwqG8Rktx7NfrIZtaeCtmcJ17SyRh
4FaODe8ka0Gp/HltlnLrPCx/QANuKEk07MjiL/Ylbo0TGEkDhmJ4EJk7ekp/wNyqo0InffkHL67L
6dsibYn3NaY090uYO/O+nSlmNQGo2FqDvJpAZVjx2AAj3hospu3b1PigwKtJLKUdJXnYv5vAlAz1
EE36O1eUWa6bm8MErTQyg3JUqNaQ5B5xCdrO5G3AoAAE2PDGQi4sIigHkFhmVfreLqjnvcRwLYlE
+Q3li129gAhodG/FYldIlJ8IaloGkmiBZT9rfyIcHF8sjeMzYhrfXsjSv1kC6GP/D11muNBFKiHc
MtiZlK4Y0++ctxHzf+vWtiFZ6Rz0EBxZ5DdOlYtDpVi3fdwbdrkm5+a8oq23gWCfA188rzjj2jFZ
1vbiuBrzhXg9fcQhP5FNQ30AIXBwC1ix3sqP3nbQE3T1vn5rZWIGP3/dTzyRGBkVPR9Phr2UXR3j
4HaJeJNLEBaOiFF8RN6+wExCDuk6g4Th1W66gD+R/HJwIrfb6Afr4Sp2Xh9QEdSS9IUn1YBbfzo5
wnh9IlaVIY3edq++5q63v+kyoxI3cKkLQFYC3gT28o1KzoTRbeyK/FaOMcfsk1fPRq2dF3C8b/Cm
Zgz7FYAMRQQ+LyRCcAw9Lm2KOLsHbdWQS1nUDlSNt1idZOFi05iQAT4+jfpfiZNB1eSxAKNagI8M
lB1OKrWLascV8GmbtBDive85Naai+PsHdHLtvQOm+WYtOnw3etxKvlKu1Bh7roIaPNFN1aev26OO
uq+gGDiifIWEg2D5q0rGqWZ+LDyw5MYAwhAeJm6NT/adrry8wu1+E+YmP7/SecIPYwvBiG1ljKiz
KkEOZAKpZdr8s839wWYl+c0Jwiz6DqfniJ24l7fyykBMeWCbNbKf8Rzt/ZREX9TbthlDDj/T5waP
vqualPgSwbXNZfDJcRqJcZFAeEx27WiMY1bsCVLpOFlHIGSJXJ4OebXETScpkusDQftiS0wgWF9P
1FXBd+2Y3xWT2fTmgyPI9fw5RTKTPAgqnJUIpjKV17d1ugo2p7cMdq6rJQieEgFYBNaaqts8y9aI
sgN2ZLkmF6QOF7sk3Qjq2IswGrJDQbZV/tbfWyOMPmN9wLxNwvjIrfUiW4bgJ9YgGrBTPlN8KYkt
Une0RPJ01jTP9gBmq9iJov3FrjmC/NboJR0NmnBG2ErY0BsJAIQ9zQNTmt7T45Hp71sMyLaNrqt1
g8QkXVKrPWJYGGFgchceC6WAB1ivHaD8Sozah4uW8DKqtSyE9nTUZO6+6IrrXodVEciaM10+Etnu
Z/jCRRHrKepOeE++Ap7DqV7AC9wn847hAMEw3EU70HizVcWdHRuv4jla15k/lEO+PvCrxhT4VceV
C5yqWnIxlTGIZ9Hvic8s/HHfTxw97R2ZyqdFxA3rRkBQm1RMRij/WO3t9T7msOqKTQ04JOjvahj8
7vUcn+itEEUF0o15QAjcuBlTMmO5GvbQuC8vh1IppcZqe03zVGGeLLXbp3y22kL/udV9utiSU/OW
t4EEQN5l5Lwfng+iDRouYnjuL9T01t1PufVP64tKaJrdaTTTH9zuvCjJ9HotKr+EXGikYGJ+fE2d
eJTjE5yU8wGDsf2Gd8goI0FFsyJPbpv+FdaV/zqL3A+6kxCWRiIx1wlbhQ/GBR5A5KPF1UDn9jJs
dBiFnAnlrY0Yi3lIDyQbssLD+NXvHKf4JiZtbMmUQzax0TIRAa36cB3AyoC3O+rX7E2pM19ZqRL2
PihENYoxCkiArmb9LfMsJ1HXbuJ8HUqOCQ7J4iCFlUIu7DxrmvyxbOGiI5qbSgbabR7BlGh8U/6G
+I6mEb0Cl/vD1+5F3YhS9nc/WzInXm3R7WfNNgiyER9jD7IcgO1PqbaLqhCTo9bE3wwqx84xFLN1
M0cEpdTIWrFXISGX3tyMOzJIVW9rOy8V+kGUTSFz0CljtXi7AkTqIfjW/ieNRoRFzEDEkJEfpy+o
Gc9nmqcTYBGwCeGosNBcPQcn/QDLwi1VfhP189qNFpQBXvn8mqWBJNypHVay4myV0jWJXgPC4KfA
PIyoueAWiMbd6GUHUQreFwkcwjIe738xjnjK4s/CJSKP7OKDOJDFivtgFDbsi8kBRhBCrR7T20/B
hM1tsGZyfiSCkIT3oqh88GIBdN9RWFl/24z9vDlmZk9TXxnUmyhYArVqCL7GwtjrjYeuuLsaAjYY
rXyo4VfXnr5CRHk7u5rBgWWvfL9s/DiiVjW5DLUTP4dkOWRrKZP4f79LX7vhHGUiKgJ6GVYOvFe+
Uj7656m1rLzFhK8Y6BbXKjaPR+cWxr5tk9P4vmtmiDcxdOIVBxjdiSbvcUBgDy5iZbQ/WidKCBPZ
zoWEV8nIT2wA/hOyG4+dMEWvFYbIOAEx4Y/wJ5G/5u8vjwdA4VLrQSKaqWOpborNnpy8TPbrn9CU
AHaBDtHe67nG1X3aa1ccexIwzCGqOIfc2Atiz5hcOf0g5g6m9PbKRjeoE5RK30n5nfnRJ0oGg/WS
ekr7wZrJELojZaLzdyQTIRwFD38aOBOQ3OFA0I9TT8uuEyiGebrS5aHEQwifyltYfVf/ZmPbmd9E
J9d6KCtkW2pWiiZc0DhcVDtfcxGM256dFujP2N4LJvDfCJp+ey2I/IkqonCUDKFpupqUKkSsX+oc
e86D8RKNknp71LKlW0nw+o+IW7hwZ61N7mhmH3q0hyGdFMQf6VbOv8fuw8wquQUUfTag3kQ5VGEq
PiSUY8E9g8UBm+6hJmvkFD24VEV9zDsoHoInVrorQU4aKjuXPjCGv+rYKb1qOCjFgwpZpbpAyezm
RtAXZKzpB0J2xaWFJZBwkUKiNklNi5EGQ4OfzDzMvZgWMKsCEevFyx776YYXQI+h+L+FHWK/Evvx
uwD56jyy3kiGK5tg+mP2/eqOAGcsLdeSYvsR/aALY9ZR46gaYk9iwvqWEaNmshCR99d0mXw9DyKV
FKzeg9ziVDBkpJI+TsfsUohiQpoRTPM3FpmvY5ajt2wlWTzaY1cjHDezS50PQ56ByhZ8GtxtUeYG
nKYp9lDKTRh4x+aVwUXxyKCxLRH8TqUWNnJOyjhlODvBvHzJ0cmtFjVcqA8pwJGK1q7WMEVVURzh
OxDx75JGM23bEpuRVEKiXMjB+aRSOm8TiZNkC2r22NpBCF0jlhqMJuyOKrIDAUS4Sf9l+zj+5C+a
qR5JyaixZnpjpb6+I23cWQuwuQIuE0HSHzSnEQ5Tf+7vhVFbWuy4eOEqQ9cVAm8Jely+lt+0pT+V
KnyOS/wf8pLHrnmYuLDRb1APwjkLD9LXXEPiazh2zKrSX1qkTQ004V25kB4S4OaH3qqr3q90iS3H
0P7uPV0dlqQ88Z5LOl6CUjWZRmRAVCfkbtc2nvF6D+iqtxzTUX46uB8Qby3keeV1F7UHbgpTds/n
op/R6pEMCrJZr085vqGt4ryzvdXkz52UkGGxrtGAhuX8pt6Dm5xy9JYRiq6YlKAA4aPZLXf7BQzW
y9xdqUAO7FNzOPqqFONbQWZm9ylPZqPGrMII/SbnRuhrXbGMP2XzpIYnJ3EZ6R1iHarkaBgS6nTe
eiuKIr9IMH+e+JSGA8vi1JO9DVwAv8uSlM78EVi7CYWf5z/NTQ8rAjzmSLkVschSWNbHUYikt+ME
c+Vkq2TdzCOqLt1XhWZkOX4VM6qyRd8ZwdMb15LsyFBTQtvDVrTgHm5vkgBb8grZbIvhnoxRVeZx
fvActoKtqTe++L2Qnyoe5Og32d0z+xCAVTSzfYGEN++JTk+Q538nybk+oMf7JyROY0IR1w+E3985
pJ/qerojrXPIF99nwbMABpSN+4uoNU82icpJzrHBxZ4kX7L0Sdjz3XveWfZkYjqrTSlA4MsgOJLJ
0d8ApRF5frF+MBhXQQeOXC+utn8VsWeEmpLz0QXN4ZJGM9TPEynTmAhDDEij+tsCQ+ziv358mN4m
j5vEksqH8COnPvtIAGFOGZfa/cLfbk2oMYUI1StgYO5Oiqtovb8n5CzCEWW6TNnZgEWcQtp+hkLI
ki0Jddk5B2g7IJ7vviSWS1RMDeZtc1+ciGW1owpiQ6NcS3pfjtkYsyQe/SPAQx2YGJQbUjNsYUHc
bNHyIxCw3af9LGbfNF4x2uEQwcuX6HNX3p+OkSECLb70Oq6QYjfVPDEEQoURTg8wkUGr/bNKSER3
nO5DDydfUkqbAyJxlM2kbozoJiIx4QvD9eI8mKfPKT/xF2mODTlEjE74pq5vnHjQs/+3VcCajF3G
JqGggPKChHsCvXKbWazdUjFHG0gNUvMe5VRszsqEeraqewFKiv0de7tOVHbj4saFmtSp4XhGRVyK
QzofJ6mTqsXMhwSFLlfgrcKa4eclfbCfRu8MzgWl6I/NCcstC49K2S0Pr9528z1LnfldYGNe2JFG
6G4p5aqXG/1PBporz1b0pDDFNX9F1nSHMW/uW0A0ISdrm7qDZvwNHhX9g0G2Kgzhd12CCBFpJf19
Kn6Vn0yV6sF/lI9jkzvxic+K17mihpqpqFyz8HPCN6E7tDEln7GBb/CQXkUI7cMvo0kZMiZdXwtt
/E6Ob6zlFiFw1HjUl5Z/ozEAb+TRZm9uRCJwn/69XPftP2phzK7rrWrLu130xIh3vqA6ejs/rjsd
IXLzaY8eHc4RlW4u0n77fbilU2FA8QKN1UCElZBzBgmoNf/11lqqRprI9UuunzpFI2lAnQKZQGjY
y1WIK0235ajkxo/WPTrjny8yFegNT8+lOXKi3P2RiBmuY6kmxZok/gr7K8pjiy8F62iskNWd591J
RwoIvAwRAsJr9sJwHmDd2W9ezhTs3Uu2hVbTZ66MgwdRlGjWS9Cj3idabfPak018Zbg+rISgARPm
TtLV9S79xJCdrQATzRN5OidvY0QohrT+z0OeVGxgFiI8qrDfvfritvnGjLLuluPsmNuGamuC924c
srstey//zTBQ/mQp29nuDoEYGibLlf8wDMtPQRFyFDqA1eqif5qJVAWavdLjKfAHeJSqRaNOiE0n
tz7Mnq6MHzvzUVmvjVAj+QvXuoW7lqKpOvMGP6UDPuSTgcOGE7NZ4tBBoO79ezY4YmwXWWO2mRvN
M5EPmmUbCNs4F7gjccrGsYUwGme73wQZE/EOTcIYS3Lj8V3yB38YIYN1h4vSauYqdQ6BQdlEB+EC
IMqxiJ9MIbhCRWXcrp33wNk00usECQ2yRmKqCMdAklylGIo7rGPFUiJ49STuszTg1jAh3VfJ7Za/
eJsmanKcvIn2NHzNj5hachtu/085iDr7et3iq3LfubL6VeoTK+NsqkCeoeYbpuA4fWKXoXs49Kql
L1G+KEuse5m2u6bSRqkmPI8W6deGDiqylRJG90rvGEqEX/5Sdpwb/OEsSifIrMODkd9tpwglExoj
+MdqxnHA7ULJG3n8F7S7vAa8Oxk0mZia9qM879zSUTP9caZ4JoAbcIjyLY8ai1EAaetN6UL0UJpy
aB9dRAy7HOJlZqNLc/VmV8qjOQBL8WDfg9Oy1D+ehE4o8CjqUd2PqlNWMxbuQJ0d/lHR9slsJiIg
4h5ZiiroCKW9Zan7zJfMYhoeg45DewQw9P8tJBxW0u0LL+ePoCmAfVvaHaE1ChJNGesp0JnneDwh
evK1EYlXW+g5NW7bhxr6HKCgvMYr53bsTBf8O58u0gglwk18zQ4FOS+xasPT+T35VcGIEjD2kvzC
kv9Sz4+LofD9ClwCS+dkoUY75bb4mlT2gaH7ehJShjOgjHHcMA/UOqmcRC0xSOQuQ9Fc7ehxsSja
TfEZTeSHLEgkfG1WEyZC0ZLT4tD4YB/ElO/nHtqht5l2VdvC6hkiwzo6P41HCxzyyzi4fyyJzi48
vqhWRAVZ03PXTmRT1uCY45SepCHotnWLqQGiWNw/P3u3Sf43vbVTXOvGOz0UODZvnW5vKJRYI63m
+Gv56oHxoBlk5kJosQB0WwetOkKp5XHXvhF+oH7IbYmOqN/hcq6q+lfV2EHX5fj2CFTA13UhkcyY
ZdtB3OM0FMY7NF+iSFoPs+qSZ/9BEqWB9WK5SGLE5X1WfPqZl/btBg3obb0LNim7Sl6fnFq6O3M4
hYrdkUFn9pYyjx6Iumo+YEALlb9+0uQulvH2VMXB3RHrNOAGLc+G9IkTvVzSmcFnq8/nGs/a8F4L
aJBWmmbjl+TUtMF4JWaGBdL1ftrEu/uILUPwYTlmy3oKi7a4ZrCpzvJA+TCyt292uQq97pljUfT6
jpIlgTWir+ETgY3x+N2lpXgWx/Ai61Y9/k2hvpGgwgf8f2UKPsObJpbUHI7JELoETVpYI2TVnRpj
re89EkGvOXIrhDN1ZhTCZsfFFN84rrrym2adgIV0v711EI8+6P4A8Q3loF2DAuCplOJDf+5B0YmJ
MrQbH4mzKqlVk9zurLdhPSTFWrEZgHribVBXMlngaNm6gCZ/Ol15AUBZAGzFNTUdz7xuhN6guZkk
Oz/ZIx9iUun86d0qjMxONewSfSvfsl06nAtYAzlTQh1cpSX5JPFh+63Ce2rtjDuT9cRoBFDNiKjV
tCtvYmFokaNS/B881+AEOnSfIvUlTiA5YTGownJrZ2c3JQgBkawpe2UXpH7Y0IsPC6XUHNPQa+Bl
h1ltSTI16lXAUlR/jcuI01juo6ucPiJDAJ4vOOERJ9USPm92K9eU4Cew2AOOiHpGftXm2MopH/kx
FiryGdEEsaK2BASN4qhD7rFqRxnlDxAdYG92f/4xAogBBh3SZJTGCA4oLwHQ61Ejg5NFmVYg+HZL
3yBfSELwVwDdiYqebSiUWDuOyoPKDUKuEqsEEcYpZ2Olz4qqT57nF3fVLRd3pvUX8ShfcajRfgUx
ijSYg7kEZLMSCig+QcJ53iUJROeljVqPc0ntzRu80U+7eZmogMYvXK2juRgjfBfaKne4vj2+sYGH
WEJ2T3tHrU1oHqNc6w8GFEJnUI+1kQvHln/ZRmDoxGUQQxc6gWBratHgk2pPDvgm60M8ldvNif1m
DSf8wS+GVazuVrQzh5xRd42g0BXFS4+CymN+AAie8HlkWueYXqdIbXVkMQ1zb87riNO9+6cp97U6
XdTFUYkO6ArzsJqL6OiAyfWasuzPbxe2DqknJNeMZG25xwet1/E02V7QUjzgHIBRjPR2Rv1SVX+0
qzbHjqpkcV5luaIkczWPWGCjRO2OJWdt12Wu2w+reTlhrzlbqif8yqxgnlqav0ces9RF81tLH/ws
kYv8uHAV7OuRQ6XBh0ZjAs+WjVZdeqd955PJY9q/Yz0lTcB7LlYC/w9V/hXZnnCX+UCY9eQ/OkDF
m3AeJoEz94hQo6+JB1LdIlOjTV9M6fJMMDR+RVmaGBRcJr1TeqtNY4FhLhgO1BVvT8/uCMsIX9vY
6fhsR6F3NgDZqpQ0d+Ik5JZDACbH2iUZXNY8defTog2Du5BWOQVtQadDHZWlWaZ5Yo61nZ5OeURO
RV6vUfB6IhICnOIoqrLYCS3BM7zmYUezOrbXTxUW5Fr1snCp9YUQSA5z8PEqkOwBtQl4oYd1hvgv
cp5XloFKSN2HUtCV5JOfqze57CbeXOh7IpVZmXO/oObK2gakozLfTY6UrtZQTcqEzBi3WTyjH93s
c9FHOCMA86j8EO+NX46HpJW0sfqIqGI/F4nQxiRCbRGdYdaiJW0qIzS8gPruOd5pygnLr1+aS7OB
jG66+BJ+ApNr5EPW2DhqkKysJ411EsNx8Yv0srd/okcxcGOq+6bws6EezgAHjQn9grm1Pnj/f7jF
LNjZysQ7Ai6E7xJDZ/a7pwqyyO0yr5HpoP+vReEYXYeOARllRfj5bhm8Mnd96LMg/H6yh5/Ivo9T
arQeGPnwactebFuNjkfEEoVJa0m2bP6MUq6AuDlsvQ8dw9JwlmdfR4m0/2KVzW8gSNt2ft+o9dsz
5IZLvfaTVo35LFvIee8r+RPc9J2sArtR60P6Q3S86pHBZIQK5IriNwp8N6lhUx2ixlVG3D7a0dra
xNZdYUqx0JphnNobaGsq4a4ehtTZ87DZRohtEqobnlN1jijkL2+I/kusa1htQXP9Sz3nE33qgTza
y4Zs4VP4wAHfyQgt7wXVY62XQEmeT1u/ivfG9YLe7dUEEQ2HqL5V9OY1TvUMbvswWacjh6DgbXLP
WAgviS1o9v5RhVZU+GYEopH8cHl8vvhmt7b57CUdMjIyr/h3iifkS3NDv089lfx3WueqQrNWnRGT
UsPvPb+++OBq89vq8WP+DgbqCbobxIGnJ0aj7fkvlI9eSTq92B+YRGofzlndEqnPOxTD7JnHVZiP
MTZJNX9m2O+c9VmNn7ILPbp6GrvBjbz38+AFJJeW0EJ8o33SBOTY+K7Po0Ml3/BOoJ3lhgJ1Bdjn
hX6hPUWvVOYoTOkOfkFncY0yusS3GnrOCyAjQcx4Tj62dYQPzRXszpIXAxRycmlnVwaJtDk0WuKh
/lGF4hNEz1CLA4rTJgSMG0GfJMgYJsetI0n4tEyk5Y+3RbwUP1r1la4W1noF3wEkA35gbFQYu0il
6baunfRSALe0rn1OZPVDiGW4OvP/ijA6ResbOF30tif37OMbTdi2coOt/ZKfjHZdM4GcyNnlpD5H
V+ayKJnE5ozzpFGP849ApYdOFzBOubvPS6LGaKiC1Cb5IDAc3smSQP6lCqYialf6Zo1tHLcFXgex
7Grh+/SG5Dzzu3nSNYh70ri2nU69D6Fkv6Knij6LHjyerdnhCnxRHhsuIgtArc4+xmFgk5gmI1VJ
+BOHswMT/4kCaVipSiIn+P3IUJ96P3pNjdgqZD/uqvzAX9LxwQsA269Wk5BSiEID4hE8cOsKrByo
Ksz0H9qvE7rbSbujNNO6KBOa5glriqGJl/x2+FC8d0NqLaMP2J5TGE1ceWxtspMMMKllQAtjq2OA
lftK8XiT6o1WjCF6Ow+6XT8fcwY6WHbL4UuZZR6Jhf3kwbATjVYGb/HRscYPNwrg6bJyuKGKSXwJ
EWhJ9eiBFvSTdTsdmEO2sx5Guep+m2ASsbKUsx74jCxDAk5WWZR6weNOBvOrtllq8KjlKnx3Yc3n
t1ttdo2ipqatDXcoTPfcawCURLpMMbkx9D5wpqv5Ifh+svSKmz2BC39EcVaq5vGJWTYOEeCEF8Z3
hgUCGHF2te/tUFTiIVa198Adq9Rv5DdHOZKej11QJ1rGjudwAslCB6IoJa1rTZd3IdPZbfmtI1C1
pBQFs85nkc5DOKmi5irZHrnhgxWL3xegu+aEBA+lPfk+iqZgTI3GfanQ2h3Rg8MMVX0usmBV0HRG
XrsyO7Ab97Kpu00/zv/nHBj1JL1RbP6Au1FI5BGFv2dr07HZVgYf2TCZlyJ1vx3cdKJ+RV2oFNxB
rPQ/6EuJsyeH6DwVfmjYEUc620365PkM8wlatmQ0UvvIdldZR9hSvUUsGHqmDxX/9x8G//OTRjh/
w4t1acE9/stXCfkbO01BNo9q2BaQPlCLW9pkFp6em40f9cOW9EOxyGFRsaINd97LGxTJUBowRBwH
8DhicZ46IgMB8vF0XT6lZ5QyGXIC13BSP/6aWM5/IN1E9uCg2Rb7DLw1ec8bc6Ece3UkuCNX6TpN
oEVW/b+tNXkszD4sk+W5jW/NsVAyrp6wjVFDo5t/DXwd9sbF1U1oaL3G9xjKtQwttU4Dk+cBgaKo
Y8cvUkhYGJk+1fkgs1GYjf5fGbSfx78neFO2TTb2N3UrfU9/WKBHsMtDdLYemdCBmH2nWO0eqo/z
jRhS2P0fw74R/EGlZTD5l5B66lfPlyFKCNLmkzsAkqfV6N+QAY9rjMbulmyRcqvreqAfdb//LbHU
9p3iH3n+uCQA4zxhpbHW0IkYd3erZ76BtPB+hKVTYHzDtUPBjp1Gv8KzgT6w7fSs1pLg26AKGtgX
FQ29EtfHF4XjeI8v8CUS1GmX6fZTMvzSca8BNup2xuNXb4uwECrKgzafqA4x9Iyo8Yq2QLspQtHl
IpUEXT0po6maNcFmJwrN91UmN3Hk/zrEAEhPwUL7ffC0LWHhdM7yNHFczcQKeA0pxJENAOBfJ2Xt
ZE75247v5vF8gSkrHOxm8wLim5smM3Stv9qCnd/5cx2XAVaeFJO4+uZynB2jTdvzyXOFLbX/WmKU
NFFEfdLBYZREqGluqO/cdqh3fOqKBFAa52NcqiHeWlCnteqQMogEJo7v0r4UopcZkng+3vBYLWhI
k9lunj3IDO6ht+5h1mtK5mLxvpUgz+wPtdQlF9Bx2YlVq3NwMNx7SsDMe+9VH3FwsduPiOFvrr3f
nbEJzrhBRyk9womzBSppztYBhaTNePyRwXeAAb+VD1gBrYzmNFlNzvEPnnHZZPTKo5XMHv2l+92w
7qnNuihYFzkSJprwOhJH1u/6pl7G+WE5w2N5bRnqLIvToOY20I5FSHUXrFhc6cG1suPd5tsN4yFl
2QDVj70lVP3TN11KJ0FS57qS4FIcsJeO/HbbHc41CVVmSBn6JeLUF/tyUHREO++ERCNilFNipUlA
r9Zjf/E5hzOLIxpZC6tBAxsf7GTaLux0sGj82/ZnDv9UcE1NP1URFr7iu4PwXVky3QdCVcp83CY1
Yx3JRBMLqhOvQlGntm/XNruPEAr8+/8RmKw082d1o4zJlRacKwcF77kFAy3k7wATGRWg5SsWFpex
r47CzgZ/HgaNt5tA4fiQ2/4EU7Lre1gtTszCNeyhppKVwpgpNjSvEBKHyuX0qEWT7B1EJeOgA3jK
i+aVJM5gWg4H2rtUEWeL6uto+a5ADkXmD2qFs/e7wCEPDp0fcZqwxc+sJeEb8kswVM3YszjPaPVF
UQc0O/glWwwrLSm/QM957bdmapsCkaVeBz3a6AJMgYcWWg4cgSTbDshofNoDjBTX7lc9TM6kHWEA
/Is9+pfX+N2nEvOeL57BBf6tQfZ/BpshHInDUv0lRYuw5W9oR618WNLyCUYbGUUfRKx6jtr3y5Q5
m5qfT/RtTzQkgrdaszGmhs2vg9D4RpFwvq5kP2Uwf9fXdrxfh+nslKJtsp8ehDWoyBgtg4/tFFlI
0hkHWHNtqtSOXrdFtiD5uYd1c0pK+pKVil8O7t7ibO2IMqICw7BfTXaDWvahTi+ZKZbA94/zR8Fx
OliaXFFDExEnaz/hSYIcqhYg21vg54p778X7dKnnUVhGdhNEn0tgCYC3/Ir21GvD7udYoDDq+oLh
zB8J9orztC+SULJdfi6oUosib72wbKjIWqwHcVWXJGjZBpuKElrUjDHkow2UEzAl3RaLLWpMD8+y
Ugf43nOK4nhCVvCBcVo5o8/Q/dhgSwuPam+Db4bE3qf419Xf5Aq6hGzZ3Ylep16xGVOGm7yTF6tE
JRNwHdt5WnrV2/kVedLyEOiOJHdhLVylFKAbI7vJ095OYWXuekEc4hB2sUxqGc2KUAMt8GPtCNBR
MqMRZ+/JkrbmxPonKJ0un0Q9t9ebKvOU+L+k9CStdGre2aZ3vc3HN17EGa67rlqG2DcuGhwSuE+B
w/6aEXCm0/Ad8SFGeeEcH21Bwc/G7xcKeYu/9ZEzCPMtjihd5VYO8ead+ZGuf2g2r3C+jkN9YLju
ljH51aSHGklkwjcxefxF0iuG87soglxK7uzESE6tcxsrpTsV51WSXYMlOrtXla6UAUwA9VP92LZ6
taTcVrt/yhlh7EDeF06Q2p/ZUiiZpXJwX94WliyR9kCKDK23IPhKAI46b0kQO3sTKPPOMRYNMZMG
Kln/CcsYA8fbGImjjdXgGCgU55TvUr/qAn9sdly6kdu0XLtxySV8j+TCLLeMENrH9GysFWna1EYZ
JfJWs8gvEuzsusx31ys/6JwsqDZYBt8eq15dc580Q9xzJGP70BLDvo/jTFzCko54rlGL0HUJLEPH
1nqYDtqt9SQorQYXMJFB16cCNTwt+OjTGI+bB3GLN9wiAYUQRPWT2xirxMN7TFmSxjBznpmBx55F
txPNODkw+q5dTQ0u0Vg1+lg4yoavaop06gvj5AuraruUo72dX9R5kXzQyOkGx+vK6OYQUnYjFaVW
W7FDgoTFdvcQcVVNQlX04vk0TEWUYK9lqp19Li29/G9z+pHD1rgSkbGnn0hn0oeYsFueiLvFtN7c
2QseD++aSx//y0MtxdPZ8d/HzwXqzMP/HJiJw5UXXaTJqXD6FlGnpjl5k+VXE4yodW/9qrfkC2gk
036Yp4fKj+d/pFumiQlD3dBOIDoxTzYiJ86Q9SWvUl05U4RPL0eU7beYgMSXcCaJrnKasarNdrnh
8a4SXJ2dqxFTBCMfmmX9L1ggGD6UWPgi6xFP3u4+O5CWTdlq+b55ZimsxfmW6v0O69yif6/jIQf9
Dzjmlqpzf6U7YCGgO30BpCFwYEafF1ppwAuKzi3nhbX00rGXW0VSgcI5e8aeQN87mOUm2EJOQteg
upCix1+BWSGcAhP9iPZR3oC0ESat37SeaBRsOr8B83xDSAsFdsfKdwLvWXsJgMv9eJ2DRRdvHn1u
sEFGYoNYMAlXkWME/4SkGXLs1G3pjk1Boo1T52yIo4pysMkMtALc6gzT5/rUOMexpunsd8MBL9fG
Q8yWJoPiyDTYMN7isOFNhnreQLFG1OvhbrQhQO6Fm7Baa9MiH2ATteFkgx6kiQlxh5N3gFDCNZjl
f0NiONqOUXNzv5J3UIiUL07ilTdC4+vWWnQArnvLDMrA2MpiXC7k/R2utM0y7vKsYBXLQKTpxRLS
Jv3U9eY09QEibBKVPvh7dfU8i8xe4KTiOjGxN9A1AYhqH8esWyfmoNcPs4hxuCWw3i3KPdC+BNji
HZfQX632VhBTWfSe3enIpGja6PU2coWQVQ60N6H4we0UP3aiuJtoYaMz7Sp9m4iqnz78Q+z5rM3f
5ZbMqYAQvrZJtUsQCrImKvuzs+hvqDgtgQphqQRnl9bJTZ8itDACwyhy/oJfWrdB10UUbRLnrKhw
JBy/Cl9lXFO1KGgpho6MgW2miYCyVBwzy+pF2hE10zvoeNVRMwILwaGEwzdIXTkagtWFVD3/akrp
skkX2wCDW4QlWrZ12mL1AAtKG5eXCB/qgA2IXtVJnMOmjZVV/TFvSqaTfAAgqn8Qf5iyN+M0O9uw
P+nnOF00ymXv6zzfQqrHc6cVOtYDlbX7Mgz0CHFCgIaRdYsjbNauOvWzIbNksHb4XbEarYJILNA8
Em1e2ijvjWfDJ2yALHw1IhnoAhbDf6iQXi7d94QmLIhKHVAEvQH3Ih0dRMMcRav8HKzNMmi8Y27V
IQNoO+rOY9uDR86h4mNbeGkecLQWX5HraRkskNB4ae785nzQb7DcJ50UU5y/9EqJ3F8qzDxlMknO
uI0sZZ7wpdkXKf7ZuWKleSKnNGj4/3yxEYkmstqkStnOmkjX/dHL8PpqdpPqUBdf/UFZT1fSdqxh
sTkTm1gxrtbCCZDcVG5ut7FqaXhfa9/sHbVHqQQ1Y+0KOzuKy59j5aEkHIC0iP9i/vfS2A0PNRAh
QZHnWRJoozSOXp/zwUg7a4GCkmb9mje2pQ+fewvRUGAtM93H6muXSVYX9kzTE4QZOxNSk3xZPz5F
fNcCPQAcBeEtCGPLp394/bhJSrGP1eWcY1mlH0bY8iN7QH707J2kGMydeEfE4imEa6r2/NgHlxEp
diYvO7em/4d1iZL53hQTKIO9esg94Y45SFwhH3YiMZ+t5b9CmT136jl7NreA63AbGNlHecPTJu6L
2AxejYc2iIUld2w80cjXeAaoEYO+ZoGUmI7La1LF0BOK0Q184pzXj1gBuepBAZO/Y/elCJ7VcLf4
d55sMQm4AP/Xj3wMVERAuLZDlswR+IRFKNMrmL992A7eTJy8cD7UFG1S152qZ6a846gxY21/l7V+
mZJYcXUQnzSIPxliWmhHnfSZ5qC+WWOgPepgRmHcpkyPjtRV9p3l/jNP/PVeC9xSAH2g9XeXeG7I
rCeQOSEl6ihWJZmsT45yS56/2zh/m/RJeOKYdMO4ZAxJAwhMBjPrOPOW0LmHAVerNecenIvVSgEm
U+6WU/wtReL4iSN+BMUpoKraLMxxbMXd7RkIbop4JkHGWbGqDkzrCaZmAywXAsRLC0ehzj+LUDFn
FG8lDZmQ5Ju/LH3my7CN/LYE79DN3htdDUMWv9Fu0TEsiozlVurIWNlDyayCZAE3+n+5PTr8DgsF
nh5fK20UOw+tTfchynqPV3uZt7ZXaQwUoEG3s8eRSbuuiI5UeQC8gPnfCx4pEyRvutIOu5hIj9ei
FfYcFaMvorbd+FTdM39+IIDstYS5RtQPSiiumFUmhd47auvNNYShFrL0f2j4pseo6IaNd5AS6kAA
aFqA2cnfbR/ySYc9VLwZY8TF1+Zb1ppd66zxaDFA3qpo2NiMFZwrOiebvQWsGrVTDVZ82v7VA7PP
9m0i9fbFbTcOyoFSfqNGtnhNopRXKbUcG80n5SM5P3GYEIgodEJT0n/8uspJ3hiKxWgjGFZCZqKG
LA2jTd0i9u+lVv3YFsvu+NI+8ZHkBajI4Rxwv0jSuoGVofcyNvfsyMH4aj1Ce/ED4X5nsnXlpozU
in/Xz5tNDQpincK+sldFKsm5JLfdbPBbNw8JoOH/eXb6hkoi1L/pOalwjfS2IV3psjwhPqWOlaax
GfJUY0nBHfAzze8qLI6K65ZnS8sLz+f4Gh9nWJ4Cx0l/rJroOJpq2LgVwlWjY966Tn8dczjv/zOe
wG0bngcccSldocTV13zxlT/jg0LrJwZ3ow80ApE6oyQGqBrH8ZER5eCEctRsoZ0hRNaVEZ3WLP5t
3gRdKCAS6M33I3kONH4PTxA8ANeZAIHvihrOqD4cysXza24ODPu64It/M+ZiT99r1F1fFUCfQdG8
4AnHUHj5qYYWN+XuCNdRiPERChwkNf63UwGlqTJ2YNdLIPg4mzSzjIxsj/9ABNpbCuKUrqjQEJ0D
rTFev8Psda3vvZyfmpET9Bs+S1f6dxLQCPKBAovOIq718WSDBKcdfa+nkjXSL8IOK9rNF2k2XpME
DqzO2726z0oPEZyF8ziVLKgLrQfESNW14fgN5m/uU+bUaGNHfJJUOyz8sSQW13KF5bmY16pc6+cD
YJB2Jo87DTfHy1ap4JriyH4bC6dYRha1lhAhR5Im61tax+d0dGy1Hcwl48JY6NmiuZmr4rseMRAV
fMZ/Ttu9SnuXDZgIdK6Gxo40kyk9fhOw6+CRZ/Mbxc/mhzoVYCFDwWieVv6Z1JC9X1B7WF6uwX33
1H8afZiYYMM7NsVdcE8r7lHCd44tsQ1OQx/65XCRcIDVq2KV+iGN3vdeLgQp3gp+i5oUvUtuaYJu
7NZZpwQ3ZC6g+tQVB/zD++9zjza4SdgfLyByw4DvMXgUOHqN7/8kwT9XmCbm/Hk/F8dXxQCbsM6k
xdLGP/jA3H/jGjFaqa+Bx/7oUYWqfoeStV80AQxKnFQtfXvPVto6HmC0Icq4mZnUB1MmmFvCbjLq
jhhR4b6oI7UmA8wjkXnRq0SFh+9mM96+qVrL6cvS0AJFl0v4ZKczrpTHLGPafn66RubfFTbwYr2U
mH2DFxLgcuhcRmEDd/SEkOT5/z0NIl5bBfg+3i6nx97esrBYmLndMKV/TNuzqHqsvfb/DEAB5rlv
xYIDL1cjLtcnBzOceR6F6BkQZ9BfZc2bGDTm7QxhIDTqQihArmV3NqJ3N7tMbeVcVi30kZX6AXkS
6nOWewckPjmdkFDJIKIQr2fqllJ0sNJlv596euUiqVFkSozo306yp9nzXppmYSiBe0ee9BsclNOe
I4Dc+wNM5nUpXcT88prquxF4eQFloyfRvwftlfOatUuRaS5u/njmEMedm+ot9SvOL92COXhryfbK
AXbdQkcDOWzISd0+1MrX+aocJ6kBDlXOjhvm3vGKT2xYnZUNwhWbAg+xB12SVwG4AeIxcMvmaFh3
lPq4q+S/Frq1hHU9LscV60MGIR0wSiLQZJ9eslG1q70bSYv4xR+KDMk4jOMjL/q1M1sJhKmKDhcN
Wg5p+aOgTG7OeN7BGddfcSRzKC4FygcRvooiCH2dStWdcZX+sLzUJXd7ALHWJsVxBMAVANvW2OFy
eHZiixB2aDYHULu1Z3KzODnjJQ7cdnB2SqTkoP2F7YiJBh/fbt7AW3H/z3xTMP+W0qFdnmf4+AIT
H2Vlc/Hydv7r6CsG2HezT0ZxYr3in3Ae2b2N39aG2toLShHacUtUpJq5lkWD8z1ayUB0hiIm0Jka
1Fq6fDqKXLmvUG8RGFA30K5uyRea2aCN3WKLiRxusErf9oUm/BIl1IvdYBToTgEaLqFRunJ9Gwm1
UqVhwmoL2K2v5nsIiH66zXfkHCbrENJPCkXQP4bJQVYw3yOe1lq4wRXfNTGee8e9PY68SyahLLcR
8u4UDkNVLF5yLbmxkRTb4Y2BGeVR1Y89Xf2UIgoafv4+xpjKuJ/mZE3DvsSO/lEhAK+4PaP6gH4j
wqsKfhG898BD4Dls2Vd/zuXrnhpJc4srrttHmOIQlr3cmTCLf7xa/qNf6FYMFBXfipXC0vjeYLRw
wotB3/n8hDwXIcK2dWfYOomhjGJo2n4ozOvQeF/q10RG2nYIQhxGmn71q2x1jEfk/XsNod8vr2SS
N1AesFlLqMbiwmRRZJ2kQtQZesVa80JZd0pz8xNssbwkxnPGY/KYmxmmIzbtNYqMx2LgXJPF7s5J
qF1egXHPJgpkq1tOo0p8z5c+0jft+6aMiCayQen2RUrycycDERImaWZeGECoE5tLaWvuKVrzT34N
rVebWeHfEw2K5CQFifrBtBVywJDlshKNfSlmIJcbA/Us9cks2mxcw0sfK8GRZD1D7bSU9jvXBqyM
OHDAFclugjQHoI6+jRSEQiV1o3siiSSaS6ZpJTuwW7wQB2ASQk79SSJ/79TMul5K/7vqHf7rQ7Yg
/dc+xqc6eDWOpVc73iARm8dOCWeOtnEX0fBdX4K2wavwovC1JdJDXtPgmawq3lYByX56sAV4swGg
BFaHAiiBWRCy1r3m9ukQgqtG5b4YdJ7QNZnVVYndv+wZ6mIgf0SFMYPU98HOOVVMKdnTEs03gaa5
ijsIRJzbJfDsp77IqDr5iSdQrFBLaLuzWaqX1nZattlHf0LebtbD0V8IQs9DJXTFmBo27N0fUJOq
5FuzrYtbXVBmVOGjVicc3lg4VTk2yN7EBnFYT8kU4QDQ+ql77wBHlOYxONAu8PE9mr35hfbO4j0G
qceyyEeRDPG3Nx8EdmUR2YO3w14dXSW2PL1WjfTYC1SXFlSYACyHdxzJvjkOjk+ATWbc7GJ+eQBC
onDQy6J+m3aTcUCrttf2cFSYTahUGbhKVAJ40cj3TlDF3e4MRj8xM3XcjG9YvI0AoxLLz9TP3Dg+
vJJ/l7XPjZBUoxkxsP1XGD/Hw0jQGWnCCJsnlBZKOqaq1Gzqebd0HAS/LQ+Zmv8L5v7eTgqT6K2k
y4wp7d6zbpMO3Bd4fgVxyyeMu1jdDMTwWSBRxFSLdKRGKZLusGTkLPkq70OEjqHeFyIRfA0pJvAx
t6alD2dqnt81PCjXzzuXJvCn4ptiF+L5LdbOMvCvAHD+ATBD0RpjQbQBJspDT/fo3W1W9h6ObJMf
Nk1slNrWVh0qzA6B6FAGy0hQ/PP3NB7OQfty9FHYxba5tzdVq9sFt/Yuwy9TDXn0Nowq2zm2rLmh
Fty+LTxNxJ+PCJhfOQ2rWqs8EYU8akJ7CLkEcB4f7ljHoD9R56dujKmdZQg2Hm2pKfsFpuolM566
nBHdkS/Loaps7/QHsLInUylvM8LUjDAyksyJSpMyOqGYBc++stgiOBTeToCIjSSXevKgrLXoRJ2p
1xU2WG7pXSsl1kS0VH5WzakjCo3sUaPQp7+CUD3iUvfuT9VIux77xece1VN5RRfD0dGLylS/Olp0
6YC9/IpIKEIP7tJnJ2pV0HX/lykxlJLXjjli264f9q4iEonvfiLX79K1c21g3aiLAemUOY3hmZaz
83NXkPvypElJOaP7u61UTRwt6D9+Cayff+lovoVe0Lxc/sQwh1MUUy5E6bYkOi8j24j2U13nXDUT
spNDgrYeAymsyrDokvw4AdLmojlZMHXGzu8BQOlkzLAGrrn5SXKjcpSf6ugQOMjQPHXJBRxtLnZr
fhJY/48bzWq0iVYGnw9wad+WahtB7Y6w5niFvav9N4sdVjmqiPLGR/61sKkR6pc1PoHZWLCzRddN
N/BpKuKB/KhKZEQ37l95Hl2EKwOGbsS6qrJByfGCgbU/zHVKEoBz8NtiOnVL8RTQPyNl0IEd+m55
6dloBVZSgI25D2JAVKu6f71Hd8Oj0g+glNbpGPIKivWyw13BUX307DxtIjnkB24DwjbjGLowJJsD
1CX/xdNzJQNWfVCOaYzatZ3E/pQuEjuY7KxCLc3Z/nWyZcngBGN/bIWLsNzPX990HBmWq8pGNZiL
vAAJmeuN3qptYohJNpm9q/y+jXxL51agE0f+q9R7xpflEbCygGRowDkXwawY9JKfW3fT+mk3AblJ
Rnhi/Sv9lGMNZqmtuscbiwwV45Acenmm6XI4beQ8uAkL9YGhzfyW6KV7PWnQRg0TzQYi2tIVZx1o
P8U/2qp6gouOJQOnzp4dUnSxW2gmbaw1+ML0mqpiG4+wuEZjZerpCE3NMGmmSIqB59rkhEO7CCHD
sX6nM+TXpifx9/QwCU2I2cQXmhljEZrQmQ1BRmoNS/4R3nExMX7OTVjSiyl9cmz5zx5W86bg/yLW
iLDjOGKj6f8mg2VNebxoKP3PKnd8fYMxdhysEt4HmYiPKeQ7mrp/KGxF/8L7Wztm9KghfSnyk4Sh
6XPyoVv7EHexlqlY2yCgfmdvBaxbqTJ849C+9MGoOh4Xp/Lx3AR3/zODtZ2crfr2DO7CApbZwcTD
thn9CvETtS4Z0A2NzDsByF7WRVMgmfJ2vJC8sGMGGdumH3HXSWlZomjEDFSaSYpIy0JsxNWzsVcr
Yat7aAeviqGn88t0fTdxh5qQ32eVEWCBxRkjqXy43br4L27gtR3UX5REAZY/PoReaqEaaawzdJm4
9ohp7kioPHklK7FgMRM97BVLHLdNBH4Ws00p9aMKIth+JrsKXjlOnONxFwDalk+HG8JG3153ZCD7
Ad4CFuUfZ7wcA9CYc074gaKLxv+zxePDECbudL1MM7lZ6IsQ9zS5NKUKUgaOMm3yt30066wJrNvI
S/giTP9z04UBZwYweiNZLYN/niLullzEK/YwhvFKPySe4yXBMSNmj8RwI+AgMJDZ7ROwvmFOvisX
/EVxw5h7AsaF1zKdYfPZ9LKgsK00diGxIHqrF5sbNncKFIxFzmp4MHR6SKIX7yWynCIJGHfPEkfw
BpxZT7bChBo3mPIHapkio4v68SevWKB6tOM8JvcB5ELiPVyj1vyqMRMN9Z4/thzdJhPbDCZqTlcC
BARfo502NyNSjniyo/rLYXIxRTRoG2KFq+VfGSH8qyJIh2Ok9KmQI/9GDZy7zxlbO2qmGYloTUxq
F0bTTDocjfnObNseEN8QhINjEgIucMBf/sfwBRqqz3pF1dfcCtrbljoUNVDahv7UoWLZhyz8zwdY
kkX+poh1MJqJtxcWhg1kQWo2z7MGHOBVwZIKGjKG9RZUZC+6+4Gy7X0eQ8IzW97aP0mIxweQ+cy9
fC+LWtIrrgQ5q/L4WWPF/i37PssHeb81IBV0pGNgc47TT5CbvJgmXfR0H2ORON9maJoMpgrgtIcX
4PGVcl4ytPc15jdrQ+JUv2wfczWAsQ4a2yz/ZHW1v4+Lbk0+9DlrvRi3lU4GFvAoSTSTbFfnMWDa
zvk9cwG1nqEXtiJNpX1VIZlvcYirU2I0GvAi9Ql1niE3598FPRkr/+OddTKgxN9ubQeTVBpl/CKm
9yyVGAbVbMawPmk4ucTgTe4+8Ua4QeekPDF2GmeWTuG7qX68jQ3bNQg5HbQRt+6UDaDcONf522Mj
v/BVKXZ5/dYIW/yod8wo9W1jqQPLEE86ONMrMViHCWWbwmKAW9HJPxAcIrU2Z/x4UnFooYD7xx3W
r+IfDPJngxNLAEiCHQ4W3+IPt+cjbjfqqqYbEYZpSm52KEHs+fijPHk8N9ufYNPJF2rBU7/3Zhkt
Oh9GD0GsjqK9wBo0xmvbwKjknIgrWIskJxE/ciaP4aPEope7haRFEWcK+W3/3yPR+A1FtjDY5YZb
LefFnaxfXn1BXTn3oZRmDK5blpNe/R3sSOSz9RmN0ESI3oHE1SS2TA3LEYGgI88Fh+2+gxsB/z/l
ninqiN8RuA3DgjybheFegCIlG66LOEqbIDz+zg49hCzaRh4pcLCYSa8wwo1tgr5R+duQALPM3I1q
BVE6aXa57K3XqLqjw6uqrNC+O4nU9s1LSI4S1jVPyXjzJxrOJP5h/55uBvmhSV1Aerqjm3tg8om7
WtlOuAaB6z2V/8REuLR6r0mtvh52URo9A0b1jUEKrRxJ7n2iBr/hdjmSdSb6qRZKSJdJOK/AyBVQ
Cxi/G31NKrXTpfh7dbNMaVuQLZIA5hHc0f/jHuChWTGowio0HEFpwlPlBPWe76Cq8Te7vCm8fhru
l8JNFi8C2LAQdejUshd8q+no/bHSnCQEY5vxM69V7STiUmJJHsMBg7rMgk6exS7WvzOlCCzPeLQ6
2ADvDvJbIoEyllffIxTxMczvGn6IuMdKZ9Wyd8TVpVh2RAlQbc5ZvNfUvJ/HYJXTtL0ENjwcBJVe
h/vX9TpV6jmAqtfo8ApU2m8OLxVjz5NRZQAGkHTmd/wUv+goO2le5Y2FBV+FDQWY0/OHBP6JUA4s
nmTscZbxa8RgGWCUMdpA/CaP1CwbDvgtYaVypVG4xsp2/Bi+LInrmekJpeOWCC2TMxw6P87u4XHk
xdgjaVlm4EAHXMLrDE+bXbHM0QwAEMj/pTIawl0JVckMEMNoJyMfzPkuMLRlTJ3//b98mgBHfChA
NaZXw1D6Vo0xr1Ttnnsz4TroiDopOOOmgu10nNCOObCwcf+yHAMNnObrmXQdQW09Gw4ypC2S1JWB
YYNoxKYvNVzItwJUTIKAHrOnmqKslMm3gyWzMick1U54MFrsYWg2u0d6SP1fAZHj+vHQE9S3Mmud
wgZkS2+VlmrkuGe++kC3oVsEPjfKAugoTdW1OoMmud5p3zlHP3KJqEq4jnCn3fJqOE4YKlI9grQz
VSEUyGjdGee9tjwmYr1U1/DZAevc5faiD/rL3L/LhCRP7JQagl9MBS3JfucujILfysysbVuhNOTV
SGM/ugz+y1I/Dm5aoAk3+G7pWos1NP1imSHFlpSCQPqSnLeW5m+rKAr3vpCE2EakMyXSQRs/jLje
rdemjkOw8IktUaGyViaVHT3kIdMnw4DmPEym3dsyfD24DSLLSKG6gRlDXqiR5qGP7XADCXhj5Emr
LSKIHd7f+QtUa3krUzvZyuJ1S4ic+H10bVrhK5Fty2tGWNAEPvhJTICP2xPPZ8ShryqMh0o+hDD0
BDReYKeIajermumAiclOC0TK5L5yVgBlIRNJ9sF9rDh5vKKf4HF1V027cWDMHGNENLcHQZ6mgj8j
FfQ3W7W/6Yzag2p7MGUksHMvRJ4PpM+nWBIswvCWvxKmYjVf/VHQ8CSZ6IwF9CvMZMFSFHh2GOiv
R2ckrUe0V0exZhHasZnCxL2vr2egnjtm9kvtQZyAChgd/nahahuw5xI2RklHBIi+oOdk/XceX4LC
eubnUHIff1SEKBYErLsGLuceqveADmgeAzg/ANItH+2FOZNv4cJpfyRZ8Wbf6jJ2ZQN6+bx5iiPC
AccAmUzilTUaCXOjgdk7PzMDOupY/O5g0CkFRgkIls1fBamoV2PwHkBoRg5gt6sBI13nmXrBt/NE
FAvyiXniM22/R5tgOoPd9UjkRSTk2jrR+5TBCNFD6rUrcSznNu+kBzryzAWEBCr2oldW1lY3ELE9
REVrO5ftaOx+i8EGs/HvRENRLCjFya/olOX+u9LggupuCNYdaWEWvhNaYKEtSeBAAmv+DGvU06b2
4sXDFI6/p6fDnENZ8Lgx/awC15Bb3XjX8fuP5zIrCB7jx1eqpfBmlD13GRUHHqnnkh9I2U3HKUdw
eAjc7hGloXIIxWrKJjcMELS9G2UFARfRx5am2VqbKXpKa+4MOQUWwo/twtX/+/4G+FngU3/RXpR9
y+cYSt2q6GvQQgkhobQ3B39Lfyi16BPygriW2HbA8OyRoig6lMNWONVi4+jR8XjczKN67sGqXR6Z
KgK1jrw/kdToC6kA3+axhtM13veJgkIdwhWYYJLQ6mri1nUe6C7XEcneJhBKe6Sb3d7a95ev2G34
OO2H5H+EVWQ2WRoQus+noFRSsUdenH/LTczLfJiWKDRgdKdunIZOBgHH4J3PzYK+0r4R7hEKzHuN
41p8pGa4mAg0SPqma5dCaf4Nz7n7SyXc0Q5Tjo5A8XV2aNrSFfdNJmCx0zbXC9IS4wbPaxc3Rle2
VU+wZKSqjdK87h5dEAj6SeZpb+B9wSk0TX1RMo6y/ID2sRjk6B/rB8x/tdCNL6sFxQAAvkxmk5RO
+fKyAAaFaw9LWb1PJcKh8kiQ1qzMCFVlBcuWsY24dDvE9V++cR4511YZQHSfDQYbSIS2TYd57i8+
tPf1gpssvlA5OdKFENZMHJoLt8VrYgD9cyc+dYGM4CwTmYzTH9+vyi+W0Q/GZEq/mQ/Ug+wgrj/k
sUOFK0Gj0RQUpa8500wmW8dfksS3zZjPmBsTiWKRDe9H0Peo/jeOAber12hQk7JMxTISryZJuzxv
dHPwRDnq/wV1LCYJfKpBy6DerLiLHwPh1OKeDJ8AJH3ZoCakBxyD/gRfGaXqfcQTLm6/4zx94AOQ
fxHzi59Cp+oyNXlz2q80uMayC33+gTG7f38y0K1WUXWhNycmPXhh9B9Hxv59kNm32FVpJONVMQvl
4nvyXUgzAAl3yE+z4dgKJEdCDXGhFJsd/PNFJPIagz2BMwaJ0VG4l4+KyuBeMuHBD7/7bNqidH4O
F65Efwmj2yz8q8zAPw12eqEk+7Uaunom0BRwhdzp3VUmpexxN27zRHu1hCzEG1GZ67RWXMKwhJ4W
XHbs0j1f7i1WjWc4eTM4GAmKCZXquK3iaObUbMUhhu+qKfxx8CEnoZ0eRY9TnZeegXS1kcOXtUss
a/iNO6fBHFDpU5yaoZ4A8YJUc4H7A01JaI5Nzrkh+eCHSyA3gh3cLtHWULgC8gGIHNESofdJzElV
p4FwOGebpimdEu0IjZ/zz5x6cp7dp71vIMsdqMtlSKyKD4VrwO8VE4nI6Jt3lLc2HNW6z09Iy3vr
nWTcmEjMJX34LKJcBlHOs7dopajw58BZR5UXybQ3fTlR1Wb0d26n5gxYKc5A1SylXCv7TNytlqMi
7o8Bbh/vx9ln2FinAQTtNloaz9G0/5WNBDHuZiuKVBHQFFNuVoDZlRVp54u7DfDIdkIJPkfC285G
4aIN7Mw69SHVc97Gv8iFMPEFSlpRzT9OY3HwjHDcgwVWZrmeHWzmiFg8HTZOJSdmdLxjfPHYnMRr
l744cFG2xmwjBtjR4g2tnamXB1aJLjLxSm5g8fJmbGqfalg++2WueHv9Mm7JLuYwZVjJYdd+9I4A
wL4nN9+P/7NSi6NTSMg9qzV1lCx7iwXh//abn64TufJi0v7Kuh92JPGqMshSdHDsGRxH5mE/7rdm
FsvR9OBCnrd5wFgozSPD5mAIK9zgAPHtXTySC3lIRXMdL1Gr97alnbeV3/5jpjneOyhXBjpFnQG1
skLVQNEnj7TlBct2D+fodN8z7GxALATr05aAL2g04MtJM6hzkOkY4QwRsHo73130dS5HQpFqckOG
86ohdX5Nzqf0Jp81+aWVtE/BY/pVm8JpHHjxzuDLkYciA7PhYz9450N8MwE8+YJev7fZ/zB7LJqo
Zi3AnLO0vnnlGf8D555f8o83zw6woj0rvDfkKBMYVcQPfOuiZzoogSENGZiH6V0VUtILLUCqL/CG
JrF5v+ZERnBT0A051zgTnxoiMgjmkG2eAn/sjkuLtdBJ8ou9vE/E2n7ebk0y73rQ5EIK4tHIVNak
SPLdNQpp+9HjeyaZPwW4OvgJGOC/xRUC1aIYQYfjd/B+04S6BvmCAZejikhYI9oHWG9xMKQGdWgK
I2rU4a3/qClaH/7v2I83Z/n33l8/dSmCosk49rG3JSKDVrC242lD7qbb66NRSW79ZszkJCaTsSpp
i2iJIRBS+QbMViygFLtuOpJGRqxdRfyOaSp3Nfu+rM3M5iihQzqwefkTx9TXPzma6Th2ltJw69Yv
8ij9NYO4AcDR6i0ov2ZYwZHBW8WMwxkRe3jp6v/MlHkK+hfPyt+sK/KylRpQdKX61iWPVkqcQFf3
FZBsiXbq797DftmVbtgrh6yp6asgmeBp2OIW6o05+jh39yYsjjetC5qYjR11quGuK9AdOBc/0D2q
Dc1aLRudI4KfxNy/X2yLZc0NbXz4x3PfvXAD4bQumQ6lMySJXggTNBt27D3GHoVZVPRdPEIk1bnL
6AWClb2aUr13w50s/BwI/+BhwdFEWqYV3zrFBd/cjNvCb8BfvgBo5yaSuyDliQy0V4SwOvfeAMFb
3g33OplQoiSsxOkhzZ6ndIOa7hgoOyJjEKBpPp10TqCC3qNl+IVbgiZ96Qm6Ug3E5g9CJl5+Kdkg
pIHrWERvxn+9HUFODxnUu5Js57FKnl/33lKWP/7Pd4j9J8E1LJQdBtlC3FW9yNHgtO108955bMWU
V2gqkZte5i/fWT0o6QT6m3pCSgylyfG5KZyTqtWn/yQYxmabzr77TBbfl2fl8JSFz2bQCiNHH33s
T20A6nRqPd1GREDMB8MEbXsg39rWq4Ei9RNOJutQQJu1u6pMdRXs7K0xaFwDbvwFKGrtnf3DVfYS
rrxiFcyTUaM0xMnFeNvIPmh8EhH9yuF2lTqPZZlEEK/IX/EbYBwSA/entTicvAoZ3dBOVS/AuL/e
n5h/TCbA6ytpb17vaj7m3ZtkOxk9MB7Fn9TE6HLqe8os58Pe9XVqsbPy+Q4bjBPHCOHpZdexgHaK
q11W4hMzqwF4eOky29GguaE1m7sb3ukjQNC1MsYRqMfwxoL251Gos/Wl4trVRoz+X8v7zR3XxlTU
NqZECzJOxtUQPMahl43puNkgXVtCz0xyWEoI9cvnRkERLD4oevMyPe2kbmfHGfgk7ab/FVfp6sr/
iqd/H1z2Mji4Auh2SAzvttl5ZuzJcqHvbqo4EGC5ybhgGo1Qg0R8ugRyCcpL5v7H0R3XN2L25NN/
kGhScMS6VZIC7L6srAYznL9uHdwFF/DTzlJ9pfS+4kDgWH3rexiQKkHIOI1LfFhbZu9OdpS1FzKA
MuSEJ7AN4ZkMkyPxo/ItoApunt0wv5TVpnbKxtFJAL8r5nEBrm3yxdUbLB9ObsAmpw/2+lGGHXY3
JBB2g56NatotCVXiQPrlqyHJut/ekOgDEe3kxT64EY9Efe4NOxGK96Mb77kNegKP7kLAaW3uHkS+
skq+/rH44qo37h00dgMlxRGM6JzGjUkUuGMZydqgJ2ohXKXvlkcXlZG5mHAg6TgGH5CInmQPYiQg
RUteX5a/0yn8r9dcTfmGJZIMypUKINR0v3nv0NtgRF5kZBWpfmPEIhguFHrtDZHCf04QISvm9Z0C
0/qfOk5RNBDFGLPadbNP8hwmKrb2prCZeG+DSb7yJdrHz6HKlZjZ/ZLe0G07naEK8huK4qMBf3GT
wRiNHqP6bCnCDHEl1Mxbup1OhzV0W8bx1mlGUOPNoqgprcBx475IIz9szyh8sDnR3TcZLWv+yIi3
QS5KTQat5q92nqgKhmMEblNi4Qn0gVO+tJFnCKtqLTdEwV7pYbaUfs6f0ZWldKtukz3oklbFKbxI
EI4jqXaoYZ5y3QNH1+5ja2tIwHkGz+b1pNqJ2xo+dyokd33X1XynAd7pt9tYtH0+DRLvgSetxFQT
KGkw2tIrCrTp2yBIhP9M1txEUTn7HJWWL8DTOnPfwlWssUOcECKixr1BqtHIsAgjHSwWWHD/T6Tg
rgEKRaZQ35AupcM4DDYulDh3F2/K9ZmxrOMCnE5VathNfuVYrRhFbI8JutKwtE/6M0Wde6ECqaxZ
WvnLHYUEkXZN9rNpxB/kpyI0v4j41wNdq6P5POmMfRoJFNfOlIUYGdwI4+0T1IIhKg8KwTCmlX1f
j1Rt9HBG8s/uxUIEa/mJn1fhNA1KnTXQZ8TB0gTaYhPhuKvdIDzsqII0rxvjSPLl3in0/EnkdYEm
qhPunNUzt2QpmMS30MmKejCcoDn0LnDyPEGCSEVJ5dgOiQgdagfefMvI4vFlG7gpG74/csN90RLR
HtrvGCnRoRe5exs6vEHUEHux7sqUHjVcOsAWYJO5vC3OJKPXRe4UEAzb0lk2Dmp1vCB7S6xsKMZc
lJ+9wSPqkrMpD/YRDHcjj154ZsgYFyoMivE/HdkKtc1EZS+AnCTQiudqdOaa96319TNMTED6T9t4
M1LetTFg0f9RA66DT2L2I2RSvRlFca8gLGCJ1vmKwn52PVvytnppJ50AbeYJjk/JpsB4AjhQjpKD
2VdIOCqr1r5JKcSJVbSaCJzJRssKat1FxtcvZOdkhPBeUa2Mbxm5XBkceGS9hYF/9UzQ1RD8Ykpd
NKN0mR3m56mj1KLgKSbEybHN2W1pZQ/cGHWJLTIocIDYZUO/AZkpt8zIQI8cC6Y/KuJRcMoiQVGZ
0osmcS6DNvuoVawwag62z8O5bBKRHc58STxTAhPJdbEXGy4bPG33ZIMgy87LgWCSxu5o1kx8lJk0
pGs2D7qgugOBKRpOXyCZDC657K4FNuSwg9ZH6l0tH3ZLmhn5n6RgY5RGBQwDlXdePoXTM7hukwSW
DZS4JLZKbA14rXAnyt3sE0qWQZTwaU1bvgoRjXusl1QLLTrcZ9iudhxornKYvINstrgCbVz7vsNM
4qXR7pf5Hd++ygHnGygq1X3dqbZdKfDbf8I32rocfQ5p4A02TPnzun4Mz0m8Q+vhNN2OZsM/jhuy
ebdgyT/uLA9o+ZycG2B6/N9NlfF5if/Eke+XsVw8Kzqin18tT9sbtCEyWom5I/Nj94cafCuXzANl
UpGL/EbdsJjX/UM6cIRXkHZWA0tLzJVnrgl7P85xC/9vS1qhl46CtODzd7zGrZ1briQXDni4/i1o
j9pgfj2dkJwRzq3RV1EQEV8LftloxFJCCbG+ljIFCGthqAXAID8YFaHxXkPE48PchL3yJdCCXsow
oAN0ja0qN6jAoJgHbE4rWY/9nuIZeZD33/tP4IjNF4OtJ/8abYayGftPw1vsqR0ExIkIc18w5kgA
7xLSMGbCa32nYDR2M2CmyhD2qR1GXV0aEjouso2t/m1U+OrzUq5ZTN4fAljINfhroZ4aLepGGBog
KQ9E5n+UkbJUwgpk/01jiEpJqB1W/oYLThNiLbkgVnfrRUZ9SW+Y7Mz8wJkPQE15u6SlG/quO6Xl
F+NcDXGdfcOcwg5b5GW+dIWMsXFboycwj4UpZX0AI7CsqoCwRT09V2MMhDdaf3A+W8lYyfEtC3jR
GpyDddznW1l/yijuawIvEf0FCn7Yow4EReiQ1th9sLnuLjGk3Pq8sXKZ4zc97T+1PL8zv0TnGl16
VJkPXRBb5nNQJbncLqdVadh6UmpRZp/3QkdFCXn38FoH3o7ZdFdYatVVi7JdSNx06uUAvjVh+yaw
2zmMW89NXk7a40myREihfIzoxLLBl1V0F0Y0mYmMPRCfGVRAjCNbph6LCu6rx+keVqyVp/0bxBeh
IQpbSn+hobjRbUqGvqcTyqnlx/Vl838XYQ+xR7xnZ3Ej83eoGJ4yJjMuKJ2IsL9IkPde2LiSywJ0
97xa031HjbWjTV4y9ihYjez6nz1PfFt+SczJ+wO+fPXO8Mj3Xnfatxxx6ACq436ElqKod5UZieRQ
FriZ5S7enOw/q0I3EAOrYLGBAGJXeHounLK1texK3Xadu5cT6WfWSdCBtuh9f+johGMQRTpBMfOl
Fp5PtVqDzi9jS6Tn8QzHPgv4wNLT4OPfhB8ODX+r5GglSdlcwltyZHxhT7Afvsh/Ui2qaJz9LhpI
Sem5GmxNFVbzYSyX2sJj+J6HXhf/QnswUls+O81Utr1PyDvYYBmoQe4OVuXEXGEv2OfYDlzcEWqM
+vs3I+v6Q9rp5yTHWHjFghAZXF2xtmCp9T61XLnRQ/Q4Sblz1R/AaCuzDdfJun476IBsfaSdxHD9
KnPNezLOV4l6cN0gO/c2IdPGFOt9No+ARLj6TyZjMBGt9Uh+Kw4RAt/hTmHOPQCGfIdb2E5PJYA4
HutdzYhWGMi31QcSqkAlWY8JGbStSbrvZuIVzBipFL39gReXyF3H4xBeEWjHIwx51F1f25dx+Nlo
p6DBBSZ3uXMIOZso3cz4zllFORCG1m0A9uDUUEVENnzxkQWzRW/4tF3txVj3WyMY4pWQmo67m1kr
5VfwqpL7SnJBPkvXND5lG1BeEihwD0g4XLeuoOL9d8k6R4vCLL3aI/NIcuqeIiNSAQHlscHszPq9
C8dYc+dW6Tj8cUg3OOyj+y49ot292wjg3tpe/Yd+h+o2aftnwhnhTxVgoBFng/0mIScMwaGG25+W
mSVOwN5zMW+8FmiqhRDLkSDYULQ5eqrWzjf3K0mk44Aag5oCPhWWQWTn2Cui6Aab3/cA2fVxjY9N
wzELMEhSMMqNc0bcG33b5dS8HI44sJVmLRc1Gxhwv3kuIw+2yN7UmxlZ7eUKugCq3pMiR/Mov9pe
iC3AF9LDf/Rgzh8pHCwWvXVpfGA36cUOpwhuVOkCM7O8rhy52Gkec2PQioVYejSBBTcz3/3a3bLM
+1jDkAWkVUpou2N39OBQyRoTPU7KGnoeqpMyNSlvJUzSvBLDOdt59zAvvvjYIgCxVBtyISdBv/9i
Px8kyVKLnhJVoFs+qW8dp03ntCDEGKLNwiUkuMvaT9P8MLM7f2o/9fqOt9lf1ya9nHKnygYZmkz8
3gxdtcZW9xySMXgqGasYIxw9Q1uX1pI03Kzu8mlVxSaWOFgXeEsnsKPRA8tQYY8WgXFypwab53Qx
kdEtV8Wmfzao9tq0es5idC93decB41HIveoryNuRWTLhXwO4V27VhWMtOUaRN49Hd6gYmr/hac7J
V0cVkD6ufUqos1ClQK8pFajRXX2OJDLsjkjaa/3h5Lrw25cDlMW3Z7h98x9bGBeKxeBl83ukL5KH
8NMTlbn7PVFa0jd6HgWNb2JkR+d4KBaJj7vcacpIELno5npuzAsnmCvPE/1PIkfQj3lnxdr4O+tY
TtWwKXUE1iihTGJ4/hQWjGqrS3w8REV+YpOAvh2d955B5Gb1/gJ3Zphyu0zO20rvhyB5kPfsefAU
8MH52iNCdZE+Q/T+VDQAVKR0inH6y+FLtKPJEaxW+1AK0xGuhK9OXnm098Os4zPkW1SZ8aZyAvh/
Hdzz8kxeWWdMSnTd6MMuGDpGVzNjKcKOLFaFgqCRsDw9Val0EjeI9K1iMeFxuWwoqRHFNKePPFUQ
OERVXWBJpevyMbzIA0Hs5nAbjDozHX9ASAUEGPeqnT3Om1ln8qOJGp5wpa/1/V/84c8lDYIzytZC
mnoVK+oTFYyg7cNlQrLiWg0omhXYBXVhARYk5zOO0rCs4T/b+gFvmXHi2biaZOXwymjIn2Pr0SPa
qtau5bQiHX9upW0KI0LEQXy1PmXrUaZRjqtOMjVboG6yuNS6Xu7Z2W/vLguxG7EM/9V2JaJNRI2a
zNVV8X+P5250j3M3g0GZI4HcuZxKhkzuBtHbZCdvtjHq8/wrR7/1M3CozrdcwXWQRz3vQjg/FScY
3cfFGhvsUv3QgNGar4mVXstWgyOGDW2dcG2Qh/h0kut6phzlUVGsdhTWqKL37Eu9j268IqJ6vrJW
W77ZyPjiBfHvW+glvWv2gI6ruJgFRkb1TtqFsbVF3CDLZ/WKt3zRfvgvLuQbk+5vSRfeSgEl6O+5
owJoXNYoBNIK5N2m7sY9KaqCpLoD8dV5d9thY9vE6GxwzP0UR7GWtjTVDvN5ZUurKsKXgIaRVJC3
zL5enE8l1EQoke9LZwPJAvqJs2NAlIMmylnHijR/GG8KgzLmR6mysOFTHy3wJOJxBHp7tbGs0sJs
h/qwCcHHVVil3TRRhkgxYALURBWyYTpoUD/Z9X0HasZNsNVry3SiXS2YTt4s3AdXxgNWCQfe403Z
PCZd9O3ZN/oTJnOe3eZpaz3jyHVX39fny182x6BzGZWHIwHFw9Zm8DtiY1DFtw4Y9jFjJnP76ARx
/Xy+eHlhRR7GtvG7rAzATSXGsYSLoCy87EF7vFDVU0MRPYDPi/NmR3NXzYpFX5ocsZbljJ9oTpA3
oqiF/MU9NCjG6/cjILXfcKyLtkE1+NHVtzSqf3s3RQDsTOOlsbq7wNEIOROYj7wl4ssRewYCdZkC
R3hZgM0FIlHdowQwhX1+m3A37O8TTZ2aYU9/foQrJgNHewzuLA5C2nc4M4ldV8BJ8ny07iM9pgrI
ItJ/iadXwGJAL0uAxyAc67VIh87fWoMDoNSfoCsxRuaoCYImhXR4HsoMEdvkKOUW/1tkLyYjUKpe
67gROldgThSJKZN72hwO/iesR3Z1djyrWTvWaaJq2e3A0GHIV/43RYjyy3blK3dxMQiLy4vjYlGa
7vRRr5+DqKTTlCdecUQwKq+j6lp7AUZ2BKu6rLTyfRWEbK4CHPjq77a67O03tKprUMngSTrn67Bi
oNPKYz44g/WkmDJyZfrl4bVfovFgKNqeUf2orkSqFLxQCdwUVYW9vM48QxWwLVzkCTzfSAJyv8yX
amsl91jEl4nlSIcgn2g1O7lWAFGZuVNIvRjSt3ecUy2kKmJtnzeKQTvfKMGR4PZoXp+MatNcFch6
OIZTJu+NCqn2nRXf96IWZwwfBZXLc5j81C33h7Xg2jiBRIqN+5+N5won7/8vB1N1LKfII3+ujPLl
dPEjR3A/iq+rKJFIuKwiMPDYGZ+O1kJz7owvg31wfyrB0Zgsoz2Z+kWNGPhbDFvayErwM2LONjuA
CpA8xT1eRRhODhI09ZyJF2zX8EeTtrqe/jVPjvpieLOcdgcuoloDN4EX9H5FFmfiHY1Ez/6mgoCG
PJYX+EnXi9YsV4LfRYtnwwOrFjjOEszi/Jrnl7K8CNpRsOFjo0MT1y04crc4kQ+EEUCvMADx0wa/
LST4Ut3BnouSBE5Tsz9q+ON4H5Q5R7Q43QG8woYhbQxOqU4vV0PYmMX4thSHm63YHNKyMDjwTYz5
qIccLYX41HS1Y1myOMF+eCVwIdWRsoO2vY1MH3Yk23kUjJaFz4CH7dY0ZXpVXDMgu/AM1AraHiKQ
DBMmZDePPOByz7iSMOkVvsVqjK0ZSimFK1sBcn++d2kCU0Pg7zp88PtRWpuzl/ISJirXY/fErWUm
u5R7B0FRoP2eGKJlxB7P7AtXxmTeQQMGPph5VDmjTn4vsS9Sp8EtD4TFNbbjb2mrsr7k0WxXj2nb
WizXevwwba1sxvm/mQsOWyBuI27cxmOtFVvuJ8oUu1AN3ou+mMBJl/4yCh7vIPnPqgSshf3w8GS8
4+j7FVC/VGsHIyEoisdIc5Rqkp0EweuFXUrrlEuCph57h6iho5BeFB8A11L1GogsUp27XQv3hxzu
zT/k86PSuRfd2/pXH/JExJTKNkS2s8B7LdkUpISlKYwjTl3VhkzgiGqS8nojHbTa0OKiGnJbzon3
7Q3kXcnEmFl72JYKYJBPPlg4fSoQ8LgkrrcpFkQhZnSquMXH1jq7+2p02yvRQCYHHmkau/CnYeQy
MQu92eV1ut6xOs99o0TjrRDykFX7PgdOYkJA9UjbXZh2C1DB9lgJztCyW79V6NzUYYAsdLCJsg3m
Gb2nluTmVCNbZG67Nxi9R7phLfyojXjR5zhncNW2R5oZOZRh5Gu+OkxbtQAZHqP51R0L5kEx9h+D
DLgU8Lh2QqvKkZevpz/wmxCIP78mkQR+U4Qdt3gWdaQS5IH+0cm/j9k3nywtkyrud+Dj0QexmZGG
JcPLfK4lAxmRJ6VH+1pDu8MCLndRmBsvyKsMUypF/s5BB1rlIPMYJwp8vN1woyb02g1xTnWLoP+C
qvrLQK4I9KZ75FsQvlTziFpqLtxpoGTt8Lcj/uteQxoAQbQRpXTCKUQe3BaUIHz8LshkuWqZdPaN
hDamCyKfpLPgQVSRqyyt7g4pOfXKHg2OIIKSV5k40az3SMykp9tFR94F5iqEPW1niEt0vK/w99Kr
/fZiRz+WPhorwp/HNsOnCZ+EOLfB60XYKjdNyfV+G/ayfslCkyeJGb54UnXYhryKs5QssSbuVywI
5tiFFJsX7CjiOxf1odAj3bTlPfC5bQwawdM9NA4DAdvR5zEnfFjopZCeTjaf2WmfDdr7AaYOaIwm
bQFNXdn618Ra4ZpRkr3uGnbPPAEI+486Ahwc2YCGVpUE9s1HqnIZMDLozDqlhrb+aQCr4HB8myoL
bIuzdPPLY0hujU2L68Kx0ni3WP0/qvEpiO7T+igNviqteKXJZSpCTB50aDw79N6ad8KqQ753yzY5
ZM2u+1yKhFmqPF+SfL0ACNzgubm39/UlX9yvhYmZDAuVy8Q3rMClKpN2343hhKK3iZ8MH9izvTPB
705DrhBfN2l9W+Ay6cpQSh/nd4kuPRXw+L5BYHboLGurONgKcNLNi1XEKkfadABtDzFf+FoTffwZ
nUa53J7J/pqO4ojryr4/sd/2KgtlPEz/fU2fJVgR7nwGMagnng1CIznlNrehyr32a4JY+P9RbTnx
+S8GXDWAsac2c9wb+lmEytfLXjWBsxqAo4doDEtjYbNjeB8VuIWhQHRMjTGsxnpJuZqIyc8HOLlV
ECWM+CUAm6MuHFmYvfF/5JRMR7iiuUx/b8526/NfvXxoCIuIXo0INrAK4NOB7QgYjjZ+5ZiVW+NR
mPRw1ilYg1YmcKS60rg5DnsrZtz61d+WSGIVNE/j84j6WvkeRRlX/8ebonDO6T/847jaeitmyP2n
SifdlgkjpuB7ACW/kaNyvr5w4SNR4LmxBfbohK4p8LaismGFjbYjNEyLBcqh7QQTmjo7Ko9wZGjA
Pj2cICKax/z6xWbc0oNYiXx1As5IcNDlpooV2BAgMe06RuswJPboxxQkMEkJbr3AoxM8vH67RQ3w
oeMGXcLecC/nhhsP5ABdPzaeUEPP4GtI4vJmWM3LPGeG+9UuOhTQhTJoN625YlDNK6lc18NbIKZy
aP/YKg3OX2tYTVKabaUAXFn65p4Z0viYtSW8peC8yVGgeaju0mrxCfI+hRIVZGU8E9ohKlSQcNMr
WhofAOs60YcHSyn6PmIEYKYU8TrJA798dJIpt/tXWJr2wvthwDd/Zh8fO3KpdXjMgwAgAi7vxdFA
0XI47SFnG0BQPt23u4WOhXfjFVcTxwvzOXsw1AMczP9plROYbCN6kkPfKkhsVxadJN6cBoYnxgbu
O/K1lLFtclGLqQcVB1j2MVqwm6yzXJa498ckmgisA54krV4ZWhqR7Y9hI3Gv+NAmlRiW7jXO8EAk
/F4msk6LWUpIZhiQp2xR5K/t9B5+ECnGEvf1pNROR7ajb5pKA8FPrrrzavoxeqJdoVL/AYmVzp+5
fX24XfztchngTzgeoWsr6H9Uy4hYWpXa5SdblJ3UEnyIXGcWpsF0PahI9EbWqge9BadntY2fqHXI
5LTg7yE/1YnKw9Ujevh8+8RiOPf6snyMH5Eki/l4UMQOkZvtXCzvUkSFT0R7MHHKLrbRjwxUWAhb
Hf1J09h5LhZZK4UkcA6dOntwT+DxALtVjvPygDG9ZvjBukYtC/ccYzewMLMWqEOjo6vcU3A/IGC0
zXrjRr00Lkv6S77zZcWlG4cpgv7+Pelie8grovTlfxxxAf2Flxv52grMRmjsPQEmlJOkve3vr+aw
4kD5KGFvfgrbcXtpSIPvGQIzYzh9rxHAkjQ0T0JG99xUysRTSNLg7mXtJOq6pcLLCtrL5+VDkDRB
+uCkn3Q6frrpfqqWNJSq2TM43vDYp8t3bobbMRk3oA3/1t1h6ZRvDU6NifjtT0SK3aBGubxcHXu0
ZV1fZbqjZyJMbJzMiWLfoQ208TPFqcHArGitZEUmAduinVgB08bjuboADRnkARIDEM5qSuXudeIM
bc43dPj37DimrOb1FP+um2mFip1QkCHk7RYVt8NDl8Xc34HvLMNbtbkqMzVqE89gx2i4irCstEhm
ljUxUyBAvTgQZivDBdIS9wr7JfDkaQgL2OqlEUXubbaP2tdtluT+PDDHzDjngWPLA24sSBOhjLN5
aAQgWYMj5y66KCtSYG954+k/gzsMB2vc1hqq1KHtV7XTW+SdGmCtzyZnXMj0yn1kSbXWwcejh3yB
EOeNWMk060PMNrcKKMGHiFzTPf74gEdw9P/m011P8D7WewVnYcDSQ6DXqWc8W1XLiNiyoY3Fzsxi
3eHN3L1Ya3pFfW77IRXHriE7Y4AgT/lqr3AVuQCoAZJIQd8SOTktrpPkVCYna4Khr4IXbEWj6aNj
FEq3falrq5tW+h0+j1YQMc4JUUFHjkUEZPJ71FI+nf7JprLLZGlPsYpJIyNJrLa5dtxVVC3dyDIn
Mo0cAY2K3jFkvkqa27hDDngK67HQZiKbw/6j3bUPD2jKdQPssTx14YLFQp2xptB1AnYEGcfYFMSZ
OgmYvHN3oTPKJ3vaFp7loSUqeTNH05ZLEyEWuQSN8+z63fNaoebee8KubccTR8gVqO2HFjOTUBNc
SrF4QF5tioLtL7gwfyW9ySMOxIfXWx+/uXGGJhG46NHQUcLegPHfjQQTXTQpM8frXnGIlGTipyRH
IgKfkHVWirsAQ4Tq8LZ+/mLc5WwejHfBzb9EmA/yP9ZLH8htM574ff323Ejb9cO6V/wtLdvX3u6Y
844ObDK0JTgAdOficLriMJCyWJZTCDzKEpyfR7d2LOlpS5QsCP9w424mq67WmRQg76nzTBdkvg79
4uPjXFbWje7NlAQnKu/uK8m9M21bDEQEZ6H9hatI9tJl1ZPiBo+41oEanrj1gPXzbQVBxhzM6+70
tInPzRijegcV25HdwavCJeDpz/AZoEWBihS/+F9X3l61xgCLB73W0ouAszppU+2QROQeQmt4xq6V
cMX0bFOjYRLE2BPevZcN4ZYtrxctW53gMc6iHG14pcalLBKRkePuDvxMT+oPD20XDVOWUSHrWz5w
g0L+m3ikJg+XuP+Lz2XS2AaArzgv+GJ86ieUqt+vwVKvF1nrN4y9Zv7IdfOEWcsrdxOA5HoKskwo
u3k1SzbwS5d2d3D3zvLl2z/YyBxq7uXubBn0mZA252IVIyFpnUphMfrzkf2sMa5s5FvPQn5mtmCQ
zXSoRkIpZs9EH0Yti+VP8ydBhKj1ja5jUAxAlzjqzd+3lBrfwx0e4NpQGUVqt/NxtKpDz9tpTrMA
H71xYFiBf/Ms9TV9YZcLyGiXl+Tc8N+n/hJWfxFMEii0wl6NS7kB/2nKvLC49XqdRaw/lLbcRrnh
rDEfZqFIeIOnQgXG36zqbMidDRSczi92e37ZjKfpGHM7eoeRwJBdyoEMW6sQO29xnYKc5NEdjlc3
vqsYtWveDqmVfQD0D73CVUckTOtKfKgNDuEXTB3F+qOwoSBvfW2M8sbZqNUkr60AuhAOVg5avi6/
CS+nyIizdR7np0Q4GqxI5jhFPECLLiEY2Xs+yRstrozEafdcpAiHgpa1Da4Qf+zIIyIqlI45kaBF
cSVkWITL/ZTFat9IBCetTO6416dqLseHP6nShdiBzGKS9RIhGm4FZc3BDksh6Or2FPQQh25jRIVw
3kaNQtV/lseRZvnDDHdqHj5wLqBZwmHBe/iyNSaPdAhk2QF7usIgiseV56Fl8X9rHQqk46cTYB6o
WxG9F3t+gakuUo9GIVQNqqLoMjoEWOpppyKu5Q8+u951Z/U3v8haxqXQJSrldNPTAoB4a99HvvDK
hGBhvNHrKHn/FOn54x08whmzFbEk8LxA1f5T+sE1Xhnk1+kbycHq4IhSwy6GBBVAXWYNa2WztdU4
o5lcJO5LgILW1Op25BRFj8dM/xxSx1sBe4KOqUiMeHfKE65qsjbNw2jutOxbf2MOmHXBZjODTiRk
DMff90XQ7Z5GuV23lVMOQyfq5zRjnQYpCPAmd6dJkHsl3Nd10hbCC8Co6bNXeeaLExEsjEKlVg13
KhzK6K2fS8nwm+yia3JY921d9OA4AGb4rZln+Z/kPt4vPtbZop7LTOm/FeZY0aNnkmGTHMz121hp
9twoIvgJrq/h/bR9uhRS+O7DtlgUVWv/sQjiEyCj8AdjTTEwyERqORkSp1qQUkUhl6LhE++h38kS
hlZ1rBvjgonHzt6cFTdwKdpz0lwd+/jWfiEvEXXGbtmlqy82jC6829ES5LlNBF/J9N/GUS93dUFw
r0Hgi0ErDxPl5g8bnB0ZZlOoNPYIBEqybGrlEjfJr9UQJj0EGqh7ZHc5cy42SfrJSgnyLmyN7Q9A
w+CBxZarCcU+U0vrpLeCAgIF06va3OePu8nOyara9b25e1v03CzN0HmUGIQi+js6Nf1No6dIylW1
q8rxDNOMDLZ93vgdoHEDlytXX6f8IBmplpVyhf96Zp+EDjvzuvfsi3qm492eE23hu4VpPjVThxBf
8wtg9H70ctsBCUgal/T34jGIq+8J7RzQRAVW+ZgmKWiaQ7elHZf+XwEEw1GdpbIsfWI5NPRErZ3C
kvpEJg5oM+Q+dtsbHGNQ1Y2RToDdkgFAxD3a9OcXVgoUQiveSOQlPj8ucPY78UJCS/mFxySLxQO0
+UMAUo3CBu5HOw1Cdit9ZYL8yIdgih0dzY3xdghAHOOjq5kPKAqaSOYFiZExwqMduIxxbXAUCVmv
hNtUk0xnl4+3vq/SagtMU1zLj/l28zzFqTzyXz9zmF38iPGzZ4aG79wQWi4GYyaqIQZlZyvsttqk
X2rPqEXXqF4fIuVgmou8gcGBxmx4dqaqUI7MYc93E8cgCU0YdvzTemcbxMsa72MMYnkcHaWJp2WU
LnDQeSlwXGN+rAyFvU270knrs5sLN9k+sYXu+4FtQvkISPFxF/5DFn1oBHChrXeR2yEQO5G9RKcD
jRzbezZMx4LDYKAR3H0Pn/0C7vEgz6pjxW/gTTZwHX3L2LAo6aPQ8pIRvxy1GDmFQPXOE5fPOx7c
C9/PnqfVDf47Z+jlAGcILaWrCIZp4Z/SoRWKZrgFKSRgkFWscBmEwsXJbEI5xjcxvMJTEXOLo9hc
7Wlql242lAFQXUeztBCGTUaM7n4SO+vJuFhNMd6UUOzEBPb+o5dBqZxS2VuxHsJdB62HHAar6D+b
WDAgZlz//4ew+zaKYeVPARUA5phUWgOupfJ2D+gFl5LWlxqL6G0INOJjr4HQIZ3veEQtvw56YgPN
DJp7P3xAILbqQsBgAJ8GwZLzWn3nOxKtnMacAVD73ScPHDVNxrWb/dlXSYZ5Kk8xpAMawDQ/GXas
uPyy0W08dL1el/oE7yA+6nPvusQn4t9mvuawaFRNkdGHRwJS4VTD2iU1X54l/BT0P/J5ZXccfn7h
eeenzHtP4oTyaIx1vmzw9JxC3jzWqsS92HQHiUG4VnH7QE/aM4ZXAe/oHfIxUt/LgLkGnPknJVO5
DowmTZ0JgpNjt6Je/owI/KPC2p3yTeePfrmgFuo8DdVKa0X33j2vsIEUE5BrivpEjlZqDKQZMl/W
IwSfbL3f/fI6sM5L1WsJdvMcqmViL28JmAZH1wbaqi9E/LouMaKagiogfMyiiRNmAykdK03tqxSM
6uaem0VR167asfWiauGZTLmveYR2ROYWO832rUc2h6u0aJI+m8DKfXi1H7qQu2XU7tunuubzSPn0
0z7quoCaa6F4kh3COwurSGGszkJrQ4og/hxlmHj6Vxrgl9qUoImgXUSrde/91HYmDttEsqDLl3Eu
786RG5i9e3NIQGXrnzzbWPk5Xi3GrXJZJepXxKmZ5DMdOwt9skOkeBx+XkZmCLByxiVg6ka8X3z8
SwbCibZ6RWEclzOQY5RVnj7JlJnc5zQWT3yjsTtZc6+iTrWAt+oxDMZORmEqpcvM8AIye5LrY89b
WIH1nZlNu/UU0FfxGdMdqsiTYXig62WIh5y6mlDqNimcMjWBRuAkRt0ydU3Rpxfh9h84eVGlkLXP
yNjVR1Z8FnumUPmqysLbtIJ54Ax5T6joYdK5C8NiiWFhmGZcbO5CRAIgfn0qDWo2J8/BgIh/69IY
hLeiAq69lUxCQBmHs7RsNXzvfAbIii3rsZn9ZARDA8crZUHDz5qvgb0jli48BkO5Vtefsaz8P1JE
xJNCkWvqp5fkPuBKlIp6zluue31+lDMR5NrGjrKxZYwtk07tfdbZakrdCDzQKO5yopyS9HEYBVRS
CI0/oiHWSla9dsAuyt9+2AG4RRutjBSMWf84lP3ebMzaUsXIhiAqfkls7CKksqlWW2z9DQmEgtHz
NW7fZVi5BM9orDG0bGdPsgkUJbL/VoSP+Up3ppxq98mAnoqBaKOgJ5PrBvfBPzi0nLQjq2gWwQ8U
ahkLIcKA3X0Qbirv3lSdWNYVFm8DK1gopxDfl7E3zffjNOApzU3+Kl/2SpYjH7gje+5o+BS4H8Ca
9un1lJBiKU7tHRKjthb9d8SgyCLhUskx3LP4H9RZvBaOSQJGc4xX+xRPLXJLYo1iv5RTLToyiLYd
/nElrY7fAc4DsApiKzew7Ci8LgVe11BL0g/F9WZO3YrEWXUXN39w7bFzv9Y05ZSJHxrs1Rj+mhKS
Jz9Y89EGTXmdxJqjTvXp4yr6ouv1thmMMBnYnghR3R+5QMmFG95X3kBtuTPbZI+LGZpD89YOGgst
ImXNKtz0VCI0SWsfShxZEdBwSzJH/Hqnr38J1FMGcgKxs+97VzrDy8b1buUA3GaPwyeOQu+UYoyb
ojVaEvK84cJxc+QMQgkthXNQ4HCRMnLXgGSpvNmZEKaAE7toLBq43gnP9wVKNC+scxnjs4vWx13Z
OHT5QCSwrYB0DUmbQee/WpsILwKvjXrtgeYmKeQHdGmxj4lW1R95VRCM6ZFoI6xUSy8hRVaWxQDP
722bqlrgTYsf/cTBnhl87P0S1EQlPKNhgZhyjgNfzpaSiCZ2vhvBINHSxZl/D8TfdPLfiXrHDF4G
5sAoLh+0FciAvzkJFsVe1Yv86PYMG1UluKnI9xOmip1NjV73m7UHGHnLt3D1K7vnV301K+HqlHKf
3+GR2iQSrYUy2S7dElc10xwDCxN150IDhkD8f28863ddmFG/Ly3+PJl6f/bHmR3k8OOiic3is8Nz
gT5RRz/ZBx8zR9L8Rx9QGVL3QTe/iHhyzV/hsx8Jhr0W7AvJrABXXw7ZqjwR2X77xaqXlFSuRnfv
kJ4QhPLAO4182zNHoq459TUhWhZVVS8X5ErfidNkPWmfxvVTLfXLVEKsxjI4VoUQiFL3FXvOnppy
P6qp+xjgLls8uosZosyzjqh3ejmJSKtRIGSc5Wpxnakyywvc/U6bOlHgO7CroiN13YajcQ8QKLSk
k2zKSoP9xIP0dilY3NOe3e0VCrgr+FFnNft2i/DyJ0Gwy4pVmJQdsSc2wQSJ+ealcSzvMtOSTjg4
Z4+VKyXEDR7a5SuneoLbzCJ7A/AOH6bZV9T159RuJsSYq7lm6JX6GqtARoruetQ7d1ByY5lKiucz
k4ZhBmn3QEraIri1MRAaOImjPo7MWC91ztDfqddROhH1aGGC2AmF0H5O1xZBmTPSjN9iwFBj0BRf
tsYLh8FBzAPKxP8xN+MdWzOippxQh8uKi66dJZ+FB/GcdrUCd4JT7q6opv6X9B55dJgpeHO9ApBc
ODQj52VJExX5NRvUECIRipwWTnKztYo9War1UI5sPd4BagihAIcUYWPEfwe9zVKVlMyX9DYGlXqJ
RgdJ9zjLmdXtXlx6hf3KsX6FuneI/7J2JXoOewZXd8WEwNTX23NBSfdOgUBEcjR/4zb2QSjp6kxh
SvBbdIpd5+TwkrV2GBi4QGAMwexHNzS5Sn5zxNl5qumPH94v380pE837CHjjMICy1vx1ooF5aEYQ
1X0FWfZiTdWW4B+1o2ws/u5eH5mc3rJyuuz6AYtCMmt+bmXyLIZVxw/dHcAL18zntv4FbxQCIpEf
9zdlVGZZpF/1qzH9F6jFeyh1k/UT+iPOgd94IBp+U+wTjwzQqXrhIPQUnE0zL1p7/HekBZDc0X4+
3A2X1XdMYKE79s0QBPMum56ujAo38qxPLbjmBv5YnNFY7ysMCSWGX0oa6uINhPRVbCzq8eS+2Uhb
Bk8il/cEF7iZC+F11Nr16eHlSfczI/hfbVCvTm4VqUGFrpROeT6LlzLXCmEJsYrYVkL+tMCcQ/Le
zaYsShUPNUfRIFLYkoRpfTVWBVJ7OOHppf0VnNnMHwCYAqGhoRIChNm04XIGUB49YG8bTcvio+8J
gQJkcBaV61Zn5OLRoOh9UQKURDvUTU73lD5JFSu2AakxEaztL183Bs+7cZ6jJE/xdMpyq/ApOjcN
e00Gqe2U3hW//fOBoyH0/lU63FByYXjiOKml0RqhCuNh+I8PzpIfadzYm0UYanVC6wxVelYrj8ww
AoCM2/nQsiRpJBNbkJHzrOq5EYFoBRfp2DEJSxjMOfUJkFOh8AHB42xRzlxg+RAr3j+8/v7fXwf6
0pNK+HvAP+L6caXjyf7k2iGoO0lt79DiTaxTp0tTIBKHEsSTPLC9tQzeW7UfI4u0/DZmicW3LPel
9+CfnCtkLzJRkdcnTWw1Ymydp91dni+Kpfc3zWbXcA47MRAdIv5hmj2wF0DNQCVLdRN8iaFRuZhV
lqwtm1XBi86/uh6Cq9O11oUlIHAQyS5tO/0Q+WSoL9XceXwg9RkDDgYPH2OnrrTuDAb/uf/2X+9R
xyJaIi9H8KxkJy2vyOi7+sw91qePPgxxkQLyGu069BPxepAOowhAM6NOudjsn+ca0IZoYxhW84+j
V5UpNBuivXZKpuvEOj+zGonKvuiN3yWvqJM4jiTRPhsVXUuMg+eab638ZCtP0IItC3WZsEtlFnos
pwIcqKVuP3+KpWgFSCoo2lSKMEeKwIfxKQ2uogIu1eCRa/+nupQDniuflgVhl95eLxysMDUudEpH
cWsGCl442mHfJh6n5hA1QpTQjrm0yHlqZPztukcuUHKYdqX1TLiFuM8XAlP2flLFHuUTAlkdCizB
tnSNhvGe9MhAspc6D0qWYGCDItb6JoYMELdtlDRlJxRjbWbgfyVx+AHG1x8D0BGaPD+lzZ21nkpM
OGwsrnIsKknfx3JpzJ4KniPJ8oWVmff2lD/wonYCn7utFCXe15mRomwSTYB41KpLBv5tkgUmSrm4
v1NMsi40P3US0z4zYeDzNaJ+JsyhyBCuYE8mkRtCMVvmojb5+Np6pPNcdkiNs20cSW3wvwuMWmmV
Rh8ISYKvRPGQPsyua0U9iVhwu6P4Tfx0fyOK6hsVPh+ph/cD9H95NA4wWfPZxqbw+ewMxxz1kdj8
e5CmRquv2E5GFyFa6udzdjtIdLruKgWgQ7vJDsxJCRkEgTD/bh4OxLypAuuPelIfCYNhpZZteQh6
+BH3hcUALAl4/6I44bXF70BjlSxxDwkIARUNu6fm2znQwN47mq1nRY0wxHQSbux6CLSEyk/HiAPy
atJTxeVQs6jjMOrYblAhZipfMByWuUWfNgvtzqiZOnuAwAxiPIkfC3E+rOUymN4wWqviqb9ExLeq
GbGJgJwBlWmI1geoPppaE2ZoeN2KOj53mboKXQyEOGlUxOY9RoG995fiDQ0N91ng1KLSQXTYNUOQ
HLpeY4ahOORCmLIY5b23pkrOv0BH8qFD4LRM+f/n7pWdvL9O0FvFPdWiZVeDQOnphnd8EaL4aWgt
kZEmbpZ/R7OL6HAqFjJqbrqZfEJaIKhFCebo9gI62NWsWb23kL0YsXbaIGc/u8P6X3fJjn5phyOV
Gnr04VAqIfREhkDw6pz1EB8YmAaFQw4BGkMWsO4iQ1QjegjDLbXETv2PFEugCikH33coPbrvhRTz
m1EiLhL33HsKajVXvvdQTY9wluriOwoTnq7SiqAkc2FDVny8/2mk2yFK+jdYg3T9Tro95H8cDx9P
jxJNlOLFqsF46AcGmiPWApzKyDyLJfGIBgZy9UmcwEgLIn+AeJamI7RmuDDzXVEsS1N6G9KTxFij
VD6r84HGQPz1A4nSDifKQmRKo1+yv6lxYfZXxuekXOcPp0fcWnKmflK9+LbQOybSdyuzJiQHjjtL
T23Pw/ZHbxU0gTJjYFXErhmn6vGaYgc3QSvfkIoei4GhwA8oqfJCPg9yykLntDyWyVmkVi+a7y5a
5O6ueaL9vhgF22hMVLBmzxH53bf6ErIRowv/4bIN9qHlABiPZVuYMNS/XvbGE0deXdfZD+Ks5tWD
+W5EDMzcdmx6fHYo0SHm2tkLFhHUzpoWs66SLdLbjmrB7FCmV191NEtPrAdObXjk+ZBk/Pu4fyxv
rggYUfxrJSi8EaClo2FQCqEVhXuiuOk6KH5a8zNV5Pp6KATqxPnT9eJqroDcdMUh2a+dZrXbRbVB
rm8GEVPAjcqbxasnPVsY0yN1oaRzjvahhMozfBlzuqoypwOCDBTDxmhjUhGcmwfbvoGbZA9AXRsX
io1wr8JeEUCuRwD6aWTaVfV1IaXAUrx6LshvJ0pv/ztBIj5bq0Cs/kPKJALBRl3cZ3BtKFmlGeNv
rt9bjm/CkdLpe4fKLZ9MRAHBqkT+pJJxsCcQU+Fmq2XGeTS0Ne4ii+nYHTDSiVsY6z/S9nSc4fDa
9II9i4gs3tYmpEs2HI/7db6HIkYUwusC3KqLnMa3xpwjQZ2q2mNiGWnPwGoxnI8skKn2m12lpm4D
m6hCt2k8JpctO8V8pr37QSmikMTZjlz1+QxQO+NKbX0KiKJbd5t1KoXdsE++6HKufxa4eB0wIt3A
MDR+Ifj1p3A8ZvbSo6HQ7n5Ryq97ByK3pIok1qkGfphhSmq0lZ23ztivOAu/PY35hZ95Ud/4oWnX
fUddE+5HXmYSPBhp7CotU7ICD87zhYoa1VcMQurrt05ZIp7pK+Fmp4T5vaAFYXkUAofOAsGCwKED
PiQVuD55McjRBneHCWmr4qDq+NyS8a8Mwq75285DF8P2QVbKbmAOB+LvFkkbXHZaoq8cyrW+gKOi
uAotwfywhF291zm1emg568XvDjQRJW/NYr08dM5/QF/auKHvK1/0B0VqduzZFMV6bOoXVhx5j7D5
c2YBmCt/kPItZfEYJLfYd0ZelEpUhzcBzml0Q/QviqWPvqJ5cMQlsmVrtFJJlOcV6M8Glhk2/L1c
ZgDUGfr2sus7Bkhfwi4ZPPf+yar3yV3vsRuI/qk4Cl8WupnRRHdYjmlGFMqeBsjD1pNOZwRcUMEt
P5c6fQOsOz9Rr0r6Go9agKLJ+8QAf6pCTd0jzMKyTyXzLn3k4HCY+cISGroMi39ela+VyFRZpztF
ym/c8KzNoY1CDo0m7YgxNWmtmDbQjf9sxQxuBb//Q9iN+mqIHY290e/pOq0kZc8YIDHot7xOcjYo
XiHbL2NOvmObaCjP79P6oGt0cmNrTRGvdP9fvR3m0i7qm+bN1SSEmOIS0iWIgRrCm4kGHDOeDeXt
p5Dv+EDJKmiQFF7nhu/v4vo2D0NAL4drsegbrzgxF60yubfpkE6Vr+Lqy0yjsEVJOhgtE8x5rH6y
fcKOB0P4NIucAPVtxwByIU2KQI8usJTuMzsssHvDw+tSEznhNYlS68DHl04yS17tzOn9TpxgJdtb
KYJt/3rzNF0dbCjnf0hlRVsmfxoGjyxrxcm6z5bqgEfdk361lETaOJMjLiuwBjf4jg+x8s0QGr8d
YxASzDM2O92yMX+wdy/scmwj2fSShl6IHy6MvHZ5VXhPriwRWG46NRrLBQXDqhZ29v/Agp4Eg87B
+MVGVL44CXy0uIA3jKEwHCbCofDdXlEsRuVFTN7pBwDuFCVdXsbRxrt0kvDuJH6L1LMvPXAAeRH6
WEbcYVXgjXpr6JPHNmBbaS1t9WsFoq4+lORb7q1KP4/wN/PjckyaxSS+6d4XDzxV0badTeYpJMYl
aei8ugEPChPB62tNV9EHa0swW/H+6G4Uiuy+kFgIW9wWvCki4/CETnyj4gWZxiagP//ftPKcp5dU
fRy7EnrQYRYzfqgZpKbBA2XOdqDPbgFHKx8AHYAiQs2datZKR4OJ5wQWpw0hiD535oQ/r029xTTV
hfWSAKi4W4qfd6smV0sexdjlpryRHI3wGwoDdtvyULmL+3QlDk1IisrzDle/Mwc+DxzqtZsK+jEx
TxLGYRRnF4D3nP7DvLasH+5mFB1acQu76u9c0t2k49vBP5PqQa6Z22ZusRPenMG/aXgvPf3r1Lsi
2F/NDI4CKYF1AGqTbDRRhQ0ou5c3iO0P9rR0PSc4j34t96ozpyIfU5dTBZIJhq7ybifIGSIh4jW4
l4Vh/N2kJD3nGzL5T2jLKtds9TisWQqoCuKSOLGjDXRXhX2DHLv6GmlnKoAkqhLleT8e4AEP/WDH
fNx9Bb2seNNNpU2Gk5LbAtPUQIsugd7um9piTMAq/oFoHm38PVnMG9Mfx6upMUhU/Vg2NO2ZlwJO
WWzqR5+nBIrHTp4DL2fshtSJAAV4Kim+t4+wCVTK4CZ7Vl0+i/ZEUr4M9/gW2t1PNIMZPNyRADnl
cfnS6H3wqdT23lnn4RdgofDjUCBxs2dQjyfaOqG+uNaYzBNpnwxeT1kMtoQ7TmYc9UBBvCmjawx1
Ed4IucJvcHEg0im6gGYmRONbDjUGuC/skEi+LAq2FnA1alWFeGa9Z+Z2NTp92PGqsTrhkDgeGVak
lxJVS/S7zHKPjIdiOsFKbMnM6nFpb2RmF+Pf9fMF1XiazpDyFDZ1haMQMdPAQ/IDVMCqKZGLeGpQ
FFEuf7kHOCyx4R/kIjGl4FnWwHp9jkoR6UJA6anorP334NvdI6hh3bfrgiMnkYxqnrt+oASA/MCx
p4QzFn0XCzoEgYYNXkFyBB0WH7xVH99E4mCe+KnDwz2yI2iYrjp8kwIHcoZdkKU+EWFInya4+gOY
W2OiHZHIt29r51wzzopy9NrCiQkja060B0AJ11QxFwDbkSW5nDt2gQ4e3Vq1qvmGNwEAF5sytjdZ
eb3pHpjxG+BwQUYTL3c33caM6rwBZYs2pOfRLGxO4/xiL8TWpB8iCys5R4x8c9xkYMnSo4k6ZGUS
CnSVajtQAvZQQuUdKjvq6vk1fur/+HjwM+mcTbNEanrTAGDPkDTIuul++AWfWVC2unIbYQna2Il9
IXyM8DJRqIQmwDwVDQx94t+bKsLV6KFBeBX/OlYVKmKksIpUYSbcC+6KDlcO6oC5+XkIB3pqNNz/
vfzDAAS68ZVL1urYaos4HPhKjfLjatb7cSLbzy33ZtJH2eKzaj7kQmmNPQyPDUCno8Zf7+eiRaOW
YV8xHsG/SiDuYZgLkG2mgi4cSGQwiksmHY7nHCThjqM27ltuA7SCAvQt4bHm2gJ/0TGuEDFPIkgA
j4AKmH98PZFCVONtnbUpq6WuzPc056iW74gZE7jJ+0qiAwxGirM0Td3vyaFvdTxZGP1UAO+hUMMX
39xkX+yvXKFkA8nBy3BCOtoQHCFxdbGP2iCHwmz+KgUX8jw4XL+6oXP+KHAV+4Y0ym6xyYk/VqcF
q+MfHEr6pnoTAEYgGwAkr4aZ/tNn6V+tZiZZF2OEQrYSUjY1ppI31hA6UfGkO8G+jMrDIRHOf0hB
b6dD9MQfjJVuYh+yijhJj0cQ0gvIZe8XK/BCra9cb6SiKD6mjK37faVt0KpklPuRWC0GoihkQ8Ex
t2MPwKNnKGsGV33B7GSJz8czsMXrxpUsHSl85bN6bet548mutNHRRYiu+e7YULvLb+SusnyYFPTp
xjZUqb7dEeowHwnAZrHNxCxr3IhQo+CDzbkKgnCUj9z51GLRlPY1vrBZDMWCTvlGXmw3XVR88U3W
cIuQq9zbnQm3Ls5VrgDZ1sg0xkFG7pObvd1tamffVS7W3hfB2R/gcq1bC3t9O1wzqn0BVINxA9/E
+UZTA4UVRdDh9KIyqQc50POv4TBdd5ahhOvL81Dba6+IQ+vtZ1pySXfHjke/7cYTUGJXa4u8boyw
sAukKuvgMHYOMwabrEmsA0V21pUoaJfg6aixlCbz+68Z+PoqVZ/cvdbHKgUAOqeUg9DgLPKmViho
CmwgSliPw6eM/hNHMH39O+xSMI4WglaAYkX6lmWgmifHLgT8lFVMto9Vqn3wJSYqVEuW/zP8gKGh
HKZh4U6bfJvn4hK0xzMoxRf0yEN9crTu/xuWr7QOZMXRfTSfKkZct8i55FwqdiQymZHYuh8LLBOy
Ei2NkywofmBUnaH54V7SCYPqvl/OTM6ByctI0AyberAAergSsD/NsZ41rmcAqeY/MuMin3VoEj9h
ffBVbYjhx1ovRyCPVhc6MqboUQeCIBDvDuEsPoz6nE0X1FTikINwuXd9HCoIL1dHEGpZHd43wVC4
3tLFC3HoIKChF84gko4TPB6c4MKepqNFrH/YfqcvZbnyGkCrTA+3xPw09AIC6Avslq5RwLfKTrSc
YdPfhR8XGm+kzmDUys69CuYlQ3RhVTZV7hy7mKAQpxdnsTE2S2wi6pptyT5YbDgwhCnLPGjxaO6f
SEiSyEDjpPMPHnLCDlitWl5+v7c4qj6Ywe3sKgo25mlqUpP/mOqw+OFYxv8NsyZ5Cb+X/IGgDSbm
UTqO898Xk8ustVhD+PyGGN19FNgxbwsJbAQahRlmMac0dQWxSr8zEC6sjUX3l3qIvOOPpligrNE0
AknuzJJTPHLkHIfQvJp7ffftn77hv85DgIOLM5hVSnwxiBSzmSFf+Csc4Fm6sF9nLVULpEKYtY/y
y/xcclE/JxoMl9UTzrKLdZ/CSfMwYhYQCQ7hWZ1y6bJovi4chKy8iZK+yPHsMzTytDy3IuILocR8
n7fIYxM0qWFH8ocNHR67CXDNgFBchworyekk9fl9PJBblY3HDQzaDdUL/f/xXAiYKYR46aBHUvBv
oGgj7e1MAylCiy5PRG7jm5TKJ/rsGzU/iC+qEI58DsYvXh1SLHfBdUez90DgdTXFNcqrQOBfCep4
qdLlhHwz/mPtiIXzGXx433+rJ0Wsyh6LEeJ+QFQRDhTQ2nGve8M11d2XCpD2PbPwVMjccTgg7WhB
u/aHW6idlIhkgDJyo7ISkM9aGC+cNh5ZxskhUJLVlR5cODvwXGmrVm3yYHwMyb5zPvDJA4gUPfHn
I5CQu4MGYfVJK/Cq73rQOlI7zqVs0/MuavL3HcMpD2VR6BSs0NFSkOmZbNE4m2B0pCIQ55zMIut9
BVEUXvoNgZwJtzWKLZH9Cpaw1IBbC/w3LP/gSkWrVcLPiIUi/QcHx2H+yd8mJy6vjSphO778NB+m
EfvW8rF5RRyoV3PK7ojcthljsl6w/MBO4g0tytRnIgB8q/n6NGvNBsmm3sbtd/3amCG75QdP1uO7
dhTEe8SzbHInVTbj/BS6PFUx6VBi3QC5bj7RlQpjnYFp+gIV8gF2zSzj08YJlKfqFI893iqpDQLn
zCxKnUbmv8uzC/6bfMEzLQtfqRR2V9Uw05ZsRnJx4hT/BizwfL0VWazIGZFI7/LES9YdDY5T6K/i
XUocCzrrJ/u16FXHQLryDvR4H2q+5X9OZ6z2o1rB1AXdxnWYXL0qUDTuLjkxlCK2Esao3krtQFbD
OvHCjWM2LEdLmnNy6lwK+h80gRoMIsAGtoxo0S8qKnwFMvd8aXhS6Ovc2LnFsAC2uLDZclk2y5t6
s0Cqq5zQLlhtJWrDclDoacUrktUVE+4WsJFHCNRhjZUAoGQOFXrNNqz1lfw58CswhJ3F4EchsksH
VXDlmUZlTpksyloGKx8MZGrvYd6Y4B8wAoNo4f2yLB/AAmLVoIwIoGHbWT0XK0XWqnBywSUqgBT4
UTn/cTDZSORgCMSxdp7eTI3jh/U+qlAaUIPFFKhgisY5Mu/7SgcqlF+uiCq7gnk56mpqddUsXfrF
wufN0PXbHSYuxuh/QqxPWoauCXHKLXF2B4Gf3xAgYwokjQnu9AqR7fHktCVQ9QBC0DbNIvAB2NMe
YiTCtbhhiM7Bpg86b9Eop67+esP++xYdAsg8GzJReP+rMZDvF9nnllB+4b3WiOBYL8gnqU44Cq9J
0t1tFdDlT467RdKKQnH+NlXqix9Li+kKDj5gN64uxeEFXNy8LhtIwcjH6U6/YwDaXdoWgO6khLbi
MWgOwPC/x6EJVJ91K6nl9YwxpQ+MEylOGzA1YnsOMELcXAj7JgBahkKJeJgsNNwgzIjABbDQFMh7
O6C0kqPwCLf4fvdiEzCAfH1pvgC2V5WeT84EOXYc4IuHzGpi4v8EP/LZ7NaeA7Odu1PRm1XnhXwq
vHKLRTSg8CkHyedFrZd7AeN4GD+gxblRHOnAbovy3MyUA2uV3AoOAXUKf0FCd9kwDcSoxV29QCdl
SEg4D3z3+v+yH/NY/WE01tH/nxzpU81YFcwdlm9WlGgjYDOMEjo0qAp36iWE123JYy37FcyoxTMW
gU9K5BIBX3VLTzoKi7bL561V2zCT0C+1bJV36RRrhc089a6jXcLcHJlZAsjnKeQsla98nMTw19yn
+vKtqbMJwfw9urMArafUB2Ykc/XelYoAJWNsTfQo19V6XGhNsVw7pOM4SIS6T5PYzdljY8S5wVPD
rU9rXUImioO9/B+wC+39MLEaRzO4I2JXG+cuoTIlGWRpbh5mKgvt92gG7h4hLvbEeBW5MnxtBQgy
sjsE9pkxcLcZC67XoWeoKiITi8uAPKOLjvroIWJK6U0yHMxPWIYnaU3zRWKExzZ9H5zIdGUWEUgA
jRqqAB5uUTyXzcSzqO7xJ0WkAIzGZeky3RI9xndpp0MSKbgPnczraeW11Cw5NV3PRzNcGCCgej0z
Rnxxwq4tb4fwrfV7j25GHwdVinYAKES+mnhMMZwPaIo4xbutbEQgmqtVtJv8pgoaiaq03Ad3CMfo
bov5xU86wXZXPLTih98yWPJ7KWws4+hteFXRdOq+s0wCQqG9zOKIsnj4PRQkYbmqYLDw/ONMrKSZ
dQAFxUC5hZx9cYycHGlwoW/Af1ckYUg2yXh5ANQBMCZL04ccHs1F3kNflYDKbsnEQKjwlsOpjTR8
wUOhPV43IluwAhyst0zDTiGa+yqu22/a6h3CHwma027ruFhwGWCHtNyykmoVS/dq0QeuO9ar7Dmf
fCiAGRtE1PDlqnn3rdtNeOcuAApl+M1R5P9foSqYbV4n7/u5tzV7B4pzqHun6nRopoAlZVzfbzyB
D53SvXc7GzCnzBbVac7FB7Li95cHP+LBRAq43luRmG8wCgbCITqnB+jASIp1IH63Sn6Vp/rSJDXa
LaioPCxqcLezzHt1CXVzuGy/xtQ+9kLCYJZjLDyWFMYzyu0aq7ORLUwFZqajmjNn+E1O0+Ye6kW1
FQ/QXENzFFO3OC0s61Iq+r+xq6HSJ5nmOBI/MEGqWUmK9dBkcEovxGk7eS8TAJV+fBb8UCoPzTO6
iyvvCQshYBs3sLDJr40DvYVmrArnAKbpudKu3g5KDLDVDmlTPrPcFuXeTdEihTi+jB7E/AooOjFy
Jy/ztykw6hOHkeieZ3cjjdvGfKQIgAJKj/1tKK/Wl9vgL5NUlg/FMNH6nrTEK5e3MZLlwWEmuTVD
rvUPnASF2BCSlKMkEf2vrbTOi+ypH+vpy+BzcCRBJQEKIvKK4E2EziWJHFhJFXVpIWDeWWcSAlOz
hy0EPae+wKyz6ZvUlGJzXc57IsU9cydJ5Ff8Y6l79FntXkWfzSi/7RWs4rqIdc1MArqW9MHzfDRn
HfDbESQNyTYUHXZkx+BGhqb6lH5DuTXuNCYoU1vfKsaiIiuG9y99N6qbasModfnhMRXBtuSZR49E
Mk+Pgnz13Xf6rOJmhyC49E0qIUhg0bbBEieYmIInyzpYfqXtiiIRv++b76Q8P45OqK9/llyT86CU
wGoXTKPqo5pc6nIjO9t9oJH+PF+b1IXdcyHOGXZMVRPVfcZwaZdotYQsvLeLNI2TNciOIZ/IX0vv
CBSD0kAuQ6jdFuqypK5g/6jIoz6Cs8+BFyuSW8NRe+dV2KWekL77vt5xn9AS6rnspJhMJdbGAnDT
Ia3ZZWBLOU9buw4WMWIVZ/8KnoChQqlpSC/+CHXZqWBAfzWwQRcgZah3KPG1X5j9EjEt08uMJ8eQ
FHETzJAaUN46+4OEqNYJDLceP4vwh8Tcy+Tl/Jdk6HhlOYORAeekJnwwS5WGZdBG7gYYK1WmKwkl
Yl0zWTN7NV4M9eIM288Qqsg/esFSd/LONZn0gOeopki5wwte/ZhXHza226gsItNErD+naflXJRan
RV1pqB3s+SjzCJYJ0fSgu40uT3/Yku3uYPKdVeyQcrQ9Dr6yjhiEdU7V/4XAv4g9JKlPM2OUxhl+
zaP93A34xda/RWfesAy8pT37EYmcAhLxP4ZkDcLS+IlrJiS0vZactCJZl3IWVgjzJAjIARBQ0Yiy
MjOaHm3tBDSkGT8VauvPCDNK1ZFa/vDDt62k7kagrTvEMVEKVQD2pEptkmK/EvGXkZbSHian9A5Z
NcXuRwAxbR8JtrVc/YrNCjPsb7sQUoWn3hBxffZTYDFUIQ1M9+7k+gmoFvFlse9Fi+ruqxbZJiib
HtW4RQCBQCDrCEiIE6/o2mhlEzf5hLq5et04yT3D5QQcAFk77qJ0LIQKbzmw/17tswm/ExD5FZFB
prTPhVfqbYCGjWBD3VnafLP95H16FqD4E5h9k4imndMFYM6WTFnsF+G/86uFPiUn0EanBteF6Dvo
C8hDb3Gsa+oFIE/iUItAbnZvLOU9GAXKtXC6ea4yilZlgbQfclLmjnPtu3fSDjdIpxmoaPWe9U8K
tQ1AKehuUWWCvWxuLkWq6qrPzfgOZaIZ6eP6122Jx41QVLaNwVblDfrhv8eKC2ofQaKol3y1Io6/
KjX9hVqx0Gcg5DywlBOGMbOcgxhtSn8peiJo0OC21A2kPqMXjmtBrRzkZYENVR0HptFenz9u2E1d
SMbiQngYWshvDRbypos38KA+sVs6kSHUhSWa2ShO1oAQJ1XpOwNqrTFCaqumKMdyjzNAIWGjzZcW
FLe5vjFCsjJaH4JC8u9Ps06fcG4Fph8x9d0Q2P89WgV+e0QudQ4pA5UfbD9ozSNT0tF0WCRBcYVE
oXygX42PDPso8mgTVgIdJmxOXVvkiFp19I9tpJsf2tb/LmRljr2UTYv56eOsp4HHaKIA0yUDcI1p
T6GgFO1AvKmDCgegDyFxe7z0GwTb4nzHmPrIKFZEw3XGuPwXjUfWJnPP9tixg7tEL3fCod77aWJR
JWRkX2Cp9s9BwdwGC1QiHh46OHXW7mXl3twjTak8nIMHgi66H6RCv/Wv25fZan7jHHuwXAMtAvMy
IGoyW6Y7zeuq850QFVfCsDsewsNoRUarFxb1vJr5og2QeQwDR3qTvRQOtm2PwwzFKgR3lpdOl+w5
KT3Q+0CfkrQ1lGsC5I0iUff/HpuUN/PgUDxL5IbXcJUZfXyXYToeQLIiWdJMJuHxyU4lJp0HqDZJ
Rsx7p/3UoXXUxKWTcTt9/Orts/uGCSb8itrzzeGYlgf+cThTNwilyhS4gU4gZW4KzO6uQBwk0+m0
iGUeWs8HfxeLOqNrzY4oImBMUc+I7sIIC20APo7FpmLjc+ZDIs4VxIbsj5/OFTGapg3URujCp7FL
OpXp0vE+y8UeyaaCBY6Z8EFBYFciWTb26g09hXSBt5djOz7ZgmigA6uWPhu3TEW6DsiVAmDyMVH0
E8sDj/pYn1YlVxQOq5yxWzXiP5QgdSjhtPj5B5gzkh5Jm/8HCQfYbwt3T1QjhVWN4nspfTqsbpwa
sXyQWsuA5/2DNCRKCGgAy0nUGHEMrymSQz4k6qdfZbwu40EfRTKUqu6aNOlsOOTgVxe/izvtzmpt
rF5vO0mptAjzV6rF0XkQP1mEr9yDQ1FNy3mqkzUOH8kI3LuCB6wGkK5dy2YKD8meQhvhru08A313
QS2FKumAw8OoWRy/HMLz96Fwh0EXJ8tKRARcs8MdbXlNF37RLSX+3s4jO9stjOubxFR/TxlO9YdS
kzmQ/EEtbh+VShkRwUyT/Hgf14nfoHDIHEI9kVuMFqKslBVIx6AIj4uF4+6nhMvKnzn+FoaL3gRX
bXF9aOi0FSf2GmrPNTjMxg4fyAYCgDp327EvVJz3URa2dztZ3pwpuL6o+79yN5Jd1GDycOEmot6w
nqJWTs8HklJO+lAHjkfs+9RLptI+mmHwBYNm36MTzmt8Ml7eCmhWbryexWJ2RSQ+bYXAVRoO9otq
jl0wmTW9qneaRBabSswo/ALuvJWjNu3eDmsQhCx5yL+e1tx4SoyOMmMp99Xj+OpUW8cL6+7vS34w
d7yQ7CON79AvJQmRgPXoSgLkFsVdYvwx26iL2ME7oRuOEDZzRypDUm4sqa3Dl+LnhVlf3qyo4qZi
NZf5HYbjJsMKOe6skY/W7u+OiQ2pcUTdo1L25/rs8j6bWasfEBHlNoj5yE7RoIhgr9Nm65ZclRYp
reSdgVkuGwGWdqlOX9MNXf/cI7L1Gdj7JB0rbVnI/HsmK/7q622/J+/pAP4djtQibZNj8Z3U8ft8
5Iz1M/kNv0MMfPLiztI6XABXDSJwuDOjuWZeq0iQWLSTzOLBVNPJzgu5ZLEHzQFsFFeSrMEJCj71
HgipVQjRUzNKaeeZzBRc95hiihH6FqjapJqXxNELIv0R70oXKh8dg/9fMGI6BeLXWYr4zB6yq+Gz
xdsfFh7ZW2Uly8tBUQBfB7yZj+I0YyfTsnlwY4lJ7LoknMume1gJf9dcxV1wFv2XogOVeidcz0ub
IBgg0jb0B1OcnNWxb/edeOD04KRLbN3jMjTWCU0ypQeqJPM68DXDahIa96Dlc1wqyNlJJFohksfr
BSLnb842Zq9xltOSUrLUt2sNrB/W4OmPdBQPHcjlCis52RjNqza6PAAwA/pN0fL3Fxr7PrqIzwt3
XzJudKaOqjyu78PwYGe22gWmxZIT3ctOtAB+R+x/HMZKTXeLe1EriqCVtEXvHbxsdwrT0ampn80c
YsTeqOVKbXGxY6tAFMzW2MrsDN8TWUXZCuK/yOXe3Or26TL2G1BzIZE93zfazocN2lMpCHMszNRD
KFnQRrO6tNLfeulYQ8a9qA6/syvfVO4GzeXhSZYj7KejyU7MEIGkVsk8WrjUWUTpizSJ8T8UPp2A
bDKKCQGn+HhTI9sScV7TMqC9koHBywSA41mM4M1nnIZYeABTOklSwUXSyJy56HBxRE4GEk/ReyXY
GYICh2ToXb9o5kC7xBk3RKjLQQV+PxpBQ8eBJu0YqSC4DrA/I1IzGFZKhDZddKZREbZ6KTllmQV7
s7Hqm0xBo8CID86BLj0qUhANYkSUXALYAF9z8SclcB4Y6GGtvgazXlOP5zd7KhTySyqfc1jsxbFz
a2fsbYd/Dn4KVuYCQgweJjov5/DtIy5Bz5Jf8jBmgBcEQAm4nO0ZBr2YCodXbmYB0H+eZ2FNWqlF
qK8rExjOMQd0I5Q2dkkSM61Oqv3UUYlXtM0aQWiXjz4OkLciSsFC50e4jGEIKpms1q1flzIYXC26
pSQXKlyZF8vQ2ONIlobkb3Is83KjyfDya+KGzus6PZ2IwsxXCafIqZzpaCMUgG4RW1rlLLTcn1TP
gjKtuEP9sYT6APS4bWISPjPym+gJ88+Em/MIP2O6nS+oOOW/+UhEJ9G0Xar03qPXZvhyN26m7nCi
d4TAR4j6aScp4JomqfkJn7CHa1dYg6j+YNwfIhWfMZlLoTOSEH9Z5HOI6Y/272XxZoCOEnlAgHmd
ZXAM85WNZMQRerEdnvlwSu6wzIHzuR4obGYOMEKpUzk+krdtoJxGXSwAA4l639sZO1JimMtQYf4R
uoDwSE2NuQrjCTFCTGPQXNOZMrbRglJ9TbRm3o4w2hTJoOQg+nEGvWtZXk3iwyV2WuXsSBabgAhX
b9ZSTL5yyEqYLaZVnNrjZhIrFzKgAR6SbiqFj6TPCtnKPZtglVjOpuMKutZs3MDe404ui11hYQE/
vi3yTB4jQTcWAyHlKsRHy8ZbdAF0QQarrwIHFykhAWUpewofvosfu4kiwlO+Vxc20IX7PGDNsnei
AmJRSks1KhOPWq1S3UMS5Fhrki270+6CDjy16f90qe1/CHgLWaGVYrk+5Ewk2/GCITFzmn4sPL2o
30aFQqRPQ10LaXvae4QCjuR6w/0Hkyz7jejqevMss0kzsvZzEmcNn9s0UaxCK8VSVdx6iRupZkxF
BrUS+8m044WSXgifMTLtTbw0j4LwgACXUG9Pjrxcp0NMhC0MGIdLnUsQt/fFtICj/6xmnbAGdQZx
sx3/txMeGiY5LaXaGM7DRm0edgjPiGm5Ve8Rts97Spu2zInCVUccLV0LQTopD9O1usFH96s6Ta2K
UWhjVU6Wxm/r/PDlL6pdImFnaaaifymdI20VuEDiNERTv30JdyhYb3v5N7BnmLf/YTRkptzf2zKq
/CI474JI7Nfak9/PkpzPiOve64117NdUBxudNqtTSFjrILDuhACGhCLoSPwTR55StFaDmilPu0fa
Ys9uRWUfZbebyXs56iBQdJZHj6ux+e9S0wJHMvsDNjF2pYaNpmneuOVSal/oK6k6hbZad8ElucEk
C6Kno9DxM7lkQRd7dFCOS1+ttFwZsMDSSWX3zYbi3OQaaZubpApxSoiRHbtpSxea96IsYLt6WVeT
Qrq56rmJ1cZCRmT/fJlGAUqY/Q0+YWhsQNcw81mjrQAmnQ3eBbh41/0Rah/179abtueA9duPM1Ie
WU/bR/ORBb1YMn5z5UaSOCm/+SqRYk40SGPhjElbYvQJxdDadodLMS4dmGWgIVDUxsF4Xwo3b1lV
k9oB0iEONEY2KqvSaMDtbeL3yKtUGJHKxBj/Kbnm32nWsEmXDa1taYTzN+OH6iFJ6tQfRyrZDOyq
VFSV9LOizp2bdV8hfiuchQzOHCMYwGgN0gkWF6RC3EpQjXPv1q83LMfnmJkANpEnu/GApn5n8h6J
QnZcGDlweEqtPyaRRh6OEzTaRZs9zdpxhu7j4oQ0GAhNxuAe/IgVRlldfuiUFZivj4yUjRRtt5GG
ShIEmfhKXyWRUOBMpQOcQxpGckP7ICQc8/5+snoaveRRpVSWXD8vCnK/AYENmTUul2w4+coGaGCA
h8akk1BBmoxfI+8EHX8a/evIp7eajLQqOme1vTiWhBgdwvh/tk6/V3Hirjb4PJzPdu88jUQ+xwU9
990kcAjQwWd79IQLkzFnCMkNs1Yy9LGoskxkiIqDiBkL4hEZdDCIx9+SB9Pi+rq6+zQPiWcgbKm6
BwtbGapNveYYX+qmbD5EeZoU1X9hEo3L4zpro4UrqsOhd9ylB1IRLDDTaGFAPw5yHQz+JFLyvCSy
EaXbRr4wXzklKzEIu3xCRCEdYMcLP5z0Xve1vg2c3RhUckfPUgjfG4Skr5uSc0i/cOpSx/C79VC5
7mOLIrqyy3IysyzwnqRRnfkItlGTpt+b9B0/09LM1oZPjj+kLtQYL85ILWq7hBN+Dkge84tR80hn
7Cca+fRGKGboLEivr3VH7CoqwAYTz7HSrDZ8AcNVyqXXsNOFbdSH+mA2eR1mETiX/TLQy4+P3JPc
z2DS12wYMlqwNBLPa+UqXoCmNe/Ck7Jh02eQjp3FVqk+uUnCYxBbnWBtJd9jOqoCIngPcgk93xNi
g35YmsWmDIjucxD6pANraRGwwbrMDToNH9ITFjTbGY2oRzooktnAbbvM7JhD5bdA6xoW9QMzl3A6
eXewGoSSiwCoE5zlJapg4er8CZAz2n/+RBKH5arvYUrW2szjL7+c1Vrb64IjlNTlvzSHTAIAySGk
k7rJfdy2OILwgwLYlTTNMa44GuBZbt/JuaXsX2/W2xhgoHgbq58R50s6p9J89C5slAeTm/g0gqxk
ZOdSYVQNK36LRXVsxN0XKORSz57flUA9uo94N3uE8XomaS7L6MFaFYAKE3Kd5tiWb4TzDshfneWx
bBUZY5GPnFf7HU+sd1Rsj2LkrfsffhsrGm1tRuweuDvv98KmUze4RQO9YO3d414lSCTO1oKBylfO
qNrcgQSn+OEFa11x1jYNasbEXVGQq7zXwb11OEA3bWOaUXeiuSyuENCaJ3eYPTH2Ht4OxNHPhDPV
ZR5O4wd0NrkTiMQrSp1hyzTaXKubvVkPPdeI74RZeMWYp7E3iQraZP8cmhzbhMC5vWHYUcV/uSgf
BX4OCgRG86V5dDKiOD6tCCPNoMBel2JKpih143wLRVJE+4y0jitk8NmFk6vMVvBPI+z9OPGYIXI8
TIWSVzTY1faoRkpranitIjjB3ROUdW0boRok5I8vEp45K/eEfbth4ZM0r2zIhCBkzFsCr4jvcEJf
0+g20VxWcjLpMTwYkxPXdLcL1UKNBRCY7NT3Jw+iJ41yTwQzvGCDlGMdjGq4IcUA6JbcFXviGt0I
9GFRNjuepBUhn2iTD2NG2v1doT8hJFBVrrqJ7RMvqDit0lacOohSD+UO5L3ryopx15yfr0Ng0JAD
RwvIHLnKcWxv0wJtvAkYnQidXSWCv9kOgZV34M9zANPk7eVr4WWmbPASEfG1G6ylez1AHkUIe5V/
qIF8rRWFzNL1e6c2Cg17ewd5ZNGiijFEOhN7d8eU2+i0sz11EoGm6CiDyCYmdI2W6OlIX3CewnKf
qrcds0aqNnKriUH75/bPxcBfZex8LMC9ok1JpeRrGAO+9fZsgxsP4U/xtg6WQAaUt+vORbeiv4Q/
81AHavBBQO18JpHrp32bP9lZUPoDOV5avBBo6QStBg1m7sBvKLs8h2xInWCxLju7I1BxffRnH+ni
1+MbpD4COBiAl7AjrMIKGVt0b+9I0MN+b4L2Tr21cx5Mb8gkgEwLopBfJpJ8x7tVd/uV5/Oyei0q
AKybTmOkO2ZQHLNUHAR3J8g7/ub5oBaNVKi6g1hqOLhSVMFETJjB9afKS2HZt/qE5k1slVs2kbn1
+jJW0avmdk4JZazvvh1EkhogwdTbWTEokQIELJg4onMrETHAFg9XIDaowNnPx/Fh1qfhI1ffQ2b5
xJYJcn9Cxelrhc/ABHyjC62TEwbSuQkbAcFmxtnmXmeVq75R3LtvQc+8l11F9ZeubY717y82DX/F
IkH6jYrVxOg+apoa5REAvMbnxdtVC9DmnhZqeTG6rz/eEG/v5rHSfGjbO7kz4VY898FvMjsueyi7
IyGI6tscBMoNlpzlITs3++jARTxlM0tYcK3WZA60EWQCh+RvkiJZy0FGo+yj+v07UljMJC1WQpms
AVfs0/ppz57g+ZP7NDpIbh4pRK/xoYLxRv4iEKBdxIWfhHmzBL9kI1yYm3yUkrL9nZ8vAWtf93mS
rAgQwP7GLlCYiL3Qy2Fj7jYsiSutW8OOH2fassqNOu6EK6VdIV3SjaY6p9IoU+JHWDvk1+9rN1GY
L8IKKbOR5IWasERufMtJWX0YH0lqk4kwlv1bPZrueDOyF9hsZbnQHOgLWdPnUB7DD6PxCER5IrHf
i/tYSeGvLuypAvR5U3clvnykzTTWO/FQ9fX5JDIBPrgMwyJtP9YTiZtGLvqE9PjgOqNaj6CP10vs
rXoyQ2rHEZf/awoTrSvhucaK1jchfFgGmLzdtFcrltQaLo4CYUAJy+ciOaj45Kbd3io8xUnihM/m
1sBG2ZFUWaZXSe1mdRBiMHxtC4T0vE82y4Kd5ngan4UzygqIHNK7lTt91lZ7n1V9AlXbhN4BW0yn
MwvMj81NKrfEiBdwhLjguZj+PhpoWe+OYKVlgBWcOr+4npRZwpRwlTks9ONLymlhKJEKg3dqP+cM
F+we3RiuB1COlkzwtFPmubtSWXHYaBoZsBoyaXdOUcMSRpeCP8W7tnPxSMFlneCpo1ZvnBWVSjr/
CMNnWfdScHPSaVY6kRtX73UstbW+48pj6t1Wzprr9MrgO8di9Yrmonsg6Dj/oNH6K/AU3D2m1Jkn
msDGz31WQjck8WXIwPkX+aoNITfsbvVQRfn7QB/zzuWZw525iPAOwz8x53GpEr0aQ6/HVJRgO0Ev
DUV2cBaWXTge9h9vMrFYygaVbAaDy23S+iMpbGHtgzg/3dyHUG7VHJ/TbISJPXxtiOFeCfkpUlUb
5T8ceiLtBqfdvzsoEPHdSWz897xwXRuQ9b9lzQ9MYW9KhQRfKFda2PPRvMGuuHUdqPkfljx4ne2H
HJPTo52zVpKEvwKjyYWFDZV2TBENuoTzDF3WBTjcqKsp/cY+uGNbd70ZGoGpPV7JQeSdHg/RO93V
PA1VyzfrB1iTfATgvid+1k073e66yCZAjbMiYkF4qEfCXaoCkYFm8KaEOGEwfyKA9LIGA3jdN50B
taWZ2eArtlct85TStriqueXSONJkzDTiRP2H67EuDL+QRNCmPt+Dd+O+npeUmHYFgQTb7sp5was0
TEeIt79tNCKyXjdVkLjlpLbfamIJxYNGwhYgGUIrx4I13PzUA+WNPym/B3FsWaPcHK6X5d0aLBGl
ur3zWy0dg2T2t3YPI3bNm/VfR57+IiC74yGa8LMv+QVhA/N6Rg9onDg8DGWp7iLmrcyxIiMaAVvg
3kH3ytL1wRL81QiKCDv5d1pbpRUHszCSRmfljEbujPVPyGlgBPSlX0dEIJuax2iGT0bu1tyivW/3
EtgF2cwEmmrTv21AH/0uJkrc8gm4l3svxNb4RqePbb1ey1TNknEa77WqUJ1AssnaF216UZ6SA5kg
dcMPlJo9PsEhVSJu+XUvySKET6shVYP0ZZmL1m1R8FhCF+49XWsy8bvMEb1qy9Ao61o6sGIwGQYA
gWJSgdTLmcOGblayn5EaDX1xDdYpEZW0UzXpz522cV3hMRHs7XoEBZKe3aCjvX+KCYA0vcbrDLaK
Afh4MN8h5n3q1KsAoM3gm5P5SP2o2FWhMIDwI3Av+qAqbHklu+nVi5qxPMj3W+A+cpDvIx2dBt4Z
yeN8s7WU1WJzQzvMg7V1SIjPOFzp/TNwHkEaBdN49lpvK6b+DUkDYUyWSVtN3e4Umg3mTmKPG3o1
Veq9bT5w6pJaSnlReXe+7oRPbydDJKbmOezObIDK4O03k0RsOggNtHqbUuw3gS4x3d1+JxCWGim2
oKqTroWPyMYkFLJE/WoSi5dg+l1UW4YTylkJ0V8oMFcYA21b45DhofQGUwxyL6P/kE4KJWcIfCAi
UnrlPz9MzQpfdZr2z4h9o18g/xeEyVq2T6n9gNHafTZogMrTl4dNJZ+F/Bxkvh6yOgRo0B2KmYLN
27yQGSEyNJ6u80h/rgw1zueODVhJXZgKsOEHg7i2nlKItjeS5phNqvoSrltkxoOa8vwLpqtryguH
p5Jw4G11cbXKFw95IceZXLdn7E/ce+KzI5GqI29d4GIMWbUa7mi6yTVl5x+ujKu/kw5cIAB3HS9v
yLk7L6w2b/HIaLMMknVEWpy6Ic7AP0UNDE8QcNz4Ejbyz/lgnqFExrEIAw6W3aqJ3OM+YuNo1Slz
7w+0J6FSiC4ZDfJRI7am9LXj8EM1hOXcA95uwfmIHKbh1JVSCh7b+kB0cSLPW5tRrCz7QS+S1a56
YSjNUIzVKIPaC0/VS09qlxIR1P2RyYuHb5N9ra0LoouzcMncgRYInptMTLNBi5HW61R6SjuAJnUZ
jhYotJcjE1RiuTwIPyxpbC3pn5EkxnRYFobQ16uXsVjHjPK+CvJsGWQj1Pxb24yUFUCfpLgpSvOA
RV68l4kA1VurWCUbNGAsdJFeZ9rccWn8DmmRKM/AsZ3Sn3FK94hTzWESBf4SKwBx1qjpWMXlZzfh
7xH5g/dqRNY4QYYRkMMa7K4l5/KX0DQj1wUCepvJF2iMaDyxAM0lMTWBmtwLd4DLdcAsqmOO7Skk
QB7Vl3l+/0N9/vQPKKjLO4dvuSy6BP4b9e0U5MvbZT/UmfcU6NvCtcJJQXVO+X/6XyIr4mZEkW1F
L8ICq0WRz5acPC0I4dcTwbe/NRKZcr9Na3FNv0ESE7XYIVNv0fMCsCzJjpSqaJkt/uk5/jYQg5CW
apVvMmuI7fyXNj+EFb0EvrOgVkT0a979MmhUQfMJZ4WypVtwPyxpMSqkzs28/1p4ie0U9Nr51iZO
lhbisUSkOZAp10FQyIQMfETetQ1NbnwmRsKNdXr8sUmQ24k9l3vlCB5T8UQaHXHFn37s+6714G07
kqZxNucmb1cVb8Np8rxaUXkL42+2yzUoXzRzbolQQ4CVb9z68VoJDikJZ//3A5OMQutibJBZWPtV
tmrC9Rna+MbQX5j776nI45GeXqNl3iQtMPXSJZ0FUCxTvPRc/tcE7jOffQ8l3IjUDGrWjiT2pYKV
ZSmkMlu92z87YHIEbUnCoaGQmppC8S9bHZClX0NALydWHpdp624VizjbQJSFgkEjvG8hy6aKpBZ9
6eSYLPgBu8nZiswDN/c3osQwGtweJKUGXgyPMuMhhJAYQMZ24iBHHe6HAYE/YfKfX4/I2wbO4YPW
IIAg57uf3hb9DfXIsL8gJ+vsrIOH5xyRnUMfvbCSSbIqsnlsP3tlxNT0MhqALmQSiC45/i1T68kk
5XJCkC8dxfzOyZpdSRD0wm3HGa1qYRv+9NsvnPuuq7BkU8tg2d8w/xMdUFK19dX4/BFGVPSjKvj2
i17sxPR2l4sZ68z5SfgGYoUYqE3lYnC34fCWEBIV/LrH+sukeLnzl7Rmpy71S02S2G9mYpac3Epc
R9F9cIYCqdZC9RLjsJejw3V6V7gTxWJ4rBgVroa88kldEhR6H4PAYPZXraZ4oT3Dvvodog4tUsoT
1581JEvlx7gWkpIrjaQ+L1VxSmc+4OwGE92wbg6IOUh8LEYgRq+C44ueAbyJ4uEN2MHslPRNq6Ub
iY14gtHutuYTl//n6x727y1W63CGbKZbkHwgVNy2ptKim6EMBhxB7VxtpO0Rtn27YmAhQYZX5yz2
fRd3eTzhFLBypaOIkZy704C/zve9Q91//6aOmdkeGOcVH033FTmwcyLkNxZavG+DGb6F2zc+tcp2
h/cQqqBLRkrcSUvx86gMM5OdMkAl3PRVKJyJTlawPjlWI0tNqtEh1jJCUd8th37Pp+WoydyuxW3T
t+A0d1ATgI7YKoLewym2cUJRrcn+pB1N2wmDFdGVelGYJWqJmGBvXrv4JN+AMXxFjnkUsSRI2zG3
iwVmi/t7AUU9exqwtkcCOHg6p7Te7KQXELqKRsB06WAx5GZOWfuVChkzOcttVpyHHNTZBbsRtww3
pvf+fCwVR6sAQygPChTY51/xLPRHUFUwb5N5ndxVLJqDleQY9kHSo+tnIaHG2vPyOEvZRv+o5Ixr
DoP1w4SYFFGeBqtbIgPzQH7fePBpVHtVIAgu72s2iNFFUHRQ14ZgzxL6H+FldwL5Ml3TJdODFene
UqZ31xz6ac8x0wd85qBKJ+oXvRiUU/WdC7b2TJj8j5ng0j7M9UuOgmO2XuowEbvj6JRBWpBkuwxV
czLTpDqq/0kEVQIUbBqb1tm/sGudjlsZAG+Vqpfm3ZV9LAUOEQDUNndAG1bFsoToKWQt2jDw9nqi
hZQHTiWLLqraElzHj3X0aoAMfg+o7qkjydR9sU/0ByOcgrJXVXhawnH2rTH+Gi/vOshxOnu2vvBl
/DMYhX5Io0bcpZwcTGiAJJ+ScR/kftMj/TF8kKwH5Ux5zVOQ+lkgwSHecjqK/ldLlxGQYXf6MRwz
fmZ+no7tCUVsp4Jdg9ZYXVOMv7TcMxhl+Sf0dsZ2NZScZVTov3hFr42fUNwi74C+mTPluGnsmXQH
IQgwqKEAPlMe61+FTkF1C/rDEw8CdkDaX3/XRtEd1gQpE2lconaSQAN1qgpYc1mfug/IRidaqXIk
8WLEgXqEzKvuuIJvOfHpCEpmEM+0LMP7Wk7ge7lPcGqhXBHUeEHch6uaBQx7kOmrQsi4DwJh6UEm
4W9KMkkdO9tXqBbPSLvCNUM0p9JWNPnhkZn22WiihXh7uCgeRiUi7CA4+hGrbgEUVwPR+NlyEkD+
BME9MfyA+/5Vbg7XVEFrdqLjwubjlEjWfjbfvbpCHtHzphCHYeL5nh8nm+8CA4yeVPXlDKleSihg
ujC5n5ODZqWrxH9kDvWijHSO/y8/LuzZ7s8TzwNbejeE5q8+Si7tpWtUqv6fIO7VBog3YMK4Rqk8
sssi367w0LTvYeojrFwvrmG+6+x5SgwInL1YHkH9C4CaKCA9UfXv7vj8cNRuR190iNFPFIt22Lb9
9UUQJ72kr2IRr0sDGnpKga7yzaRjPJD/wgBRs30hy+0E9TfJaSGMT3Yhnk84+pWS1DX3b62SHPAJ
Tnynq51S8+sk37N9BR1JhLUPnNKTUbf06jsY2wL9ybtS0o6H9YyVNx+F7/EVR3UoYSZaXUSuKhmZ
ObKceVcnnN7yUSXoid/swPUHWQHibpI57Co0E1ajJdUfa3J4XO1TvUIRvoAlm1JzYWrsl9ev5fVX
r0YvmWiiBNfysQsIXhX7/4WVgQ7yKwWZWs7O4KqFVAA8hP+aJ3m/eHKQwzTk5g/TI0H31CuU7Kig
G6OX4gbRdOPbBOhDQfKa3cpvbnFI74j3FJDFy/cjkCzJQV3k0e+jMiu+bdfYj0ilnwfYN6LYPCWk
r9PPwwDqJGIHhTc8Qpqu9ds08Vovau+cOgkJMTwG2dB7UpK2YuU+PH77THlpBtf278gaVimLhHFh
CXP4lr2aYW7DUp9gqPQ3twmrP+Nd3Wqz7Ms/F4iWkqjxfm8gZm4yS8Uk+sgAGJ/pGyAOwOOkwocd
8tbS+Lh0N38laRzkganU2suYTu7onCXzOR6bJORTtT9Pu/gJPA+D5g/KUAmbZ8zs5mMoeynaETWW
mX+doLRI0+JjJbUiy5w8xYmWiCYLKnT/aUHZI1Ckfvs5K8Zt/wC4shxY+r4hoCWD/1DXyP3S96wd
wzJOftZ61Ti8Viuf2cCUYVRGpi+qJFFWSGgrySBoF+BZOGQyTrfj5ffCP7EGOvzNjvgSzy37LOp8
VG741AT1psVuIA/CJQGZaMHLuq1xk3Wdg1hc893krZTMF8TE9xu8oNESsuFs1perOxThY0tqbpVI
9003ilkEqN3ad++nWUqk7L69hCY+QtGDfWURKpmtHxYDiVAET3ah/6ySzYLXmanOWOzlQung1Wp7
kvz5ny1S1bJAvY5KzwpjXTZf+tv+HNzws1PC4TlLTRhvDIEZkYmdrHFVANn+p91sZSlakcGnk5Lg
z+TdrbBBSSGJWj0AV7izNgK2mYC9eklnGw2N856CdxywJp7duU7NVMbU26tlFrYx0X5jskNb40Tm
5q6jrkXJrlb59oFE4ePRYLfMdPVqNPOZIlTcjarHvg4ghFtlWUqm8P9m9EYrob2u6se+YgzSVxGl
CGiGtunm9A2F2S/70EGMUPBXWroyFC/7L8QzFAncfQd5Qm5TK3MCDK6+0+77oxcyjqkFXeYqj4J7
46gonLUlMX9t9BoH98FiKuKZNAdAYZTTpL0zZgd/R3lzaPAc0Ld6YlI4mXIJW2mihp0K4C/i9kTR
9UX5hDAGY2RA9U5llRyZxuI2QSr0vfjJS4g0kgdsJ+0VPNQO8ARiK6JVS/zSW+LtNtiidNYU0+kH
tbr39U2BSRAWhvEh2ZqvcrGHxC5mDiZn16bPSE+lgs3jff6iwQvYTDz83ChBQruXMtGcJ/MF0klI
jVf/YwayVXjGxZGV/EAicokrLQtZERAHbEdszqiNjMbOXCpKJkhVgetC5djC+6vVVbQmWBnE7iwo
fXlU6qC5daI5lIl17Rp/s1A1iumfkbwVk84Q/9r+Zj4EwjEcTR921gpTNJHeAmyudIoKHI8QUzIi
rnfGSe0nW94fOIMbdHKbhkFw3ChSwqxyvkVvrzNds4d26cfPhA9UkgxcQbDZBF3INYa4WBgNdrtC
wTr9a/z8/ywlWI9UQSaxnCkR3NG9ttGsxlvUEfF+BYhtpBElCqd4KYk8nx7cUW2zo+/KyMIMA4pw
7Ri31+vo6aG56tnf5E4T9mEbcaw5pdYSF0W41GmLjlKWpZRZEDJndU7pCb49CpjJmuB0o/Iw/0y6
kNzPcoYoLChR0NTxSWI+eVGn0DdgzfFImjgBMxxIUddn2HxZ9lpFoFNGjMhNfbXxVOFhCBRUl81S
YcYHSnfjYng6/hbU75bnRv5jC1mVM9/LTwQ9roBrWzZWaKTA37DVWVGIbr2ahrSGq91HlyyZNEGY
nAV7HM6iKS5kkHxQotceW7B/wFJN2lKvVG5Y++dFXE2Jw1/ygVO1YyNEPW7rJYvOOFGTDSIxWAOG
P7zju+3p+50a4+sBBcyivu6oitvTviNM8fkrDztCuTJ564nxx+Xb3bKYwjJzxoUlIwjq+wZbKgPE
TlYESAaw1nI9bwmOSt52dCzB6DIaymt2PhQW6eFa7p/POO84tC2kvZBNCZyYufm5/Vr+0tdT+zIr
zG3TjUjPGmtujgGA2LNvqh4pWujkMneJZd7M9Djm64gFpftMH4TnMZlQWrMdjjFu8LrHb/s9M8+a
DOoMqabGfGUT42FNQTcwMWKqdyXHI4soHt0fTnU18UTsHcGK3ZiXhc4K/jCYZxr5dDzLfXTU5iQB
1VOT1QfFTEmq4pv05+0TCQuTpjqFhw80fy8ug9YIk4jNt7IRrZODL0WGAbuXkxLFIhctNoLgWvu7
kW+M0poLhru747wStPwQz3mKio9jlr4wsbTXVaaO74soBqSMuPpNihHgLeHPhgl4iU/ectUcgzV/
x56hADzTmd+qCtPHxwlxjyhOBwtQEGa1EEAxFlmk62Cf/SGD/WuzLf5XxK1Ir12ItPVQBAbUEktJ
I5bIMvgpmUjCFuDx5lw2Gtj7jUMD3XvG4zvO7nG7ZoiGl0NspmqfzmoPVEZms+WHZ1KLx6ENwoa+
BJ4Om/maUN5g9dnIi0F44Ulr0FVzdHOlqnzIAdrvK+wibNe6E62O72tw73dhu1n3rhWkETGtli8B
rL5NWmZAuHU7guxMCOIh7v8dq51nTdfVMiVigjPG47FmizPlMvAV/fHqWiYg7LrQEqhsBRKRFVni
owAzjnOtRvczTLoWPiDWoCeVaEpl4+FZv+3qFKfa+YVcFoExTx4e24AZ5b5dGvOIbZ3nL08SgzQX
a/clAxFFuLTXWNjirCpIEUK1Ksj9z2lYWZOKGVaYd0/zGtwBvXv2Rcb/HGzrikyhyiGajROKSlCC
+t+ieNy3JMRDcUeqLB7S5T/l8ztBqUiJ4TuseRqLbhgeQ5itOkyt/ry1wW6ZZAZdsL8Xnv9L9zK3
ZbavnMRMKEM/WI/5+SfCn2oH1xhCjk4mTnr5gHO1RoDd112yOZaLoFpVllDGEWyN6mL3AWi+zpMi
85zGM4qfMc8at5vMOGBKSFMYtny6jq7748ZObowBawqTSC3pFH7JLskpxyqzAftTey8PCpRdYsha
F6bbdWN73CVzpwVSAjb2kc61/KWfSm81Gi93nRtwQ1plwkzsz4oDBsOHHLUJyq/6/1LOWhV0kzeZ
W3dKrAyMAKCm2Veagck86Ny1eYIDhnTKuQmWxFSL8ne1F1jyTZc8VgR9t6OmZBqBSLYannWVEFHV
eJjiOX3HOzqDVcMgJ75yb+hCi9oqpNL28Mcgtn1MbEbcgEPOE1cy+dSl8FCqiAN2afCGoyj2r89x
XJ8BI7FeABFoEkJgQpGrLsYbjEzgMYceMAxORgbSXOVOoQFatCnoocUf5J/p4OGXM9/Q36IkMR4Q
Q/xWBAxbRM5Nzn7l8LIEpxAtwFPy7MoopHEPFI7nhNMjE2Kk6zfcXA4eH9cvfTmGAe0bEE8hz8Eg
pRrrPEvDKbb/6CBZR25WTNpFkd6wRD8uCM8c2Lcmx6f94aYZs59seM2DI4ODxaN1M8tYbv6jAK6I
/dsrx40dn10Y2YCH78Bjqz+vBJ/W+M2E0bfIUsnnllxl4+hxl7GiXQLuk3si1p+yxihT4/bIp2Sx
OgMczWyhgs3QfPgumJGiAZpgxQoQTc17ioGF7Zys16KDlwOPEq52AedB4KKIalhb3nYSVoVvWc53
qPCcTtlDF6/19IA3tcLaeWDxCBtj1vJ+yQogULdWAQ9g55FQhceH/c1mr7ojhQj5klzuQZJo10ga
KU2SKwKlgXCj4Nx93Hm7iGT3rnsJBl2mLI9LgxMHyvddxpjeNkOJ+4fV/7eNKEhGiI/Vhx8HnkLq
78TL0JgYo+lBcNfEDB0I0xJ7eHhhN1B6SiW43i2bsy4YFXJCtJzCFM7G3jXpxklrCq+K1zmiN1TI
B2VvZRusnrjwNMtYge8WLEiNUDOAa65EJrC8wS/V38bzErnjahzyw6kEUYrTy3/yjs8/nku4qkLn
M7a0hKEhDLWwZbVPYJSkkqh2mBaI2HnR7oGbxq9mMDGXwxselGh7pNFe4uyAGpipmF+Z9JGACcfv
KeulAQQx6f/ZrIOIdFZ4zcXnLFZzgZCDDxn9Sqp6LLAobaxluooLYETd95HlBJwIV5S/gDPLjo8e
mbiqtMGs1S7U8i71p77Sgwx+aTdBYxbcIBfdOrybKj4EnbHgu10A+gY4yveCKNbku/+u6hRHKjDV
0PEh9RNUXM7O1iBSinfaGCx8+qtr2C0Z2jq4th58jJwD9SjcBFgk0MDiUYR+KJqgAv9zXGrnZOAj
5XNaVOpogcFmBXJAH7vf9Iuf8xMuGHNY+tJnf7smtOTyaR8uT4eGwOyEYn8gcU+Xwl8NjjxN8o6a
P3cGUfm2QR+PHfDdrFg5cCDdeCxIW815bioQ6dcM4Imm2WLm4lzz0LswxVQjUmzvgetzVik/BiTy
wEfiHCJ7m9r6INK9J5JdXx7586iNJodAmURv4V17NZ2tClAfM380KQaIDKC2dBmAeEzyooLFk4Pl
nA3wXYNvCVIB5jpCxuT/ULwg+BiDO4NrtUA6Sz30VtljTHnmJ9xWW4qpot8ZqYaKWQFQdrHCa/x3
dl4v7g23MlzcVhfJRJGFHX8giG1wiLtEvZ9xK6auTIJmAnNWLsHlc5nC5ZbAZOWJtPu63o+H4LvC
YMwyU0KMKCKgMVGCTirw3ARxY2kceSho5xKLpVC3hoNGRid2X/NFn6M2c1k39nClQwo8Uh1h/tT+
MKBR1btVe67dEGVeFUe4OvY/vNeyY6d/eSI6bcwWXMCg1PLQuKJa6t03Ok/XgcUmypJpVuJ98NXD
puRawN2bvpX/7PJIrq/muBNceLwlfiDeicwsgkxSNFXm8RtNSup+VmC+yhitM7CbivAxJW25j17Y
AOn816g0rdkB/TrTPEIfjy9Qqf8/dgEVqKY0MBwKZ1MkVX+YF+eQ4crmbFywH/EGHwR8af5oUYIY
1GqV67uj1KI6Qrm/Arn8FO7K1M+cNVPCKk+iRW8QxyYxKLKHobpTmS4/XGJ7GDsyDeK3wE6PA4QO
rQw75BxW/VkKMwT14GRCfuIrLsdUu6ah+EZZsJK7bzjAE+HeR3SwG3/XXFMYQm77+/4ix2Q+1p3d
Czotq0ZurrOIccN4WUMHzFknFYFQS+1giFJwGdUIze6Gq5azuCw6vgnTbgNErl1h+kQIpWHQQNAe
vKDmNQ8ohJAzgWccs7xwX35I94C0DlRioJ+7cJqq5NpvZ4MJIu1IZ3JjP5cO7NjWxSDNFZO1qh9z
cMqtmuW0bw1Z+3/jcI0nAYDSfQtoJ1LPwoxO242Sw1MBxDAF93JsjVEvWNzpciKQz1kLoNa8uG+C
HYn69ecJp2MNZWfrv33lBjtJIMVzPkEF8dkjhfL1ga7AOY918L1OTAtUHruKBORnc8Wl+EQ++qk6
OhJvVAFqxHgc18WfBhwNgVp5vTJTwuKtp93Ok9fd197mmzjFdQMoJtTMU830gNhec2oLo9QIfOY3
vHYsLlWjIzhxwQPRIjOzmvwWM/MjlT4E4wfq1HHPaQAP8uVI1Sh/ka0bdtWa5Flh4HHDVefpNrqk
vqKanBmek16fhv24AyXlS3jP2Tq6z2vtZY/iWQneONH+BXZjzjYRyaTmUBfgXaMHgQQz57p5Lieq
0raXTXoB5xcsaKjUgjRHig6/kUIq16ZjyHmbggizRfwKEKtuTAqNrPuPBWXrnN/piHv5J42OCybU
KIvOjc1hYE9FobRG6T/okMH4oMqCKSBCOe2byTiJEmPRMe1fPhG+voiZCDYf/Gn2JzLl3RZ0QMXa
AAZJzODMFS+qE+sPNw0aBrLPc+5rtIvfAPDY5VNFV19mYywZVirLjitWL273vSOE7DHLvgHeoaRR
uFrmQC/o9hmZnVp+U4hiSorfNaHg9WIo0+LmQcKX4/HeNCUJ/a0NDyqM91yywta/BrbSHyoGPpm2
kKC0ND8CVfytEsm6LD3Wq+WeF8P4E+cBCz5rJ+vWDZp9nRtVpedIv6Rx56vOCdwS2ErgsPQ0zbd7
VNv/0vEdFK6NYJqYsEjloU2V66zLzDzGRqf6CN5mNi7WguDaG2jUUzTIWT2fYNkxsyyrigBd3foy
suwxJDdY7cVDEXTh8yOmSm8ZnvD+pQVukM+lnaADB0L3p8tTeV62Qc/hH9wW8tMCHg2WrKvs5qVc
ic5699cmRhK1przoFI4GnC7DA1zCTinDOdwjfAJzKMKlMXqssJpw5Cbnl8rhTCXvaO8ikjvUkazo
5YcdoniVKh+WqHEiCDU+MLPNJoZfNRFGQ0sXNg2s2ObW6mRNmrAQAJ5iyDQeng31R8LzDPRhgiJ8
x/lxDONdt1EtDIY4PJd+S+fLGxqDOrGW9gxjCLrutauA6C8v2O3BvZvZIGcnHE9i3i5T6QmThkZ4
PD0i2b48x8EdD30Kh6/LLI3gy4QyNilXqtB1vXURhDYhuQ6xLHBkWMi7ijUhBh/bzXSmRVudUEnB
+lbixRpiVymFtNV5tLjeth31SMn2MYLwcChaIKtiUdq/bs/rZjSzT4Vxi9Ci5IeI5EI17UdGdEZ9
YJTkU7Afx38NrvkVmLLKLR3L/sucCo1s+DoelV+ENSWny/7DhKQ3WUMvFpPYnGSMbu3hebLLbGtV
uVXSy+kVzh+tSqNdEbjWScGoxM5SnaaJBPEikvpCUI6bM6YGs3YBwQDiiBy/uH/2EOzXJtBy8CYb
kKWldogawsARQF397Pb+Uk2yi95khXUImQ7QZt2sQowhTYgchcgGlppQnroA+Gktv/ZqOGD0eFVn
S997y08EP5JtnZEqxvsVnIV3lyXo5ccARjZe9nQj5yqsv7nivYjDOT8S74ut1doO2IL1DI8oTzEA
tkqCzBjC/8ZNkcmjzvSAW7gWWRfs0KknwGSV3dV0bvJCgK/s6isEizcPwe0U8VKG/1Oamtnoja20
nORXYjP1fQIsfnscFiqbnD9OEfq/C6zEmeEdcnB4iugFsYaQbbFOl9yXHq9ivOqrqgHK6AMblFhk
0rLaThk2lLHmzYY1dFpg1StCrwyTqCcEp5TFn2Z7NFqm0wfQ+eZBCTfOctDaZNqOL9fa5L1JwSM0
HAlOUM6gUVWT2e9Js7BGByo6Uc6BCtU0nzpm20T+jaj+/kNjmOWFnAsmw/t2hTPGX1E3FY8VhXO8
IQkY7B+6JiwA+dAwvRQa1X3AOtL1ang0u9t9dUPU8n1uoU2HYdZ0hYgbvWJN87wGCpJX1Yszhfyk
/5duzEspUD7JR3GpBZTcglj64adjDw+V9wR0WtXdAD5y4RyWQfCPeGEJSqdEXJpSlR5ojuU85rTV
v0oA0m6X6PIVaTkr20LvfuFQV6dkxzLNpDwFkU2pEYLzxVhVZ00uWFq/dQveD5BV+zBFlvk9/+xh
wzJeYtoLok3oXTAsVrSeLlwnCFChV1ziTukbGDgRHjvFevghO8NTRs363YwL+37kyv4ZaGq64t8/
xH+SyDW7OhemgaV4ZeSRlNcEnDfYAFC7hl/LPqi6UEBi2xST3P+z3dXhT59Ha79syBhZqzTj/8hL
HQHfZOKcUbQj8LILC8C3I5lfTsdsVBcez3nq8OIwg8wbMcOVlzqIrdM1s1i6HjMIPwQCJgajIUW8
5eL2OTukkXv6ZFKOKNdnuLk0gmqL1y9vYddggDFyyBZ7WUWrDis0em5ZrBvms7/VGUKr/vWIsm7L
7UCQVTiq2JzVyzPmFTWydKFG+K/PHRX+v6qj1cqbFjNBbfzls/GokY8Pdmlg64IPZoGoek+wRWMx
kfqsxOJPLsW74wNuUN6Rpd9OF35q5E1l3bvzLQ5Llqnxzc1TsGxRc7ZplGqB5Ti9ot7kpk89N7mU
MSnckGXGRkpTul08QkUwldo1LUEGwHWxTaPmHKizZ7wz/pi9BurpWamaOLidD5q2SkK/kCisF/jt
q/T1PNjgWzeFhAHqIXD6GZcaqPlT8UdSKhVUIE3LI3d2JwHTvKphGEN4BUJIKleGOYziCjWNHKW/
MiFNFe4/tYHnPUQZV5M7si57lWaVmSOa7PbxAT4cTcPQK/ULAi2j1/FhissjdYUHaaBdvO+mZrwU
g98eeC5MTnmiU2yG58Lkn1Or0y7p2A864/pKguriDYAw/BpxbGBc1OW9halMbWU4o7Y8W0iid7I6
gj11sdc2eQSD6CyWuXRUYJXWuYtMWitS/h0bN4zKKYoHyN+Pb26auyiqdllX7noVI+nkNYMqG3Q7
u85cvl5MkdkR+Ur0oQD2oRVw9fm2wibdeXmpfHoRSTn2UW9rRFI/hwEsPslFI/+IX0IRa+9Oos2E
DExWjv+R3Fmh4CWcT0cUP34g41pTBNlcHu9M8N68Ey3SvEUWhAOXPCjD+sYSOIwnPo/2MgPzMVgU
KLKk+7lsgCsFK3hyKhrOtEtZj9OwTL4hPKJ72dGqFVnZ48SHeO8z5Z3WdkRn1WKk8c5+D6LnGUMY
XNmYE3H5NWI2OfwdHEUl9A8sYk/eywRnm9gnRkCiR2dWDXmUNhj7ettaWkjGW3cDFD1dV0OCM3ey
ZrQcxdpNFQRyXLozsy0Nd9ktTUNEsdCNLILPpuSfMZqkehQXZChD6ER2cYtRFnMFPOaShl36PK/R
mkLgyTkvEPJD3NED5s57mZXFbe3F6vy6AJMDEvl7Na+RBIUSPYUV4yVcs5PGrbNyovc2H+ELiJLw
zyqK29iw1wZd8HiKZUrGoiMABVyPcufnDgLFepXaXUGleQoofXfqpeVduhPRPeDUQq+KRlOcnaAN
7jPvGrB0ch02qhAkjqyirQ510ylnaq+PN007IS2zHAA+iCSYZzhxnormLDnGWOlXw75qd/s9gD+g
AaO7JJ+UUqjPc9Eem47RSA8a4zLLjq+T7JLdOGSJ8rf0OkSb/KN7lmAznQWE4pNekS6E+ZFuiUT/
asN2nsgV5drYLVt5eg8SO7SnXuEQxeMCmxvw67IIyJoRDWUSpr5mMlXmvmd5Xt+Lp3ZWjRikV8Dw
wXsuGeSfGkKfZFy30EvYzqScTYnsOoMiH70ZGrTar97ii5CVsIPYNB71OL8MUTSfUYHCuT+sgrDZ
Fooux9MfHtEiNHvvA52JT/jQwBYpd0knHfOCEkXAPWe6zwF7WU3ELwThPGEOYN6y505n9idXaeVa
Z/S8cphKf6miE4gthx+RfNjETwOOLANxOUGZYjScfxUdLarwTopf0/GGdmsDaewKuWBV5o+2Wl3B
1386V6lGy0sAb7TOCdTXVeXEl+zQOJwnPH49DkGGGkDI10F9QdtPGaQVWUsShm/39VnCQtirBgyD
WAPFxroggZtU7A/sE8GjWPmtM8XHaXzMDyd5s9nc+NcCWIpeSQcvqHBCofv9FT8iUOuLiTmHNEDE
rj2l+9oohyvgzahWhLkGg/3+YDio9mCfCwgmLNL3TEzCo+2SLuRLKTPzIRWkZS0RpHvYwU/XEG0a
ap3Uppaft29R1+PdBYiCR572t928GmJlfkhKgY92muQaKTd0A0T+znNR8h84Kte3P6HhI+k3xppq
XZuId5ZODFzjCwedspAByDQPkZtomzpB0a6uqDUh8mhPpbUKZPPC/PGyxQoTlKdhKVD8PZYPICoU
1UCBxWeLQKOL+CDggK8/rrGKZ2OUSMeH/L6jNrGWrRmT3ebzi4VU4fkVhVPorFvOUhqubXPu/5UU
9aSErMth7NKjstJvhw/77Yt8PjjIe/G7MnAp7hArYhgzT07l/uxUcZkhTvrLH3nWNJhapUzThDaj
ZY4TdzokqF0kpmnXMJ8XQagg5q/XnkAigJUnztXFUC4WbT/+hjio21W5ol9OqgJBwLE6RL9XQaqx
eoQFlVU/X6yrDczHNT0mQZUJ65jgfHiZwyMFTZfiYPWfbqSDo0XpXCby40ZWPckVt9Fe1wcjq1Ji
wPh/ABMICfw+eOhzeNBOK+V/YU939dvaqRrU6Z1lo/Myj1rwpElQDChWsbI2TfnTH7BUGOJudhD+
c4jqF1V5ZY0bds5486jF1CMz0rjuFIO3JVEiplm1Ptq0crqQ0AahQJq+H0o0MFtd/wUH7VFDmkN5
i95Os/KQG9NcsozJwpASmbZCX1Y8m8CLH7+k1hW5p6kDtRDb1O5l90UFciWjps1X1usa8hZKx72v
v4EJHlIBkL33s8ZXQYxYFPZf8UOIab9wiHeAQFSzDEvGsHkFVLr8DJ0dM6JgIpK74w5CgoulQih2
IDo4f888gtg1/qV/CJ2FZEhP4TBENt+nro00IH4kJeqMWQleTFL8gysnEGxjBQ37Pche3KHTXMQ3
jRFMfLmup5k9t1HfFhnlyD3Df/zCbrWIgBLdZ/VsCqVle5aS5055HlNQaxLwAT8F1NwKSEn/O0nT
+oYFgePtSMPUzLjJ5cvcF63DuAMJoAbY12nt3TDMMSeu1klgYAv1YwiETm/izCXwj0cmpxcIkCXX
ykZSk60eX9MGsYr1TgYl/w7Fd8eAjM4osyJjM7uRZQjEYY8B4qYvQBIowSYZWcoBQF1Zy883zQAk
Y0cgHPXQ4CKRjBssHFwPeXrI0MBdRQFVmfG0q/3x+s+d6CewbPG1aiIwlnsEfsxKwHOQM/UyjPqm
0apIYkWbmpuG7CihU250Gys9aEzwcMaCWbMxjfepM77lZjCyUTzlF6bbByqL/cOdcVvlkNrmnIXn
cvGUBMwP0yfgXWac2nF2L+N7lpaS0ijvLP3xuuULuNN7a8BgN0FhZUQYm+4+3rN+lALooL7zNsbZ
D7H8BcLSAXlfF6FtvyadeUz4YqmgYkqm1eaU4y80lMfWIDwNQJnp5QQ4HfqwfOZqZWB6BaJJRBD8
/Ypw3gSRF2AUtlZPHYdF1EYbfTTOPXyh0GkBnVB1BL8IOsu7TvFPpQofCv9gZwDYo6ODXLswh30O
6YtbZlx3PHialt2zoFYqKovQPlBwek2+/aDZxmOJY5jM80XLTT9HERpr8jOTTf8GCKO3noxOgANv
alubgwmiPPf8Apeugsfv0+FDtOuS45F6vFTJ1gBZhx4pJ3L/rw17J1O7JZ/M5BkkJMuQCV3mHfYk
I4jjfIT8uTPYEtkLQLjNKYO4nQfL1RZ9GlPCxO3+jyS0KCawH3N/NUnP8mxKxHMg1LWuVHO3OX3p
/zO5QVQixChtRXyOxP15Pc71nIq9Y0rwp4iK1nBRDrgLR4YqEA3zomiH8IPfQFWwBKjlIsBDpKHK
wKPDfZT9zGUmubVcoAzsl/QlkK8pvIWyO117T6Fy/DaYTThksuSyjUdM9q+QRgyXiY4puWdSftS5
enn1jIMrhdWBqIuqpBbo/ibVfVE7lr1YSqjmYXC6PE3MUwQs/wm/jPFkSnAoku5UeY1r9qI9xSLH
JO9dSl32CVsTDp6Y6mlqbTV3Mda5Z215KIQalAHldfitUQfgLed8Q4fdVVdjr5sfsi55gw8zfDzl
3YRsuKnv2P7uEqWcsS3TZsUez5Fg8js3H+qausmOI5orgR2fFOQje1V+3C9BCTdtwCLI6DT7OwaY
08/R3CqHhBtvNJaAAB5lo/U3UeeBNrlF9ltN/4+pvqcPCDt7r8NZJbuCl2QHzStm9P9srfZ5UbIN
0sPsiVy5kJjLOQlzkFLcOey16EPfZpHSF/LpheK0DIgml3Vcr0u2AQ+48RyAh3be77L1F/hPKdM7
4dvZbFuruGjr9Zj09xwt6ohdyQsKLwsUolko3QKwXoAZdccwKRyNafRUABmaeQruDn0KsiA943p5
QnpevdwuFjTk3chvT3S/eRK1xFTaEeIAOnCTnb9TDwpK1XS1HXSIf9oNUIts3z9cTBZqR752CHvO
fFkJKTu2dSsJdXdCuLmCasqo/MKfrXXDfATD4Q5zMqgf2zEpzXEK+mODeyuWXZ0ebUP3o8kay4ba
gY1B0h6qFWgewAUrViPcMG6izjMkB6lTxk3i5GWcvcw3zUYWomKepWQS0h8bcvjUA0sVDLJn+cVT
JXcSrDSA+7ikQSSvNuEPKNhESb7V9xZOzM7X7hEQRx+FV2kmZRAQK4tW6aMFMenWpk1I25h7JXlx
rQux5tb3CPypvMFMR2ZBYQ6zfm2zqv11jDkkeAMNNkYU91bgPoVzl74azu6KkbrtHC+SwijOkDOB
fhP9GVTNYWE+AK2cq7iQVoSc2UQKdxYLLGlcNr1zzqhmbF9XU8L06MV62qJUC1LiADZDg2TGINQf
7jJolBdsUqGfx//4oS0MF9ukcVoxK1s0y0/9GjSLr/xx7gIadblg/EG1duefqveu9PEGHw1N8nGk
tzGktXYb4I6NGvs+lxZaFqYId3Gg8JfNBy4dU67iUwZiZxUfpwIXUP+oA9+6ZJoJkLSSWZIH1gko
7ftVo0LYwX6cO2chIvgTbvXsuKVvwHRI2CRH8XhZv1sHGz01F+oZV2TWapIToPsn6gRz40z2XpNC
5QwgjmHaNbliw2mlbIDv9GO7PfMXbLO/ioV36WH8bp3toTuSSkWK39GlboZVMqsXm5+pmxhRw2/c
KkPqc+gC6efQSzlQcUxS8dGZTc5RQ51hB9uk1MfPLPNN+7y9V+UOqJQIFQhzEUkBsSeAAr3SpgSa
noS72nVZmdf+NzR6//+oePViqPnXrQ0HiyQGYm8KLCSyokndRHoegNiCR4EW9arMy7ViUX3osrOu
bCUt1QtixSZ/s89kivzdo8DLRN5UkPEm99j2bWP2bTKFxrXlSyUaMUqoyGswez02n/Az/g5wBf1c
XDdDQiKrbvAYTC4MllZHilzm7vCDknxy0kgLmUiKgSZfocGOlFSF/Fz8I6WXaSBrcdpHeYo+yyr8
IOEdc38/b3nNSw9UyNxU1RKxsG/HHRhZHtM8sTHVaQzOPV+K0HwnyHJYRECqJduNKA9KRWLAUK2S
2IsQAaLpzqXYHl4m8q3mO6qNSxe4oQY3L9JDX2NfndZxRY4BVD75hE5wkOBKPAfjhfwqcx8+9WCf
qa9zJAR7H3BIMli46+spninAPg0QHJN9CQjjGCy46IwcoN0n0C4wgqXF52MD6jXqSMnMOHxiYeum
zvobWXqL2h6kZbksnv2hCF9a3ORZxpHYDbQ9aT8Y1RFc4CNXsQykJX2sfSTojf02NbK+XSIiT6q/
AR64t1M0lrY6XR2XvMM6UKfyvuIiQYpae8Nam7QgxTklydRtK6UbwnS26trBb4CWbjNEWalYGAKj
E4zEqt9fN0hSM3RJwK1E7oNJ/hc1MBkgXZuKoNq/a5q+gE8KBnB9rAwWw5fq5LHxPE4LH8mGz3tz
gLoly/M5CdrJ4Am+epHDgJBPKvFvTsTLbiwRipZ77rwXsTGYl/UZmyg7AP/+xNkbSKCQqIiwvf/m
622Pw2IT9FLasa54n3e0NFqV4X1B/k73e35DLoJ8Hsa1sZ30cChbqPS0v06B2eEajOgc34CZYUuc
MdMFxNQLOkKMR+M3mVhF00LyiHvgzW6PbwgDkUd0REKsueFQbWLqOW31V/80Y/CC7TlYzal64TK8
pe3QR7NdSIutMilQPsQSTEWbC1/9qc/Q/Ejtcwv+Nx99NOL9XBcQOiEknBUmq938HG0GqcvJlJAR
asFv54dXEwkCFv2kQvaJ3IZnVkjIGqfwGEAz7MLm1xeIxMZ0qyJm0f8cguLKSxW6xmrvSHBqwfj7
cmlZGYPFKTbpGE6JhmT4bAgUutgLN6VhpyiIuV+wm5oOABFfVQUdJ9lC6OH+gYmZnZPFU4mg2+tP
k8net/vlA09LEJ2nrSj3QVhitIApvixbMFnqpzRAjctDGaFjR6mhPkLhtHgyd2YgUj5psoMtbQu7
VzNHqebgL/Yr12eG0NJmv8FQwkbnbDnfXD6Ves8ASyp/C+fWHJAabwO2X2n9fUoJSahGSeP7e39G
B9s0DuActPOL2tfT2dH8oiDto/XZtyQ35PBglUNkeJirCX44dhVYWahjHk9z1I3buMWoWio2RDPL
zBTtfrzvbk19Sgkz1mbjDchSqBn+9hRgX4pd6r+1Wp0cg/pG/Hbq7Das3Ucde1l20Al7OhsMWhHH
X+jF/2tX8tg0cTWvHw3g85Hh7zMTeLnt9i7EwgZm1172ePnQ3MMkBVGTL+wwOOjYBo0plUtperRH
3DbdNOo99kEECDXgEZkl4o3L3NgBWKFYFrmqIh/8znz2sSZOenExf0UKhyEvuiRunVanxtbLIP3r
3McSeGwgaiZZM5M9yz2Zv1x7DLXzcg/iJCtUa4LSOvcfg+bt7kU6gDvBCm2wY8ScpQAWlAQangiq
B5UDU2Lj8PrFJTVaA0X2webP9NKD4qtYiLOR+lnduBoP9bNZJaxEKAAA+EgfF9ieNYj9/hTapM1L
zq5Wqh7R3oTcEnQ8aw06pHAZMRW1iHP8lBv4m6C5IC/+Dr2Ym3RFMTdYCcIhqYiiY+E7Mu/VoqOM
sICYa7R3GaTjuu1SQHjhWSbJdn/Wdgb1TekIT9tYcjW/Gpt/UI44AtwK10GYx2EEO+77p5K4E5/Y
/J1aEWugfyGh/T8i4A1HHgQ9zn14fmcBblyBZZ03Jg0qUPVMenMPuqdgMeaQTJHe4JAZhJQ5DEHP
LoYCQSWMPYWP8u/fBc1gqe1U0q6cYX5zML2An4B1TIT+Ki9nb+UMOsNial+bEmyRtyE8X8NfJO0X
w/YPTJlvJAFoANFfrwPiYdMfGxY6D86duDb+OPItGxLR0T3sbNdAv5cFyvxmoY1HOMY9dhYyv+6D
MDcEdpXt34cPVjuAF7tN/a2GKvF/fO09oviFO28wEp9jS0YFkyul8EQzqeFXEODkz0JMWaDyA5Rj
jeLrb+7bxiwMv+ikgJWuYnhTS/T8S1uXMBPQ1IxX36HGudNdlyMDYWL7p676GkIz+7yJHmBIxsJH
IebB5MBNb/3FBeoD9kMWxFpPUbuU8km883Zg0a8Zn1JFlAaOxS944MlB1sfdiBoFdaWn8BKiJ5eG
imPI39Nrk+DkB1rvhhgi4x62+Th/Qs19ybl//eSczcXplAlbqJJJ1rCDWev6EsM/lNrSUOUmBfvZ
Z1ECAp4gavdGw7M6m0+w24CSXtbFJNynzoKPQuJzVSpyx5WI8BsMLCXvcK4o2jooW2ZYnbyB9cgK
gKKhWH6EHcQpNYPEhSbkXkZe4MpD917N+QejwhdWMPUduEuAOZOLwvnhkX/vO0eRMF4DGOyNcz/x
GL6fsy07z/epNHrtGkdkNQIjrg1oP87xL22A0MVsMgl/OkWf98TpYuQnnmPL0Xg6ir0v/fEBODJw
RmlZJqbGucmyMeTeO84lSO9h5HcE4rO0kPpaevG4WMp9PR6DL5tIFGA8yMxUjNOR9AOzpHR2xC5c
vWDo4M1di4iK9U+1z53co2tDTwjQwhfrqVc44jNKdasR8Dyyp21s6hlO7T1uKkrP3rDAT44DBusL
kky90XyCnP0rPiqPbggGjCdW7aVNDcke39JUKplgnOdnLobNeFwHFbXc30H2CCMKWSTRJBkaMEXF
s/7NyK/23xk4Khwmh0VNSYHxjXFKuVTNpdyCCmkC0lTagYTbvqSyWJMzIgs4/M4I+T9kvZYlyUtg
wfGW63LbfWqxO08YY4+McqO0fSf0gpOsYOT/aryUPD97IqfNtqUrzgml6YFlxASQu7G7GvQkL5vR
QTsxzrtfNy3GJub9fHM0G9+3L4uBg32lTMoa3rH6fU5y1rzp88mNC7yQfLigQOE4op9Ee+SZjArE
KP5Qz/0DIMZpY80/auu7QgGkrmWERQ6hoLqNXUG6Cl+bRJJswPVEPXC1dj3837gzLATsQ5YHChWL
uJSUx9o992fyDNloGvT9xdXzT+Nfvh9GZyYgSa8g7yGNertLPyqP40S0II8v1AgVal6Pt0l1+FLq
0oGmr1e8xD346RgGDBlOF1bYPFD9yHDPCh6aLBInHBeVen342eSYwOMONI6E85CIw4ISo0Rnehm2
WqUBQZKtLDuA6yWtq8vdA0eJG0ZzaVeKwt27wcOxGcWSkoHtp4TpnuvgpDOCnHLqCNPwTrlwc+UJ
q1EHBMssF2kVb0LM8OdI1oC6cSkCbLBvhy8pKOt3ZmVWTKcs1vd1PxHKOPcEVhetvOtf/5wJrLEY
lOexC+JIEE+XvbwhgJ6XhMuf73QorU9bFDo+ci8/b7q3iWs0tbzubuNWKZIHvpJkfilS1lVGo9vC
ryKdpvwaeegfKUEZspJGQg4FTVtxdV8MXgckIN/BQ1HneALI+7ZbOis2nwMs0lHaNCQ1vw216Sfp
LQe7aYoAZzSNIpu4+SpVbstCV6hoAN7mhFkUSPq4sz7TLBgj2X3IXaDrRvSgowSvQZgPyA9oONIQ
Lb7BTrUivQfs0sXrlZuozTTLoiqsTEvRKKjhpvdYpxuMEphDrMoRgVSNUYiRQuUGN9D0WzeTAj9Z
/Q8JJUEFwSlqumAcb7lC9QRf4NUxgd+TojS6nB2kYyf3siu+9O4kpPGtDD6ipSiWajY9pceQ7c8S
0oO5fTF8xSwI5ilh6HCGIi6ZpHTrK16/1g8y2LEt4Sjyxr5ZzTaUlPgoeSyBghShRDwo+PBLpoUM
FHo0HqpeJf5E0swIDjEl1WTAHFBbx/QDERcwynduWbsKdrsiqAY9YNcZMiHyP0sp4T6uEo+FPVnF
G3EEF3vWODeAe3CZVxAyy3Be8DQH3VS9n55VZF7ZHm8Bd2e0iUplsL/yUx2jlilOfNYqzU3VH4Pt
vjuUtujwiiNfmIm/o6o24F99cfNIEzFk5splIV4ClKRMsEu1gyx7zXfNx6YT04HiZwfXaRSxrO1V
Tq7mMZDU23ON94iRQMAl3Jlnz9Zd81gAaVqlFoOZQd3MaJgs6pGmhLK9mxZNKIYIS+bj+ZTAG0i/
qRb0GLfCJyRL/YESvvq+QWo0rWOl/bQbqL4/GnZuY83H8A2zrwBsYjQHsxbml7P/n4yAKuwXilNA
wwhSfB/OyGFs2xQaOwRSX4UyAXulwDOx9bCaRgYaUf0cQr1MjEr28OyougjVzSeCUzttMJ3PxkEI
jNBmd+j8EiYImo+xAZVZSrI8cAPIpnysLPIBJ095diFFWHZUYXy5GhojIgM3AUXcHAh0sIf/0zxw
KoDcCPCNVxOzw621BsT4taT3QP1LU+HlbTxd+8bX9OmSlA2wVLlRIw/H9DaOCAJdGRGhizH1l1vr
backjqH0iEkxolUZtqz9xv5NkwK4u9VNXIGcE8mn2CgMV4KUpzwVywOZxRIbp5evg9B6jh7HcS+Z
Rt/wqY0WQZYhwbptSlGHU53UpyLBzdTPK836vOt8vPRLnaRsYZsAoLISKAtvxJSIl8pPe7iAOKVA
UfH7QGOoRTHL2cfOClcKTm52YHaVqFVTtitbYClpW41UexIX82tziaoRY21D7q/2+EeFFEIJcc+W
39E6gogVZcRnbONRld1/HJ5Ge0QFdQ7j2BlEnLXH9Caany3gVGQoSetA/DV1b5d0vyJuLru7glHX
TYXVpONWA7vuu8JPV6/5FlfQ5nBqdM1qLBqIGEiWn1cu0q+9UuQ6VybSb5heNpv4NhjTkeJsCf0k
+EAq8A6GyLwOiyPGyUvUW0K1mH+lYZL8NMQsHU1MdhV7sarQvL0OMW/JKAkKmxH10mWXBuqbO1eF
CXRksB6teGjx4EbuHf4P56IwMkZuisYDW+DCbhSoWIz0sl7x6cT7hIHqyUVFohIZ9bjyk4jfxa+I
Mt4h+Qg2ymuZKGV5tMF/ExI5kYMwBr3bL5htqMc2HD2b2ZEhVJhb8OnGFy/eOfNAMhHDb/uM1KNq
DK2A0BD4Pld9z3DANfCgsctGnAe6qn+xYGqMTUg2LEvABMA8AtFWvkIyzRAeqBpFEK5Mk+rGBpD8
vhAaHw/0Y016bNhvWSA1oEBWXlEm6+jnrB022nhC8Bgj85Vvh+UBN6O3uQqf7gSFeEJRqf7trJVo
PIck8xIdQKuDuNKCUW6+ThllBpOTH5AiZbZ9HxspAbJqholQatmETN+/EACHiCA2mRbUaOvwT9vG
oJysaUxyavHbbuEOsIJONE0iarB2AHr9j0qnyEqh2M1721iMwrwd8vdJJURjw8r6dnghPa76uW5R
WGAQRGDR96rn+srz2ikxHrziuVBrR6tTqC13HPhaWVxJAT7wb+gCPzDOgonEqlqSjRegiuh07hOv
CON/e9aUKlKPmnFUsGr6zjco5oM24cFDUyAmdaAIL/noVyZoU/jEgZziYH6dPDhEwS2th/DgEvuv
oZOEdaYlLrBIcDrLaaiZacMtnbgoMmAcRtS5U3DIaTN/sSc0towzeGZsKBmS35Ux9fAle8HupLus
wfzXsG71dzBI8H5CVD4xN+xcuFBSLm70YhtK6P4cWiSRWbm7oKjq32+lNxL8jn1sPKcjIt6zddv/
f8a4qx0lJyZDtvh+vzmY5WVk9YLxDheMG+B3eNOiNh3E8tkDn8qaTt7wAfwCd25Nl/L6z/AMRzvO
a8goU+AJk8RxiTdHYnMEkRuX439ZdxN3DBA9whjfi++W6mwStuI1Kn0S9ZPsOfaBrsSrJb4JV4uH
i7QmIv8EFWedrXCWEp71N0PUNOT8alCnjccT7YOG0KJmArCpvWYVgbJaCwdoE79g0NgfbwSU4OsF
459eW9g8x/Jo/mguOEFizFvdOtnhudRvvfRYidxlHY4EV7iQfR5sgF2hUCXhqxaW3ElqSwAZq1hq
qvYM/xg9svVPFnJUt7g60VivcwwwTu1s452E5jNk5XXjskAvtuGTYra5TGUvCx1uk4GPrK9bHcFq
0wosTMTjT0+H/pV8QL+z3QqfjQmDnk1LbMPsdyLs/PIOOhm7gtONOekf78K5TFGRXUoQ2kW+rrRn
KhDaVR15HJIEDL+++i84V67Ck9vvF/mbQqqjcP4jDoKRrZlEKDKcqKfg+JtBPgUfOn7GVJzajA5C
uaoHIDSbiN9g0IgzHymZf6knZZ4l4AmFmcntg8G7AYyAmz7Sq0ugHBTE50vRcDBlCmVKCFQTOXE8
Y3KGsOkG87Ehef2afpQegUWzOFL0Vwe/7qYKuad54zwRlfyIEatg7mqLO4atpGZzytmgAOvEqUyn
XuVg28JJxNL7BUAHASyA2bNJIAxF6LBLzxJVgm4TU447tmPoq61KViMrl7a/ZU5hwqM2399gX5dF
WK+U6xqLOZszBWtYg4G1WhS0gtMlI+uUDj0ejXQLeBjB6uUpnFOEuZBGYm2ebNMdhwWtkDuBwga7
/7Fo7xo16TCn/SzzN9WEYlspvbBYg3ycPLxM4iDrTnaiTYuU4+rQBMZoEreqCRvFWdGaUZ7HW2M8
HU6h4Zhz0lIGl6J0rdZOdZ8o4o0MNj07VIBH+7V7R3twuCgdRXJjGYoI9X0Jmrlm2UwJQqdFYXiu
U0buE5o/CzvgGrDusEcZYB5Si/seC3q3PX4rxW/EfeJ8ghrmaFEo23M7wO4IvE89OTkysfEuC8kS
cxbZ1SDNF6S56pjIHFW7B5aG2G2SuSPoz1GmWh/Vgpk80Ovf/jxMSEwJ3TVQP+nHRd7TNHXrqhfw
VpLrZ9eu9O1wKrjjzN+37pZfZ/Rl9nrtOXQsXH62cA9xOl3XqV6EGsWGwiUyx8KxrYp1h/JL4bnp
GqLsfYE+a67XjQu2gunrn/qkgIR+aFa+wBSp/isWzhf/PlHFfZp3z9hQFY9N9Ly3IhIaXW9vUL2O
tZolavQzqN2UcEt48j1/3RdsyEWUTeqDaZ7zNMn/KxHu368vGvYCMxhWykIXzdBsAlcGapnuHUWe
rJ4dHzds097DBFiFpu0QswwdBlUJqM6nj8wZrFqC6RpZDetxVRfBj0q4BA+1xHIydXqLtY65tauL
+V5tMnJewLrtYuWOaoXeDEQQ6/paqlPkG27FxkZ9+D8hU1MqQodCS8RLFyNKiMprqVhca4uPRl0G
bnmai35JUrg2W0UxQAFb2z7P4LGiSIvUi25NA4YiHUjI+uMgdfzKt+T1SHFEKa0nKq6+BMtNcznF
YIevuAYvbUKYWlEwCxzrbrSgscFwNaqUCJqxs+/YsVqSfn3/pBJu5cI3GhVD4FgAnwSwfnjaFCWA
T66VWBvX3ZAjPgqK14ZZ31cu4sDhWoIJXCIcunXRKypnyjyNzuCqNI7VJiR9nsCPK4xe3Faq7vQD
BGdY1hiOLtLHGMAmPfz57UrCGEFL824jek5TMWieCC+9Mj1JZSS2uoYgj5AurUsici8U8C2jnEUj
6ItQXEpumE1kCBpK+97LLDEcK0R6/UeGQFDAuI6SD8cS4L1veKRPbWa9jahvSvjWIA+XLwY1dLg5
Uj7thT5FbjQn3ehJOE6u3p+GVSstZEYMDvO4LmE21jUx2Ggk4C/e6zPSojfQkubVx307d0Mqe0bS
Ph1dMrowZVZ+DfcEny/aPassWzffqW3bi876/1tkcQiUEryMv14cxx99y+XeM23rLeyDWjr4hk3+
tBLls/yjEYbdLbEkZx9072fIpR56YSLSbLOI9B4Ojcf3R1ogWyKIrw9EzaBaDX3HGmkPTXf5Nqpa
JO1DtO/mhc2KKJuRksobZeWYr75AEGPZNylUNODKT8ctLThAUC9L8dgGkszPKwFWqP6Zt0f3Rqf3
8z8XZrQG5lpSjFsIuyDAik52rIxpJTuENOARAsLQAfMWq61uCHjPmZRQbnOvVCRrY2qnmqwFBeLq
ROny1ZeJbk50D5pcsmF/9xeQM7hOcQS2Claa/KACDPNOMc2sUjSdxO/dqc1U7CTu6h/QQa/txyPg
JuSkQuglN9o8aeiIcG4/BamG5IIvFFeiQLuIzVXk84f5vK4L3DrgZwKAQviY6eG5l4XAl7Aq2W80
nUJL21N6knr3eLFF5Ps75vq1SKM4WQ0wN0P6WV5Wxaptc7oxylJTJYw0KXYN2JiBeuwpR0Nk/yTz
Y0E+Qk0ievrxhEFq3SPl3m2V2DEXRGbLL4DbNgGg0BvOJvt1f0uXuiSEinE7bHDhHYc8TbZo6t/8
4dtJuVqhO1IJsbbQIJ1tzQglM2y33cbBOie+U7byBbSqkwSn/1E5/6/gqtuKFKgdSgaroi4CZKxr
dE5eb1DKckB+9ycSkQyoOk0vgIPucLCkI/aW2KKX4BuYU3HLZrgPqR4men3+OXUlGp26xrIg2/JW
Pn/ysUC23csNaLC+jyoDaKIj7QG6xQoAJaAKKNtjLPZTCbUTHq5wqdd8JG+u6rN6ea95VAWhzfAw
UCch9RFxOAKnA3loWBdplqQTpk1mEt3X7aceMFZ/XssGh7XO0pD2bHmaq+CVCRnBVDBC0zkwKPGO
blfi/q/rRUYTiq7AE726iOVa3ZRh/9aUYyYPVMJhUIMrpbebRqVD5cona4AnI2rNiqX3dxSG988l
r5TyTpUDkvQgboXZOxMp0E6xAKgcCVl+brWDlg0wT/FdZOBA8htox7ssidCIV6vP6Whu2tKlHjoZ
5edwzqI+PXw7I9ezYouQtWiqKL476elC9OsnEZ8GyJA+S/c+E0YNezsZogsDet/C70LwjzeTkqcH
yjgmyX8BGLcXAflzWup2vVsXVFj8AeBMl7cfjMAkyPMT9fKNyTvE82bEXinDu2X0QUoNoN9fgo+6
QZBbQikcmXojpZFP4XlPI21D4Oe+q2UVE3ACNK/DYOKGqDxEpffiFrbmGZgCHscGDIZxgYmvPFd4
I4wiVr0Zsm8Atv/zwZ7V+NZQyNA3zElNkglzF+GL75ecpKQCoNtl4YrDiLdY9GcMozXfnNYFHaxZ
XW6VVsXIJr0WkPNz7Ys+wGjWfRiwF//eypRjuw/pxxnQzkCzydK3oIcBdyxAZV8O1MDO4VyAAKTL
INQyP+DMy9QNuWc1z669UQF1f28JsLd5RqVtc52AMM0ixQkOTymNt+ks8cTDS8xy37w1/fIenm7O
IXtfW+X8SKQpaiXlFpgddus3vBmoh/H7XlPuXqQr939XcvOBgetPIT95xvfFuDkAwr1IJEz53PWd
xlsVyARiSucbI/4qkOWEKjEhME55CNQLSwLXENKpUUOXcQ6BFEQVY5MEZ2GVe6KLlBHVSR+8glTK
ioHdGzmGCaDETwVwPq2K9LmDuF0BG85wNluwFaHgrWXEd95vJDZE1OPXv/Qk7ioXZdLvJ8cqb0y7
d1ewAlwvPNnCRmFAArU3M3To3Qai6eldTVvNHkurpY38XoZl6PQLpwBN+ydHdCumW8ciMXAHBOZO
u/q+vH+d+eXoJ6VCaaYpw5sXzUHyBNEONFgRuK3ifuXjXx1DQ1Zjne6JUALpVsgg3cO/UqugyWOT
Q6LgMv8lPti/qRZYi4bQG/C3acNHQo/7VX+ahWHVTx4xZ7mDyu1jHwFPia8nkTxogx3bFvd5Bb+K
FCCXSj8kIrBlNBbwXIefK8JvGLSli7BTBl2a3jYPZfH9E8gs8IwA2F+cHBUZDOfgZNqHxB6cGpzJ
TMaxoqHX5hql4gMuo7QnkjTFZNrdZRS4P0rnSLLFhgqCkgabrx/jcGI9cIWUEXt3dx99EH83LXs7
hGEr/5vxJqoKqp/PnzF+Jq66xHFAxXfg6X1agCpV4i/NNo7Af/yRXrIWGgqyp2IRWaNLpCceMDWJ
iY5ZTr5a/JIGyA0/NlODQaXXK24ykv/nm/YBcCgZyBqedoKqvWovV9GBDImlGQ5r7TbE+QR9+Hg7
qdCgDZ2CQqO4cGIS05oe4HZSWLQHlQrx7wzCvpu82BezRnD6pZxhQm5iTI0tctN+EyVMszeNpAs+
o/VAOTV8kZstWc4EYUDl7Lv5L3TP26LyVrxV+ObESy2ay6fWLbFwcqjdFI1VvWwldfCGZJOmGuo2
7NB2c6pXCzhEB4gjND3nhWftOq8jS3Xw3C69hjoE5vw2xFUwk9bTxpiPAZY9B3pts9WgT6AeNnuV
Z8G4htY6QHYA7X1lR0eUWCEAWccRbH5D7tSU1DJdqCxdlvwWT91Dhhc3bV2HOHLfRUI3G6VGuoXD
Wje9+IXswAy8gDIEPxTkSJeVe4fdqc0Y1nd3mYJnX0Fbc48Hbwbi+PzbUrbnw7ZfWNdN86ygXLjD
09uApXwuUo1RHWcc0Apei6eaaO6vR3lsi/juTFyEtASs/gjYlllt8r91wfmd/r95hpDdEk40lDA5
3WNDNEB72wz6HQX7d4KSFVmGd3U6KKJONkrF0cfmTYE/10hd5yFvf4iRRXNmp9rm0fRAg3ma4Hkv
YfSNrstiT3nFdImaboe24rgDkvGpeql2FckihNgQSU9afqIMhFTGxGB/D6q8jvFiwp4jpTmF3kUF
SUG7/uii3xfROpX2F7uFHOdhB2CGjNB4Fy5S+EHqdfJ6Olc2a21MqzbCgehRl46sw7XTW+d72KDi
IiZMM49R6/IlfDZ99u+28LtTRLOXDpAoi5iAOobGb0Eo7Sc1S0rBJ6Fhq5G7hs+qsRWYOqud5PeH
eXGte2sNMrTEn5EgPnwyUzctvtXs7yV20EAu57mJu/8LNdeCddFyk/EzfOUDWW1s1msmvpR0dZXv
U4Yi3E5yfARtguzAKDTSA+fqN0J7lknDMMSH24q832Yecph+Xrjb0Ww+FTJ88VoyBbWjJkj//N6Q
JhDw0Ze67H5KQmp7jmNtkvYCocpNgzp6eB8XuwdGR0IQN4QPKFd0CeB09vS9kqcLNke31lJ4PIlq
XiC9LA3hd6rroxzOg6vi5LjaobQSWh7D5kCqehG7Csp+ggCPMHAN72p+CeZTkcxnRWnde4kJa8eD
amptbVdqKcYoj6uzicbuqIxKq3ytfu+p2AdSYzv6lwNvhtyZ+F715wW2MSMnEJTwMd5S8+hndhbW
kzMraS5yxhAPUZWT8JF8nCLWs2fU7Uu/duwfQmnvA8NFXpB1411dh1+inB5+t7nHlvHqjT6BE3aF
i9bbiCoYWG7u+M2hQrte5WckRQYMzswAagu8shNJr/ico+29oPZDfa+yTHtbpkDNfNC4EQu1+fY2
Qx4uU3NMJSmjG83yx+q8L0iOwu7UvXTQe1gqi/Q8FNG+zcRVvbEqoosg9fQWOlKVHrHPfdnq2HEY
jf90kXIm6O3JLxHOZ8iZU898l0393A8uE2GufXG586XIAP8zT4WAij7t7E7FbKw43VfdIp85LWC6
EG6gXNoVXp6hKcePmai7102Jp1spx4xjVuD+wClySE5BZnpcsA1o28Sxu74DP4d3f12kztUZOjQy
AOkTDZZKuhAQUnv4cal8rh7Mib4FqWMkUqZIe4YHdZOFYnmFJtykNvhdQI37a/7MnZrb3eaKu4wM
fvVAEvx6fikVpudl6ELgoOwmKWs0VHW+1lBCBxiHHPPGedj/DrWJmYH9gV76Vws459ExfQ2ZPFRc
3QL4xMiZJazS7rQTzBNV9zvdbyqht34pAw+5RzLVNq0zVS3d1Yxe4yy0uw9KNEGrh4Tx0c5DIVxO
2P7bGaPkrUIh9kHvfB55W8j8Thgdr9AZdn0f31LjX4ynQcyrevOog5sQsjqv8CNxpLOu3Qxs3NLd
IRA99ZRrXlqyShtyZGCCNQeXt+mdP/Mg3/IeFez+W+O3ck0Sxs9uRVzr5sPKSnyfv4edd1WT7HXQ
hF4kwaglZH/0+6tZqbree1UUfPH8gee0rSOx1WU9dz0/xeTyaBNNd0bdWQNqxksH9ZfYxd8J+zXC
2PZrlioEaUvw7pXsLBXq11NjNcYJOC671L9egCx/bOP7d4lx5cnFVk+CXtaWyDIMoIrOzBetDBw7
z/HHJadWMwC4s+6rtqak1IgVaOGEuw3us3IbswGcfTzmKxVxFSBxHQ2OHLgxQ4NGcPDXSYPxtXXr
C5iRP+PT3huVf/PN4Sv7tRLQEUSpnDZ2zQCOyOEoYXqJ08tFBVeVWR+iyQpy7NmORnK9FogHxqd2
swXUeVkrPwyq1MPFnObw0D8ywJsGgZ7klLXzfTXTwd9xo3K6nx9U0A2Ps/H34s3Z5QiTAQqZ/EEV
aNmshFgKrx1cckpKkuKK8ORdz/x5OKfwMNmVAFqPMJ0QF7sXm5enP0kGKyQDZlGmTWXxe3tJO3ut
A6mrl+3fkagstknywu9pk+3305zJtU8yrIa3P/eAZMkCqood79Qr7C4k4HOz/qs9HVKrDIjEaS6H
qD4OnlmLCkuEsxSujvLFQgrdm0Q+yVrDQFYQhG3C0O6BUFFyhNgRPYQwWYHqLrMmbKJ4hLxsSdqv
KPD5WYEw4KvE+B09A+zIjNHnL+GjnZyEe4TNsPpS/NASrULvxYMQnDo2JTHgix6HcELK/lOW+Rgq
JKJU495Yne723pjz4JoWTNKyE3lF7nT3yLuG2qnw6O9SB2BT56VJ34cxFWJ1ZQJzHCXRAj7yaCDr
E7IQSIqRCRgG9jO05RnrER3DjUL/E9c1aTmAk5Z0ybS7DAeJhAgmj2jbKxoOr0P0ww53vQIFmGUk
nj7TCJ0TB0iANvHrQNRg4+lgD8gg6/ePcSl3jig4H+PunMykQqhaKr1PaJtDbXPf6KWNG9rwslKT
m9t/ZWYchWV3cbZSYdb7YYghFmWJm26bVNcoVfoayRjNT9xfDjoem3h6UGKrYH3xiSrXpzBz1Hk/
u0TMnSuNRevlfxdPG1kIXEuK5qQita4XxZjb+k866lUDFu2Ne9Jnjmd6W5s8Vyj0F6xU1hWBg0uU
BHnPnszSvsynrr83RQl5xmAk3+FXWq4ln+xdtLtczwsS6Hzg84Ign65ilYyJd3JRJomA7q2zNZep
fROQ2fpVOnacbWmfnX45EPMJLVZsqGmnSnha9QVRbdciFm4eLTLJW+668tFiY1DV9YM2/Q72HoLU
p7fSxK0hR1Kero3FA5MYzvZmbEycTlmoseQu52alnkfhPBKv/0d2f9abE+7vNzw3eSKO7xWNXmLD
oxYLwebgyzQOWM+Z4zN47vhqDDKLrrFIkvs5KQCPiIcyCybXeEpGykT+m9FzyzAKE5IAYJbORUye
QkM3arhCz3XgwSnrP/6ZHut//nBZi4Z1p07qRHNOHPf2XMdhE8LBvsoO96EIPP+T3NJqCY7AkOlP
QmmGYofKX/BNa0cqFHsceR8c4GxtnvrqtgAIzh0l6hFS2bTKTQgGvtAHrcPM1ff7HyzZGzcmhB7E
DjkbkpeZduIx5rgzv+W3hR06igNwtOUuvjX1r8pWPdvMJ7Jt/PqDgCjTnfsI8Z31Jpi5CMj5cw7k
kpeGLLv6kGieSew7l9+OKijGTcGi03CowkYvzM/jqi1+GeIhTLj5sndF+fuHOTbe/akI2PMy2Luo
kZz6wXNZK+itndZA7q7wmW81TgystMnOExHArvtqoaitiTa/PUDP37OpFLccmYsdIyJscyF9O9nQ
IDLjQ8bYlScGPuUyDNT4BaTD3aSzsUwu3Vt4eWle/noaIXwt3wYPpTB3GB3/meAMjmzVXZh5zOWG
eRXhHTsEQdG+cdmmFU+CiSPhPGegEz8TKoMO3rG/H7BqoAkiQoWeBTzqu+qL6bxt8p81A7FEHJha
I07E+8TJlCt2phzo+x/SE/vwwgr4MMxtn1lkiP3T2iZ2jolNRoxgCxEx6QxK5izURaw0cM7O5MiW
e87OIHnr8ckDfSMUXEkK1ohIP7mdntLKtGmU3Rta0dvNhaf1f3sHOubTwkcApfJp2n6rfN0m9h5C
mKtQhTh0nDgeOntLZkRxdvxUCxoXspyk0dBq9L47ba/gQaN4mpT7pwPGniQK8Jk8TJO0saQlsutX
/KFZs1Ue9blaBrn0T1SKsH5dzjwf0zziSUOE7inOPPtxaEYnOcq6QdUt/vOfAtALTKmlPND4Ziw2
v4lKnVk/hBCHOEdXBwp26hAS6u+rsih7W34zKsTpfdtX9a7c5EnzfM+8QVHSKxvz+Mo/aXRMJPLz
Ty9iUblNyz6fDrLMPUwr+9FZbkvcMgOBk2t0FEt/ZCV+CpYAfEFSGORhzJxlOLUjFofw+6KvfADK
wr92DahUU7Umx8DamiNWMM8ezXPonUR9xcjH8GqbK10LlIMV5bhzmgo1YPNkiuHykGVOeu52JnXs
OJhBOTiUnCCmcF4Rbyfcc/3l/Na/hhScR1gU9ayTy1gf+DxPEpLOi5lF/D+mQxF9oyb+3XYtIS8Y
bK4xiXJWfi3pMVuHMnDRWiLKMVU4VxlgR1zSqAKFIHUwnzW4zJT44qYlWSWIP8Aq+jpJkbL01AbO
pSA/kA3xGNfYb31N+6f7Ynr7KKhwF9xQLsv6ZZ8lfQtrFdU57Xhe/Q7y3uo34yGO+pa+Qe5Nd+rd
5mmUm7+j2Jl3oue/7DX09RrnoQTcsCvayhyV1JpvCM9rzyFAMZNdTkv3UjfbJh6YhnuY1TyTMLMs
tOlK4tAt1fld7A/2ONk2GKcNEPbazHHIFhJfI7Bw/k+j4xHGksAWAo3+g7zEOJD+NI/6D6SqZpmi
kNayDCfr8Dyhv7MoCmfPnvtm333+Cj6qcQ8NAuVG2IcMosQ7OHuFRewXS7xyRCdcRYmBruMaa0+Z
K6x8oVO1M85ZRoPkJfwUECGvomtg/aqf3sulfP86goEabS9IWelDw7LqrNc+9kvIG5hvkTGmiFto
GExhU+3BIF9FRmPcNrrpP7e5ZpEdf0pKM2UjqK39Sf2hifWNaTxZQYkU12bJ5F5cQo+ths4TDCMR
ab5AMNzZxHQaZe/vR09Xw7kAAUJyOcB8RGWn/fFgzZurQjYLbMKdC5bPzVf3kr69Qr8upa0B75tv
+7aaypDYQBlhZVw6Ji+POA0/7chVBFzCiX4QblRduZgaansfULwu99vTFnYgh3xQ16k9dXi8+nHw
UYe8zufHuYYtDuPxZ6xIWuyellu+k+Vzx0ljbP88tgYAn7u5meI58r7aXTNAGLKBAg+fMX9Kczqu
x8oOpxNRJbBJqpjJAr5/vBU9lWlGIspZ6vW/lmA56MTgDUjsQ7KnTzdC8dF6+LMI9ABwIsyiFQpo
LvbMoAt1gZUfnAlD2TW2r0FCCpVZv758RPurL9V/RaZfN4hYQnXR7VZ+fxjSJQU/S8zbNPIdyMET
vAA6+Qj7WXORhJ9sfegZG7tL0U09hYrIkM2mPYsJTpm8HHQ6yUFvY1azVhkzwQjpgGxuuSFtJje+
b1sBJgeY7GJES+rpDqk6fM0j4A/wW0MLZYr7eLffC35otctnbmyy4strW/uAoB3VqGA0BqPnWDQX
1rZxKIJKWPS20if+DRq3tzCLdsI8UXYAbASZg5dQC9gTmxFNHK8qcJaEMzxiavcLU0Yzq1NPIjK4
ymKoP2x6dCeoODfzVW1I6MvLgEVvu/6KY7ICVIyxoIifWaECYzCFHEeU3mXOWQX+njluMGh6GtZh
pM6POiFNKnmhaoU314fvrvV5BL31XvDMCeRX/uTuV6ZrxqWYCItUL7Tllhn26dc/aNBv5VriQSYs
c0KzzH08XLOrFJqkXh32m5AZZJ46RUaXBK6P/OmEXDk5a/CLyQyiFyF2Krl5lISDvnIdn6QCGTV6
VHSGAcTwu53lYP+EDpj/mg8VO4/BPKnRIiMrjkRHrac0f6yKHa1fUNtKUZTFyE5pK4oSQHrB0R9f
Z3qs24Z3oqdzBi9BhTQ0Sdv8iFzoorC3hq+JZ7HPTrjk7YpuAfzZO+r332n+yP3EUi5k8rhTOr5W
+YlnBzeF0rD6/H7JqqsRh6vJPU+5R8BMnEylYrvU2L+WxPAM5IytIqIKPI+bHcpoqVPht7XxVU9j
GHFJlP0EP60OjSR1FG6mVCHjdbgFxbidk1qi+OFBzhLAkGhpPuByWv58pjM6U9lfDptLCnfDO6/c
uabKfRCBW44rtJmCq1HJQcw05z20DLmEaIxYBYGWJxngvMLhOZ+6lwlsg1TVMxlYVjzJlBr9NGg9
90WygrozeCLvDN1ArlBGhS/xZbahsgoul877hLmlOKcjZhcXcsX6dHUyMBQs6YySFQtoBoTjRI98
OwFVLtcNJ+4NCw/Iy8XsfJiVljxWXo/64WwMY25fQsZEM0n8M5YEvQotsb5arRDdyiJfqF8vDGu7
eclfGBb3+s0j6Kcu9aBtgp79M7PrYDFsc7ttEOeZI/oZcg025uB0AUyZKWBh3iSyY0XEhzd6DQdQ
qnepNPQtSQE2krqK2uuDaukCELO4Se1/PT7P9Q/n1qEjDLvF7dcqyYj+f4vyFpi+zbyTFQ5oFGD6
6+7OT6qUUlrLDNKU8Rj7ul9MC0xrtN68+abDSkAYEvCzaf0euZ9Q3jotU21uKbPcIt0IoKePBrVA
3MXqbhR4LSSKBz1v6cZwIyuqVZPR0MantpitdtYakUOhobpl6+zoQaubUeQ/CpOLda1fiJVFQDNi
HCcs4ygM5FJ3BvjQsk1I02WRUNHY/BnDiwiLFhipOROcKUB84JoyvK9iR+MUE47Bp50Npx5fAgsw
knTQPc4uOmrrALUUZ1hAjLiPEh85St3rDnKPIDHCLbvoKxSyLIdpKu5PFEBv/Im6r/sKX4F7sy8k
rD5kYd8H/qf1I2fRIY6LfZmcVQeJMlEBcJWfhGzm0KabDYc+a0tFvVXjGGgQuyifmu85e6ucReYv
Pul8GtAIc5REPR64xsYB4ZY7J5kvGVVljG5JoIdzBI73eWtZOjpVMjwJ4GTskJ38nMlm4+9a08WZ
d9hOn3wq1pny4KTAjYR166S81NPyWd6PiTxEq0SX9/hJAXB++UNH7N5VKy3pWs2S++Zyy7Icnljr
/M9/oSdbgLeVA2A5mGwrMe8EO7vos2Mh9vDG4KHpY0UL+8HrWKiXHvmPJ2t9v8pyBpouKwJGK2nF
MkczDUDGquB7TgQP+9QDPBR+LHQbncHY00OnjzoWpQWxhWWaQwdBfVybcUNeHWAM+hDWfxi82LAT
umPLWoM67eDIAQoT4W2G96PlVScc/k5kfqhhDXCSmrbiEbUQjvRsRYfpa+CHvqdEr7j4E8O4tSjC
CxPir6KAmyd2vAqultmLPKgR2ozHpFydSvR7+jeyDtmXA5BT31y0gEbUstDceWoqQ/ygY7NPp0uf
uT7ZbJ/i0b9xRCdUMXxQxWIsVT9aTZOS4GWKdg4ZTdGffJIEq0LZuTUBlOoWV1RPy8Sgq+rYUYjR
FpLItWTqFpS5p8X/frXVDzTJwXYRVutF3hz0NFbGZQRIyKy5j6CzoR8vZhmhuw3ObJGR8DWnz+Ud
6Og4tF3OItOO2BB4DdoIvCf8zJY1Aj8D+zNCG40f7/yYy7N/QR/kFbUMOijwhdt9X8/NT51Yck7q
ejZRgM/wDcEE2ta6tLOeLI9k9URS9elSOKW/UjGxX+81S2T/w/JsbAObIIgLSUEJXHSsm+2TZhFf
SWCDEFAqOa/bKOGaJygOE31FWarEwXmtSjgPTPbSYYgku0XrMZOKXJNzt8r4//YT4GdTx6Jwi27G
NvoL5009s/MIMqS1AhHfETXyyQrlkZlI5ntNCqtLzNyjxfXw5CwYSRy61VrXCXFTQmzine4FqTpQ
oblXFB1/HosOY7VWWFflAprTBpYWvmGTZGWdV7S+Rj23WX8mdavxpFU3LaZpPHgAtawqTno072Lw
O6nJViA88Ba883mPNP5bMH8GvKRPhbIBYX6GWjwgYkuLkZ7X+8GXZTNdUSYzeCK327GaulU4/stw
OWHq6tZUjYJYuWSpz+BnEd6hS8X+a5dht4U/odENcyTPUvC2X7S0yz7wor9lxtKu6L6d2+upTX2+
oMEAM4GrWEeBJI20ay2gI4pNb9RsixHY+Utc/kT8T57MPjK2ZKePtZ/vIBLMBORq5UTTyrzNk+6Q
xA++dNhL/D4vEQyxzgkJwyCATdAFwqDuZPQUc1N13jeNKIZGVe8o/mXOHdUqXEb0dquhtinaCnMI
1NPVpScUv8+Q4mM0pvWKhR5uIQ5gwKRT8yiIhR4skuuo3IW2LX6ifw6Xor2qFfwfPwwxTJmg6h+g
+VArnHGU1LlacMsqFoHlszzsChQT7TuT1qZ4/B5p3ZOwGWS3AcZa4h4b72NrD8xvLR257TYbhzh1
AyWsZJQLGs7+EB1JinpoTf3f1sNMxWkn9cijO0iAMyAuR6Wd12moCqYXeG3orYgzpT6Wh4PxHMM2
zzuf1+lMbGiu2y6hiVx2cb5fTjYjYNzxSTTpUYRYJ/IGNEN+xDTnhrVXGfubWxsbwEd916/OQCEp
6mEVLV+blAtPP8CnIP/DqHSI+gLJ7rs5u+7TIcd3jXtVGqSt4fwikbdG29d/rgMC6FglqN6WTeF5
9W1CeVL51D0QuQaUYqn+e1/nYc5gL7XPWmUfpAGW/DoTTllPRpiov2sDyZkUXEjgmDgLNKx2EEvR
pv8NGLB7pocEXwduN264WGjvNYOAZynSO6JCPitevS6fKPZVFm3NfoWx0uo35h01OvwDRGJpkDLN
CFqFwiZRA1d1ZfI1zae4FTv0YLoywTJAuo0QyDuHVKfGwWDbyAUcqhdyQB3AwT9eJYXM4ymP+dyy
IVjmVo1hb3pwigwSbjCrxYFcdUB9xYCDlVvuTMeIpAVbVIzEhH/2ezVX8PYNiDvqheN5dZSLSyA9
gUIRdp4sIO5zvmIilmbK590Bci6RgahF4hTiJt9tkZxU056xSo9rcErc5ZScfktg8AMl0rALdKxj
oO3KbmL15eQFbCcl7VTRoxPVXtWTXe9QJsQUb3H3r7OLZSOIyhtfLYVxk/RFtNh1rvl4L2HRYTAY
sTrvAXOSyUe3mtr//+MK8j7cCuuvyAdLL9b01v0g4W1DLIJXgnOkaoRrJX0uW6sYlhAUqeRmmuic
APuhysqqSr+PMUKU5oPA05rrDNy0MlUGTDF+BRh8EIefAZTjKAV8BgS5BjCosMIgdLsfjQrZJshe
64c0rZEV+tbsYy19f4/OVLagurnvyzX4NrePgkvnfe4O7oVYVPFqorupbrMvQAsCMWxb5uYZH0ZM
u1mgE9eMrWyX+KtteHDx7jr/XV2vU1rc6tfreBoNr50NSqkATTw8XfTHFAiRaPZgtRf6sNlsR2vi
Ztqm9bv3ylOCRp9v0pDnrIkPvPNUAcenE+A8mM0Znl4vXQ433tJ7mkBB7kQRXlK3tiwH+wbQ4iUp
wow2nG+1ijCihlkswDKldZEoRg8ChSvyjdOETZvY7GT/V42VUoIdwb7bocoV87q1oYe3+LZBPsTy
2A4VLALgzpSnhAczvFo9gZj7wWqpRgwMPTqZGX7ySjjvQX5ocOmTLta2CFdZq00K6pMvGatQ4mwo
/fgDWLPhEyEouDEcB/fAVXx6tQDqvx+R2alofdE8Cfed13RJ46jLLyHDcsgBackb2LGjTL0DPIe7
U3EeNRCNyT+OxD9iKkv2/zPEbhIUSOQG2f9J018BP597eQMCBMC01xql5zspmj6rnOd1uDR820cv
iRQSlzfKHzRhDTuWCkn929OUJWXf+dugQHrMPlMZ3AYGgzfyZ1riDBL8qHRWe8D/4xd2sYfIdW/9
8tMmjYWRBPGyRY6fUv8XOplbgEqsoKLiMtljIELTXmI86ycJrjf7npjkrp73ciYnx3Ng3Lv8REo7
ZYCsfwQ3snEPdioFirV5PmsnkWa9Uujr1m+BGpehoDGmvkAhD7YmV1eTzD3BA5v4KU+AV4psdqgz
vgOPCK6/1qG7Vak05CQpVjPLn4m1h//6zUolE3JBBMYFMFxsGSScWpZWIQP5NjLup2goxRPpYDfg
MMgzeKyBkH4OqDj/81EVHC9uGbIQVhpvmKYXxYwwxzokUjo/POYyTmnbbaBOrrjzRyDfpHDrnZlF
0LGuDL0IvUFkxJ00RcCFm5Ri66SrfzFnF7MvyqGhNVAWNSeDT1Lso2gFufo1I2aL8585v72RYHRI
C1SEFfd+o0AMhe5XdUHSotOY/9xuYxtOZKQE4LUA54ik8IqqPgNDH9ACO7W2tCoFBS+p3jEyw40f
7UAQFh9/FashcvpR9H+hLA7u2Dval7aR4vUWOISitI9iVkBKUZTNgnMFg3kMLphhAoQ2HRtY3/70
6VPEzCkTMIsUZftD9PlKFUWNKfKsl5XHMhm2A0KAdtBMhkTmzXkXTmVjldu8A4L/E8iWtZjT3sOn
PgkK6m7Iec2PUdpSEYsD4HFFZGbwThFlwbEQSPxX8pAuE6jebPwGp5jc+eek0tzrH2jjssBX2eAm
DzcKXU7s5j7OMUp6bSpXjUTOp4rf9MswGBdKy45RupEuW/3oiaUGJBkQOiczADxnahBYl4sU7G20
cnT9FJ+2JVwalq9QMQ4rErm7xSl2ESbKBpldCe6CdXBsctl0oShIAvlxvmN+FHsFS4ULlnMjNdWB
mV9g/DlYoXq/d5/8OBPm2B+mEaXn9YqlEjxW1WhFWAG2eX8aFGntj8xJVM6a1zOdXSY6tGMunSNf
qvNVgjORRHnJXUGYm38vs0cNad39mRrGAAR7dKQRn7EKG5qGquAkU3VsYwurib06EikiQWr2lhMJ
mlx+g2yHnchC4Rzwilj3D9dFUpvk9jML1JwIY+3e1f8yzuGw29+2zryo0R7jS+YJU7nv4B/XUlDm
XA/lVeYkGW7XRfNXYLAfwrph7Hu75g79NrGNSizKGFauPdZn7JXC47U3YkoH3e7Im6McfPo9BEFy
AVu8suXoE8kt1M9M7WHeUBkrF5AIVl0hoj1raF+JJSjoHjPLlmfyAdandHGLkqd/OVX6xhOqCehR
iiPsx5IFY7par8w6uHc+mFkvM/41NNGKICUdRh87hda4S7cDGFPBIRrwJSO39pgucIdw7ZkN3rFO
8I8inzjfiWOARjNZl+60/kjavVZCx6I+52C8sZjY4xwwGCb+UwmvxaYzJCYc1gYCny7OsFrjSSS8
WgZG0vQ5+RSAIR3Zhw1g3Acvd4zrt3H6jjxZjFDrM6/SI7gF3VqLklJiIJRS+HPEJm+TQ5hSODiu
bbZX7Lf9/oEGI1BWO0qTlFsQksH6hkw3QnwIQRPRj8CCTnLpFHpAnwg9RglYCjV0QgpTaTg70k/F
TwpgxsH+8hIoAzTEw5mEi2mD7Tn4C9E90LbHeDWh6KAfin3AbZTjGXTfErsjxgvgOkkQ++lgln92
90P3B8lBBUvm3zDToqQ/7oEa2Wy/YDX+T5ExyL9wdZ/JBlzELx4eFhfQe+1Bp7NoAYG5SPtpil28
dCBj1C9Rnz/zPOQKjHGJwKjtciryFW6JtMgJPJW1y+FI7+H2Zkj+eQqAZLUFyN1ZxMdhBrd9ve01
4IaRGiQbDeJBMB0nb7i2WacrGQ6oU4JBcWHT9qXvvMy2AKMPdNSxNZtTbfimcZJho7yrJRQ5QJtL
VXra1IF4+643+au4TpRo1W0R0U5q04a1wptCI5mlT4SRix8AMHFkq7isX/PWh7QXA+NpHrzaI1aA
lYOm4H89flYoOkYLnR44e2CYIWYy+vY9RngGH56a9MJMwECFj+64fFAlMsnVAHZtBBIIef39ep8K
L0kP8BMtxETr0t3gEwH69WkgiLwvZa5xgcxqPGM400/G2+WHUOMGz4IE5P92gRlJgYVF3S6LKpw5
0moyU9pOAn0gOD+/HG9YUfIgBio7BqAp06TyJcUXx9uxIXYvhCUPYTB2+w8P7GbOwD4LyzGpo+he
W2ORdwqKOafxDE0NpMFjAs5TkSsV14zJq1CqVx8VUPJL2XR5RmMCTGnle4zCHsCYVyKs8Ps4eoW/
rSMFwh0IJvs/6iuDw5fTFr1WZQFTYSjXS2tZ/wm4i8HvDpdZDVHAtfODiR46vy/AYtXGxlKhe17w
/5zAPrBciA7WZ1GB89rk5cHGNFMV7CKanWJ6Elmt9zhJrmlbUSg5vE4uY+lt5yZwR1UPGypGh8zU
bjrxIjrzgyaNZyGJG+322TKQTCVo8VhuBekbfCKvWBLdG+C5Nfhlr/mx/nNjxAGx9Y6JJyUXzY3k
zSo8iUKNU1VFw1xzmGEFJpk5LLRP5yoiuVJHHqfh+hEccR1gH25KrP4lWDUEPZWhy4/5rZ5YMhZc
i8AqPjcuYkfJtkqmCgSqsoDztUUu+FgNvc7lRGM7otyvjWLB28fSUAWYeAsGABxlIU2eIKI3FR9o
gaEHLbG/Fn3u6ni+gtD54QomT7CAiWY+3IS2mzMW2eJ0Z3TV3/haSEyjWieb5AgtVpGJEXFMtMO9
fq3jCsb38/0a9wSikzZjUCxd1RQO0uijNBJFursfKydatU4B2mZxTSfD3LK5EHF+lNkX83RdSD+P
9kDUkv+NQ4u4LZnV/XgnvDPj/sEymVQNdRsbFOzbIRwli22NSblP1N6Ht5HQ68AW7a4Th0sDlGVG
Q1j6vVEhN51UfRSgu74E5CvethIvbDE1CFiwUC7KUeJmy/DQrgn78aJrtnQswGEuLRVEFLRfCO32
NrZh5mggrRyVAEhLUmydAFpes/aQPBfah9CLQ83STUGqSh4ZNW7POY8G/v/ODgPqtoc50Hx/9D8a
/nIJy4E0ozVW2K8JoBV2VMnZBJ20KLIRMnnI1jCMYmqYGOLDB/jJ0XoPIMQaLWtr3QpYJx+Cnq8V
e5axrB0PJ4cbBWbXMAw9q9wNcN92nxlthGueG88+gricqaJ+Pz89wCMmb6tFkXzEqq6dM7TiSPdk
Vh8lDr9amfKAEVNRk7P+qMrA5pn1LULF0mDALBhf38P2UmSv1svENpkXZAwMiOSlV3zyDkpYCAXJ
G0ntz+a4gLP6eLrN+qGqKvuQg7YZp1FgCJcBf5vsMXkfML6xWl0a8no7oD2Za/nv8cxjw6vwlKSa
CSf2adRIE6oSV6N2XCzmwtdo4D2LDrLcjwPw9Ce+bIB2vdxKNmLFek98j/HZH3WY+hP6s9r0tH1k
JfSNTXwXuR6NT992TI5hb2nrpshZ1Nia7FYK4hgKY3yulFTF7VP0itoBLRde/vDQZR+9QGEtI7yy
Gqh2HpiV5XBPd9rbQ60E8nzqkpfSLiAS9JVlpryf52UnPwWhFUsYWr2vZYfo0CmAvbTQYo2x7W/Q
/iMLtI67wYfastjItW8uFzPsskD9NeuNC4gcOwYP1qf8I8TpeNhCbunPkd24sIMzuZuAJfX8xTwg
M1qmgAjNQ12teW8O6iY8szWyqMsAUqDAxL87HphUNWdyBiUCTRbCZfNLTymakqD6kpuIOIqXfAcq
Adm6mXybx4w2jZIJIEsdtmPPxrkOCyeNRksmA2SrmOR7L+M078MhEJwH0NTMSuspFgCBlAWoR30x
Dc49zL0+d0UVoiulXzPfx3r2ImiMMxPcA1IzCJneiKlOzGjL/ZPNHj/BokXLE80g3Z/c24lzzkbG
M7sZBaaAawXZEPc4GHDc6bftv37ie9YgvbmDjS8GB19sTrYt6r+FD63zkZbI0+8RnOl3aw3Go9Ut
BjagEgx2nqDQnKdfgxpEKz75OUOSx2FBMjddJ3iAFqrRCVBX29Y3kE+vZICFMPCTv8hmiQxwuza3
gO5HbESrpGErYzTRQ5HrkUJYjSSN26LPsspLCTzeEb2IaQdjxnkEGL/aPF9n1PXFdbikkm9IdsTX
ZUfQM0/rhhVOevqgJ1bdghC2qhFQvxJV7tycnO1xm8KJIk5SIQj5wxrIdaCQ9F18Djuxr09bXOfG
u4htIfUc040GusBFAS6FWtYMQ2W6VIcBdB68MuzfPDmNplA07vR/vZCKJXOMplpwHNHmmsj3B2CO
u4mLIV4vpzXskQLfWS2cc+PmPkEd5avGUN8h0zw6W54fP6uliqN3DQsG7TeyBbr99o3QoFihgbXx
Ox90Jf3yyTL75BGPnDMr4EjkIUR04PUF6pXlXTfQQtltSPl6yhZVI9qF/9b8tItAb6U7xRilcqxk
ujhw+Aof0JTAdLNykSMs+NF4oNFcieehJnEi0lwm4dH+roocDA+e9C0uy36u9+vJ+eqY1EFMM7cp
/URTsyS+Hf8rB2AOyx6hXsLT+c01LCkLKg0Q7ky3o7Uc3FlAeFbRvuJoArRrplcr8voFE8SBHmOi
36/hbXckkCkI+bVrsM33Qpph1d8t7NOeYXWXlveQcYPLhfdLEab5+pBh9R0+S8SzULPIbdJZzEmv
xxrGkpsIZJkcrgi+MLp0I0CN1XXw67MPKxRB0WkrdtquqIhry9DlA17/QUORttm3Tx+1gKZUxdnC
x6Hv4aekx5Xd33cg0MiSivy+XVQqkJUNldX/qZ9p+1wcvd7IUijn0eabYfU/TozBrUNYTjQBQo9t
OY7cLBt5eqyA/mWlVBVH4Jz78hTGWJl1qETpk7p+1HF/QOKvoqWff6E8ugry/am/24HmVecod7Aa
Corb5Fsix1YQqa05YWr/enRZBIEJDHezDUSQ+sEa9uxtB0AgB5jSu+SGRDC3rHLFZk3TzUxJgIMm
YnnNhA4HDTN6HJmdV8T56SzNMCcTvGyLjQPMcFx7Vi9AEnCbIsYOZb2KMpWm+NH7cK90VNvkHWPn
Jn9tgu8jyjtwlAD3c1rpN+V79/ONVCHkR7cMIrxsHy1aerLqafXFrz0eE2aksuQS1EkYg5CTT0bL
6opDv4gyCfRf4lrAZwEZBnfRIxPKNG6CvlFPQ2dvdAA/IYo3kqxu2Lab9iSQYHFWOLIovb7h1c5V
5fccu5uzn0blLK7BD8a6pPsfb496gbc/teGegVo8TGcHr2riLkcdv+Al3Z2Wg9oiynxmRlgZ58TK
0w+xVNU2K2wvEnsExDwYZvg8H24oNHOk7sCleC6Wp1b4Ch1Q4F25AnguHjhIHEF/dM0M61FmjhTC
jEm1jnnoDYP9Uwst0mTMmHmrtcFzhbjpKQmLRH1sBYkNCBUxwvjhUFEBMV+5rpUY5Rj6nD68Ros0
fuu+KUjAuF21BuTlL7FA5JJkLLumNRgMl655ZGCwbcyPcKgQzD8dxO4m0QuR86AzST+DEUfO209k
fseV9YRVydv45WzORGM9dmESDudGar0lr0d42tfMdza/yDg4MInE5NZE65Wcxl3cZQzLdcX7IpXe
f8aeGWoZEUvFuhzVLhwQWm414qesG5woaunJO1D9lfzmXSWy351hK/5fkYNVMKc3+wdv17LTvLIp
YtIEAzhutstc2bXWPDDfj9LUiP1Sa3mIs+TdpUFAFbnJTlyklYlev9WLOpQHRPhCq7HWrXEamyP6
rmBDG4qz7/ZBsPMZFSB29tbv0U6GFfOgHE/UFyBiYlvIrQn8RKJfvQf1rhaZ5QHNggGJY/MgTPxq
Z7Ta4IffiGOeNlIhTG7QFM1i9N2ddMlXtix+W/Yzw4WADYj6KF3+mu/siWBEfzcS99+5zG582DCW
RMR1o4OBhdfGAWAEok5s/mhO6Xz7l4q1rYhn9LoEf/sSHfERzu64wWhP21BQ9SdpH4vVNl8JwLCb
LQCFcXsepPDnUzT6/cBc+HP1qLezdxRWpDszVDYm3/SF/g/LT1HtiwrvyAWWLg5c69cmghoXcb6K
A8EK2GqEBomwF/WL4sZZPGWNFJFhvbJXsR7HfyepAiiGqCgld8vdXcmz+FFtpoOuZXruXacUwTfC
x33gXNnjk3OPwDkphubFB9lFA8fEGR3rJyLDdrqkzWORuFU4QlVXf6isYF2dgWhyq9fJr3RbTjcr
9AQPBbS39hz0pQIzCGsKXfN9tnRLmmehruhaknobRqByhZ7A1slK/UncT/CJ2HrnVRlljDZfUSUG
uD4S1HOV5gna6/0BLvUa/gElg8x2SDDXK4/LcUb2qbU4sj+EWECL7BGrzGNvFN1rKFY/FK9Azuie
Je/tFmLKwMffnDBoFj05OJ9VckaTZX9I+WT20Tg57WXVoxGi+qXVnok2WhsH/dAOp4nhSTsV4oAu
DHHsBfDXw9NJJLa+e8vdV/1ydHIbsyXEf538VUKR1TskddD5t0vR1Umvl6msW2ARIdAvAcHErlbP
XjWMonEckGCimxmT/sRFIJwz6SO88Rs8bNK49Oa/SkXgw8zfT8ATqbbcN7PAcqurTWMOkErvilKL
lOylmBtyO/Lw/Aw8tQN8eUmgAxrFQxPG/pwoEh+8Q5e0wyj3gb7YrxhqPSr5+9sp1q7VHLArNZca
3TQ4buDixd7Xy7/BQkwldx0QV0Y+2nRA9RkIfoInWvhfDArt9Q6H8LkV4V4ffgYaG6vJ2JCna3ap
3hnJz67FKHlT0P1tD7YzfRdY1nTQj1GYHlPIVIcSKOHoz01C/CNYAqgNT1IAX3Uh6aIRGHg7vKV4
YrIvM03FHdCR5GCx57tsYF6DV9WNmPZ1AqXRaiEmdLhHYRiS+P5X6VoKLfDM7q2c8OD0wf/ViDnT
lV4aye25Inc0rkFo5MpR+ziPzPttYMekRIRt1juDusdLBNJ1KffxuJ+00VPGScVWoSMKk7tB124i
L/BpZ5enVPqpIPA7yYVCjp7xNnJifD8t3ugDZV0hDzpYdHAwgaJ5gTLEhK1+zxEjPpWp/3OWZMBh
fMhOer18Pd3U7lHJC6HgKFqdZuFvKmm8mK6Gd66AIyt2Oom1bvLTVa9CFePzd7uYaum3oS+72aa5
uoWXRBlEZK9BCdUF4C5j8xMX5lsocJoMwWtxUm+qd2y7dFlw1MgJdwEkYCbe4Tk7DRIJ5u5bjuXu
n+AFrxXZUUp066QfxnKXXz2k0SG+LDTKlohunb/OuBCcQI0dIh+PZuUuRwfJTBhIF1b3v71LK/kk
vgr5TDB6J5T++Em0kSdIvheYV/YjpBb+ZBU3Gjl8ShEn0P9yiOwWNvDhQgxyglxdb9iB33b3pbh/
cLqdFGqMiPn7mIsMEMit3JONsC9qDY+62jg3VvPTUyfFi3umHZ2l0gfdVJydts6pgm/j49DTotcJ
v+UZjZYYM/TM8osUdX2guPkzzZhBT354GNx3SVKTWPnSmwsfZkVOJt2BQ6i8grCEejLmf/1/BYVv
kxWfOju+iqXdmVahvGXeZsfejPnqurbbm/nSl28a9De2oXcNM7UfeRcm1PfvILcBs0dRDdOGcfdd
w9Nkn8DRA4sN2IN/2ESIDHYbz9nMSbhCCynbqzJwGtpvXI1KTWJ9hI/0iH2Mqxi4tam3kYZBKOgN
pgEUiBqziG/BuOHAwYmcjnibseG7t49sqqaaLtw/FwDMYXixkql9EKa4mwePM7LtC0dm6ooSeITn
thXMx7OZpnbEz2lJP5JbxJ3dex5E82/EX7t44h8dv/paY50Al5bhuKAqFxueIIhRJOZT50H7sWEu
11ZhZIHqKkwM9b+8F46HUvVbrAepXuIHfcREU3KxCThVtlbIxvvBpFVjv7K8VoyRiBzc4j6Hqwe/
QVF+rGCEGOrLDeBHcWzpjKNCb0LVLGN5oZTveqAqGl7lZ1DuymEJ/YkrxwbstwctwOQ70eYMkefI
2e9G+wEW4sdOQvuDUGJ+VnhM3uk2/TvKpUtI06T0IDeEA/ZtXpG35cCLkszPpl4KjwXK1NI2osSb
PYd21y+Vi0JAxKUIquseynBu1UnQsmj5wqx06gu1UDn9zWiyHC33Dqks2dTqghmVkPHNHWv53dDq
2KYmZgW7n20GludTyuTUpWg7ub57YvnmeSTN5mIaiWTGlhZzQWxg9plvwGMhS6W3oF4xN1pQv1ZW
XW1Hb7DsYDrbI4yBe31aE2QZRmBg5QCrl6aunIEScajgFS+4f/Q3pL6IgZqo6Pea+qMpydb3nqoT
fD0W0R96te/YJkkQMiK1nIOO7m1zp5TlNjDlmFoiHTILVE80SOBTYi+KNpyoaabBiF7fEnJNiE0C
PSF54q4BgyO9p7cW1GlkR3h/3eb7t7p/He3IGs4YQZGNTsm4Rilzsy02g7K5CIUUg3yzizP0hCz0
U/xJ/Ps6bCQ51hqoVY+UXwiWK95MtU8RB3VnlFO+vJHmAD1yB0roCgFZ2SkilO1MROTPf7ZilF1J
8Dj3L3ga47i4F6F53vxIhJINgl+d5oNTb1Z6ggrbSWUhhJYUPClb07oPcmqoY4ID7ay1nHx3OE5J
RnGeBeHeuNT9oQHuwl6p3+rp34Qx1x1Logn4CBWhLWsPIaHE9oin/wBGIa4ywrpr8V+aiFCIkx0Y
AlAXk9wDx9i6zbJjn9pP25QooMDnw8ipsfu1f9khUSw0PtkQO18mqZfNiLQuRKlZNBKmsutWzXyB
5T+FuRZq0bhZHYKTNDKUPRcQO2Hk4QY3vz9uANhInPIj0XkUMgj0i9mC7VBrfUoAtD7oYYB86SLF
hMJHyt942NRG3Iz0EYshks/YvjpyY1xeSAJ0zfaiqf96DC/wN7fmqLIJjOeYIjvuWeO9G+mEP+NQ
LjqzS7HR2uLUJ2Wpa3myTTiF3NgNuXMlPIHnF9MMiX+smVbtZLqwEU+b7OMp82DWS4AD2rMEgt95
PJsfsmsIREaPmlsv0Wfi0Kc3vtHXVP7vTtcwT1Lb+h7R2oKPf3B7EGfZ1mPLlLVHo0s3WD6dolN3
3a0MpUcHQHbKkqMgRsjHrShU6ib8cIz2VB379o5bsI73lft2SlkGZltiIuXIcheWNA2bjxKOp7Ee
CWsY1tk4mKd/xAL0mB0c15QhesAUHfoo7YsTELxEvC/BEeNG4AhXLlSPSlLtzNvgqtW0+JgT/L0u
altSYQ94aMhNz3I+6VpaJ38nj/eT0Uou9FeRwyamjX819OVqyxPqA6fLbTOcygHMQrhbRh6SqX9+
3lST/p7qoEpqjHkiDIOeSwuwX+l4w44QLT08P4BPk54UwOZXnHzdL7yM0wD3M8RKcpePFmA2vZOy
Y9tLngujjwu2gdbCvX7na4Lt1AztxkF06Oev1zDoc6f+/s+hgXohlImxoPokUBN9WBX0qlZcrjXy
A67pul3P6PuNOSpVz+jCTsvFdDRlVhZ+Jf5wAT1JBdwMesfYGKdoRCoMsmc201HP4DJsJ9wWfDkm
hWMrPGkPfa8k0O9kIx8pEx7/3lpwm1tZhNjK00KIoL8jBFLo/GKmlQ81N05JYjlyKYJi2Yu2/buZ
q7St7rDp/IUXz2Q2YSzPMcUaNAedTpbwJXcAOwvU2CRsEdYljO2p0vb04prdcQ78321iqPUgvUd1
KP6EMRNYMvw+/uiNz5xRyXW2PZ6TC7Qnxiw5wesuANtRKA1mPHdNXeq9MXty/FNYjT3ZlDyMQXzI
nFb1cfiYXSX4nqb4Z1azDj0wXuAfxkwj0H4cHrLL+2Sq5YyrwgpZUxLoOrM9sqk0riDdPg5nuEeF
AkoKlLZ+iHFfUKPT2+9/ViMJn9++6XJNITiF0i+sdm+EYY5547Tm6hoe9GNp3dUrfLWKdPzXPu4u
dZ15WhsQwI6nto4J1N+4u63LDFOOOqpmcbTjqK5lXhaarH0EYHEl1EGL/hawo1aSnJRXCc7L2RW7
4i4uiatpYLyPgseQArG7YEwM64rkiuj2/mWoFVyE8eRBPkpk98ue+8KBnjFOYd3aNyD8903Myygr
f1qaPjLI9XGFZn/bqaVVPPp6MlaEhu02mQgMBEE6NhLNE55g0bYV2jTvFpDc9ijzGy5L357Fu09o
Hv79K1R9B5k2gzyAOWO+Oat9xD9FJYii6UFY37yl6/pFmKe6WKBfGxZaepM3UbEIBVVa3Cxae6uz
lmgnq32JvcJU7ghdEp5vf1q/GmrgG5Wfab5+KIhUj9X7qrxbiyoRpAm4nkeU5Y6gETtR9gZduoEW
Axc3+vufdD0m1RPQod2xwpH8Szt6X9XPIDiu18yZq5fxwzbme+KqRRI6UR8x8AJ/l/+3j+zpB2uL
A3HuNziGOlQMCQnEjfFwbndt/oQwK36EY21vH3gYbiCbTAsAMdXdENh22vXmtBL3gArn3lLhs6/v
gFl49z91EMjRTbY6KXyYWjQVuxLttShpkKy18XjUJOOlOiOirHoTfz+C47W2RrQIo3NgNfFuMtzQ
+nzHw7mKZBlN5yDeJocY/vH363qfwHSySbroFLoJbLhWrVwThjcn23g+JSh8UmHu/iKmBsQ9MWN6
ix96fk3h3OO4BbvZcPEDj8GpiAKdjAlcdpvMq5UkE684C5zJDD54oZ/BcBDZrJNU68I5nUU+5Zzi
/lokVLATKdIHziqqH7GY2fHltegCaCBZjmR5EEtqV6LN0AC/rSttasM0j1SBPqesaWm0yUZ9HgCu
UlRySDE75Crop0gmALvZkip8m14T+m6dtCS8dN3lA/uo5u+v8E9bmNqTl+03iimJKZ/isiHoU5IE
4VZb1QGNZUVHnOTWzTiKKb0wwajhTFJEA6glBlqtv14qsui6tLN/BJU8wBiYB1q7VdLu9kwDPWZi
9hy0sV20lV4xVQX3g7qq5ePijzpwKVPeW4wL7JOFwB25/ePpGtklowvvBytQQGKQQElQYn4m6V9q
NbOm7UhbY0XdEipPYyIrONsZiE0Qqkd/P3OtlmuTab2DN+ChLZ7JbUxf53gXGLR3OdqLrks0wDrm
LCehtWSwWxhnqxLMesj9xUgI05CksoI//LIZPdrEt1kstNMPGH1XaZ7S1BWLKbW3l2oy/T687d1M
kIA/NgKWGSHgCnEo/SinHz03JNIoPya3nJL1qF14cxi/zz/vEYwjLkrcDoG2eAXGcQCK3EmtOuao
ulJZR9sRIYWaWYMW5fJn1c3+GdgtQZBEJ4xc8Q/hqPiL4BPF6Gzu4R5fd/XFYoUUzouy1Np7aKYu
/9UbjejuJBwMPkLV2bWpeFTs1RbpLF9eNO0sky6fjIl9SXGnU6lTaRqyAjPX6svhVJYYMLmTStti
0bgO0Oc9QG9yluJUP54HkC6rhPhSABQG9r8wPUtwhok+2LaxQfmvuwamPUgw4GJAqIznREN2Khdu
3+Bvyrb8xBpmqtWYsJb8RtM/x9MDxE/OWyaTdQLsJV8AjakqP6tKWqwSHRggFqq3kcpnB3Tepjk0
OccAX/VUyLuR6zHEWNC/0WgXKbIkkVbsnrAvGpsUfV7HAWYAg1PTFwI4Q6BeveRjipH+PwFFOI6T
wVgi8bUmjGjXxRSEp9yXdyQC5Bt4DdTk2Y1PURDGEVtDWsK2V8ISBCqCl7tLR8S6hzkQFvc6smv+
AU0CbPqdwSZLxf0NP2+n8LKNGfNyoUbWy40vGPALGfxJK5wBMqTUpnbY0fB42HShg3F6JMQZQI/B
sA5BjjCPuw8eOUGWUj0/rnMHjwzQkrvvasdlEAG985yk8gzam+3VW0E9aauCWMwK9pAY2VgB3Hvw
U68r12BmTkHcwVAJhnI2trNcTu/nFNIaSHeq0JpE4ZWrM+kx9p2FFBg7/ugbaFQ9cC7b+vPQotOk
jMKpJq5PUARUanOPI5xn1Eb4QkEQbOLlimm3Pv6N1UCJKe1xyJ3DodRjqEM4siLtrrFHq9w9W6cn
Xc8tOIBt/qxH1KAqZCrFleFxuu+FqZMs8tLUhtA4EBJ2KZOfjLzx3nUGW2pHnGFiajCG4DC0t+ZI
SRfmKUwVM/jyTRkqnl3xA4MOVQaOUnwkDo9ENa/rJXNkeFYHH12Pg1GVaPoyMg+YrQnZHdOq2aTI
LGJNYeGLiptS7uimuYLlAU+t7zjsfG32avQccDsc5hqFi/XhTPHR0dyfMhvdBNsKalX9LMRzZAlL
tQVkhBaKd09yzNn0kCU0OTzTQz0GyKhWdjTCTCeC5Km+hXblBo8v/SWicz1uOXAFtbftvTTC2lal
TIJng+K9vyEiajBkidZS86XX4fF/0SWg/vdwl7WEtm3dSNyu0AiTVIgu8WEsQab2qozOZNLSwVn3
EB25ndgwt7LY2uOZZjGYC8anVHhvPbAsCigimj4PF0cV1R6y95geQ2+wZjfhIpM/Wt40sAnr0xHZ
Oox1jovJkShOFHWQ4aMbGASGyVZcbBxkqKfRmE15veScyHli0dU7fKGo62nn1ps7i/OHlZtj63kK
l+BFxXDa1xZWeyS560yBVz21eG9GuiB8XWsmumuXmeeHBB1B/rdhWFpjnv+Ct5KDqsie2QC2hAs8
pXDJVXxlDjBPcuS3TXCJGpoJP2VbfSw6y+ewoffJbDwjJbRUnnnPhwCtG2kXnRJhfncmMUqh8gD8
QO5acplGdZjB7gGr9DS8scGWAM3MYR6Na+O++eHgRbGYRF/qv7kWkiCmaO62qmwN1FYuI3NDH4W5
2/F2C0lnDToHnDreUB6stcWIf9U1nia4NiMNNJdaEEclPXjSUATthc193ezN3LnEQ3l28j1H6Z24
j7ruPx2EYIP/3O9nj0hZTpY80Ngxo30jvxi3dPeIsHKi/wDTEbelK/rrTC6AbDvYU5xz3km5kFgj
3W48dZSqU2SABX47hyuJG3kQAQT+IrwrsDo5akcJDwde5dQVE1OxJGFLej+3UUSA9Ao6b/3yYm5T
OStfO8MHOJ6bm87hXZZnxPimFD92nhe0AY2YrHlothaimuWm9Oi1t7Au3BL/lw0o8foFJxubkeoD
bIARz1PnID4Osv7q5AOl8H26bDlJFkhRC4MWgQx68EsVAeIe4jE/9sLV2pyDpLcO7AUBmjtiocVt
90YOWJV0JwykFdR/GHTVj29Xe6kj5ihrxyG30uSX+IKM+3yU9qh/rvqLiUJrD0X4DMMvFTekZvqq
o3ieI+VtExId0ckJtDCe4s8ebJ37wXsP7EiQPYpBdsDJxzqMfp6TsvP0nt8aPsIZyZHg6DrgJR6R
fIKnQ9/fL6wLy2McUbHMwIMc6ng4fAbgGWLY48rVHHl5qQ8fNUa6CTOtwe9gZKP4OHSaaF9sAeAL
unhVyHKs4kGwp1bsOzuKJs6HCdwznPAHA58v/8dP6w18qeUlhQQdGvcKZXSVivIhg61QNPAi+qX7
cyj32WRK655EUNx9kYkotgEEtuTncqSxXuKHjlsLvNB7UGsYUvRL9eCxlkKttyWXmAjFGFooMyaR
XMHZh8X2U3HObOyY16etvQE2w9bsQRhZNPrOZMO/FkYwVP9Yc1BaFRgiy0XHT1hcXD2sVnR1kIwR
W8DTtiM9jlCCt+K8NhFBXfSND8THAPn+WAtb4ZGzKHIK1mHbfnf8wzmu5QqlDcLPTs7u4gtK+I6n
OAhfDKTiXE+MIPNXBHZhhugf6kxT+9B3VkGWo8nNrA9PiED00g4PQWfUGW7ps8fAfuhOQGX9rtqF
9sO8K0CD4twrh2+LjXqnOieyGb+bLG75Wes/nyd0dJKsTbl8ZKYHncjSWn0Pijtu5DZNl/qs1pbg
dIcyA6KpyUQdLihUF6Ju0xhjQO4ljbSjeOy3xXskXrFJrbglR0CAlpYjN2LpeNa2koYUdFKHfy9w
BR4lU3GjA+f0YplA90+yRJ8piV8HbL0g6oYlc309OHk/C9/eDu7+WlJccFIyyjf24hcuIuQyYqmW
QEjSi87QoV6fenDC4+GLD+4o+3Z6D/QcUBzSvFsXWytDFjhl7Gbch8X6bkwt9wBVbGxXaW9sUvgR
b3jjYYHEIy9a18zPu+yPyk7PXNPvstnWzMWxZb2hVjMYQh41o4HVKOlbCL4DXKLw2yX+C41OWHpW
avqBl9t7gutQYDX6adAf35pByOvT8TkUvdgq0r/4Maga99UaMpo0DQQfgYa3xdAfUC1Es7GNe5a3
C1ZODN7Sk2ITLDL0a53CHe3x5NJk3ZKApdmFk8vDL6M9WKp2w0/vQ/vsQwqJ4LnDq1fzJSFaPjWY
pKzmc5AC0wsyKfJnFs5/pW10FIW8YEb0Bb6p9B4pEp447syFqRIW3Pst65wnCDxssk3NMfgUTJ1V
GB1aWJ/gE43iYT59bgH1t5kZszc/36Y/8ijzEaW66XkY+MDI8Epqa0HuRO6lWo2Blc3NE2CNpjLP
MTFzjIKRJ0gDIZFSHWu6uiFiEC4m74yPzZXPJDQIXMeCCOIfbJQLityH22Se+BL0bKEYNrzKVGoV
YeHo6N4YhY2CkMAGf7PAJcJhNckJ7/pvkqAUL6ApFaq70YZ2fbKmgrtG3G/+EYlhuFmpHsY0VYxP
AGCNGRlW1ErJk0NMcWofq9jy1xEB4Pq5wUo8yf0GpJ+NWmAxfPR5j9bMdc+Ipqd3exVB0muq0pOV
ywKLmv4xnQOw4Zj+lSnzRvE3X6k8WNvMFiIZBq3w9Z/i1koLle9R1W0C3BxG57FljRiGEDSk7dC3
MJEWezMHIlCf30NQvc1wfi2kJr8F0XFyFNbLdM5FhU0TbspIDJkV5teUkiv/n/rIBXPH7XciVl+Z
VMPTkSTBLi8VENI6VbQpJrqh3YslxpS1YB6T8nxD+peV1pDxkDqSuVMrZNOGgzkqnF8fXWbQyaME
HwFu/rwUmRdnXU7gNzI5w1XNlR+QzqY5yUaTGcZmedrL06ljB7y3svbrcfZfTcoXB0ZLFZNaQQ6P
+qaiV94e6UA5Y3sa0A3TVBqMytWjGlaoBHHMA09j5mxOR5RsoWJLN4qxjsmJIsFXRsu89PjMucZ2
Ja0J1VBZEWCRdmxFKZWIBJX5dT0zisRDTcQWTjEPi5baMLgrH7tFVDfOGxyYmSiD3CowPiM4GIeN
iVp/RAQSH8KYbU+sV9OuTxOS9t+dSAavG9kk6DEz3pbLefJjPLand2ZUvf8PW86+hIhdRf+Bpe70
ssyB2j2WNn+aKpcM/NYEEigSNHNLLhDWZYiGIi6kfXK+bgJa7jx3jidKl5WiSR729f/3/4TJya4E
YFcGZ774kchn/38vNuL+7zJy++PXgjObTpmf5RWjJKF2IBeex49EBfkoXMbi9A/3YmX12Anbw734
Fb+gwyitLFXXeUkW6WfXkQfwKxAGZnf/Ci8+rwcObOkEVjthwKkDMjWDRSNyEwXQfbY4ASGiJW5b
OZFpwpG7LdPfv9A/kc/HVAAGRt88E7V3ZUPIdD59m5AuAv7h+OfUmbOcSj8pl+Wn0tcv2kLwASh/
ywl2uauJb5puT7ygKqzivFpQBmYh82jfyfy4PD9ZhnNBZIegRiFMG8qukJYFusSk7+vu5l1P/l8I
vosCVShU/ocHf1cfo9CZjpiRer6qmFMYP8/EZlIGEVL1+ECKH8c9QoxJd8sfonNI5/4CrkMtb+J5
5JLlr64gpHvZX6FZoEHLDjwjEVLLBKALmPKcp+RLGTpFkW/SrGy0Un4I/8fGgtxGBqnyFM9sV6Mb
GkHLvFlSkkgMiNAcAmLrm/iPjQmCvuvRzthlSHhkVu8wgOvCQhWufRii8reyaRnXv5Sx6V4fv/BB
fZ+Ode/OTmzC8J/EAun7LXh3kvvD8LaTZQ9y1U7avL1bd+3bh5xlige19qziRiB3fk1cQMQjx/AR
gxsZ+t6fHvU4ERoK/EOs6D8lYV0VFXD7h8qqKUsk8EUVO3pCF4DK0sIAG3qvsY4rNBtIsHpANEZN
tCvMdOZwiddIY//7p7y5aEmjGM/OJAQSJfYTBnSLh4OSLKoVFRhatoqqTDhoXJD4UItd5I7NRm22
KvXaTAy7bhHY6lB0nVn+SvP2ADlSbgxtYisBHayHlBb3W9b1N4HrGkvQhU6UT4yXikS8iRqLyVbt
0tMChNIc+9mZ+WHmx4bFrnN9YebW1rump0yqgOPnR3x+CibMh/Tlg+Js1IgSJcw30+dJRZhK9occ
lKyMk0lD9iyrDiFSn4qc3JQLq7RintotUhw/mICFHzF5wPKdMF1VoVrc4r23QDXdTetmr4RRVR9T
wss+ofI6XiCcEMyOPGPw6G/IMRI+s2voY49ioLbqbUhsP+Qe4+9B9JDLLoET3EEzwePkbfyLWQOF
9/mquSH4l46SrJCWOwn+ZeiD/O3B+6I18sZtOwDQPAp4v1crjdRmYa+2xcoTIbCxcRJ9W+f/VWjg
dWs2j3vla6TJbEwgKTVh4awIXNZK/gMNORepyBUK+pj7xl/H8vfpJ2xwGo8vGfPdQ5Yh2iCgWLm8
R5akfC1mvWAsJGnbw3Fon7HPKkjlxrnmn+i6gg2QimbUxuIbbQX/2s0UdgCOIKztcyuL+peY5hzf
WErBCx3tdgmtdFgnagPCLz/o8jqdddOMb5BxEmJplkZG2aJ2IKiuJMZkPg1mv+MkQpi5MBtGu4G1
/H8Kc8zwo+eKykoGgmhDSPhmjpgXYhkhKrCN4ipQPulHH5/SkRGRiv16egZ9nRSqE4PNmUFCSLHO
1UPW0WF7PtHu4lXvuA+Tut2bhZ+HdOZq2GsN2EnGyhMguggPomBkFTHXwQbBfay73deHKD6URF9W
ryfV4qbhKHbQvnI3aBfdyC4lQ3U+AHOR0GvZPgryffLIuc/vbgxxSkP9qFOR/K+ONUF1jFk2GyaP
Oo4A4r0io8Q37hStRdMy+6yKOL9I9VcutpP+c2VKE6G69mRAop6ETOpJY+D5C+uM+09fKGmdJ5ry
MSRQ1xa9suL02mgIr5MQmy+4PqcVJ9N8xxVwzzL/akiv2xqZ8OBXa7SptrOlNnIzQmhq+ytACBqa
qE2/py/G1Kb/aXsMV1Vr7EJWhtfGlMrQMqaSyVwvCBZSOkZVjkf5s/hg0H/D0lNYVPX7o6/kaumY
w3T58VawSe+dqN3BVpo/9FS4cqzEWEMscOeEqSVcePWo6KkxWDOwi8Zq3ekzSMF3h+q8JJ3bKNru
qQA4UvPZzdh+UC3jcgQWJHAAJHYYq4Yo5YuAmnDeXjDHyeBQNloqlLIDNsN0eT6EVVrp6d0IAG8a
nZN/s+EjGG2tcN3zneoueE9pawxdCzPDwQr0q9leM0yoAnQnpESPXxgHMZXb+CeMO177plY0lL1n
PblZC9IniWpagvOaWX663do7rJtJzAO6HJXiqc6vuMOMiWVrweT2JsavkMKURmIVTOzxt2MLMjT6
4nnQ9DREmDALqbpcQhN1gbEvbeWwy2Pg5wqpL6DWjwA4cZN7y4dvNGi9DGbkDL6Y+EQA1+fzImKO
V9fXQTCCrA559fBZmqLbw+eFxOPFbyGxuHXUpoBNoME9TttfjSORd+iP/ZUOuOLq9fkA1LrfXl83
N61jO90fPdy1b5bRevsHV+/iVZZf+KvzedKm/zCEkAl0hcOKkYxhcnhvcoUt136tLjJdEpfeNb3e
V6rlQJfWn0Rb9vcJA8LD/KPhloRYC7/zF7VRcEfSFcEwgXYRtnElbFXERHZNEtcexCXa4Tstebz2
vg+i/11tmNaZY2X/ibLOqf80SlOKme9LCRLIwkLtHXt+QbQuOuNl9OY/uGU+TPMFob5kkY0fXvVI
ipYuHEWrJrKkhjLbA0uEat780chLO6EBm5tXRWSxeNOIlPWvGowbDQNc85EkrRoNuALULK/dJvGb
msE3SmHWmj5pREefyrEd7hQvnJTmqyVDE4Oq3tNbFd+P7lsRD+kNJ33nEdruRGB/B2LNtRhdQYLk
42SmE1BJFZuDi9GCqJNWKs2aHJcoGa4VrkDHKTmsliMGkCL7z8Oery8T0y/RSy9trmxY/STAbwqh
9ChAernQv9SWJF+HHuPRL7dUX57vGBDk4S1wUr2/IBwsWQtzRqmkp3HgxrT4/7D3Dz4e6wcZzGOS
FbdsxypWh3wCQUXwYTaZSauxJ94D2YvX0eKUTXQATIXIyx2eKydMnlTB47HsgaVel5UZ+BU90//x
Tgqe7SR5/TupExBc8JGGINFT0I2pklKnGfiRMq7pjIFmTNc690eTHvoOlNUbbBIsaq9aFdIqQr6Z
0vZM1nhZwGz/weLMKJaZeynHOanYlc3CBl5wvOXfDBPsZ7OGnRhtDOEkSGXE5HpEogzfNYbKMju8
B+1lvU2CTPx3OtweeSOksA0msroDpj6xtg10MeiZXxNvCJ9+uMaldK7OXbJb/iDQ1RXCZuibtj0H
rw1VdrlGTOXkwa6YeJ+oncvejtbksC74Hft2K0hx5AbGjN3TtzEafWV5OzrmcRfdBYAh17Ns1bku
pk+/9xGdVmhkxQUyiHzgsRSZrrSODCnc6MCC5hSWRK9cJvOxdi7PTqME2Wo3mbarZJae3QxOUerg
MTN/QsOBBuyPbPVmK4Qt+aGTtyfFVgDZO1AD331U1TaykgVKq7bsBmJ5xNwsl9ViwCZ5YDkp9oML
xBZueTPRiIk42kLAblWuA9irwDpdj8sz6yZ1bVHI+69ouGh9I8sk/aTel2xA8LC/xC652nx3vTdL
tU8yMmrs/QBpFSXFiLyq+YeygnH0ncS5rMlsTQtk3eqd51BKuhw2znCHwLcpaM5FDXKnJry4WbEO
h9Vm8v6N59oVDbJfYqU9csUXGSqH2yIzG2bNxBN4lypg/aKA4grqmVWtjLdFqbDSo5G5TSeWWdRp
resFRsI+vXIv3rHKhwfB9a9moM5No+YV1KEOuc68AnfPyFmxkfPkboBY09c4TxysJhwWMgx0UGSQ
3pXM0rKUqIkRG+FmF0FB///YxLr9Eycbqa8Ev0HcopJIJk3D7ikrGiQMMdmxonlCEaU348EAh658
ptH/BVWmIPkuNp8NJtWGGrAxmGfwusHtnknCBNdpomDef2jNHtROKLeVom4SvVKkpEg53+tXKKgG
KFrlm19mGdRp4SLuLswaCj1gW0x+7m5Wd5dodwE/Zx+SJYkvWnBlEZ+2mKujvVgN9zHQBpJLKV6h
AIDO3t9BDGAXHh+g4/cZuwMbM7ytQG+1z6dasGPBfYy47zI7vh7mnc1L6kT3fPL9yLHZklN0n8S6
AxYN2HD/PP7zBHPIgKqB0mBlxelG5HoWbmYbatgucWFsfBB7GNRjgBVGXr7CjFXFTBIijXyFic8I
kBaA57S+80SOah0qKlHfu86hiDQmUyAmlJL67Ukn5yuleKxjaX4zPb8GgYIemsP+P6tbUGmdqucH
7ukgoRuDpxCc/1XazAGoUEn+PnLoggL7m28LeqD5ZuUXYQSqLwQcfMyhJB8EoynxFnz0lm9Rhx9e
BofcJvo9phHpfycDeXd3ztE8mzK/6bPvogdZ70iGxc5WCFPKl6wmOmEtppt4G9y2g8tSaTXLy7yr
vKChiEj/E8wdB3oppTT/YNpjcArf2f5pZGa+nPUfL6EmvLq8U6T/dc9sI1COn8TpY456GtcMn5uN
9fptnhHg8FdEhIONK52N3zUFrRl2PJ2U0Ozcqve53qzk9Bib663JxzTG448vU9u29BRafEFFt5ji
34zCBm+zxif9kej/ZqrJteezr8Su3BC3hhh1pHbachBnN9y2hrKcDxVx+6QLSAmNGuyX+TQdjSN7
3+C8oNVC2uwbvDSZlBqEjm8DAkM55sgYAjl2/gX5TNlkN0NhrSfmTHPah83AzAqIiEk85uUwCE0Z
t285Jo/mtSX9MTxekU6ioz65FHF+ju9iSrzxyJQ9RvuTDKsqPaRI5l9qKp75EYNG+aAjD+aWV7Ia
ssEhvNYGg9l/AmuXyIWUUXmrBiplI9A6/I+9vJxLqYXTc9zf72Cu/FnuD9g8FfW8act5axw3go1b
EiG+GExAuRUG/CfWqkC94fVZLl3vbTRVdSl7r2gCjPJdaUD8eaQypYurfVSgWI3CLonAdECfBrjP
pLgqYYeg1XDs7LFK0SA63VegoNwVi/OIBExxQbt3pXOajiRwqdguoCEp/1EcEFQnvEgYkaPDtPsi
ztHs1CMnTqpBcaj59fgacl6V5++zW0lTgMGGl2zJOEqdc7cEISlvyUn2YHA/IhpQtXkAw+iYtSrX
xIJOIFInm+YAX/ZrTNoSi5fjswhZxtVXKVVELCeyIzk1O4W5FKsLtEK/9WOxznS4b7FWgPKKY8DL
JFhHcQ4s9NFdgci9bcdSLNoSv+dQd7LKPtdMQ7i3OGTQfWuEnc0u3nkLu4lM58HvnzgB/jGYtlsc
xH3XbRhW1ECqHXZjfiYbBiDTEfnso9WnJ1HWTRHTaQ80zLRJkNylJaQof1Tt9P6+EfXFIBU6Tnsc
U1wym2hTxopvTJcBW2uxSWtnjISKsE4Ftq95UC0iDDGsp/d4/Ujdgj3Dcl4C5iT0lFs+9IVQfW1J
VOLbUiNzo06vy9Yt97lzBfRMRzmp9M5HGcbOgc1o4+NEP8uPgnDIfq7noHSR7kpKrr+mAJq1bEoF
ePmC/3bwr5R0+ckfnWEddUUthysT1bE/BP6zMEmpmpOqvAvCNhJcmL4bQEyE4BSNy5pELzqF6q8i
WsB4SRTWfFt+GYVdWEatPvAcTRSEIOWCX2qH80evzPJ/Eg5+NWn0VVtbREcTZzoCS4sflzu+OUFN
n3gfRjhQnccFPM2MJnOHKpvTYtD4cLw1zye6y3BhUTMcAwQ5Sb7lMHZL+7SReC7zlpnsspiLcnwI
NTPqEALcLsxIonGn0sPoTTsFDB9Wd0e6AQ+ZBjdI63bWBmgxcoynrvqk9q/Be31iuqEwBMs3tsNu
FIa6EOtCskdA6sI2Mk+0ChOqLgz8xx40bPV+d2dKF6isrOxMouikqLP5WBcjgZa+w7dMQ98PpThb
MBb4cwf31ZyaqeyWwpbUJ5phYrCldBj/nIhj/Zogn3bSe5ATxGD8Vq5FgGkLDIcFe8xB4aoHKBzm
/E3uNSbmThBpqxIRd36SwqyCFqidM/tqRWTVTdgF9Z61rZnRs9B2GOoMWcjhj1nWEilwYLJ/ye7J
PGylsp3uAYanONTIEX2YMkVvaq3hL1TFG/SMjm6iPLIqfdM1bAeSZNKs0BJKH20rvtKEh2iAsOt5
a/CpzHSBTPpH9VrmC6AYgGhmKBqdjSDWSh4hNhWF2fqdSltq7wjQr4Ln0BHoYxXLSNt3ZmhD+3qY
cyxZnHiOBUewVXvRK3Cx8EAzVqiw2vUN6SPMNLaKYIri/0etKN8pMmoJlBttgeCRZhaAr5VqwOIG
Ot0A0k2Xq4fVV43hEqnhcuN5KkxbtKVBaO8B3rInvs+7ofTaEYUAnT5ulRUfEw3+bWMr5VPwB9vx
5HwBJFK9NlkvfTrITDoEnDaAu9awiaU1rUXT8zfImvysXsmDFEOUAPierm0F0WVmVMmKMg/c9BtR
fcifn7HRuBqjq5IyBiTFNDWKD+XUgIvXqFN7Pgbpp/OvrRdnRHZM8Clsv540ox2oKXfFgR+bfM7y
bHybLgig9pidyzg3swguQLWqfDqAjJ1YgvOOI33ajwgX2x73ZD+Wxu3bVM+8t/Z9iEL4F7+VQq8P
ftIExBNQ7uR3gAmBpzG+nXz5VNg3SUosuyDiic29OjmLi5ff+RhE/xEgSGBuQgdSc/Bjgue81rIB
FaliXhI5RT6GhRbiwDYDVYxeS9nNI3bGvaIUabJiNT51Kmz4uSMqv2QQlEVNfzaHJBUlyyJdvjzU
Q9rDTUQgC37OgjB2pOyCWmaROIbn/a5Yqpt099yETWibanrAy4WzrVQqCJeQo0keMhvVSXFAVP8M
seYa5TPiDrPMITLYBXJCoYhzi2irBtr5i3EEvEEyF60bwaOopYW02vNSFobNhUnndcSgTo3NoK4c
ef4RL+DPA3rhm4fow1p3gGoK3Ir7V67YQOF3b4S1MFyX6Q0CdZGTZjWFAybRnolDWjwS1xKD3rrn
CWv6xz90vE5RnV3RKMJ5dbBrY7qP+hVuhMY4ggpngGVYzSAOcKMmePL0xcIcZIoX5joGQkpjp/Uo
24AyT1qzoIFPUHMl5zEWQWc102QZD+H3QI6DD1VU7qdoGdeROC215x85irssA/061lcuT392Fnrq
el3wK1NrOBITxGjgTSM3gx4TVTP9K87A8s/ExSeTgkVE2JUs/9U2jcy2SmLW2uGKl55mZVg9qJVh
JUAsB1Hhe3ITYLtoeqmw65JgAJABFGf77LcE7cHNXhjK4ly3B7G1MCgIccvaMJfqGt3lQk61CmVB
4sgkf7DoY4QrhvJ774KCH7mjdYC2CSMbrWJKSMAyb6Gjj/YmatIEc9tXcAVsRmUfRW/rcA6eOve4
oqN0Wt+cpmqJ7aAOt1TaC5HG8DsTT/Y/XOVDeKIB2cZM3rR8478Anl69Ds89wTnLXplNDwXM4W+R
3+uksPTR/+rj3KpvyRhwgFcfOs1WVsjvom3gEe97UxNADNWWR4WhadLJECQ+qRRPyBYqPmJeecro
ab1F3SL4UgVpocJK/hhPnVCmvuWzbQVKburbmpN8MepGOV73M0ktWNGMyUNHqdtmNm9OFiAbnrKb
b8MqHYJq34aCkFCsATnySIYHYIXkB8II+nr+DLqxwAEvrjG5EjQoNq8NzDkLPrDytEjeOWWB/Vhq
T5hd0ApwOdaZ+R72s5X0Nzhrq8LN4ZoTvR5DJDoAB6GYsicHRwEUqExsPf2iPCHbIC/84+4RFn/W
z4DHt5UKAOa7oYBhoLymszdIYWsNXObF/hRM5nJYqTmIk1XzhTVotOPvq95X2IhJD3Hnxd16zGpG
Ij4fL5xgRRrFF6x3v8o29DrqGO7tb9urLEL2nNNBJOdlrCpieu3rdVBWP8HsX065KsY1BTQAOqBA
IvqDyHqEdAJ212Xkw7oVZ608ungXL6DHFRzJxzNCSFDrmUSlTtvynf69MgCkZ/zs1XWhmgCeO4qw
zxYz4IwWlz3lpSChIwjsrhtWD/jsQhnKjyvjZ+IqATl1wqyEBilToBFhpKPLqwOCmz1OyQFUjBIl
orGM3BL+D3eUxFtEFzfd1I+GgX8/mz4/3MiDpy387qQVRFTJMOL6+mmDyOvUr+a1fWMvLdlkfL2x
IIVkpo5DSH0iRIqPThEbsbu+C+VlxzFvkE0xK5bbjTpPo8dSts+DqgBiG1FuABA7F2cbdITin0tC
0T/X3E2igTYxkTWynEDCgNTIHe0mr9azBoZqQ211cFyghO+A5NwXAm9EJOofAbcBRmGoSkR8GCmq
KVVyQ4DgVO9vfSb6jbCQQ37H3APlGZK/TsvjB9+zEM5u9fxmysQ15BOvUmqIca9wAWE24deSYacD
zNFHRRPE4eLuGDKT9EPq4iSMf9g6SBQEfooRWvNp27YloWOWhz6Q4P6Kc510wZvzPla2USwkMMIr
YK3fsNGlhPB+VCVZyTvPfDPyZ9ZC/b1/EJBpnDMJnJ53rZ+V5VpRfbzlgL7NLeJSuii7lfpWp6i+
lmQVj2/SkgxjNyeSROaC4X1mMD4thPqseKJeacQt1XqYLo161kPt4Oz1SEsxG2/y/c1lnfBWJkoD
Q/mD/eAW9GKOWIf3Al87SPGQJHlvJWkBXjAXZ3WlPWbWPVVtfBBIzcxCTC40+f9lVULznBUujgi5
ronf81zwuSgEaZT7EzOMXv24OqMOJ1ndq+XDE1tHvgN6uEOjxK61v6Y81IwUD9W62BSZqdDCVVNi
PMWKmFMVeDH3PwuV2HwAUwS4UYQDNKR9WZIi/Qh9edyILMXe19JfYBIcM5BXgYpa8wTnMnGY30YQ
z9wCbgy8I5p0neQbnf0KBxpwGH4wbFzu+pOXj5aeGZSlV4GSSDhGWE8PnWiRuj6919Z3HptKy1lL
AvMOTW86/egVnUqBRET4h5ELxRMW+L/dj3CbkcwQ54jDux6GJb2yoRNhwaxwtfIBzBIbLGfRaxGO
nIQesB9Tl6hClis5FWYPjWhzH/V3ihqE2Kncwc1WTUmSlhFdievMvoLCfTgacV4ydgG5Nav2rXpl
NzXqCGfKS0ejgkhgsP/TKyLodwCFFTC9yuPy0VzsX8vYz8beYrYJM3iRnvnc3NmAxlB9Ei1ClU07
giXYupmtmE3qB77dS+C/ohjOCYuLNeb8G7LkF5oSrY+hqxYOp36Xr0kfjHRyAV8+/bUqU9J6Px2G
IT2nOYXs3eYVwiFpEHpgQ4agvbqtUMVgwmoyWTqXypOOrie2U0JKbUfn0lQXtVwB6d/0kAhIF5Po
BsqA/YGbExosYDbA4SqXhY2zIAtcR6Rnu1+0583BcncQfhC+5fIWV/AczuXNYBkvJpEK3SUDKRD6
b5bSkZrO3YeaITKrFc9/Tt7biNrU/YoSGlJFB1LpPdIfhXmPO/Qb6Os+qmyKT6B8MAJUse5ZVkS/
EmgflF+6EGX8zeRyW3tZ5Q4pgdas/MoBEqCoT8238HjCLUPUJ+21W2N3sTYVFAaEIa+dOdfVpWQn
l+jIcIN6mM7jOqRKM+8olcNi8kjo4HCaLonQHvPIdDskKFLbj+3/o/TxxgMJKKzjb3zcQnH714KB
tMCaUIu9sJr4TUQgCh6SjWK2nogmnCzQExJLjPy2cnuoAJt7kxbx2Da3blLT8eTeieHM355TiFBs
bPOKFh/xKUc18eOilVPiXw+Dj3q9UFCiRJx35qiIgRDwqeT97GuOaTJoUdsZi3PNHee+jsePZ10N
ZFwCwwXvDPpIPt/R4hoLGL4JLqT5FI2+egYIAEh1DhNZkYlQw/eilJP6vSFwVbElyhqf1kDWMsGY
0XwQAPeOEJ+SE404coW39A5XvJvlAEAN9f1kP9J5x9A383J76klFxj/XtLDnGKo4kUl0GxMqa+iS
EuMV7J3MQ6E3JR7A0/ESw9AM7rvDNL/Bu9kzbGIXRVI9yx5HnJtXUjC/ZGAa4s9l1XPKzi+BTz9L
gRp/jy7UxyJU8URbdZ1FMrU2YyvKl92mw3Pq79tI1f3WdjkphjnqWL8BNVgGsoBZV8wLPeg8Dsb+
xtVZj92ldnKLo6wA72wUvb8PjgmvQ4o5P1ugLreiiyqtNbl9xLTdFregincCwu/IOANiZSqoLfhq
vEfhnym7Zalf8duWTWOBo5bQwiYtrsEW2FR1biCrkfqxnx/sA1MXjb1mXKf2dDg+Xzl/kgQ5/OU+
jIwaNTo06SIesBBdLfbksucFdF47SeWMB8opS2uWjOYme3p41dS8K3pcgRXS/FNWjGyr7wpHhpex
9LT2q5/pnyzugoqz77Cyzc11VA+O/kokAhJHerI0BKuyBmDfc0WOUsgSmUUqdJhYqA7Wp7jQ3mvx
F84AC/TMzpz5NyNShrhxsyvMJSbVv2YLnpd8dDwrpQ19h6B4YGFgUEvvPp+HCEVIzfuLye9rxWcs
ci5hg5aslOKbyOtp+AGuWURqv9LBQaCO3CNuzx71HQAK+W5J0SkKjy7iEan85epoocGW8tS5K1Sx
zhOlNekkgf9QDHw2WCGAj3tI4zX288acSzsizJLHSaTmGqGjZ4fdD7g548mUJunoqNiCmnh0nsvZ
Mwk5/O6v7wVHZXEFaWJOhEhMfJVLBwm1OkokAiNxKQjI+23OU9xJGgo9TNHqgFeC2w3j+blDplFT
bLM+ciEdnqXwn1WQ5zqOr5k2JEYhKq8FRM3m8gwBnYKpoqVIHCVhU/ahrLNSK4JnpnzbghTrP3Fm
V1DN7fLQZO2VI07eja/AhuftjRrLI2FBmI7mGsOjQcC5RsDBZcxAd3g4tKmFHXWuTT9gwtjrrg61
EN0B5eaiJEZnJMUiiAOERBqiFZCyUqOG1bgMItR8ARVsdUiLwGGjP3Yq1mHfppqlaTBS6M6Br/7y
U6CS6b6IR28oepG5Ix8Nr2kt1GQlFQA4ySTzaCAzmg3R56BhX62Lz1CIZp+dxMQUl0ezlXscYG82
XiVsBWSVW1wptIqyJxDhVi6Z17UQny/GHfbFHP3lrm3p4FAHYXP4SQJr3H8ME5jQJpDnfAS7+rgM
voOgCSAmSsccAjCsFswW9RR5Kq8iJi8IC3FyZd5wYac+NZu9joGmD9yimTZ2jtsAHZyMeSHIAX6F
trujAcCr4+hdZLdb6CwW6Cbm1FAF8oTv7qpp1LRfO1bHvt85o9DmattIOMkNuf5QcH/4sfEelca4
5otY9FWokiOa+WT2Ls0Vdxme6DkYBBjsrGlj5Gv089uKhsv8iJgDC/gD3tp/Evf9vQFRi7GZeLc7
nnk2V57NtxIlWpV1+SgUPSJ/XwWjEfbtP6CCQ13CwR5rvm4cW2skqTSkpbrroBzHO3yaytN8Jvk9
XqKqKgtDUfVPVeqP8ipmQ4CjfDP9otDyWe0rdlYL26xWg3VbSfxmjTyz5deccykeqXwv1DjNwYCh
m2hJmRJnZKhdIXxoA3pqPznMz12udQpZaMIbCPOfBFcmum32/Pjfkll6b05+Wk9Pg8RpDrPqiuro
voAO7Lxy2XSQuGjt02oFBVJecboFvd38fkQ/TSniXRPPmB3LDriE2TL5+TVwwY7O8zPSTFzIsoMI
pOzbRbgaDlZjQk/UzQW+LbfMNPqD+DT5PRTKCL1yOvmdxO+Z6wQwYlZ4zinUrh+TZ+HsiuEIfxgw
GWeY0V8B5KR/E5jRH4XrdbVSv2VlZx/h18SBwLtACcpA04qwg/ukIBNIHpkXfVB3IJ1fSS/pgy14
XYK/ozvoVTRo9Zu7bQKErh0nv50owiqXgZjXkr4nA2Gf9jvm/CwRkZIzmOhkaglSyxQE+s4FOeAP
5EA5aPxDhCOWjBkIeYaDjH8jkHbCfRIF0F3qTjC7Hsc0Ed6P76cQTEX8vf7V+jclUbOS8tinBaob
PA7pPFs0nihJfzw1NCXx2Bk+tfR67Hc9DQLCMnosMmB4GPij0ARD4wLbisJzRUZ1GYQxHhThkvmR
xkUmL2fRqZqK+KLJ402z04CtaRtqbXHtpD+EzAiSI6CiROb0umvUeIhqg6deH1ae5T066L4+DLP6
/gdzj6Oe77m/E2jW9NrJoKVWVbqWPm+/sv8p09eFhuKfNm7g5pwL86PVtHC3/zRcEcxmOKFbwHLb
yb80JG918soAkmi9AU3BrEzJSmgH+sTZlsau+NE0v2bL0+gS2TZBcvIo/lyCDoYE+VoECSuC5nrh
YCAPzvjEv9E+NH3Le0hXtbNGPkU9bA9LfFeWBx9YuXdaKgYumu4yYEM2KoDXjup9/4nItW52QAYg
Yo24qa4yKQ3UaUN4HmksaVb90p104aZW4LVptLhXk5vwUqSqzD+cc+ZVhxNd4ASvNTCrzdyMBgAV
b5ZSBg8AlQw6Z+uW65Ej0Blrqc145WYNlnhD0bHVtwOe9J5IqBEWAqj64vQinaER6isLXAJr/C/U
A0wqj00e4XYI8JYTdoqEaciI55ivxc4Geri835qwAyOOQekRsmghm+8S6DOq3WkzyntjXJV4QYyE
2QWKZfAPqoylxLxtImp8kNIyWacVF8RoAsuTZFTeoxMO7kptd520vb7rF3u97EyouehzN+I1/2wh
Qnrhi/f0bM4eF/6mO/RqjDnuvW4jH2u3L3bxH7zbUYH3Q5WsXbNGIZ4JQHmpiEOMOTsuD111EXe4
QLf0B4jAkpGulbYsUPjndevEboNdR15AThezQFR8GWQCn/GWydeiJddonLINnfpLvUNGJkZtsjYB
wInTAm62RmBighw47tMe2v7FaleIO3yKx8xeJ48RxSoyRAPYe0VEo1tAfIoe6s6ZAW1Ft76f9+h7
BrhTcrTN9HAMJ8UyNNRE8KmXjRV9ierDdSr9TezBLpViKMuI3zkgU8H5UuOHa5aEZ5xFMyM1/Wa3
bHcUo1Mr2wb5Ph43JBMasA4qa152al3uxFZp5LD+RviPssKwjTfwvd3YbGAtuJXmb5PHmegvM9pA
B2Rgl8bupFEOF9jjExvS09oWS87jks9eHi9ty8LsnmTCeLykT6W0ZhOhlGHHl1b60bkvQ1PrL6fg
kNSbtsYGJXQi5y1iujuH2jWWms413GyQ2V+4lvG6sdtXuhh1DZURtls5CLxPsJPDBd/jXJ0Cdrpp
jrdA0r1tDUx3ktOrW4c8rA4metTQ4+PS8u+y2MfWWswPAMgoJnCyxnCN2y92iG6qBFORoFqO1KJj
8p6uJcBB8d4AzY/yJif/QtYwO3Nj7h/2QkmPloeyKfNQjdsS6As2qpbQixN5csR8bFqr0MP2bUkL
FJ1BkpLz97/0P0E8wgwtRNrm3erJEsIcoU/RolA6mRX1T/9DXQW1hT+P/V+NaIiQWDerqk2LfWJ/
/4vnhYiJdFfqhks1YC+GrPD+X7pep6k6wZyIFsIGihpl/V41C/USoJkmm95WehFd2RDiJVWVSAEu
Ihr8FTlNkKBRaNm2YWWl9KjgnODJJQWvdnXDG45UjEC0MalTQHEsAeKM0HDcCO1GZDDMyaMU7jLY
Fbf3Z4+/Wme8n9XoxmGvn2bNy+XRWxukhJC6iRk2peMf+Lq4RYlHihydS82JTmdSSs6yTC56FEOn
vTQLah0SQjERmLmyDBwxSQK5ihQKc7wr1YC7P19CQRyCIDLsImacqR3Qv9ONer11fPiNEegYac8e
HYZT+oK9WU5FxCe/3193rvpH8XMifRr3Toaa4td3l/JeYjcESMNeQ8OU/cqHwlu9whJNADr05eLB
PPkzkchxNKaGMRKqg2Ww29qr+FDB6WBqd9GQQ/8MOtkLLNdyAK37KCTI7riKlIC9FXa71cnexqER
tzTKM6wJ7S1EvS5MW7X7RTu1CmMxOeJE2oaRQ2yVgXlaO+Qi0Sk5SbJuzMPPxhMoNvjiJnrquIfP
59Epas/uKRo+lVOn8BjVYlFXT6FOA9f3SH2TvIcLxMQ7m0arn11QZIP5SC7UYp9sJFjklnDP+0jZ
o1AIHoYeT3mOTeMJ0wfgEquTJx7fuBZ6UlW2VMap4xbbdjGJUihoIfSEYkEu8vxgSmz23fuXLUhl
+eDqZZj52VDaonlgFtKyIMdSf/41vBOuuLafCFz67JkoNEPHPfd+csjeGkzDoN2wvHOeSf6i7HoM
NDl084JB/KzpbsM+wvdzfAKqWhkDoXGMOrO/L6LCaymdiYU0gKk/QWKcIM0pXoEObrjfKxspp188
8oUJE05zjXHnKicXcdKAEp2IIjIhJzY0w+T8rOx2iuMEsf9S1tOfVdaCRZeazxzebWcS/kL7QV9B
gHCAAfpXs8tP2AyaYASHsBC4UexeoKp58ly4v73/IURoD1e3pFnZ+q4lNR1ZloVnJIcP+CMncazx
h3YZPRIWs8UfDVUgZk0c5ylNq3q0r0gdqpelO/4X0cA/Lir7F+qVKgo5UZgEv6PKMP7ges2zO6cI
8yKWvSwMenl29e5YMOEOuKy7Av2Gm56SoumQL22hp6t35w0DJzaYi5CxC9B06lcVAE/rcoT5RxF2
N7q9TJciFkxqmJRVnHcTOQllusrIzwsbeomyJ5jiZHJ+yhu6X6/ZA68MB4YHq3Cz/lY2TBemNdsF
SARr7ycJKyj8785FMdVNv18N/HGYDFq6hSB9xolL9Lid+hdL2R/j7dHe2JBpGdHA9j8BwwlwVX9e
9w9B+Z2zNPNBefXmQevxboe9PCietGvX1h5HFIj1NFzDFNhABCviAy1+r7JFVR6nV7/DVj3dwXhj
CFHfOZMH8K38vpcTr35FXTG5TlC6Rw/QeEkLSmx+ssdsjGS1LaWF8jkOwgNBNfjtt/Z3Kle2u79K
3Mw6z6iEV64wxgvDQaStf2r4xqZlUAUvumef36FwhU6WaOLKAyJ6Il2fHgY1NilRQ7b0cp0LisG0
gz6zNGxOuufGTZbzPlvtiBGAXpM7mNLT2L4SRM/AH9DRaJu+JldP5tnjW//2XUWqJB3bri87LOcW
ZPyVqb/5BqublPUhLfkhkabdNehG6/ykiFH+4Cbmf6KBHWziepmMZcjqBXS4SC9JnBfo9I7eHdyA
8LbCgqpeE1aR0g/0aWQ0VSuOZpahY4QRJ+TeKDAtekwZa2lQWs1A/d3emSvPdTewMukmDxZTxJYn
AiE0teE5woJk1e8Fa3Uz+4SVHqzh40MxCYdtJeAfIGkhEB/pwUZMdgFRNRFgL/5qQOcy/Oqo5bIE
lkLtj+cUNrEnCKtp4jTgFQcoYQfF2PTu3SI8b99uQSdj9F2hX6KGa5HxDfGFBLnlhxWUNDjU0o1N
nNVuwUc8Ini+SseO+8+TUjdLIR/vn31L3DqcdWn4kgH5zlUaO8KITvfU4wFasLwhQ1uieAf7YxYR
6NcIIOb1OPu+4Wo90twf2MZSEQoqk9qJ5TAv9gSJwQSuK24Qu+pdbw9ETVwGixsxpg/Y6umGphLi
YmsC/6+BAI1Y3s5X90Hk42cztH65gSHQ0ZS/ymzNKsGUrsGtbmf4RcKp2cTCKWLMiaXFXu7nRvWN
U7BsGMyG0TErjBADXOGf+GlnQVd0hYuhMaFQsoO0UE0D2z4F5RdqnQXg1QxAP5J6eYfZ2LGjajVc
s7YJ5xez4GnJQpDjJrJlgUmnVjgCQXXZTqFxyeseVUukA6CP3IPuGUlOLZ6Hcm/Nh6QbRKBdnVcP
XUwN3yi+yh/ntV1mY3Nitrk+LhnKu3p+ZH77Lj1cMguXqd2IRgyEgju7qS18qlTPTJoP8LENQXUP
ZesnNNRRWELHIzrMVXNYrvxqFM1avSrxjY1Ir/hRj5YiGe12v+UTAJBfAhV/buOG9V9UHDxVsG/V
fpDjgk+bW49RK4SYIlrZGo1FWWvwWLm6pdelh9pcAkh0a7tXuHkJSzzRm35E4jT7u+DVQMJPDWFn
MkgMcJ+bXkydRgtBXx2HuZGiO3EvS56/Zfirk/frkz0OWkuUD6Ix7hPovciW/JCpvevCCcHwDBdV
Uk/ZLm87jc4RpjeF/MgHXCKrVrPi0YLC6oiM81K3YfzvUKA5GcjyhhQe/ZyH0S6nLWTG8p6MgMrd
TxzSdjV2AiuZMO4APJ7VQFAVsrXp7YzILggKiqlbsD2LEEpRC3LUUlFbbGHaYnCKQDTLzkjCgHQj
NUtlB3muI+PYKwCa5seSAV+r0NgEO8x2oL/QqBwIm/TgWv3FMyE0qsEmQUfxzpaPh+CK4o7KtIN5
KKzzUBpAEK1qYJD5NvBRYOC3meGLa35667q5XYtmvHglvwwwb3mPJ9DlC7HA+6jRB5QQ7w4wXVO9
LzGlyIT+B1Xx02S0ntURsDo+WOwDnLeRMciIiV/WF/Ik3BvQMAo/A2pTjuSi4rZqiqK20L6ZkHx1
zBa4yvhsKhMDB4qhkjO90fURRxRZr/wTp7DImM/vOzxULRMkAhY6YCH+1PFJHtplbR8V3A2Net24
2dni4n+smNOyxIa61oyBWgP2kJhRigJIGmqlA/hPtFWm3Sf6ezd/EG+umogkNk0xysZg6j1josth
hdVqnvo3LOnmKiG2wVJ6TEVg71sB1UX2I7c7r/Z1Z4FWyXcUKoIL/osln7INtSDiOjqoxaB2gIAL
LFNqiCrOVZ6kbYUdptEwiMXLkn7+prH6UpGucaAD6xd+yB/qFQSzlReQjfAjBT6beiCaUyriccqx
fYJsGT2+6L8GU1IWT1O4Bh56AUUMCwAMkT+7ZL78XX/mzoAFYMoz/iB3UYJx7nbaSBj1VLmPEU6g
I3VQzdj+qntAyGwjFZCRpsBBCZ3gVbnVfrN9yCheSs8YVa2d+JkHVJWuZ9iouFkvX73ShSRysTu/
QsMlwkusNFPkw/hHu3W45HK+n4SnKzaIMZigpkJwPlJOOXqhEQSLfIYkl+ERIcnvT4u0e+d109w9
u+nl5hXQjp0kqERNCJqJvQatn4VfgouVZZ6nHG5sE4f+sVNn3inazujwEebpqwTvfubY0lXeD4oL
VRsAW6CrKhDIo5Su/C98qpFYd7PUtdRD52laKv0sGhnkQxXQOc1468b1nnRmWf+qO6z/cgjQmICJ
DmDVNHcAAybtIsK4me+JBHULCaeyXAnY8x9SqdRo2LIhqR0mEqfytZ7+fJxgJvvkYO3grO4vbKHd
oPz5yr0V0SqnKRwOjLM6zw8DhjKozwNIzzLq6yTSr4YFHRlcM5vQGCT7bsVnmKosgVpkliW9I5bj
MfVu6vYpU9IKmGrQkNZtMBxIjSVjYQcXdISWccVZ/ZYHC94WyylKIE1ruppWXav5mr/oLgA7wCmv
NqSxGRKy9eKx5D1JPfC/i+VeC2sCjM1BLWN5KFaodtQdXGtLoeAYrAqclDDTBz1r6xCOMAd58inM
4bTk0yP7Bxcm/n8rvEOBtGEt2TxMtn8KI3nJmy625GpnQRoT5ysMMaElv6TTDBcmL4LghAsE9yRZ
E6RncXzCriXLNa45qqmKY0K3BDPFegFfombDx3AVuyQeRJE0V4ThWWPrzgGPDJYX2V+GDmLLQhiE
Kk8m6snp7DZOSxxXRvo4sqjuxICEkEbwdmg8zKI7RjefC294zozHEP0jSsF7PL4CKTxNMrhETf6r
mY3s7jDgq4lJxNIv32W6NKTtbPz/nm0g+Z1Fiq13H3KVzBxMZpGf+e4MeT6aoHJRYNB13QVbuSCz
HQdZPagvTNoSvqZqthV4ToirbTMvXHCU5Go3xVJbVmIipxZiR50evoVDD8aCSuiZEDAzo9uF1ehZ
ArZ9/lGMHX0SqVWp1HElmS3/zkA0eYAI+jFncssib1X5LQ7MmWByNVVlSjD34h/FPXYs+DZysriB
t80zt3fLHjs7GKstJVeOOL3iYgI6pe2B0gB4tXR65knXj3ZzzQbylsAaR/PdAYTj9FfJt7R0GZuP
yq+QSG5SGvAbXJ3Ip1be32wBGdx3ErntCYo9L37596J3qWeAJ3N4bRtyC3Nn8a1AcHiY+P8C1hmQ
Smw6MwFpS+tFXcO+9beStyK9Sma5irzJlQnSwmHn3bN1wx6YiEg7q6W3z+2cvjlH7zyYwtgamnbO
gOtKjX83jly4YRr6p6U1O0YktnLGFMPnkJkAP2nnA0BTScArlM0uGNU+GyS/R36M5ppZfjyVdctn
koAHJ0zvZlOA44RynGjbD+r9kZQPj0K+QSzsy62ZU6QLukj4isyE1BFxh0WtyNgtiY9AaiWcbOnZ
wPB1D8plTC9+gvEVUk5BJ8ayv74lPmRAOzcdKi/0Re0lebRXaHTHSpDTn1/lCkbylx6TmONO9u0Q
NZw42uQBpw15S17WrxwiVJQZvKj7uMs6K6/r3gVn6+j2/hS/9WJ+Rr0JkSLa4fMOorOA9hZtT5YY
dhriS7ybnClvZMYsRJuBqLf3ClDMhsHhvzvMiDmyk4bMJeecIBCqv3UyNnLeU3lcqdUGToVhfxev
eRrI6UvD8OfX2+CZ4X9sFecAhODWz5DiZaKbxj5x6LW/PKQLetuyeyqi9ngLbPwF8uXuEpH7IVDs
Y6xpZi1PI0qRu2VrRoZhJKHKsFkybHJWZCmNj94Q5w7d70WGOCb6r3Opm48RGxCVM3gmmxOmVSIt
/yEggQbxJAIsipmX50piHdg2+t7fitRw2D95i6olPSZyylJ1dER7VQTNMbDpqvCYfPi+IfRihxIl
bvNNnjFMkoG3hEk5Xq7o1DWDVyZQZfuxQSw09E1B8WOp6IbQJVLJEc3V8vKBXNFj132JowIVkcrq
ks1PRNvB5CocQ6zCOn3CHULcd8xhg1kKAW1H0hTv4xNBecPXnzQaVf2EDPgCjYjXgK9/YERrOFK5
QDgJqEFeEs7FOBLF53tlRU/GXm8JmHAsc50rIjTYLOUtUXMYYJHpszcikFvCVE1o6f0MtayoN0aE
N6lFXWtK2yv2FCOOfu4poK85cGm8Y2PWhqyWTDehNaLijFdkp0TxQaQB/Jc4W8fYIuASGHFkyh1Y
UShgu+2BMNM981ZoQ2TB2lg/MxZaimwt6ORVYPaTredhGb/dWJaz6MSYhj/SJvSArFohyL7ceRfC
UaZ+rNR3LoFjpn3gtfOaLC1XrMrFnEr1FD+AsZi0NfUOS0UgUB1eweAArywqFSGW4++B4o3sz2V1
Xx6Kp/rs3ibTNDqeo0bi4JnetwLxH8DstK5sNeFqUKgBSZQa2sno83ra9etR6xNR8dP2CETcfj4w
ry9ZQGE8XxicP91aDvn3f+FgfLd/4EKXhqPKgQQJQtTG+XrYuC8A97029OtTNDdHYPRdbzHETO9E
lB/Y2uNvuKFJMJSyCi7cHTrwZO+NiaVdbeKZPVZ526Nw05x6kR1lbjw7bY833EX5BqZ/3GurXbSI
36fvL4Ql5QS66pLWGn+kK7TByFrygpB6lZNrWeqbigoUKBuy6q5Sa2j9zNnCsyXyRgCcVH7vmefx
H61qf12IS/MUDlZFl+7+ztRZQCqY2yYXdliq8QKH0TGaHDF/sWmxg2HFNFwPG7UX7AG0FypLDNxc
xtA71CkbTo9nYiTyB4Oocb4aY7ywiAEzcBydT9gbV/x+9PzDsODiHl4d3tF0D+o0z82IKbIKsnkM
azavx68nVvgTpE8LRySslCU2Uimk4vukzGwVrQOL6ZALZQzfp82Mbd6N1PxVI1pU+6hWGdmvEXa/
UsPZCM6BA2S1d1PV64WgpweWP+xsJcLJIrqh1NM2PTBq7/A0RH1QEXCo7upZW64rBltGKDKE2pE2
9bh/xqPodq2jow9/bEW9GQgTDiEI8613O4h1tU47OA6+IpdQl2ORYc/PmZoBpKSI12AkF4eSyXq4
FikKdEt4NDPtMbIW3rXpab0/8S7TgJ8HMqHzeP6e/LWH9ntdCoEKyFFS/yUKZ1ClILNgghLFXMei
zj/7FG4423SbZszHLLVPqX6UokTEXQquTQ6N3rf5hzUNA1A07usAQHH2GYvaJgQ8rMlphfShvSvP
jDVyAqnyUiSf11hA0ga29QcP6/5GtrO67ub7rAR93JC2f1XbsrwycbCAGnWGBkqovb26/9GUndiL
UZ+Pe1GkcLwZmyD8Cf2Jt2CS35kTwsxhvJcCklTNxDmIlPLwf65TBpND0BhIxYe7EHtp8f6Gsll9
Wnm7uKkKEC24fwsQ+6Bxt2PgRRU9jP4NUrC71NuJ/Ifiz85rvgs+EE1sBGjbfLER3uxMvKqLWYkm
/KsfdsarSBxleuILd+N+sVh04O5J+5qRqChk5OQamYdu9H6AFm+Rn2i93VeGIVzsyGEhIUSjaiTy
Lkx9XcZKa5JuHR62A+qS0smdGdwLpL15LwHTA7gd59OnCTXBnjcXcVLU+kEs35ogJqjJStrTGBY5
MDNiCzqUXGp+5DVDJlnZf2WNPxQbCbdghT8d/TcA2tykMRTwC8+02GCg/fHuuIo9wfSgSlBcjsNN
xygJranxeCXLKlgo0pHWHgBnKY7jRvWN5d11uMLWDWIiDvhFOLbxCYNCQA4mpQP5/wunIPcwIVqo
O3xpSdczruxHwrG+TtdE0qsvDMhUFXbq77PizYucCbYu4CpOM2t5QusIsTvfclwolWwlEV3DCCiM
y6J7Pm5rDooVHNfOAUW5Kc+gjoEcuo1xLAEX4HvqeFZ1I+SM/Gpsu3meMxEt/zv1VNHkxBbSaVOC
HOKvnS9aukYMSPuq4IGbrQklx0pVOVzGCr/4/S04EwXshLFCQ7fwXQjnd4ljY2vzAXdF44qhkMOz
TiDY8D0bLHwPNOjazRvW7fEBBaoiJfeC54gYT2jiVB2f+c2UClrBdB3cmhmRC9i7/Rn4ncF0nOyC
OYXnw6lc4rOgrO5EwvdjQdRhphh2kNUm0mkFvDo8x7fz4l5rX0j/TLSovxJQgr7yRI1A3Amr8Zvi
9iJ1KFe/jWG18jbJcu6fe1l+CYvPcJRqbpDplRvnAE9NmzkhGZMjwgIkrqh43f9Mbk7vsXKzPjrX
y1dwRkZv2OokyyK1VnzBq09Y8UkgFHICum4itqXEfRHaJq0SIdHUlbIF5G+4SkqRVqt340lSaxJm
/YjQn/RFxFS9TTRyWloiHioEkFbYoSyFkr3mqnUomRipIo7nO/0soHSM9gFpvGqb9uV4bldfkH02
82QMadx7kGKkiVW6V87GpAjffVUkEFxR5EL7t3tapfiExnlh2+R/PsjMUf5KczthzDQOnf7PKxke
Ocd8W1Lh5xrYsinCnE4XVkzss0GUbkH5E5S7spINiaEpbZjSXQzFWIt5zxvolp/JYl69nZ6UEpQv
7Xh6O4ToA6q9VSeSjmmcEzUgnHHx+KxXC6ySWp5+kAnBQIHol3y5bd3OPmxjKmcIkh08zGJsohPs
v3eS0tOQWyg+sDeC0cQsXTcXRKBPsuKIpykM6J7zbOiH7LNh7W68qYHp4R8BZJ7zhHjpG61cHlXY
xiBaRiBFIfo9Lwxa5bhTuhZM0QWieSHRcB1qfhFTNuHuTyMNC4NEp6Vm551d0H28dJy8VSdmISba
VoUXuNlAYsSJCJuEL7mpbr66CeAN9TxtgTU+Oc3bPPnJ4a/oQ4LYGmcfxedpys/WI2PaTFCYhxxB
jhyPqGHUaiRvU3E6IKvwdnBJ6ZZMbXWvXY8jwrO3fTk5SdywaW56Q45+71eo8pEMFbryg83tTO6X
3D0lsf/sARp5zQgXeVTDO3Q+w1c9yIF/oplOrNO29YE2CcP+MA+DTE5o6QIjYULYAzJ/Xe2P1zw0
Mci5IHvqXsVWSqtXlUV3g73gUS513RBUXFT1A5ZRZ3HZd4Urr5WmUvxv+VqJGqfHhqUOp/mUPTHF
yAIMf+xpHDNxjtKpOYv4t8hQIYvtatATNjVjqfNsfcchT3t0+CGZ6vwZl42gv7vruGFJAR5nQDr2
Y+sxR3oOcR/ml1Us1eBXD5HvtcDklsIwQ8Yw5k4CZ5NzfaNp3AT6RKbppi0lg1HxuvCxh6dU++vL
luqqFA8B9UCNXnZnxnFdjeVctUxGkKMSsh+h4zmJIu//rsCpiDAXPzntpQ1tyg5+IarbptWDFG1S
rx4iz4FmS/K7AuWADa9EGJxMgR8xHZmDZ0AOJotVsxQ5NQtpr9EqWXaJywgdRwNSXAjEgo55ARN4
Z1/kWa13c8wbxN6QgQI0aCmNEyqiM2MzKuNO7fhROkOZ3Chx3k/5GJyvxMZQ1FEUixT0s5s+mh70
DMei3xG3O1EqAAV78pQSkLKWb1o8APLEDINcjGg2QjmRYHz2h3z3reR6R03XvyODGeqWmr13tz0A
dG8HcVI10qL2KCw3QWPOqDkXo1V6WSgZfFuPGXXm7pBJlh2vURkLICps3fyLOSeQbf+CGNRLQmHJ
rGuVQJirH+irfN9Z45yz/wdTqBerUErXD4ZdaclvnRWThnXFpM2waUViB5exKJQJu4KXPQCrs3Yf
4YpFCEKRZ3hWhJBA2LceQGgoFAIX15y7h6IcwckzG9qEqYAoSFDFEehQRZZ8j0u6iuQJ+YpA+B5h
vtGokHQF3UgqgA/SuGezhxhdZZJIzoWtq2txdYVBDzYK3SFKNT4eRNa4Dt6ul66IT5x+emUBL/AR
GlodIoecyUcbJ5xJwkWBSiSuCUHntfLNB2FrDpLRBbrhLLWCZz6KDol3QdUjawwMblkzn69Gpl88
QZriDK6Ucpb0qWVndC7ZE+p7hpgmGhwsyXHm+qJig2bSethzX/FnIX+It8TDF7pLWLtiBVAIdfzs
pqhedNJRtJsybloqFQKSe6Ibg5iuP1NYrlA3zFmL6IFDTetSccU0OQUa+/g2fIYN+Rm4xwCMEouX
oCsAAASexpoUKwC3Qkd1PPxj1/b3m8ULEuz/60j0dRa4amyX9hycq5lZC0F3si7+/pBAan5J/tkR
0v6q7NN7h0HZ0iF8Q7kJBwqFragVs9GYNUXU+NhNOmPgpXfdk9e4ttISGNwT3jBwwyHyqDsJgS0D
zotqAqNXTm83pu6TOhcVrPGzveb9HpxYqERmXR0WYqQicek5AASkMpJpn2RftXJRyrF3R8i4LtQt
Pj+S3pvYcvNefOzuoVT5oKq1A5BdCDoEl4VBehnfU7D4A8tJ7zwxpYzixe7+Z9WQtWd3TzQYf72q
r9HpZJhqZuS2tyxhNhfDvA1piHG4bO5NxNSVlowneYLw7w0cXS4cNeACaBAkRwQ5Mk9L0/YCQyWg
W0GCILekvOGLTpf1ekGCrbBXT1kQA3jNv30JDcbkqvDvfGy2hHY4N6iFMQXKxvxxw2yu4vTlhYxr
eh6HSs6MLEsC9nAz5ulxhFliYaoE0pbQbWpcspinEeJHU/gXbpiI6EN+ITMxgRIFiNXOB8dQOwSw
aYF8rduVJdF3JSBQQsWjPeqsARpiDlaNU4wKeOSnoV2IlirVQ7vY143onO51LpgurXzxV5/IxSF+
bTg0b9jCOqXPR576TUPAYx+GlQyBczBKfEb4Jxl4M39y48bI7oaIiLXvzg/NmtGW+d9TmBx6AQHN
iWUra7KKNkKI/lG0MlftI/gJtH4adkOmu1JdFyL5qSHhz8fmmu68w81IF2jEEnBCbkMi8jRBf9b4
D1R5cGlQCDmSh3nHBwWEVjA2INtNfhjJDA/E4iKtSf1BnMxx/wkoP0XU+ILtFM1VuMyhScj3KPDp
cSbBhwfbkE/oOMIxJn7d13afd88bwWTuhgc9v90l010PFMU7XYFXRfWT0E5UsY4+XwW1ZqHURaGk
JMWT+2vk3nlTk4TXSKZRWNHGozPyOH36WgRfMgkHKKh5SepejhyyeanrwJoYDkbyc80T4mehEU+r
rfFwGBBfEwG6DDUsbfdFD8AoZg+GZRLr+jHeNkuWSxQmbbWJvLSFzBoVHoV4cxbYKdGpHXUzbc4d
A3Zh8SpMkyK6HYbTR2NNQV8FmrZvOy/ZkpZKU+VdWoj+I1q+jOmc1RBJaIx5zz//jIDcx9ygDkwx
lK2TR90I5C9rOQS1+X9OI/nWqpiqz+C/JapVEK5uTHpF2+cujX89LV7egpJgcD3w3Jrsd5UIBqY9
Sn57uZ79tokK/HyiFyQspdIzS9RgDFV4XxIQozUUJa/oVL8tlzP4L6f1u9qwlr8r88Owbg7mQB+4
izOFJ9T87trGXLLHmOlNvFJhIOMF4OWaebJICuT4fvnV1dJrEty56in6aaE/6LqE/K0Y5L3JvuGb
vBBGITFnEapubIFDQWuyzYadPXHYvBFdevXBtnPDUlWLh9m9DFI+39ji5K2noXPfkfMOvrKCvVj8
Xv+K187anUBLh88Npd0mR2blssr7kQwwLw10j08k4KWOYqDc9MgsBcicXAzB6mfQM5rOj93Kewfw
wpWLtaSw/0GLLQX2K0yQC9oF7H7ZZppZfV0kgge1y0Qh6B8GfOSlNR+HxeAlX89DCwugEEwKoSCb
3dDd4tSHRl22Pa3JuwIQeEbLDVlEavoU/VTewOvh7aVDFsUzl441MVz1+GES14uIknsC7pwI/iKI
/5nrv8wtDKGhN30PcK9sco1qk8qoES/uKSuM4xdpTldlc+a7JOLqdJhSk3AKU9dfsUoUoudfBtNd
MTNTE348Efq0wr9A/6J4LGtj3ixU3RkRInaQ9bZ2I/Xwo/upxq4xwC0X0nB+cgMiZkXC+h1Iehyg
LuEkCFBU1tCiZTtg7qf0qXjXyml7Kf738KqcOdVzeF7D8UC5R+TqNttDYJItnl4tH3nB3bw5v8qA
1wKyLxnUWXntKp51nHcuaFpliyYGAI5dGA9UCEJIfH4kX0DIpffRSnTBQ1OvRE9WGncB4YMAQYJV
gFpTxe1qCnUIHc1+Qb0mNM4H6tjjUFql9tt7uXxuA8HoAcnwBlzlMG4i2eOw1dSppeSKydERiwbw
5ucL816QcSP7gIIyVi6r5lv9+KukZ23R9jviioSYwlHCweiQb5Rhp+1CueTwFh/KGj/86M+1IdI1
jcKhrG1nwpFkfPVcKAYbsGy8oW3gZg4IDsLXNBlceczpBRh54R9tQDnUZZKJcfv8qOdpsPi8FK3b
tc/n0ox5BZlH/Sc64qTVZMEpFMyNzXhJ3agx23fd6lwLODHIS6gZ8nBqFCvL0YBiWn6z/fm2j++U
h+blcXmWmiKTzlQ+TPYov7CH0IxxpX5rH4eg4HJFrZPoK6kO3N3uZVvzFXdWpzTnzufVA/nnq+jq
ydNYPf5IRK8Wd//N2ZJxhDhCbN6acpGMZzZFMd+4FcsWuYhnnitHMyW56HK/lqcTl3eQj/jaeMzK
6zYV/HUIEr2QtmecCJc7gsgM55lg3SjXRutFu+tfcttOKpnTepR/TnVGzeyrPPknGYyb7oEMX8mC
o+f+BsCFQEF5BukJo12IIlQp3XBpGmlVtz57UbziVEkAlgDpexCMM+LCDCAkiT9iip1APjikSep0
dx3osl7I3aBvi44XsKMejrMG91JiO+XzN7mwElOWmgCpjB/mevEB5rmnAE/y6kA1bss1ikSimlV3
3RtKCciWACVP9tpY4dLYoSfjG249wDn73KQo/2qyEUYbct1Qxyk+SmhlCkTip5fnLObENO2ZVymw
kkxE9K8wTcRmF3alCGMsTk38u5WP2vsx2DfbBMptntUdjTcmbmeweYxeut5crMBGHnd3ZbeOX4zZ
LhltcFoo+ScPeoBn838NIp+V/06UAA5rW/l5VlOPnKypWQXoncaOL1rLImH2QimaGGC1XZt+7wJ6
61WtzdcgGyFiTbn/8DKoljwaIv3dDrj9X7v+cT5SR6eeuBGQT9yoCXToJ501SowqsF4WyDya02iD
8XnxKeFv3SbCPS/JldaOBOuYp0lkbxIXVYTjcPf+fya2++nBABYRAZM9kxH5hCg9pLHetjX0SmfN
VOZoem0eqwHZY1p3RkGxgFIjdwA9kJrCQ8z2S52C87BkwpwArM0/AO+Pn9iE8MYPhgwjepH/63Rq
09HWW0dwaeyQTJwsJoaDnMXq1S2RNKOD2b3BORNmbnnRm2Wkd3ijK4fInO8b+cj4qKsYY26/5FxJ
t085RqjbEqKHRWTeqlP4iBH/To4MNrw7lIJqY2MBXOSiFGSdy+QYcrlTqcmrIHiY0ck8OqfPE0fC
oE7F56hVL17ViTy4lxbjsPSQikB5gDcHRUItl6x+GTimAolmCVX+tgE2YdU3nD91MTgDOQ/WHtYB
HKz+14tSYu+BjogPjghQ009iZI3snGkvGu1OZuQp1eGMQE9kOxVQsJvDb5yS0DjXWLS89rM8KsUi
tA6JiA3dT17e5lQGcL4SwA8VJy0JxQRF7XfWyp9MhPcO/5RL3abK4QfHg2UerXLCNLkubLKuug/x
EqgWNNtWRfp/1xGSDWEaai1R+m3F9DPkmNystP5agXESYxqUJ8rYBo2sC43STdqNne7W7J/Y0XJL
L0VQOMsKo4+hIFgOOOsvXlzIUGE4oYsLam1x1kkr5GoSCCa9dQDS4IF890YOv63AWMbkJxrZIlPF
9E/8mTSXk4TQOSVk9pfhoQu0Gr6Y8PeIu+xaShCu34U6eVJHHLyZO02IyiX5U3otIHZTufHIbCNq
f9REgNEsuH8/0rzISs+sfEezjAnq5tHpVKcTcnRJ9FUP6htbdzlsYO18+VQ1MvPLPqjCVHeYlJaq
Ulo0AUjp+X2hdl4Bew+VkTniOmHoSBqJn0MmrC9g/pBUuTVA5XciWu2AwQH52yz+MvMfR23oGse0
ucD2RS238O21V9tLORT3TvDqw46FoZvVKv16256bHoXp6HL1gUow3GVjj+eSNS6hjWCnOcCjI3N5
s+VSSIfw7VpwpljOwsOizZinD2KMf+k2N2jSVSUBCVdZBhKQshOL5al8soRFsRflDM03Lb1DjhQJ
uFiZMj/krImcXgnYB7pHp8y9PTto1scBzEewe/Xo9pHX7ghij9Sn4Tyg0hzA/ttMzg3Vmj9p22m6
iG1Oi2Bj5Myzsfs4AoQ72L8Y9dJvTeQ/clv6ufUIuB54JjI5CDahS+MufT6ie8DlP3bbUtgO6au/
jaIg0fQumwBNj0bx0FMqWBgiIMT4rwYNCzHFXTziu18SM3a5AqPpxVhYY9kRqRT1OjxFnTx6omEw
GBna9/j5/S5mTD9g7POk8zZCu+EDk5MujpoNOGiQZXkRAarQARG+Fguk4tNa2hRD055gHeoncR9u
7APwuOllMof7GifSnHGBwDXTMG9a2/USKNk4SQxtm5eRWAV80YVHzLMn0q0+xOBdFSjC8gtb9299
mVTOGemUthg//rQithbmoAE98B8OYYNHlCsM2XdSUxbldf0LaofNduM3n7NwelnbxGqwFEfyTjq4
IbWm8rSltdgIceXFkptsHYP6nTSUNXAnM1c8p6lX4YWlyYcqfrKbVg5lXIO4ywC6tYmJzFUi7b2A
UXOUxnQVfINoWpfNd86FWEa83R4WFoSXgA2aQZEblAJiEjda3hxta2AP0KQdnV9ISPCeiOrOE0Q4
+5YAyMBso5zUDc7a8ESnbZ9XgbanZJauf2Ti1HVB/bGJxMRUxMKpBrWqqVh75VnRBGpV//DacvfW
ndGexBdVicyuxPHmXEaV2EZNw38Pj9tOaPWxliR8vz286py+DnHiveW7VeGj8xuThWTE3HQTTwmw
UManusw5RgGSnd7e3H/m2HS0/NX+FfI+2ZaLL9bSq5/zy9E60uFthElluznMhg81BpKOohT546kH
TgfTt74SNJWJFkKzsXH7aBYHFWtadWZqq+r5GhMAalSbuEbbEMz51qwJq12uQBL8Cg62h+rJgAj7
22B4Z0rapBOdQtW1UIZwHqZ2wN7D9iOw/fQ0tfEXvBWGEvBqki8ai617aAwMrOOD0bzkIr5bbfGH
hVHTM4ztbs6/SmalMC6nG6fA7Q90RJ7tLIr7MJUNsrqK1DD9mqjSMYe4dKNp1qvwRtyGLByN/M0+
rcFO/PV0UezbVZ/71NHwKYc0tqs2oaPwhAKrhrGomUkQHQbusxcLMyHoQ1GyRMWHwBE0978ZIfQy
/473QIgIUrtqaG8/97Tb8udIVOO7B/7ohjKvJAP8to/EFFBO+LOVsj7ndiNON8TMnCmf7BeQTgHP
IdZ0TjRLSC3Of1N3de5EGm7NvB3LNgKse+vFbHR+YZ46jdiCej8EZNpRJjGSp8cICMihBq0gaWBi
Qd1aVObOIt+hLkVuEd0L5l8h1qGeekEnX64E1+B4gZRPLyybzX1hkODZudmoGAseIRFoU0lTBsCM
v2RH65obYIVtjXvw/JqG3molciOeJCytPC99ZW5m8pLIIS62FQ9X0mv2g2nP+JAg40cLJSeJ1aar
cxIRVtw+QsURVAcpm+SXvX+iAs1TiVKlMxoeX7U1fRiXNbAmcfyt0jZqv2YdSrGhN572lyPaYDFV
GhmJoLdCAJPNLAQbvLMvHfldnrSblLITys0v8ieMD/1zg29OKStFnzisxR44NfWIEeqvf/zg0OSh
TgkcdGWa39n8tIXkWyMmNObzDF3cPkYQqHbhQtXQy852bClOGY1jadq7Msxjb0oiiI8p0zCY4N0s
1ko3AKKWddJSyZKtC0Yvns+2ync1htuaNMHyuinnoxLgi6NwpzZWPppORtSYdP8OE4703WyW9UlV
Z9PjBQEkhhUg7Zm2abXyVnS4bhdnC4orAZhhkKBxvT4FFtri/ekxhzjjXwJb4J84D3kJ77ApDj04
3zDmVLGOFtFx8C4UwLrnGs6guOWSgwxURuRLewgdZ5Yg5xMLXeVdQWzscb4lC7S9IZqW6CSa82+f
o5iymxX9MizqWzmFICg9dA8PSWa90tz8yzx65I8UTUiOkvKJZTmYoU/1lO0oUETgT72Su5A1tPIa
scf7iyW+QRQvVMyZdjKzEevmORx0+bOl816wKKGOpOlgr/B9n211s8qxkUcWcOJstNbsyQdwo581
Jod8Kuxi9zX8w9GrtcCCTIvuFl28T81cBomNo9Wn3g1l3tKrM10wtS4xABANnP3tw4nko544JdfL
uK4FLqmf0gbqZR9jD5iKBk3VPDCPb6nDFMBbvplnYPO1Nt8QuzWYpvp2xmi+U+dCiba1r8hnogTj
31w4wfWwewkzz7uDoqf8FM6Ttl/aCQUjD/C9CTKAiQwndHx9pNjHMqwLVD2GiHNoBl/5RZkccJAS
vV8bNBK+8EvOYefRO6f0h5sLiwsjsflPfKrg5zkO/aqV1QfYOc6HyPwMogPvQrX3fyBSZq8+ZTkO
kQuHzyzVtHOo8z+TeUn5QJsO0cMz+twVaSHzw10jCMZefR1kEVp8oYfyDiKz4Tu/6iXJX4NEbH+Z
FF4B3R7NLJ7Z6RG/b2C8rtRPWqu1eTewhRUKfOTg7+miryPDbybEEOtA0qLVzY4xveuqkvK3/AhV
qVWYbWvrTObtZGylG7uC0FwZouQv5ZE2+t3/db76amm2r+Aezv7hTFeiFf7GFzf8Z3BhJt0pGJA1
Gd3/0q18tgd6q87610w1ZPVuhAUzTHAsF8EqheHkQFlt+hHsnpkwJ0Bw5ze8WKBtG3RQ9kmtWuwx
QskLfq96Y4FjMWYftcLCkEH3IqB0rLnLVAmu/wNPXeDxx5OjIoTK71y7He4sFESNZ9SE94WywENG
I9zDTmVUzZ89wgY3DhqMidRD4N08mN9adBRf+3sSeKRnSX9/rkETkAsIUZn6g+Yec7HIG8qV+c3y
mLFPrwTOyJikPl0dxs471FDwAepa/I26VXHddPgTIDge8Em+a8uCjMvogrdtxNjrCeq01kNc08fJ
7p93nENG2N9mc/IZgxzH0/FNN6n/Su1jpKOUj3S13iQr+rVDv2aNf/4Zxg1dIrJZbc/LOCsqajS9
mERozxwFeRFLlP5QUtWObh+KxttNic6cP16wFscLnuAyON63p3peg9jVIZ8vry7KpHN734oTHSCw
kjVfClq6RI0pSool8dpW66fXhmrHMYz8MtqUbj/uGPUHXH9upQl1pqt3eXf26vQuDY0MQTj/D448
uYYpa090MAdARFMzduVef3sHxaBBApiafkn6q1oSUP5Mc/fesLlqZvRMTE7VNCtZqqjh8EPCRq8A
aKCGmfQNx1GbXPDcZ9icPmyXcsbGR855fvU2ZFrFR2w2nXPoJyOMcbN0r98C9mQqnbsKBxHWOcP1
LeXS6pvl6PUVVHAAwRjUyB4IVlkr7sRqe40PDnw2FD5QmheQg5rjTumRJ8WaBc/a418wZHf2blzs
egWWVwRTvHatedk1t205PN1OxzrzyNd50HwKHOG1Mf3Mw9NT1Se5zT9RONEHpGvzAG5ZOBGhLFsM
X9feWvKYkxtG6NDuJMptzK6HhBQ6Z339a0WPqwSu/40bI+UbGHwod+ii75OXlc75A3oDXzWuCbRO
ZhR3WdN1fS7hFf81w6WbV8tMcVVnydyx3y/1LU7DY/0B1keVyszIjerQSa3yVLHcT3h7aBCIbwiP
FPji2aIowUWNyT7pcvxeNJ+3a2UthphdGxUEpFv3SPO+DWLeVQxfwp3W+A307ZA/zHIQp8/XzY3V
8rnHmcMgTBXDqDQ4nZwirzwA/9uLheKJXJxcybkMiBGXGsuoSwYm0Y2Zpnz1vCBIHjEF806kkyeC
tI9IalP47WEgNnD2hgPyzus2/3NIv+yydaiqFI4kRnpgcl2gr9x1tUZUFvQkdM/yqG6esm1aeJK5
NENIFEjjBpBWt9ONpQph3huA8AT+oIBlb3QRZViHFuic21SNqd9PFTjMcHaHdBrZI+4ciA9O5v7X
bsxjLQCzYxCwJu4j5vEUPcZnWJwOyN6zRFkXhjE9U/iAS60mL4VwM1xH6gbuDWXt9fUkudQ5WbDD
6DxSC5vI3x50k9O3dDmo687+GevpEdU3zj9rCuMS754a6WWBDnEKows0+t9ComddnDx4wxIR4KC7
M2D0wgDiqJZKBYZPgmwNd12is8lXABQAdVrHf0t6K5S/jz8+vxD5RrOPVu31EAzQfMdy1tsA5P16
+hTIA5uI8Dh5B0u3v4hmVxUAg30nq9ehcWPtqG42MKfmiBH/yBBrRDAWZXecbrkiDMzZsEeTPuft
qNAJDEHy2f8+ePx5a49S+7ryMqraKob78ZM0H7Xrc06T1wAVr2LCUdmJoRd3rouQpkfdyYDW6fv9
qKNL6IVfFR+2jXBATynDVmUycTyO+2nck7ZlrMLRjyuMVvBwPjDso7eXRZ5KEY4kTpj6QSYw2bRm
crRvD4Wee+hZw0TvfwX/PMPlNR3S7yfD+dMKoXHPgK71bZXYutvp+PRNitjPk2SZlVuLNoViCgHg
TA8uNoVqAZGSiVztWjbxvJD9768BCjBK6wFMZ6HblLeJX1xBpoxxW8C13XPvQJl/pe1V983E3cqq
ZAsRgD7shY4wwJwT8mdHPr8BVFi9iPE47Qt8eBHiY+l5tjdWZ7M+S3i+cvellLVJ3YcZki/FkMZj
P4H9yEL62om3LgRLzZ0TA+lW14RCvI6fBjjifnFmsApAuhlprgqcuVuIZ7chThdisgGz0vXOTBkA
gryTdagqT/x6PMjlWWtWHjJpK5GCCTDeFuPbcAdy1HM9tKw9ZElSB4eyMT49sfU1xzGChEb9fy0L
nnHDlXHrfrBx5gmyy2BB18MgKvoLK5ZL82ocAQzzRCayddeXCpCnpnEsxXXlGmIQEMKUoRNb6lFK
NuvMAvuGxvCXgK2F/A7qMZYECYcCnKkjmegMskBUDEEKvQW/1eE3t7YGDyCMC5fYj2nX06c8liX4
z0lzlQV5+5X0ufFIOGWqOlWfrJi7IqRdDIiwRh4eSAvLlny2bJQRB5WDVdyVrGaV2Y/ZOhXJ31vP
mNsKgVJisYea9SrH4pTfxUYnx6MHQoAsEhf6PZscr6xu59MXOKOiLRRTUl9Ak/DJDqQIuDQNsf4Q
IGVBA4zqAQe4zIIc/bTjkC5drxyM3BJukZs1XndSmwCxuX43l9H0Ot8UqE7DifiF/SkAoJ9/n2J4
YNJdSj8WqLFSSP07MH/gMkgEe+4HuPUFDGKZykna8AGamnkOfSQanXygD77XSSbCgEn//PltNBUA
4zKh5RcxeBadA3BTHizf/xH5Bh+icnupTqIGJB5JewYXLrnZYK84AiovMmSyVLtbKr0pFVZFuXL3
3P7yXSIO7eXOS8/fCdp+leTlnluIKW0qTeiNlSs1Fc1pl0/nwERWGbpJv87yayA68mY83SPA0R9i
GHLm8NBSvyW0dSq9v8AcGStumpLgeyTLXp4SaX7YNI6tJqOhO62sNWfGWsHL+bA5i2KpWQ3XdJzr
2ihkpCjIsuALUrHGjomH4JtaTKyYOJVOquA/3OQonFZkxR1EQuimGrzRCGmTd2gMSCeoOKvwQfHr
2QuhtACu7VqStjuK9aDkxSgYH5voq8RWebqxKq8BoA+8+7uw0j2PrhCAW4PvgEHtEn+nPWENvv6H
Eyj5zpjPtJTCkwASDSyfYd97wq4jZ3otRLKtO+PRbrakphvlxgBorD3QxQA4qtj7H46/kup/xod2
O107WVDJ0fYiHDMEyhuJLioEfi3JuoNIlIunB//YLAswGp6atbej0NO/Jbxb51wzKztQD80Y63zR
PgEFXUpDVe8CARNNZ0TvG0WF+mkTCoOKh8pOCvzAj0l3Hchf0BSkqnGfupB0/iZVecBfdrxaP56Z
yghHMeLhSlVEgYCGrmSePPypetaNwUFE4k8fGwv6RRUOmxc7K4+3/tiS00PCjYG3vKMKy9mabjgg
onHkGtPzjJr03FS6ejUJEgJYfUEe5UOSvH0d0a0TsyULBz06sqNtgJtEliEG6Ipv+GHOI/3hAtBE
OK8WIvzcas1xf9CwbqG8tHHe2t4mbbyZel+TslCVgTBzyWbJq5IN6WD02uh7A2S82nTcI7wWdzAI
Tly2TrsgbMfnycOz0lp+QhLHmTkDPlW26S4ZsNbGdeTW5N9SBScvNSCMMZUdMmM+5fonnImLIZYS
628a0SWU0YZ3kkXwLPU7/tvQ24VjGFHh+VzkcYBn/iukL5Gr2TeQA0kmpbSHionOs/00pCdtvEGQ
wYuDRkIZtPKP1kN3cmSD4Sb5jJaGugsUErllMgMmTX3iqVf/sadtxYgwQ/LC0xOGT0P4XkL97ePS
IAoF9bIOfpmEHPvmi8nTyaoH++RaW6Sgp1jlsqmesrugbK7Ab6VE3plgoWDYinNneXShIPulWn8Z
hpTD7tbCYoyno/tF7FFGGIRUd8+eejjXKGujv5jy4axSjRrAOgjWEMShLtF/uUAiLCsZkd9gLQVz
c3MQjVHlhn08VbVq964RCX/YXR4nDq5JdIisdAXd0/SUnnddJxRA1K3zZRI1h/AIoS0FfFSV0wdL
YFUi3F9QdXY8OSA5/mvc35znPnb9bEGzDOfaXOu/QOZqHKrL3qKeeR4f2DN7jB/uKZzGRQ/ByLfZ
bRbA3GWkS2OJOk2S/J0L4KgS7cA+e/ZRv49PeOM+rmYYWWr1ycgHIRBT+6iKk8sROsYbkO0LM97h
9EXUat00NeHbSsbJ8dwTitjCGun8mUPCFOddrOGRheH7mHwRm3KTbU7hTffNbJheS7bQW6zWJHa5
7+q7CIrp4ykNdkHEB3IjKmWTyltz399xkQSliUZ0wvwuAidFIsOVCc4s0L+f7jTx+nomk3aesjH1
lOoxTK96DA32EzNW6YFps6bGbIQyTcHg6DVALYjMzTCQILkbGwCbG5MkoxCTbaxbWBZ9AM0qcSf1
2Kv0Fb+aYOoK85NqUPvQjZ4PQoHazNeYwFKrc8lbXhlBlaLuxZ84ZEvr+m+DCyNThF94r7HSrB4j
ohvwR9cxZ/05zg5XcvjydUNyD2IWUdecpUSsWEiUKA+kXPTUUbbSCVzMaAQXLt3EO4cuMzjYRWBv
BTAq6p7fPwO+fzRfM1C3UYYg7gV9DzAvwGoOOGcbnGLro977upSIrGOOr1DPl7slvImCCgpkdG6n
6qYtKqaw6Bi+mVnYokkJ3GFbrOYJgku5iIlDcmJ7rWHByUjz2+seOFB1g/zBi7k6eyRlZBX856mP
2ES4QXjZzXuxv0Yf2jZqJNF4y/yzvNSsXbnbHekoyK8LGugFiUcfoiL/R8ggau/UsvFD4DcylHNd
X51lIIETkPCRk2Tf4W1VwwlZDGQrPNKIwceB5+AeVMd1BhXCMyozE7ngDgpxU96wE+HfPNRqUAaY
jTCQW2KYa5R07VX/OUYwG4dZ23ufDG0WSlyp9Mroiw2tXxtwHSRGhZF5VOkr5YMi/oOA1jGJL9iS
tkUC2eLUo4u6iqFFXaG78EFZPslNBZeqzFZFiP5cB+J+ajZ5nlrqF/KbqOFRQLXhUQ3X3pALddPI
ZFhEUW8v6V6Kc1bmRLNDRyqMRMTdOxJkTfrHnrJ2AkrGjj+yRPzIpwu85SDrg7fnprvyXARYU8qg
Vww28AS+PCAkBRTvKvNxZ7lZcCfunHipdKoUXt1GmN2vL3iesd/urKKj2bMFbZaF3wI44an65oic
EOjj9GSrMRsucSOO5fxhY5OyUr1F4RK+jd5ftG0xVSMlWGFY9w8iX/qtS8Ftwlk6WzaK/7CXI9EI
ZjHCupeBDwqwGq8BPYL755UocbP7rWqoA71mP3wY+Aed2ndxIQv00XdCQxqfWQVslWxNx6DsWueI
+WtINMkVeagjEnY4Gr0/EPdyBXidD9C3WF/Bi4VbhXJ5IWb+y/2yRMxkhAoKl8MgCZIrB/FQ1Toj
ng0Ahi2PXmgelB59trRG2Suf5xmBLNbTf+lBVQx7s5h98Orm1kJvIOEF2jdJIsAvuUoRUndfOmYB
MNWecBYMEN8o/DOeAQLOQP6x3sZ8/tL2FYOTKnO7ArzPNs8DyBLh6yVPBQZQ8QbFzBzXVR0g4Qvo
FdlCxTYewqonAJ4RhTDWKuIO66z3h1MBx1sAmi4Hnjix+wRbokBoz+S6VKgYko3STuHw5ePL5+G7
h+rV0UekM1BAohzafwbvDDFffi4miduoJa1B1V0G1mAlRCjjO8PQy+QCtG32zaC2RHdezE/nSYX1
vbvTF9hV35CA4TLoj4dNdJEG7gbJ8NCG5SyUwg2n/43+wPAejw5mp3tbKMXTRDc/t8jGtpKXGp4g
+7lHuy3wsdZf30AsOefKnhOst9mp8vpBwKJFVL8QBspy4RkV/PhbKjnvjJSGvt3xcwau8IM2rG9l
EWCU7O/wrvjGTkE10sSAC1Ao3bjxsW48d5WJPHg9zsdYqFD4q1uNYZrGCTKWWhizqtlezmb7XAa6
T5ahT5zzykQRoXk8QNWhBCa1BbbebOecNbziOiTVU+1fT38adRW0OopORy/K0J42as5gUYW5Yxjl
4RZ5oKHvCRL44EZj109d0NLpC+0j8PpXOoSUMRp71H1lzAI6YdfBhmUwhUTGM8r/HobU5ovHLcAO
UdpkOkO0Fp1RYW/Z6AO7SNOXq8pWLqVXEsKrUq7kvspI+Omdve/TSzn4v5lYtNPkZLg6RD/UGnbM
fAtj0ZSOy2PCj1KSZbJPBs5eVNDytO5sCrB3m0v5kReIb1br6yKc2j7mK4Arrb7UAyIXsvhzYEk+
ply0tTgKoPtBeFTOu7LwGPYE1AUbwOQZ0sZOoUAHdZ1TjRKcbBUM8567R1wf5pERtPRCaaTgIasL
1PtNKtSEfL7VZD/C/qml5ebrUG73LKSufqZxNLhjoBIibNNopq7Pt1DCLKoEuMkQbhMJLeANTj7y
ny9ccds20ch/2gc6WpLx29HtmFMZ5d5uIVQRULgcqx/neebOqPKY1RnynhoNTUCEIUWto5eSCJsf
wsQktPJLVu6T3FXg5b6tS6ttuVBWQyICLAi5qP7oYC4f4cB1H1M+5S1WUynF05nLgJHEiw4eSqDH
qd02Soo4Azpkrmj2MCO6RFNRnH8lngQKLP3xM/iHrKC9kLuFfqpl7M7TzDAIwVVu5Qy+OaBt2CMZ
DZDXC9wSHso9/dyitFZkC7citw1lyFRyUV1hymKwnC8dIN7dMxx6KvZCpr4K9teie5OYMqKJKgyM
51Q9EHRBD7+9Reqvl05VjmHkSRpJFfPO3nZtGu7tMh76V1LD0/JfpptQ5t5P+aDolquDmJqp0WG1
/h3bu5DMUaKOqAivEAsWL2wz+rsAgSkbTsQzp0yb3MRz7w2a8Rk6EVlhaKfhsuFBHsmWc7icVksG
NuYig2efPwoCetWu50yeRyBB6Gj7b19LfSZgit8cygB7fkq2xEFrChkaowH4gosSB7oaE7WLK/uI
GaKtFNZ1qrIGo7Gtg9uJ79s5a5tyrv0kXRdhK24GaEDNfMe6mfVjbbbhs/jQx3LENzGS5YSC3VfL
6TNTLPLoMhwPW7NbXHwZlGo4/rBwrB8m9SBga+rAvdjFvZiAIsZdRSYag4siFYSEzcyM5HMIobLG
6ISM+bOkXHEx1hgT8CcnmWcWAEjG2zdbVIqxyD8AF/GVZzoqrOhpsNP9YutMw3cqd852VLcIl30v
9/dJRmKVBT+HkATu6EUNsDne9K4JupkTfJX0nXn/UjFLB/EfeIwSQEsChG+4AwMOTK52zpCQlDwC
GynC8sEU+ANfVPWYZwvRHkkzILYsRkrvs5urbdRrbq8lY6nJB1+EgUi6Gkq3yz84VYINoiQDSK63
tl8lQcprO+aO2JYNb9EwkJhcv61Fkfc7picEtf+cN7xG5MxWoQVpXwOljYCq1B5kVcSmcOjF4GEz
PWQUTy4MezXvSf+duquLbWgftzDghnvIIMrf9Gk/0/RvHckxOBFqRV3tpYoNy1IWquMaDfE6moq3
LafVcmelN3hyZu5s1QNNNsKb8Yt/jc+G8URnmX2ml0agfWS0HmgtvdczCJbgu2bNDk4+1ATEeO8G
n1Zp35Qj0mP8FDcRacoBNmGeW/SVye4r/beJEMK3XAQ+OABXRqbDcWCoiNNdj8ltzf2E51uJSbtT
mUAhu+YPp5HwMGG1j0/B5u6groAMll9n4eUBlS1EIrYGSQOo1vBM8LUUWgjSefKUNZvHuQlMaYSc
rboIJ7LZoXr21nMQbrA8I+In0J+xVCH0lmMFNGfLBQwIr+X8Z7jPLvpdeZYnmSIQtPJ6sHbs+5rr
om1wz9Bc2O2qcU/tsIvuqbeXcu8KrU/iEZRk8YeG2VAABOU1VCCeZxEKhSpTGEmxQu2HpOh4twDO
q+88OUw5sewROvfvTGH2cjmFSsNnR+ei+d+9XHrkMEWR0LuzP8Z07PWYIv4axnfn04L+IplVToJ2
jCDNPjv37HDHpfuGk18/GNI8+pNoUYvsacKCkpmfHfM5W1Y2lnMEdwKVlcDu+9w9cHgG6Xad4sJ0
2epz3vGDTfxMnv8s660mxDKdkfkPHCS3+KHgx34olhWO4pI3r0QT35MvELDTQgaWpMhU27SEPcBA
bMHXE3dcEgpp1RJLOkpnQzUaqkR0cLxxdetGB/UgyWKDEV4kXBmUuW+LkCWmnkaQfGte7oSB/DvS
BRvpLm58wt+uk3ixUk2iKfkz+ekUXIIx+D+jcMLg7hhKqOf1Jwy2f5uFMWkoVSYIIUfuSOVi+0Rr
Owo3AqQvtRd/GyuOIxMHf4Zew1D35NoWWmLBEawkKZmNgUn2pkRSIBPYmLl5Euzm5TOabb7bL+Dr
6xGm9CVFrLp51S15kPgcl/fL/l3fPYnTSVTJaoTMfRX2u7gM88RuPQi+1gikEQ1BvKJG2w8mae4C
n8EiPPRW7ZuPwWvUofWU/P15U/68LhmVY4fy+zXGuohd61LNloGhOJrmxdmlBv9xLS/DqPlXsENd
nMk2VyNG250ogryzptjY8JXR7o3rD55BaPxW95Zg/c2lHgL9u+5mcbWr4EbBSO/9Jy5de+RtijAw
T73vEuVP9DQkBnA+hB5jWlvPRHi3M8HA6KswFR5St0py5MmyFbsV3EE200wxEzG7Edj9Luh74YDd
1SPZGif19COyvnEnO8IG4c8Fa7+QZmzW91XkqDsaJk/0LYWOD7/Km8/rZtK8Cdu/836WpGde/RLR
EApPiQS3LDXemx6NmY1O1f/rJg1oecK4gMhsMfYY9GC/zq8GqHj7LsiRRmUVkcDWdNRgvPFqmHZ8
JzJZukplKcw9FbdfxbmJxQyZPquhZW+iCQlJ3coD6kK4JB7wInY8O2jj/aXP680ILP2v5JYIQsZt
yxmK5HoRNiFrnq5fIewR6EM594SuVnYIBOhnTZ3pi8rRXSWftzPDmoqsy1PP+8UCka+ezuX7onBE
BDFgKwezW+cQu5JBmpYQw0I6FbpsZMNDm83Xvnq/KfSaA/AJv/KImdESf2mf/ckBwjGGc8MOX7/Z
By68A2ZUE2XAeZlzslmz64f3IPrXraeadUWQb8ERa21FadSdqjV1OFpwDDEy8Qj+IOb9jd7FnmmQ
yw+iE0ZaP7ljptFOscpPCTZi4TnVXTp7/xrBlggifOfUu7JDFM5do01ux+Y/mQYaZ3bGFKUevR2K
lgrmCy6KbGDnZlLGgEbTwRrAqGY6Y4i80cOOtZ1sgT6ZB7rSDQ7pr/DPWugZh4lCdRQiquRp5cCr
nF07JdMi8z/MwP/MyYQ6IuFT2YB2FnQIN0l5UBsfiBdSRzW/txGdeN1lB64v4K9VEzjYw933XiiN
XNX/s3beqHE81a/z79oNDud6VsZEunX4tpGCTZCJoif6gmx7ENgrz7zJMX65rGuUSGzrbxy4L0p/
Y+iCa2C1mlqHlKS9uoMWQwJYd9s2lgH44JGzB86GytSR4meszF1c9h6Um0fs/CzQnAFWHYdiPPGj
J7OSCbMv/RCkqLBMaW7+NyeLQZyUV5LKalSh4Q3jEPSWxWYpI5JgHsQtMs2gGlETSKxG2mf9gser
80v0ph6b24JsGVgfvyclvLKcsPBY7DaY3fnPQQ22QCzo56WuKNiF5nmV8luaCBmpXxs6I0Han35y
UGkP0r5/tuBQfHMx5Vq2yMVUzx4PRdnN46zQz+f5JimQvbzdHlO+wat6MGRXb/nRCp/NiLjpQOIj
wNe8URbb/cNKmmBP9tQXsssQHrCI4xsKISZMZ8qT3H9RAjLZItFsM45qO72wg2AlI4iVZZY2ByiE
RfbBmS+gysGxYM5QwmRlQvMys3fAtlQGz2dVIA1+BmjWKNznzjMVbpF14NTouxNBYoWZbepbHY48
8C6Zz1pxNiFTYXRxYXVwR/ikSl2p1Kt2Sp/Oa88UEZfnqEZIRwlqjphKt+8P7X0WGoOwjUsdh0Ny
W9UcWtkF1XbYp48TktrN9rHK1PRKmBaHst1ieZpyO2tYFTJnInZRu/izoO3L1y/A+v13E6DdkK/I
EOFJqURvdrqTFNR/4d7PCjC74wJX6owVdl7zlEE8OAPLvFDpgCsiqTUSaqHSKRssAcnbk+U0hu/7
FHBAgQGAwZTllnVC3QLprvUoxdfrQw6jlpVZ4KgExgS07axQ6DxGUPa2eZsMQvrb3b7pvt40/tpy
SJFKycyjrXBs5Xs4Ams1baGaInazArAq84StLPkLcGr1OsaxjdRucl8eAenoMCce5HApLkPpkkMP
ckt7Z5hYaH5c4mQK5KiSMGbBM1USJLNEXGPJC5k/TjaOHZB/Br7NvXuFlp9B7Z8CTqxOgIHK3lBa
UmLCuiVDxcsbxJ95wQZS1aHq5qBHnCKIDHz5n7xcpDNffOf4FN+hC5lutah30gTB8X3C826lst4D
R2e/dEsW3RcpE6qMVxDvVxa3F1mmUAZqi6MbqgcqqJBfcERESeXE3wOGvTlvtdxJc0EcjmlmOzWK
5c5koXssEe7prSahZg6e4cepyZBSvwIworEQTJtIeru83+uKQyPOPUTQniZvsChDeUpI9ooAx79D
qLSEVI7wVox26SM3XCK96QOpU1YhTRD91cJI4fLduqw78iIHj+YiDFZKYSBl7+x5GDlajlFbyXLB
VVv61LPC+XK/dUQ0x/ROKm4aLnd3x4y5H9+dKF8EvXfqaZh1zmeL/GAwlJ5JaoDFQ7KgNhj+LeXw
elaGOz7nEKnxioTie287L+SDV1G6ZKWbKU9uC01NPEG34tbCFXH5qPAyblINPK9b5VAjO8auEeL/
xFK+855d1bpyBEKAJs/A2XSq5+0gFpzIXER7ImV2Eot5v+/lsGMFRzZciNsd1J6jmaId7AY2rho1
ieMbK/In5IYjAX4hRPMcajeqwhof/XvsEzBG9Wx0P5ZNq5UbWP9uG3Gvd1/sbJstfjMx+BjAjTxb
8JRP4JtfD1xNgmtjAGuW2dmBSAuT9XXbphGnLdOC6Sb7axV9EjgODW/TTGOMW8o8Mh2Ps5W9MqQf
Iah5vjaz55krX8H/XhqbeDj5NAs7ISN1XuoZ3NBM1BBrvtmPlueVlV46RY0DAkQubzGKHsoGmXXM
zHWOQNJKloxh16lLilqyJUdURRsK67vuvb+CoTGVnG0Iq/qE5Msb8/II086j5EDPjiw++Vb8hGdT
rCbyRIOAPfclfXpwJYzWOvBjpbfA1AKGLX7q/tjl4CcueFl/FEEUDcjqP59jwC491rvm1PYHxKrx
RTB9G1+sZyGSwhpbjQSdmCHoZbvW0iNj+gIAgrgmHKcW4ns2/SsHqK/p/LQqS9ZJXnhqQUm46BKv
DjOY0mXt0d4Mti4JzDUZCH1qEJUzOO8shNORHqzXQlIDuiU/L/IDm9utHlh0GqUAOta0j04m3Xah
UrEA7v63AHDU+PlfvAGBKtF3EL/vUkHxEQJhrwfaKHKTo4HVImnguOWnX12I1/AgRhsAB4jG74MF
5s1gYX8EaqXJga1wFpEwXdMisyuOchUoJErUidCh/N2Biwp1vpUCFP8+MwXte3IKo3j6OVEaYpzW
d7Qkr6kIsZNMMCWq/zt5/67KkB09pNvvzakwIxm9ZddAs70beeqhEvouaOvn1N8NDIFnjYiXFc2w
SGwxe4nZUj6/apOzCcvofEwe2R6BN/St6XLxuOo/rllBrsg2x4iY4Lh8EgUU9OKUmC5fkZ1Jqw7E
k4Wkt11mlNGoXG5QXKrNYJbg3AZ0VxYvytsM71Nn+G8nvOkX4+YCXcq8XwAWS2h1LXGOBdtmjuL7
sJmQ9le3NuPksciePd95fZIKiw6UqTCbeNT0HjpQznedQfgUpYkQaz6m/TOkVc50WZWDkKmQ6EZo
gmZYyBg+J4WhTBeyiGsQbTdPc0d+qXcctDOqEKdyD/1lS1vNTw0sljosGuT3q6Wu06UFXmW6To4g
YOlgcDBtxGGcW5CMO+ARVJtTMT49bfO3xPoRmfgHIvrdEJE/JNIa5B6m5Rl/lO3LMf7DEPccwqik
o8idpgsAvJgi1RotJxbQw/aHAU7RjefqNXVjKZDf8yt5ei8g5YiPk/lY3SV/5XZAxtlaLcVI+wmv
WrisWM2jrZTs1t2uMUm6vcnJco3qt8pb8lcdCZXCS1+tIyFTuufxiboT6K9Ygpz+ODReAru/rcf0
ewUJ92CfcpflIufNgBb30+/R9chhdQDzjfdezBok8mnjEyO7VIy0OGIa7Ofv3uyF18OGGVaM7upt
g7S+n7L73tsPed0I9tXn6RSJemgmZ7c+/dhmqD286HyOK6fau/zt9RZDsmnun6ER429OQkJGLKRW
LZ5yTYxx0ifuAjc0EiwvnGv5wado60F1hkhpgEldd8LRlWI4g6iCu0RomfkusSwyJ4y8JkJJbOH/
XrpL7fobK2seZH/E2M6t/TCPM4z0xMFsY+VszPjjCwgeMW0SMltUD0VbSZczt37y+WEQuDM6SDIa
1c4XWa/EDXd8QNE+gdtp+tkyoHgjpbsK9/9q3MiVxukOvGscNjA2xfXfhh4d5Ny3V522MXfdVmzp
eWl5mNqrGg3lY9Y1FtGI7EV6en6UQb3wl5sQgZSX3+paY+9jBMFx6Ec1gSGk/kOJcWmT6QMehBvR
7PjDHRzFwaXM/nt6vrSkAQYd43iGvcEDy6ZN0doXjO+NlFOrvZ6IU2WREeb2mwPN8GaF94gvEvps
AB0wMr1e2uEhDZQUnsHMJbSQpEYF0flOYl1vtLXRmMH9bcC335FSuaYpatV1MmIUU8B9Zq8seEJ/
514TwVEKLA21SUHloj4c6tgDVQSOFSi/bWgJkwLEF6q8Ut2ZwKebNGIH6wu7wzn3SYJKjHcWoud0
QNvLijtbH84VA6rV+01JWwf/SXP16ZrYW30Ff65OJJUGEh8VLMFvNP66fWGOIKXrtvG9/C9k4496
+O4R7qwI0zMOrcc3pw3UyGkeWe+smV1SmmKfJ9Ba+aAqWM3pIIU8NHfBqTLXq1w2c6eoXhW7mfIZ
NobxPK9oCHCCT5Gg2DVSHCiXWNAbc3gQo5JohHyxDcYZQm6gk9fEiO53LJC/RInulEfTEUYk7NXz
cvIJlyRMGstboIQ7cUfva33+DWQ5lqNcbMFjFJ424DNnSgQeOmZHK8x+lBoPZqgjRbNZb/oxdfTp
mVhuRri1RXXEFXX9b+8RRCXr/aMbPd0Ay9oN8STrjMTaUl0nYUC2cWsuu1aV08VpKUq0jnXyfGMv
ECnMuC12MJKfEkPKEAR1gmoBZx3H9W3RI6V6lSV8WF7+qieiK5ro7hsVEHpJkc4AMs5e5IpAbClx
22dg9GZBc4F6xuxw47JLpCs2LWsPs+tTLGTBc2W8/n8PkIbBIS0Uxok3aS8Jl3yW5TeHx03KelmX
o08kMLjxGKxUhr34FHjeAMbgEqMGJzoGGjNRuaeR5/WQFLlr1AkZHlvPGzfy/A9i21Rrvfhn6yql
d8WP66WY2x9BT7D6KHEvcdQNxCx161ovWjlHkXkuxYtQv/85AnPumXJj4o6KvNdCzFJVE01YzFqP
hxYv7GwdG/2szncZAV/Bh/Xs7pE9l+Dd3FgMCrPxh6kPZBmAZkF91s5ApqdrT1ETtuYBLrsEBhFx
U97GTed4CHOo7eSi4Z8b5t80LYO7XI6Af+9+fI4FfqLQ05ZRtxpz+DN/5Lfl6KnldDyBLwV/HUOk
o+qMx5Xj1XeTZvSNhE+QQNvLcVM+tj1jxGlqgTIYaA8ZDQw4CTGgP8N6qFqFttcPvZhjgpI+VNMJ
/lDhkB8Q7lOHKhrhQpJizVzIGq3tj6uQxBxOb07E0vbcLDWwsf+WC8oOnqDVkhueh0Mxc1eYZtMP
usxIBjDd2UTT3A8uOc6eVUnaFsQltF10A/TVmwatMDA+gOjs2vWCPlPJAkgC09WO4OA4I3hX4Y6e
s2d5iy49qX+6HvuvMQBq4AmjiGSJ8pHXIxG4q/ZZNunn8NeDKO29gyxSL5oVTR+QX0aobGRutG7R
0iSIk9Q3VxncCxqL6ODq25Wj1mjPXivcJZ4Lcme6jJy3oJsRkm552k/w6W0AgluJB74QG15kExz7
wGFbQYAkDIqqE71n4N6qNdFGjLzpBs4soPzyL4T8o7ULjsllqv0x9YNfoNd2CUASECGFuYWAE0np
27e4xyuQVf2y6ElflEJ4Zpj8P01vomOqJYz3ovBFmAiRJJEHo8cmqR2xdtyIeYHorZ6uw5jHdVe4
L1BebfmWksCfc2rNS9grwsLqz7taTvZewMvsOCdxxkqH/SDgtrjOMjX9uSojTOS1YJYYl6qZLDqS
rn7kFmiMlFsF17V8Iy/8jIBOU0vccibV0Zr1bTEzj79TCq9vMPYGrZNiQhIe2xBRoRnARFItqIAf
Xvgx6Yb7dG3UVfyVEx312TSd2JMhKuGONRV2jenlJmLjzbbtoBvHsOmbugOwTU++6bGxgA60531w
a6Ry3qdBMCIR7f6vfCOMIw35Ws32IVA6xae/DoIyY5B4l9DGiYaHTmOZLEkA3bXPXHXvSIGVBRGl
kdccnGGwJepuQttW5JIi4t9xVT5x6UdAiVf1R8NSDyjpe9hU+xnyD8yvC5qHD44xhl56Hp5iwLiK
H4OO3KxUN21TuYJO/a573DyQj786Xb/0Q/9SpJBdxzJ/qL3vAVMw2E60B0tV6vzQah9qdIqtdexb
b1ReAnp5gsbJcRZ5FejjMKAx2f85ZDnx8GJvc/qotCFGgmcUZNe//t1SdIooSmECr5PaYWEXO1On
HAiCTiaJsxq8/6CElcPz0oV1izel/X1g8rX2Ha2or9uZX9z1fZSHvg7FKtYFs1MtKWjoCsjn/h3M
Tc/Ia2FBp6VkH/jQ5KKgr51VmnSdJjEruOTRHG1VLW4Pw5/G6TDzSwjKf68fy+qQXxG9iU4v/A8e
o8/QV7LJ3yPwHNO1P4A8AaISFCYFJi4BuwrCl6mXFf6opTwmBkyrtNdaedwLi7EOkVu5S+W0U+Rq
7L/+qNmWBRzWYEA7mWE4e+gNBrOiIfbQ+J6HNSePlepEA38UcNiMLRItwwoTSCF7Hh6RBNLhuyxL
Q4XrTNTK1VYlKdqAAiIiTR7U5Jy7WBKuaHqIGMJeY8TsSCBhW3ktcfwfnd/JEQLWWVsWKpIICVFP
ZFOH5EJjYHGrb6VPYgHMoOKKwB+7jbcyTm6psuJK6C/OnO/Yq9PNOnjD/iYjggSmhnxsmjwvyA8Q
7SxXv+zzOd8SkquOXN7/mYKimxBuHrP8asyZIwhnT+ss1ahri+1N7TijzBI3WlJFBH58mDkTG1gr
vuGwo37XozFK23BJW3yFEdmYsBJ+EbL0vwSN+/oyZ4GSB8QvwSRA6RQV9Fvhl15WixisED2rWnVe
RHauoWnvS9V8nKJKGLWGR06FRBtCcRX2rVsnh5Ud4a40ziAkQegKG7iSTPbofA3NACJU+FePHbk4
NaM1P2PtfNHuGFzoNxVAOKWtv4y8Q4z7PghKfKf7XUdbyUngtEo0lNxAh2bACXx2Rt3T8ojdI3HH
PAsDqaiKzB4SL018iCrWy5vuAG7KRY7qrnScjZKeCfMJyKsKpFoCSf82yTfZM8EO6VP1fYI0cQz1
4USF8ShithLOs8oZcfZISjo/oq/DJhDbFxBi2DVAOEf1+okaaflbIuZ/KpZv2FnxP7Kou+/6Di0b
OErgxOBeA3Gx6eemAcbCpkyT1BowDGc54lqhHK2ZRq9rtuQYO0UAcQqI8VYy/eVt0cmhy+TnIxHf
YEPit0qmRcqYAhZVjBegwei4QAgNsxiMsakri/ISlwbA7HOwxaeU/sLN9VJywYlA1mlPNXS8p+Gc
Er0AsvbHvNzgH+HVdg1B5FT8p2EO+XFuCEqVYtjluCanR92BPudCGpPFfLTXwlToB/JMv33/ttYt
s8Mw58rx4JZhtQupggz4XyPa5caF6zaQmD8aNVgmiBxcCoNBrDnoGJuBGswjSwf+Yli+jMZ4T0fb
F6MPmrZC9C2E7d5XBJjGkhGWDfT7mtEFWgx1wfLuYbN2sMRyhNf54qRB7uzN8lBieWSTRtdam6/Q
7hMbGk6TzQQp7d4evzpMDLNl7KG+nr/BxCvS0081AW74msLHh0wrzytV9WGre5YroadsJyUA4KSy
3ELqPlSJGqNyRT6qGY2i30XECoSBwAzBUplpMpqYEG1fQjfaT62RDFhu2ENlGM8emuVQX+IuNIP1
sh8rR4yjBqV+ZHXA7qncRJ4BGvGd6PUJLLP95SBBkVfd4bgWXgO3d+P9vFz9TV7W4hsQ42TfJ7LC
v+FdjfT8Eiu6o4quZ7a08ryGdnW08Qsr2NY+de9xdpBLg+/uCINnSS0gQly27y3TtnTzXcscVKPA
pEB+TsnYKoYNPxIdH5hDQPsfl2uP6mRtA93nT2BtZ1CW830tzVuwkfDNX6ZTeWoOX/1l9A+AkudR
ha6Xu16b1X1Fx3Hoz7IO8aeHuk9JX7oHTM5zTXCq3SIz5YvJ7Hmp5AyOlgmk1R2q04vbNPUINSCw
eH+KyxfCblFyiaKtCbgHno5lsBUH/aUmYpn6xTiWQqFPmy3Q5jn8xTCIlFRDHX/Bn9GOEKm4o4Ii
skB8I8OSc9JJb1D+jGmTpNX2I9U5zeKjrI6BngF1PCHIkOBeaVAYcOK/Wm2PcBmQWUeCNRPPSbY0
ctENMklrEpiqff+M3W77igBAqvYzb5lyFq4d+86tuuLU40PAf/AIfRUWjIPk0J7sj44hvwEziS9c
BoaYM/18H7CjbtLoYhf99mnydGNXh4Gy/y6Oc7bIbbwcjLs4hIjmqrsi/ZnMTBqeQpdQlsYrHmJW
KHYTmrMh+bOc4+l52yq8ZcuzzfCJHDW/9DQ8Pix4XoRDiNYlPVyNkW/sKlzUjVtmKGK1/J3cFiKg
A8x1ISrPPSd9N0y2eCejYGPIpMtMAPp6K4Dc6hJPg2BARjKV3RfnXeUPMFxf0sHMNwL1StvAIVK1
oxTlDn5NbvzDflEGaFHpkju5Q3/14dUwDDQErEOnSRJ7nXxsUaFLwjWAa0R/OBGZbKKVk7vCyecK
WJXKOdT/9Kf6ZJ++MBkfgs0fHIXRyPMi7cVsvwqt+ED+vJAqnP6ZqPXaVx3MW2P7j1E4m/78oPBT
tbFhQXF1XebiayFtfauZM3yCy44oX925F+uWzW4/BVv6X+cB7VM1ualEsKWPmb0YP6k4o5D5f1Wu
S/33uIzYKC+8XD8TZ+7h9vFsiZDLPOuEzfdNi8UpcFQQWKDFPVRlzct6cX0UfX1LXqUiP9oDj6ef
AMY/ptlao4kK3D8c51Nqkpe9orRQA0VKFoUSY4FF6MeIpl/jHWQMufWxJ/RdoeW5ZWKxZ8T1Shyt
yAj6eRBm1DUA3g6AEtKyHiA+y/4GHe4/lcZkwyGWz20mll4bri6oEhPBKb+RrIwpnpeQOnIG9+NC
pQQhuKP8vg9Tiqn8q2+7ha8dKNyOKLg4BIcxvaaoUXVfrSGR65ghZEL89UjvuEZipd+FJp6J9xDI
WT5oIShpKIIIcK35H4yUXv2DzsocQqlUegbCndMuHlIIKiK1Lziw4TKSia7E13bKkPHK82Y6E+aX
3YGV007rBIdHQhYzMqfM7q12P2QbDoNe9ye7qWO/On4gFGT++gXDeWOJ0GB8Acx8JF0wQ9LZMTdG
6RaoxrBW9OS61zDTa//sKedqLNhLSCPu6dEbMctK2In09jzyeSh7zzPprhuHDIdwjPdc+D7h4RsG
buu6RjdBadYrr7jrTJrichrkZSsXggiM5vW5ZK94hM3yQXTdPBztP+nVFe1drdgqc7Y6jkfbLEF7
GQDo9e8DO2mk3Aa/jrG6fL9DIChi3QD7dGNiMVScIsoVCtjLCdDq5W2opzwGIckF9z8tUOZFpBAe
+PNPrPHqqjdafKNdnz8htNXNE1LMrts+I+aeXT11gq2ovmmG39EfihnRD3t+858qIlH0Y8Ths62r
jtys/BDBXjtFnLJ++gSQ77QU29+lc5pBFY+kYHukkWFx/6K808QuO9XMRK979K2nx++rjKn/YVVm
HL86goe33KkK/r1PjlqX5o7IiPXnDobdzjGl5ll/MLYrIb0Mpis1ViEqqMLu5d0FyjCk7s9L8jEb
Sx4uJ/khFujpJZWUKi5n/REgE687HrNzQJmxEqSbfBnhr5LgwLfIZb4QSg0P9/O0LaarqyESwSQZ
QU20mBEm/HzABp0jLTuUgapGpDUGBax7mjkKbjf/LkzG9S+Ja+q+osx96WgbrF6h9OkPJzlcF9DN
UdSqxPA7EvwQf0rCmOsX7EUVKJF57vCg7dSJWHfLOmhkuPenKHQ8zF40h2AraGIB9IOpkP9InJjs
E/bZZwLX8wmoUIUcaTPhxPkpQDVgh5a43klPTUfo79AcVmXZU97XVgtV1AzWypbOQOHScjS339uV
U/HW06gRl3X5S0SOOM8BTCr7HJ3BO3hv392pBHNa1IRTVhTnzOLqwkLBnAcECGk81bN3+v48qRHE
hY3G/JpbNqQWAYaIj3LgVuwf+RUlNupDRmXoWWP3ATmVZQt7QeIfvZL6YsetW7N6rNr4LmSsmg7e
fV1aZBnAlmk0MDlH4Q7gO9dcFS3NGoZZ3nVYVE/m5aPbQzdli2i7HWFVwfXxWH02lzDBs3cL5yml
vmsxV2Vv6lJb6uro6UT8JPB9yqW6lSfrwd30lYxqEqNEqPX9pQYMoqbmWAi+oknCaCOdsSCCdivO
vfGTrCpAvPxdTMNzQIRx07Wj/6zM0PT7PfUw6TyhCSwr+SQLWgcegq4/LoTHpHjIV/qhaDBhrjA8
k/XAxM/mn6XfJHhUHSMDiN1L/klXV95U3a1gt4eqGWdyPazxr5qwkGtEoS3yciFIdUOQgIz+nRbf
1kHWqAzn4R7ghE4sV91gUdK2OIJy1dxsUScQjX6NFW0owuplhiCMlsmOBxjW5taQ0206P/zdv82g
sIr5pdJsiZKOWIZQzReV7kWAXhqIL92LB2YMJTs0oqap/MymiQ0Wme69hczB4t+CyDg6TRpDqkho
03XF4erGjUBv8NxkMIJZgVdKjgVU0A4Kgq/AXGU0bCDP6w68P0IPcf6wEcTE8aOtE3gmJMtgVCQA
XH8FYQIB5ANt1gb43cORH22Y04cN7tOyARnQO0PkJvDNtUCyyEfPlcLTu5hK2qGEdFX8AXoHEBCj
1tCt9dsxYyd3VLHveK8ndQoVe9ZVvteH6n+5d+KbI6Q51UWNg8tCBn1+7x0GKkjvaL8PfjSt++HU
lNBveHoS9nw31xJNxlsUmXu4cg9rSXw8h6hxB4so5T/kwDbZM+LhNkH0s7cdSIeAEidoD6DGFMlD
W77b3dheEtoJ6AdXaybg4UMMpS6b9yzkB4UHUV1N8irnkVlCCPVqcS6u4b0ZxEA0BPyMbZuyuMNP
c/+ndzoCfK2TaEtR+fw9CTUHliTo0kyPSM3UBL3QJDE8j2tdcrHs6z8pgKeE3FLwdw7zRqlnr87R
ZWim6uWe6eXI7upI8iJ/kdx8OFPsX5oyv4EWxcmdJJAMd/Lk0AW4YV5mM22UDGPNodrr+2UF1coa
WNP5LHmF+Eu0OGwKr2NbBHZpgxqhIyCocMbUjvdFxJb8B1nvnrh/Z2nNRFxunwROWVdQReYPso3Q
eOffDUgrDqCDg7IIwbqkoRzSOLOOm1f2H5jbtb8cRvEXM6ibJldaLNeWGNwxhGxz01kp61k6uAi1
azgqkVE5IKEQ6hmnHnuD5DblRqvetjhzvaL5Bkj88S3M7dJOy+8gJIukqqHGPcV3rVuOUfKC6B0x
LjEBaHJB3nDfNEtOi6BYTVmHumpFCGchAJvTDbVFL8IebM3bMYgL0KCPpoUG1n56x733aOp+IH33
WQw/NV6Uj9WzUCL8AfDQied28Wmsxlo6czBEMcgDurDhrnzrb3W29Ai8KHbWG/uk2tEGomoVkJwG
sZAlFcdfY3p4VeI28k+79yOGicJBJbavEVb8CyjboDi4O8jwbNAu+ZB2iJ9WK03PG/AuBMGI70Uy
XknzmrOUFu4XSguOoNsSyXigQ+KXDvrlCsQKwbGD7E79O8Uy3fZDTkc8bNBOeLbIGo/5jVNA6tD4
F4vLR+gTLIDXY/BPPPVjFh/UsW03dAoBPey3NV3IBpg06Cp3wWn+p5lCG8JaW3EiTJ01fIWB9BSf
mZJmZKrSzisBWSS3Rm/HPNemu4bLCTSG/Ou/FKd/EsfMEeR18G+0h9SCP2CJm66Ygbw2LAXE9jUS
xDdmeWBVxLdSHC6O3oz074Tf9+t5EmxrkHxuWr/P1b28TaSlj8a4fUtnNeEfMWDksla9jV6syIA8
rpv3hZM5Hf4ApH+M7JMNLGjAA7e0yddG7CEoi/2SYtkaBkoifphZrCmt8y0S2nqss+DHd9uxUgVR
kEyNkcmmtO7wIqLjPAZ4Aw5FlzQ1Ya5dc6l3zcYlfANgoyzhrOt3CF12HlE+XlwPNy0JWyKdUeF1
I4vILI1gm9a7Utbsluj2IbI3biq9PeRcBL/E8Ree/hspa4/yAptno/0mbItEcuWr6LJoXwo2HM/7
nW22T/ZtlIlyoR0JtybaHNwt14eMnhigfVLxtRgtGM4f+XKg/JWtT4RXw7PxQkfIupai3Oth9jbq
+u6jNagwVJQ6wjBzFLHcLu4Sq8RPUWmA6N065GLGy46SamP8ByO8DT2QSD886sp3UmuoX+fGZKnb
+gpS87N0RrQ3IPtq6j2jrjVcC78T2KqOFkoFkA5UnkM0ysiTI7LB0fQFObIgsX1AbEYoQM4rluxp
o/AJRa6tGcrMYIPAyrvul8NlsUBRwHVyVgA2pznbqP+OtPEGsXsk15wtrP2TB0U0hK87GC0n2ddW
7ne4PPitOBeRp/qYyCgP8uClhRv99e0y022w+kBW2qtjBG7bkVs5eB3v6nDQk9TWspFvbH2pObB6
uVifgKN2/e43xwmZ7yDUkibUEcnN99r0OUD2iTLa40M3/GWrqzrt+FMPQA8JyINuOp7Jr7In1EPx
80aDX9Ps+jItKP9fK799hHWkcEzBZ/T499s/74l69sxXH0DMS3IaV8W3T7w9xoGe5TUN8xDkwaD/
VkvCThMBvsB6UPuKTRiofFlyNR8OXNS86QDzSjAmFG6gzwTnS3Gu6LV2iWo6xK9psHWJ4DQPDjq/
Ed+OQASdVxSAobH4Hg71wmGXs4bjfLeSJGERwx9GFewzPLnsCn8AgD79rloQZ6mOuzCEdfu8qGvd
8uyB+3+N6Y89GwT/PfzP7QFstsl6PpVbFlwN84CMT6XXb74sUjTdH9gPBhcoHv2GV0mOzVfvX+4j
JO63qrd3bsyZbZ9FIEDRNuHnEdU03Q6Wh4ZOZ7cImX58lIvrXg/e5hL28K0Wtm9IbCsHO9LNUqnC
TbADpYUzJ9zIW3yFdWvxrQ5gTg0Gnu8cJ64M9e8Z3Ww6Bd+btN9bzkgZDdq6MWOXjIWXtv+SSPcP
IQop6CqLQMgl2U8yBymodSJD4VH+F+ilvSQ6VD5W79i8bsL4ie4j8X35sBmWqLh+UXaBFGzBuuwv
AYi0w8XtovW3296zokweY2fVzkL3NKkHLWaKuK8rI2HeCqozKaGsQ8h9rwXJ9zntTQxuhW1RsiE4
fnxMokFISkUmCzMiQ6pXd7IJHZYIbufdmUfs++37QpVh7mXccAXwYBZ0+5aKbrhRGlLUTr7ksNRl
QwoQPlYKTeMdTSMhnHNWo+ekuDcUm0Yofcpi3/1paoJWegmjCAscPR+54yhpDMzZnKwl1625h2a0
vF2Xtfs5EZMdOryZNY/cDfeZs9FQ/f8qUWOa1FqolOWHUdSTDroFDNrLcybQ1men90VIp8E8uleI
WGy0cJqyJNFdWgnp5FQoR3Dzv+v6HgpYDzNGb1bhc28JtUhpllk+ELUwR69F+Ol5596kqpS+yco+
k72aH8jFxgXvgCM7Dnsy0YAgXpW8ZXLrayIYOQx+r0sE2Vw+SXaIb3wOblOCSgzz/03iXXq8yVtD
kc6oG4qrP+TMGVmoAG/awTLPw07vISbjXY+dsTSdS2B7xBoyP7h4MYVJGBTuTE3hXKJPMauatp08
3wdibwrYdL6iYavIMAY0XOs96v1uE1FwABA901f1gS5qbmPdVecdC3AEXE8e/4e/thgqhRUtHCoN
8i77DVXpZTbrV7MId8W9jde0dbSkrK2BjvPIN9AX8dmi78rPApi4+SLgYNfxYRvdI6rkf0bxA5TY
yFcLTBQ6MYbZrTfcrJ0x6aVp2FJEhwErIFwdC2PSvcDiz6ATcsDyZwiLp7sSMH5DSy7afLmRhL/N
V1V3rE1sc1P1hJpinc8K0qvRATrXLkyWt5QO+kL/sp8Yg9RO9S15rOqRR6VYqkf6xQxTbhIA4S4X
Y0PYuVHFGLicar+98bpP53F//rY/ChaG3t381BWb1VfIFxYjnYbWtWIRR/9fsMIvFZDKGenItW5H
9u7YXWiYYxs3Wxv+lCplgLY8+dVWCpzsYQTnq4GhzHccysbDFDqVjuB3pHjAG6qw793s8Iij/ODW
WlxcYE+Oub2v+UQFjEt55FEHd7McI2cOJzjnfRbUhp2TTtOX7Yux3gbjSp/XAYwuqY/uGEIqW0CA
js1KYp0hNPrODFethjxhL203IjVAzRzxOQbcOCK/rMmR3omTU80Z5Opgy0+d8alojTPewBbzgyOd
CBu6LLriwxLcmSsxq8ANS96PyIGHOwAVIk0atPtB4kqhRKsg57DxmP6GcgDa1XBsNyBBWsERUcZN
ROyFe1NcMGzGaklRu+syCxMTCsIa2yTsDjueE9eOb89HpQOGyzAS+F2x7ed5eD3aSGlOqXkKGiNA
Z0dXswQeRphs9g4hkSSdgknkb1/psVOeT6QzGHx6UHk4q7CQUCDd7lx4h1sqyTIFK01BYrk31lct
8aNIUy5CMtPv6g2JDk/0BWaUY4KcEOEq6JMO1TO3DC1UQ94IdvJdCMFq61VWDlWKGeYLs47c557C
jWfTy5f2WC9c7lOhzxmPskbVtVlrVA9aQ1Qi/XJtbbLws9oj3mYU1u0K4vx4WAU6AwY2nGtlf436
OO3ZJwdlhiST+Ajm29zpcizAR3B/YO3cXhIGQ/tpD9oaQWW+6kARMQxLuk7k+8dzH038yh8XluZd
z73cPrLum2TSag1lt5e32lnpWMP3h8Fr6i5X9O7UidS64jJkfkfhz92v+AOGVJ/eqLpE0J4RD0Re
ffHVuX9oy+hRuBndI0iD36vN/lu1K21bp0JCYhknGrIFcMpBv9iQhbo7bRAAQSMAUvqFNuiT0V78
E1jgP/sCm7NoZ/8Ms1++ANrk4vJeuBDjBkMbSVw1nI1xvUxHY9s3b3xQC8Vs705CKvB166Wk0rWM
O5RW+YihbtgOFQbngJ0osaik2yYrlEtJQtYbZcVWj0BOj0tL8hcIEXbpixDDdz4EA6doV5Dykw4t
rp/eh6tq5NEsxq+kdc9vSABNwsSPeQTN/UysEe9kt8jQfwAkLTu2SiBiayqbu3AQRtUSYSsWEtec
jB0b8HV3Mw4PEi0y3oyCVDHexmbDaTPTLM6im9JxNn+5iWVWWdRSX/9EIAwNrmGbIsXw4XYrAvNT
9PIpMuFSir3V6UFZaE/Lk/wgrBvKBDR6tN5sJz1X9W+U3Je1yKJ50U/5JfDC1d8+NMVqpcqSqjhw
a652l1qVA97/S5raV2MU3DGdAND7FtsSIbMy3vwsZDM7xBN/ARgDp3uwM5IAyPHtekv56ONglCg+
ZqIxS+8RxIg3kKzlvsKO7leFE5/ZS85wsXWNySOaYUMdsps0yKvsq4ZvcmDfcr3uXYE/cf9SmTO/
nyJ23HjLF9MM675vUw7uwN3/Vm43fdDfKjjM4MHH9tn8tGQdrpc/yqcrBl9Ac3IFobvWQN8Dud7I
8xi/KvlQ1RFtPcBRShwtfr/4uCvx94rDcsQAEjA2Q/3VfR8HxfCu2vnHBKx8OBe4mTSZHduiRmvz
QA4fNDhu/Uwz7P3VHJ3atJNn2f51DKzRm11skARfMeQEYHZK4pM1mowzkAq5Ozpqff9QtxXuTQTe
A4hkIfr7tu1DnnT4hkeMbanbnh97PpE1oKwKFuZESvYmspk5F6sgDf2MnLhnXYgzy73QPAImT/8t
NQAG9shMwrYtHZrA0rnfVXaT8pJfF24TLDfgxYkW7Ck+PzUrmhc8w3ewp4bVBjzZCjgec/BbQJra
jOtCH5zghMEqfSV6t9tEp93/+pkHPTiwH6luef+YeR6vBS1cFm2t2vr+6SrAfOYLBlpQ6nPpcTBy
VCgu58yRdduADz79tlZMAHkF6hDo6lrT80CEKOib9VEjldOCPwHH9hqDjfeTN7ARRVPVK5D7cwNu
uFx5YCKr+R7OMxcu4j9xq7539lt11y444tQw9BzdaZ5iptIWFymtV1QInW7qc0mbCe7tEmXH80gN
7p0Vt1kRmGL6t4jYDHTkzAo8AirRT/dsKt3W0/Xq3qYC9/kjtCvLXX5DO1O4KyybQ5QvENYu4vIL
IKhqfXoHYmrzlo7c+Qgf9aWsownlt+LuPUxlMDiJoLsB2HpstEzBeGvDXLIhdyDQd97wEqmc9il9
rO7ClzlTOGWrT7y9UIHfDMwi5/xV2z5ADGS2qEDytQltWWf2oLOrjRwYbgrpN0A45xgOSb0M1/c6
gmZWxN/auoaTirhnLPXEHw11uAIgiswTwqXIhPYuXjRy3kSkRpUhB7TIgDF9nneNpalBbmj5L5rB
IjiIEV6kj0JZM6adksRUkDJzFhSVM9gexL6GvlZtJPgvWe0FAB2AoDj8bUfrM4Fieu64dkrUw2yM
n6cKjg9TlsTVur00pgpzVA8deMdH4ROb6Wv01RsOT3NY3POZWnzVQ6VwVqV2zLgQ2oIxDU8z4hks
mtW4bjS5ztVUgtJhn2tk+D1vJSIfkqxnmJrATTl/pgnqdVn7TLihN95yErd1jNntDc+1vl6Qu9WB
x26IkO0r2p1Nn7cH5Grezlk+rvNE2pOXzQ2XIPMS+Lk2BoVO2RCV4EbHVwsK9Rxj0crzL2dXa5XO
Fy8kCaAcwUMZYH8nksOq7JfKovMXZcpn97L8Vec+r23PptHl7ZVGLlKDBggKZ1LWePjxiuqYB6I9
It97eDYT0CcRSBlzWgwmCwkpTaoF8YCLwvo4ARc5CeeW1eWal7uq7kSz35ZGwtpPr9eIEE6iA85G
LMW/anN+dtlfWZlopEzRll8LjoK23BZfs5B0V4uuNDw8Z7JJS9OsatWws/h+pdhmj80fTzfBZxlX
oiyNk80CKKV4iPudSo3umpKEPs4k6svw7142t0VGfH502rguqCdnsCoXP/qLLYIDMXZX/FOJ7Dbk
V6WPlWXbOGfX45Ge9gV3d9A8AmavzCSLw+gomNrdCWVytxOPKxgYEEjWJoxb7QpZSexwRebGhyK3
5Hw/hfCqUGhWlDBGqop0tU43XoFnfH5j8I+2lQ2lpzHamm+P7ps9zU/4H/XZCfCCTJjS0xW0V9YQ
0rLS2ZFip3XQQp0drhUDhW+59SsG9kKgoFrTlybMltEbV6RKKp17PY0TQBx8wXaQuD2/A/GKtoDt
axNe0MoPxh+rViGASgjVKnOkJw1W0aYCaAPUa6ZMFub/r/q1A9P/LMO3ttkt/zRuKGhB94HMFYZ0
0VNe4dHvLC6CMg6WBYEe33Bhe5auMlLGgRX+Co91EL4uDkmOHxyUhtz0oEHCkYO36thbMBUF9uMg
tNPUGwRBvFqMh9R4VIg6ekaVRgFo7+FZB6yJyj31rqLqB11MknPcYqJhHDIYJdowaxNq9uV6Q1Lf
cUYtlOJjR7ZOuWI9Q7ob6Qk6RU3xwN+W0gBcP2hDEbEno7i7+ScpjQeyfY3zzQHPB6hyqBbxQSxe
0p+bazSBjhHhzDQf4NvAXdRwtNWdFCVIM1dgt/QuGa8pXf+P0zemfgZPaYexiOmXMeMjQmayAfNt
2v4hhAeUDo98OcS3Z82Etb5UIkqVbpR5Do/B34LEja86oC9sS4WNAKMMlV0Vl80qZYn2rmg5/Rs1
u7kajizwWBdIf1uoZrAT0DxV9vKgHUHh1GH3ZjtvV7riUXjlwQs0hHnJnCfD2dGXx/gadOQFAjmE
Wq0b+P1Opd6lrGShmFk2JL5yGoIe/yXXsxT8vCJ9zX8KvD+N4EoZzp0qNnXvHvTi/eAniGoN+5gU
s8htqmRhrqot89NLE+qvAROkdSbV9W6+k26Sl2HRtRyz5s+ImeTCS8F6yzarZxIaoKM7kKd3QzP3
cF0NcOoJ89o7cwMTzYYWD+gHUFADk4SAK0RSdupUa205rARelfr5VXv6J1Cw5yZcJfQUK/YLM2S+
9ClWn4xmps04kzumGZdpxDN042V7XK69pdXf2jnidviQbPDH1r7M0tRmdyt4RFoxbTPNKl0fAWih
Wk50N2V4rO580DfEO356DhlybNae7E4CvozZ5wv4dy/unvQxgcKy8v3xG98jRL+CXxbsq2aEuMqZ
hBsdUK8GzC+pDyiANkjPA2MVcc8ZbGu43jTJtFLDT2+9m0tD78B4gZJ/6qt0SFohMPO89or9ZJg2
SwuwZUkOPPHYBLpw+dLGWlFMvGObCP/SuqLkCvU4yFC2HBJAfNjINr8qdKMmCZ1LNfGtChehwoGY
yQnHl0Uxf9gi+eznmhByLJyjY/wcfC6r9R6mOL7FHizChKZo3h4CWpu4nLjUpyLYoEAxZ2SaLVLO
YhSnwHrYvP+l4zkHA7tSO+m1jaeOvSkbXl4k8hIv1i3Kb3OhfnMNetMMaVB8XOiwh3Z1Z4QJGd4/
5yF8cr6m8/M9Z5vNu4hgYCEnN7jod2iP1+og5bGLJDxybyA5h6lNDxecrdgo6CAvPodAxUcS+076
5Y04K0BXN/ndGd9cQny8kEvoZsbAeslKQPiP50PQ5nkiH3BnKmFJ94vwqdYWTCQw8m12Zn3+EGBx
REPhOj04mVeOHQeccjJLSE9ZN64A2CYh9qpKHKUg0CVUt8xvm1yoTFs40AV+Q3K/NI41qloAmzUD
pKGFc5+PUk+UJ/FSgy8Zc6lmyCZ8oKpfb2iCAqDelwmADqky15puLDfblPuxOMpF7M6tWQaUINvE
CLaULUdYSvWE/rKq/xueqNFkN6ab2m69oNe32K+QHOB2/gRW+GXL72pmN6ZxMH3eVYwAI3V3or9I
YjKA6cvnwY7wRXoBDIBvLlsKtAWSmoy6MbG7sHl/4gFcQGmfQVmvRt7aS164VAkj11SHmSTJIQq5
98fsLybj/86o4ugGB4L4HWrSNS5M4VDEQq0yCrZZ1sgGmBi+KZP+K9YXCjuVghejsb3sMijzXXGc
+5JSo4iYwfiTo4gl4MvJ5YNBfiwqX+C45AWNxT1cWwM0VjfrskJ/8xOCCWNGiBN4XGh/TJO5acj4
TFzuaCY6ySYng1vLBHFRfrECugrxLzfYs4A3yzKKm6up+xRLWu+tq+Qq7gbTgQbpCKLSq3W0CS2p
jNyBKeht2WYZ1x1umSugpiyiRZnRcyi1IGGgRMCqvFOxVmVL7sjb9lWgsIhRXefsXUt3wAq1CYbD
JOGMLd14RvuEvESih2XZYHec5/8wA+WzGLEXmF001TxCopjnFQDO2geqRTuwc5WL66X5gBeEAozE
na0gCEWvlaLeAJ0dfYBx44WiupVhcrvmdRWUorjzIn/z4E7fOui1vaNut4OtAQJXncmpXHYBQliV
0LJPj6jvsJqmtzqqX4bdKH/kM+cysKsSuCNmcHQ0gWzaUIvtrfcWorWDxpTWil5hFvUO4q5O3bB9
3+Pa1i0W2tPftv+SVG/3zqcNbncY5bvi7YokIUWe/33eH1ITghfcVCfPsJF4NKcDnSwQMZpAjcur
RJrfEWxToBkOI6YxdIc5fYA1uz7aZe2qoon0WfqOQ/UwBMCbifH0KhVerb1WiQ8ZPWDxgFRU7NgU
o9OEOOWYn5cJAIrNoez17PDvyRSl40xKhrD3bY98sPHE8j5MC/caaspORSDLVRwUEtEiroBCunos
tjkX5lW2fgO2LQWMSVMSsVMjN2sHWBFQUunW8qnVuClKkiLMv58G/JpiyDpAy1Vq4h8jrxc4hrn4
dI9XEfxTEmTpB+ycXBveysPuRq6m5jmzS6hgGKeaaIhtI40IS0fShg6/9BS62xxvrnk9MdLN/sw5
NdwdKu7lUJivWiEDgOUv4nwT1RB+Xnr9nkOG6vxnFsB9aFM5nUd/U00X11O7jkYCfOIlhWzkT1sB
rnq4m5P05AlwI+pjnVB7Uho//NgwRshSPV/dT12KMi+v2NjIB/R5TV+ZYfa9xxDNMrGsuv0VPi8t
oGlB8Jnz8zCqOyq3sRCZd+STIrwnSOHptkeFb+QCQOrrG0Bm2LCeniMDIBX4byWCEg7gL/+rS+th
qmopp5lZd0Gg+XgezKRPEkvX85r9wQiY9o5MIvpslQtBYofQ4v//tMen0Tvtx++wyepGQR0MQ8Gc
6dernS5BWYptKurAO+px6APaJ9eNHXQzlP3RMcXCJwaQzo+vKcSasDUuK8+/2XNWKB/wp2pwffQq
+iCW3JqLs21mc9QEoOije2Ti5N9rhV/ZUqrxGC+YaAB0k8V4VBTnvvEZDmtR8rFY9miC3QnPD+wG
7KjkaMVsee2CuGEFn7NX4oVZTmj9ekVhhpg6dJPj4YGDZIDZ+npwJZkJcjY8nPYY/udNHSluBB4E
FVMYgzOwDJKYiRolKmnAcfSPimQvo1iZKT5rXXCcjnXa3f5uVpMlyKkz0Gv8tcvkHOTghSXi/a9N
FG3ZcM/FpAGdSoFJ2cEmtp/kNMudqCFi7Wt5vQ9z9pY+IvzZZzof8m2w0kI2wX+lJmPGkN6o0zfG
BfOClpVu/LDCNA2KWnIjuWQLXa5V2AAJFUKPLLJUCaCKYw7tCZWND0/723v5ZwyODgprtTjdh9UJ
CS36O5gST5ZJIeoY2eUDsljilVcvxZOZfoVBd+WAg/vnMh9wJ09niitX/EcN9SM1z7VM8norTmyz
0xd5C6FX3TT7I1Pt3y2qxdwCf8+/OQowQWeOFBy76IiKh9IXFeDbGuv+hl+OsWzEoFzA8ifGUubC
BHCFqIerYUM24Mo+EsDZQR41673Bi/fwWeEEKYRNEOua1jwcRmD9gXjPZzNQ77Q5T0ZF3V4/GD/P
JBEB390NuP+ZfXVLjvRfEoB7cxz80jMJKBMOChQvNcfYbxUrM6SP9644HlnbaHzibzZAFp9rWWcn
PkE9+dNWJiOKc3W4l0IjFfYGS53fJ6o+gSPV4Mti+CLHowV+Nk2Nwoq4m4/QMZLrl1WNItFZJqpJ
DlEySfApkshtQ4atTN0UGMTWqsxlTDvRcBn1ibyNIIz9jOjqpkLkiaijeZFwvq0Vzez4s1etWnH3
Jo8Yja7HsiO+YOzNi0nl0nvQpBZTYu8rLBNZELm5otUC4IEk+7pva9RcjJiYfYuWixpX0Qfawmz/
XcthH+lgyc7FkBXTCYCOwHUzUKDqmKI2oCgN1GU5ebPaVwmhZHz5gagF3T6ef/3F3eM1ckop8S05
JjkaIfo21C0lZ6g8f5LPKujdszYsm4YX9nO0YdDav7i/FDepivRaOB52f3yBLVsCruUCFxGH4TIA
AafufmRc6m++RNsci/IyTE2kD2qRcMuP4U/n9pUktLwtdYptfK0lzHSW9sxzP+XbAG3sovpmzr7Q
CnvUSTfwE9dtwVs2fuJrbm6fV+pjnrEiB0NfRmZGEGSUkf1eaqckJQ2vuSIQ4k4EBQQ++Z5Mg/2I
kBCD7YpVciCunUr7fvhlSrqZSmLzB3evNyCi9kDRiELnOeXLiZXtYowIkgEhv7PJ0lfmjwq1UtST
9zPGDPm0qycc/i9Rh7q5/XfhzbeTWr/YQxwwPDwUVDU8/cSi711xPmSw5o09BETGfcwYi0BWT9sh
k8Is8DmfhIhTzvJLXjES0kb3Rqcc4inE5n21fSeWwJmGiGVDPdBIc5yleOb3B9XEuixXNLewA2tO
5zWPdVdfA8tAIWL+6AGlGSybqVZEfbWkK8/buc6l14kYKl0ZmWgMSBXfdYAopQyo4EjRIum7el8B
fv1fytE7J328MZ+f4xcb71yjoEKJGkzI2xc0nvvV+J0PAAf/rYSxxBLI2IeS4idUiJfPuEo5xgq2
2VMPqK8VC0o+l5unFtEt0RY0jsmh7LBl20SLdsaQCb81dpPRFAZddjT+9E2IYuEX4IgXcWN0H8uH
qYtk7I46XwYE6x30IxJSE12GD2i5Mon75YRUBy5E1aCYtl6ExKTWcwZLengLIteFdpAmXihkPwrg
ItmtUlNebsTWAbqiBVEKm3BJTuk9p3re+wmdC0fp7aJVqFyhlQ5nzjLSPZwvfrjZJF60U04VCPGY
QN41uDyRFKGVrhz4vBzjKV+PwtUKBKGPNaG8HZjIet8ZBOuK4npoUJxYasMI02npj5yy7uU6WO60
uVvBKo/6FOnhNc56funVkOyV/B5W4saKZ4S0bsWKJNt56bORgLP19JjkHNZJlLYfGrI69kfGN/4W
wyhlLpHGRyZchJ+IIaEV/YCPycSblz73dlNELG1baOxB1Wxlide7Nvm3a1+IgaaV6f6+2fgsKpS1
aYKvgdDlmgUTe0cchdR8S5XP0gBrwoUBgZEpkHds5e9sS5vyozwyXehEziFoDVhrnzmaqRultomP
e8x8jSP4YB7mi098aTW5K37dYZXgzy5v7XshsmBZHd286b6F4diBqf28CmlZMGdPb7zPvTZVw0Y7
7M008O52ZWOWXLN6iasLOCeqJJHXwDHIEP0H/bk6EMikkLU4Koe9iLt0mMfyifELFPyE0euvqPEQ
xbdpxuy3KJzhNPigt0CaTEgSBKWhOUExOVtGLatUczDIWNrarSfBNKxqFkaxaWGRjRQQF1m+JFoH
UvjBLcqqWgznjTMk+xpbs7c61vSXd63mcDAafiW/Lr/hDCbcEM1wg0TT9KkvwqFmle0gQEnn4FJJ
c7mLRx3xolcMRN0I65YNE1qyAnDFGYF/bQcJCRIIntkMSCEqtxxdKrMdrGPvr0l/sSjO96gTidke
QrsCBHsUeKEaXEISsEtAu1amni8z42m7ECRAd5YefJiaN/zL+Ovklk1XDiCzkSWa91jlJYvN8kHb
CAmkW28MQwOK9y/1KRNSqCwcE2q8Jyi6T4tL1ibZ8NNooo8epO/VATfiucEpgd4r+QLoagq/0/AA
pOInx1t7wWTQ8CNjjIdspFqzJLsPObArTfSviUZliwaHvQCd5nTdJN0iNyWWd9hmtswTmCJgYHts
r7iadfeCsgH1MhZTrx3kIuYP03o8dsNcVCm3XNhNKpTsXQToar3brIY9VaZcufdQzOaDhwbrTgPV
d2MvpiDjz4wtTETP/4wtN8+PINRj3gz3EcmNu/qw8o55nRFvuqdT2btQhzRnRyEd20Wt03qv1ZzF
J5uE6pa9bXI3V+FwC/RjzqkpTct2R3Mf6p3XVhU3LCfsGVjoQYQUbAT6FfhVZ13JBXMrh/TucmM+
fdKJdB9qTaGZBmbdifVOtez+SB7Vj39dwzbur7CH0m9xffTdFYCVydBqpXq+oVWsTF+PnpxcQ8tV
hN+PaNTugtnPQSCl2B2Zabq5P3TsVsNoAUO1zB8bgGJx/B1y500fD5k32AT+hdgkn4yB6GeIPojL
KYj+rIXn+Av3nPKQgF4gk1fnJrUGeksZyw38PR6qwVfCiJkZi8FMSeA5Yd44vLms+soVCXQOmajH
eaYBXLfaUBis+F1/QSI4o1yvOSYNHPAhz6XiV2HvQYDSHR78HGzfNLOnzXHFIDgCTsXXJvzeXMyF
8Gm5LnwBy1pH3n9MXrnrF+gJGd2H0/iaT35EtxmeDNYxg/oQjBMMUiOjt7NlwDm8nCuIzAZdY03B
1gHf4fqHD6+J0hKYTbl54vSI0MFszsjNKn/3Z2W5Z9BZhVkEqDZN5TPOGX/2S1CYQyqtWLqzuaLR
PjYrdlufz1c3iD2DP1bK9t8Uz3+xsZ0ThiRW6F5ZZiUWZZWHX4IstwRp/lj5pcyoWoCs4lXhGCLo
O6NAlOuSiRFs8mK8i40o46Ec+i+OTGXKbYItHOJedE4fmFNyf/LjUdYEG0OYLP4xGxcDe7dMTpP3
KDnqa2vj6OGsv7LMH1jZWKeCPX60HiWJPc7tna3mGQKc1Xq/Oj2NUtGpiUPYIxOi4AyNJp2ff+XX
2pCSVcLvLfGPEXlE7yCJPdxXZQhzEw1zDBssXw2qS7qFJhpWj9zvnFdi3LkEbMS7q0EVV+DY7x+b
yEZj1N66z6v1geOzR5mdD6b6O8QJZdcbvvmx87mUpD/SeyGh2JHbLmnnjePBwJGyOOOw+yp3UKZa
IKgbMCokrQ02rP5UYogq/sSGcWeJpmNwtO4iU/HXf0j9JAVyoqEaMqQkBlWlG+aZgqmaduhz/7Cb
y42x8jJj3iOHs20fK90iB7QXoXCCA9EidqWQx80XStJ+1xgPgYxSIMv7BNDVYRIQM65j+9rG/gSc
K6t74ojJ+4oOxLFKuNY5tjiYW0+YoO4XMT8re8EksVaEkZyP32+kkXs2GAnlUsTEe2XfLvVRjyeA
wxhwBkFnebQXl7hBhK9DQsPUDgIllm3ZT9GzupaAUKYltQQ5dj56qbl/lQa7VJWGsFoWloK0GJ0j
d8trXn6hcGkWggt6CiJA1wCBvyyljMa2Q+T32vTdM+L0X0QhZrlsUW1NYoA4qPWSmFn+cYVPZbEW
HZ7+EZL2xRh+lhrTgq9K6WuhN7uphNhAgyJh+WQq0bC5gLnAKmv28XicInvS3cjnoaUvmEFjolTl
x5w1YVUDRvJeqA0/9tSlvFdcw5eVh1C5jgvKa4FC4WlXc81bu0iG1zkvchGeef00JJ8I5sNBxyX6
Nzfl7g4eaH1kK1sNemeaqsOo8rM82iIY9Qucft73+f6Zm+r2CpT0KNuz0PRWj74rq+gu/TcsaxLM
nOJWBDkbhhBuCw7WX5gTvutYY1xKmjdJS+6OFw7IJDwDdGTIMtxAbo1D4siM3uP1ry6lBJsr+jm4
6QRTyOsFCCj4v/ovoXAWuprm2hhtfjxX2tinpOwnFM2XDZDZdFCs0Jq41oynRshAHCJhrOV8GmqK
GziJS3fEzM6DPMNoRIP+bOXVHjkX2MQX6J5tMNX7vjItBqmpU1ELKmhwVX4wLwbhPVIeIQsChkI4
N9YV0pDCtDbTOxzAmw5sxYaYN2U0eX9Iw0inSly666VYvh9HN335Ghx2jU7UiIyGnQdxAOcMYslT
ncYBiDWsbXpnixF/PNos10aNm+GzAXcBy5MtuYFThAa7ZD19JM+Wrzzb5BdKdifpUrtn6St4blXI
Kk1L6IgKKMCXrsuUeiN0WPX7uSxCoz7coIlIjW+54DQJbn8Pl/NShraGCSSC+NvD5i/okPSoQrEV
+PsZT1RsBb46GPuNN0/glu58xZjgZ9YPZMnBnkJh84veT6cGqDkSaGtyAC9+7tUXMeysakerHn+4
tF4ATlYEaxzsje/bYs7LA4RYojvU/CV1l7Rvsapd278LFb8v/soHsmaLOx/d1642in6onm1rzmYN
HxPz1aRgnlrzOat/lAYpBmA1lQJnzZXs2xzz0ffwluxyx+h9Fmb/0UPUQpodYwHDBetH8b4EKRUD
DP0B2zNM1tflKS2t5gHaNG3Ieyv1QjGitwe6vkWsKThiQhTZvtPF70OgQTGOq2i4wJjGRjbzd/jZ
2TG6WtG3yLHdNk5SgorARPWdp5yR6DGfF1gwbsggs9jN3w6vU2pfpm+XeMO7ERK8PxxNk3SV1Htm
pUqvdN5LyJ7PQk5TH4eR5PnYSxCJX/Hp1xTLTpH5BxogdkwvFgr7dWWBuAPdDgMYSh4KrNd8xvIr
IRXfzkHSQZzQ2fciUeI6zf6iWUz1iqwSTv0rEmMgqF6cRyrDTlDBtWYiHp9SSgFwRWXCjcDZ/LaE
auBdFS7CebifK/zXWxAbMQLldXK2l7wkotd/1wHY/svz/x0WjUMRFO9bObeVEZdVmD7U5EyJ/4FT
8qvu95Hp9NzsHYef+Dbz0q52XB2tH0T9eS7HevnaLRwMkckjXcCB5D1LQY4dIKi0Ja1qUxpzSkbh
XT1avMk0jl8nAgsyKjXhW4mP4u4mjnvPjex+OVnBYSAmUJTeNrHmZBzjXmlhiyub0m7V2NWyMJu2
CwKgZ0srzJBi37q7A/qm9iD5lEQMYdQ048z0dq125GPmbSXgH9UdfQk6fD0SUbTuQLpn70VUYZlj
jY95xx7x7tdkQSDYVlEQcPB8xqz/fWLMsVqAmkE1i9bE/2Fs1F8yjdRFKM4eKYS/3q5JIdGdjrM3
3E4m8oz2fuI9x/C4xs3khgrBr1gzCCH0SIth9cgF17XmSQx5OeGxLFeBvAY/3fiGCwqgkpdMmlsI
ALpb1ZSeTaW8hdE5ol5YpIhOA8dslHdSmRFZNGhEYn82+GovfJW8DeoUvft0aE3ZebbmDrjA3lBK
ICkD8X5W/e067Jf4JMNWw32ubBTvJBWHZ3Y/dTD014F6ETPqlPkbmpf152RGhUHPOtUxUcWxrVQO
Pr2D/TP6hxzZtrofxn9o7XHbw1UtTrdDPkPbhWHRtIviW0wveygwaBJ6/ZF+8wdQo4sAfYlm4F2A
s4HYDfOk0Wo2agRsbC8xbcX6N32C9A0wRV4U8Eb5WkL4hOhCgdM8G8m72xp/yD+mN2CmGJceVuDJ
2EXnhFnJ+z2OnL/ZNzEk/3HKDHLWjQmuJEGdWrlEg62LfhESOsvqznttifHk9MDD2XOp+ws49TbG
1jfYkB1Se4VZ3w2k/gy52wJxwY1fdlSL/+oBS5y65vQUnrZiuynJxIq/ruXUzd5c/eInpAihIgHB
QSdAm7TIQK18p4VCso14mwSoUfwJqEWLLhsioJzATvI4+YpDJoLRDsLPAoo27CrXd6PRSxg42l+/
cSUNyBuNmJvUhpLfP6j8uBq1z56sX8WViXWVLOV7deQ3xeBFW+JxcPlE0wpG56/oxg6r5XTTc75q
PKVVoDqhybsWZ8l4vjDBCNeIncDI2TywVEhwGbL0fWDSoDwLWZVQCqJi/wSLAWelHFB21s4oy/po
IIY+RRFk/RRNhSz9TED2nVwbDbaLauusxRqVcw62xWcHDD4/6WVOExkv9zT5Ipq3UlgRsuDOTvhB
QqCCilUI0VQV3GR8R/erEMl7BvJQm4AxvKQbWmM4UtMkFkr3QV3xeVVa6ONMlkN+PUTpvprYr8Rx
Ko+8cpms0WjNSzDQ+OWjL0eNeglh0J2AmvX1fr+FQeYpuvpKJpVXMd4a0Mme+EjPsoFT33ANH77p
ewnHA9E0FuP4Mz8VghKsLvqyY1qQYOPJiowZzsZMH4lDbLFM5hu6Uq9HcuFbibuYB2D92oltLyif
wwGtEiojmkmeHVchixC3D+K1ojwsFMtd6wGuPSQpKLI0t2AAhyJbDEw0NDd1NV0uCqGXX0FcCrvF
O70NIauc3QS1f4IEaXTQOtqSOdxalrP0KyGHIe64wsWPn8iOBxbDpjc/7dEpJ2Mc4xcEKA5utYCg
BKluEuz4sCElxurgksAab5pQd9uAov08y7KYiTmFWiouGhVei3iqWkKLcFimNTnuR29fRuFLGr/I
7l9WXHHUtC8eIGW2hOaiqW/6fDf/MjrC8U3qtLslH7AYaoGNJwjVy6TvyKEg64SvcJt4qLnXs0Kh
XjOptcU75TaLC5WXK6Ej38VFpIEr3t/16wNs3D+BKE0bBngpi5gBs1wOESGipNOJ1HryTf7USSNu
hrmmDVQhdmeKyBOy0eI7LikTkYckdKPbVq+7SlF7PojpkX5RlKyN2ql7F31mtHuKCLaFHOn60S4L
3hzryvB9X8JHFewWVcdkmBHhBuRMXqNwbaaN9eDFTvBADDGkcTmQj8tSvE/adAS8wsHNRYYB52yx
cPCaIAr574Bhc0iapCAnr6SSYTuYbPAH3nv5ny16GNIj/oWNcIEZ4Z5CZa0FAPaleeNkYflf8GBn
zaPtAmuC05kmDo/oBETAbk2tKFA9rqqYKL8iJNIhWBeKH2lVo7c1WP4p1fz9skpDMzgOrvi7BNg3
WYwSN5dH9i1+bZJOYWJB+7LwIb6yJ4Rqp4NRQoNIYFk9kd+lJABGitLWvEcMiq8R+ko92YqxWV8f
heXO6f4sv/AMIOJiSRZylggrcm6seQ/EgnEfqWNtM4Vk8DtSmQKh5tTdRWVLGgcRiSgM48ViP8HI
VIJvZZ4lG2xTQQCjjf9g8G50dqD3LWn8UEKdKzEnfVGuKuX88/WRj5GXOpYiIsBWN1wSeis6D4zM
Ed8DvwdLngDPp8GaGFmIl3Vw66mqGN4PonBGrJ/jVM/3H/X/slRfBWWGRTCEwDl6LCUAr/SUhVql
0K9KzFuY1oK+beFIrUOluHjtCm/Yn9RRLgD3i3LxttrO2MoB7s42vl5pDkXheRKheQ2obdzCVYpw
W6w3hQS+OEn23EqxKYMADIkH1Wyi7fH8SnqYe3NBil+otsAtNN7His7/Kd/SfdP1b9dQaYoD8HrH
HKmQUHTn4rkJzTd8H1i2DJgat/FICXDoIzaqag+SzMWzdIy01V4Kwj+QexyCysj19hsfeJH6pvri
izFJLr6R1P3klqytzaYOyyfGJXfBThdsBX/nz1BKIPXpcheXOGbnAlEhHGP0hl4brFAr2jkHN9Tk
6l+O06lzeJsjjHRLqQKnN72x1PKDbGohxALSkjrhzLy6aICAzlAPMSwfsKVYzKtCuiJrXyvSdaRD
M63eTrof78X4SrkADyrbniQW2Pb3ojoNv6s36uc5HeXYWc5BS0fftjF7G0Y3MR2NzaMrFYdMmljL
JsTgEqDxu+wrwea1ZbDQ5W2z9Cn8T6I/7Ma90qiKaPdWvfIcZh2zt5VGAQps61vnNJTxEHLxTA9S
Y3AD9Tct2CvWwnLu6m4WiVlgZ92YzQy8cECV1NpS0MRKihf3z7MfS8g+5sR3545qRkQehoIaA9yO
VR6MXUw2Y+jJjH6TzCEUDQT+Rn1ie/AkBThc16EX01wiaYHuVVxgO5nZcKbQMMJYg0nm1nAXFAdu
gx8MahKC9kHuRk0yKh91iTp5MvQpsZ4h+Dqa8uGlMOsdh1yLv2zZl44qVNjq4v1Ue9Ym1XquSHwx
xaLmABNqz8fwu9h3wmw1QI3DBiE3qdyqh8CAXsr6uNb4ygZ69xnDuAlBSVMd+zUSiziqOP7VJsJa
M5xfXRQ7150KnWhm//EsiSS5WrFKMxsgXiNG5aSAAwIfuRb/2sEKoEHtG/qQCFUikvrkAWQcjy2C
Aep+TxtRaj9Hhu2RZUBH/wICPATC/kl4ZjtVHAhtQKCoCy+VyuC3vu9v3+4wIPAPVfi9CufdDiib
Py5AwDOyEZEjbUmEAW7ypAIkfzZv2CXXMHTJCyGx2AeYK5TZSHrKku9rRvqkUJPjD2+0cjlFGgZD
SEIYbILfbJhWT5aGZvQg0N/7QfdL1AG0l3Rm/dRrVT8aSasq8d+4Tg6nly8kxqa7Il7kcnOUbL/V
5mE5gW6/Dyyc2HFL82toFmuXt3XCxrdRvC9DvmjkQTTsfV1TMZMOEoCNaJmUgK0he49YiQAOLkxv
YCAIjTnCxZ4YZfdldV5YXSGodqzAVVn8CrmfZJ5d2mzUe4DpsFY4Twj6iFfLKA+2RekVzLyJxeMS
LCAkwvxJ42mtx9vIe8ZDdnR0/R4pWiKvpS5eZ7nH7DMY4GMWO1keq7tQpMpQGUVjMFzavzB/yvyP
KLU1b+E9CLGuBgEsF1ylaImWVnwJQR9KEEuH/GJ/rf3kbx7ZPLPJU7GqzM2HI8VDxHu5weCE60JS
ZF5sb08blj/1FoTn9D1YHTy5Qj7SOjGgiTkHf5gjHHfGyY64VrB4RAl/fJOjGSlIjrO9Z1ojRFEg
Zs8NBcP63GKSLOW06a/KAqZZQSQrq79i0eWZQXvpIR0guzlweK9fd2MV3ZX5fnvpBLWsJ6EUd69Q
i5s8HM/UPWxFiy1AA7brT7fyBlCgEyBpNmPAYIO8XGTgr7DHLuujuAaMC5VzdD3R0Va3D/VUygyv
gtTiotAFwOLmmDjAekrTBS4w0Xy8cgdtt9sXhtttpKBY2zF4kakVuOM+W0WlZOTIfiNNI8E55oYj
zeDve1CCoVvmteybBGLJRzDP76D9680cEJfXQj8SIgKQEu323Le01zNi+tt6S52KiABptBtYaM5i
o+TJoG4JAutnbFsmpudzskpr9YtQ4l+D5XaWGsqnDYUKaxujyp1hhoNL9hRtroZgGdxDOXaUY4NI
MzKeC9h0jnG/XBromj0oYBg9ZKJOYYip9KPYYdOu+i7bSgD+wZPU9Dv4/Cr4ue2C6xYDV/9vBV4Q
MgsAqm9LkThfbKXbAu7G1JGI26pozFRYvnXnV64buOvRjtIJP/95UfENW8/Wd3RrCqxru7+ciQ8e
N4L3mUdz+hTDMqcv3Ul1mM9zZcbNHM52Qfkv+vX0yWJ0EB0xEshIhABX/HTAH2yhrPJNoNEZEYIX
0vQLKXQ6XlPWUER+xTUOLNIsXoUQP0dgZT4ZkoH6mmMYJtfirfMOohFuR1ncihn3dke630dUAlmZ
hgUwEOtNiHsTvYlgqHSFsO+AWZdZ9Hrx1QHeC8/6lPeeTXuc/0O9rSl/nK08oYUbqlSx3kLa0p/Y
oachTri5uyNI26Q9x5mj8BniGMVKBk8fx4fjISeSzgCLf/bEZF8nnCf6jFKk5K2X0L34WMKWQk33
rUJPXthqagxyfpUXMe0aCUI990fuHNcipdZ+y0VxGwChufjYBuvGHCKaXi1DNQGlW2j48Y6lnViq
nAatzINmTdWTm2RFec/9V/6w7hodzMe/tF7PxNBRAnhous4ZHK2VUT9NCzAhLRtrlzwhga4K5yYp
JHM5C4EEq0YxF97IMceu/U8msy6jbbe2kgeyIyfD1MqbTbRoI+IPgbQtLvFNeGbJzMdrXeoWVMCu
BFZIflsrSncmRN3ka7uPSkh4dkg5+Iy2hrOp1h7zEKR97cF2xTh71cvQkX6BYHHGDzY2/fqFSxUY
+1NsMdOo9k/EGmp+6qdE8z3c3a6Tuh0zsvcx+PhJcb4gHkyEDjLrBFB3dV60EGs2VBBV5W9+c8Tf
o5CCX8Ahrm5oS6Cs3DRnkxmS44qsXR2pFhw7dJBh7BVO6qdZgfs9+0QMBS9IiNlybxuE5FOZc++o
MrDieMa8sJ6Mgi0hHA+Ax0zedQBBYEqx+JBIZJEVrsrz2beQW4HkjcbBPmZaWrX9z1/eTJrd3N59
tBhO0tPnBYClaiQ7XgCv5nyU6h01VvHOS4ni/fZDva4ykv50QJ5+hRapqFPl7KxvkEVH7CCZyQPX
fWwQCCjBs7uc/K3/Ycb3PS027pKKiRKdz5j/GUfK0iB1jXqTGsJI67TWHUIAX72s5oUv/dKPPSdy
c8f+IFfH9NeSXo7jZcs0J4qjsWQgP9HhrNdKi71QmXcRYOx+ptnj9/xktgoVhOkbKRpqtxZR8zfX
Cg/ZY1KWaQqb87A9aLjT+FzJewtb1GkbWEXQFtEFr/2cxY5Jiwa79Ampp/I8FWJOdTgFh4rAU+9d
weVTFIrteLwtgx89n7es5lXWJL1LZSnihFBOzlwHtMivls0NH1Pj85bKsl7nZlJS2gJ6sd9eAwFH
R+xLaH9Jt6H4iPNVRBQV5DOYNFq/qSF5ftqfTBwt9pC4IY/m6wuyG5wJ25yu5lRdQ0oLhcKPWoeb
2wZEZxG3OOa+kQDz6PRm7XTneARK1t0svB5V5mj1ep/DUsFCy2PPWqTF9Kkblprf5VH2ZvEFV1Yd
ieKZFeSyezDXmq08EQnX0uxLym2eqoZvoPO1Dht8VtY936FtjDRR98exlsZcqGn3Oi6yF3NiNeRf
cfYjbHaxi9lGopPfsBT08ArwXkccBuAEGz1QSLKylH9SfNOIStfOmzrVi4EJ4XVK0vXmKfGu0IUa
tt48R51VF0nQ0lbdK+xGupiP7j4JeUOCM1x+Raytwhy4qNSbZgraIozy9FzSuTkp/9pceXiKZ/jS
DcJ9s1uaHha2UVnTBV1HJEiFH4A+8uLluEODD2KRYumaX3nOkynfyv447JEDxhxsro4CU78/3QIC
glYgywJRy1DANozLBz3GDcd2G2NT6+PTHej76h3xzzQynh8VSJvuHNNy0FsOvA3pPXzjl1nGs+Vh
A/NoOaMKUQcDUPQSpz8yPL2p9WpnPnaEMy809/NhLa1JHULTYMLibl/wJrADiSbX4C1tlvRScLEr
lfMCK2oqAYJndgDvTlrXbI+OSmaRxgRT3tlpU+jv70AVGfbzVOTC0PXqgbZZsPPZWXDFMr8OND69
kTYefkZWb/fvD3knDO6kraYn4c2dFgOXSWP/4ZKQh6VqiO+eor9ldFCJA3D/Yy+7Ewo9yCbZSl8w
nh0TJnYkTLI7JTcXW3RJlKQkRhjry5cYzKxo+ZGDoPyn5bNl4VQiIolUUfI39YNBe5yhEhCC2Zgw
quLTjhkJqJAUw5b5j9tl7M5/f2qGeSsbigkVeF+Kkf6siuiwC2EKdAbWtF8Bk9pM5Uw8YSUAHHks
vxK32rhOY21P+YRouj3Q4BbrbfIFoa98y/bW8PdQ8UoZIO0Wz1rTgruQFwzpje8NakNoveR4InaY
O38xQct1+g//V/tzaLEHOTTzq5sd2y6zBnNlHnhGUPTr3cfFaIpOZRkWyBrB0+JNItjapInQaoMd
0NEvHZ4ymoD0KgMrhWiAeveFEgM+FmxMKI2uk5TRlsqjKTrC5u0mlVldCedRmt7O9DGpGQ4Pla6u
qKEaGm8Z1955EnhLAK74V2RQNxjCnBSFJv+W8xt6FM7c0YRlN8knoQSGjjiBzuMxsUsFsHF5eKQf
1ko2nSjHQ1S6vic3sqCReIXarKyUep/7KN0xrI0H26WG5wCNfqHLrKW9scJIq1EcdV2AwW7p1jv/
rsVD1Wgv4XUMRfdAOzE3svBJIe32pREDGP6lps14Jw9SGIhophRg/JCy9i1mhDoJX5UI4cdci7J2
IpiiUiPBZwvUf7fRYaBKvoGDQrZ7vuPY7/CKY9JV96ZCmvTqkLUjn3qZYFJ6RFiQ44vKyUDF6XDf
ooF4AA6UUDtgrK+yFtRACPw1YUQIWpbrmOa+7FDs3KTH0WldQUWDvO8gE3BFzvZJ4JXqe6daVGdv
P4O7yKSaDKU8exSESw2kassXRFoQK1aecK5KhFnMX1PDubOVS02apa7UhHQheWbB1B5W9/V7NO5z
LWcAKZEn1MJOq8SWoxSdapCV/RkYU6UQahKazsbX/kCbPZGDvbs8UhlAPOmsKOqZxAko8yWvyaIe
OLhi75Lhz7DeHRhp6h/rKrhXe6S4eNGuQDxk7lTDZCXyrawP/2Kgtgzy2UPNT39DtNKAb78BGq+k
JPauOgAD9Mi6xySFCFxxrrTlQ0b6cvLESP8msC5fFsM1k7PQXH9XIBNgYvKEzZl6x+z77w0zKVjl
FQqNDzUVfS+/9zPBziTLA9ZWC5tF8VlMAWLHESpd4U8l4m4dOxiZuHSRKYWcftfSEkgdZZQ7ZcxR
VBGOpvzYyygdTO3pcjlaodM72Y+dPBjjVj1jPrsGRg3jGPaF1N9KYqCeHLeRTDZ/Nr7qWgGkI3WA
1KAPpdR7svZJ4Uuh7u9b92DglkbGypst0Jir9k4KapqziGaBHaCPLWZrTkU9SC8xaKJ+bUu5h0RS
dwUSRuLV/GKu4icuyYoOiNLrKjCkWTuYl52eZzkBPtbFUdMR8YVK7Ss6EXjUpbqln6sa5GVUZGah
f/vDa9kktd/eO98IojWtsxVwD3SXhoutIay027NcPRycOpJT0z7JDekw399okmvJw49mPIgFut5+
oPusJe9ShVRFupMZ4mZyBy6YD8Ze4u3BvoQMSr5xUCs6XtPEEf44AB0o6NwbDhZgL1peFPSgNPkB
Zi8/wpv0kRI07zxdY/GsnHnoIrLKFeWaBb+Fh3r1+QdHLhTex87QAvynhUArFGdyYd/9b8f5RNNd
sFaEFBj2pHueuF9yvFr6Ut7PefNN6DkggNU7YF2mevc16Msqoju0ffqwAKHylTW12RWmfG3NC4tY
mLXHPea5A2JmoTPT9d2ktbxFXLsd4oQyM/w+vHfc7JZAsgVF9mt6tRVzB7hjvjF8H44Ub369i4qc
FpLBUZVg+g/NxgFRmsp1LZvKbpR4/JqN7BsP1XNpo2GP4Uea6EMu4X6SkMyZxfsQEedL1b0PHRAj
cvE9lDySgmR02ztZcJgGz6eQezH/8Mv1vjUFt5UF+n1/Y2/OdvMozb/xwIxCYer5yEQBrbR12tF7
xDiVCyzmei8uqnYXDSTODGhr7sXxfsuyEUM3AY3uFILN7SBvmCiE/oNTquoFTYyiscEf29qxudVN
igXp0A5Zg9FOu1UHschXQi4LQbf/naqaPbXnhZHcS8XldCF7ntNv/11FLVQTyv7h4QkrWLXrBMRq
y9Fvh8hn2SP9XaOJKiiFiNImirAE6lNEElOU3+RkwrIIVsYS9GLkzvKUnJAkgNovJWCbV/obuIn8
1l5nyOMEe3NWc1/DR/VxGdeU2fevYaDwK/KgkBnrDhNeN2Tj/ZQQPgZ7GfZYhLE/QRbTQx7d6WeG
T9s2Sy8iHa6sI4WXhfdamU05VkRH8MTP4pUJ7g1llUpPo2+eD2OayoEeGn0ApQN/YULb82yA4Fim
DREMnR+9EKureZUHkN0OSoARwfI5Yr/PVE6Aj6fLWFw7+iIJjQtWEfIH9UPJvCO+1kAYtZr+VvE6
39w3m+HyXtI56ySyWdVeuqe9EvuBJZodWFFxYfZdANY16nsTOyDcuKBSq0mL5JIQWDJZSdtROEgw
e/Pbs6Dp0jSu4GGFKqdabQPiAuerBqj/N04Rc7BBwc7W+pHMbzAzTd65NbWzqp8tVy7TdVNpaMNE
PwlBVzLfS8kAAUdKZz4KcudptTEM791FiOw0z8xuRSSItzKBCxiWU+EPrgf94SEh/rX+rArSOMcY
gwAQg7cc7k7QcPxKxWKEYz1/XejDoctP7gOBBT2zwUsRfd6v9txTE3pv26VJfWFAc+uIKNe3Czj8
NMAsDZhCzXHg0hak/ucGH8+rvtsG9i/25dEBDvkuJ5k3d8OZDBJT/RyNo7gTJ1HLR2R1UBhsr2Cz
CCD/UqwOkwBFNOXklgePBocjgpV7gRbA7LatkR9QQNBWfhIgLl6/lxM84cLDrIobsR2vtj89ZNCY
7M/XCjmMM6raO1A/GYMuGiKuNxnpje+eHBeKt878lwU+FKGbZ2O212kKAWVU57AR/SagB3WoeyyU
ocCRZEzq+yCywjM/XjtnnY32GunnC7Tp/C7uiyU1yuOF6kgBiOAmQ39tK6sajRfHC/uZGvAIRU3j
8lV9i8HlKTdyhDwTz1QNqiqdx2o5pdnjeaWL3qiMlg4hb1f59VtXwzjHYCeFRu2NIW5JuvrlvwXQ
OThdd4gS8GRdwuIpvBQ93Z/7c2BFREioDdVwBUA3rJpXWvuUZ3aSHXaXj68Tn257/lJXQ6r9lJsI
UMw/wbqAFdsGBBUYCOOak7/jgFx7bhsGVnbeey9AMhsMuDJcIWpE0jGFN9ibcLsj/jbbyc7J+4wq
KY2r9SYtG36FZXXg5Q9COlAHrqCL875KcTK0eTsgoPq9BBg0ZZQ6E0K+dB11Om+RreTCqUsCuOAn
s7B1ocGAnR/Tthpz+zYGC0+K4LOLX1G959rdg3fwiEpYY9hDm9eDo3abeE0kOxighvGnwA7Nciqo
gjCAsr/rZ+8VPJB2QnxVhYpqAFQOsQ7ZycsZ1cEOVCvK1LuX2nopjAYF2XbVHxhYSlu6Rs05UllD
+xrb/oYU51plzOQnZHpmGkoo09o0N7TQpzfNkut2KP21Z0hvfR3QGV4Hkzd8N3zS+CGDIo18VmbJ
L+l1wkNH7uCgx7mg+CsVr4CC7QELlPtd5STURhdaY41kMVESqfuw4YEnAefiXDHcgfQ8BkeqX5Yi
y61F1ZQh8EZzEYCtmz0h5iaZjNYVuARv/MUYq2vpxgSJ1zy018BNxCkKMggmj1kdauutU8MMlECQ
qFBumK4VQF3a29llwZdfKKAI2WiNU8SojDQqENZ2ttNAbrmm9OZCpJvgLCKPvFbacyVSne2s7xWL
OuEAHWjjzRIo6eIZ/o3CqWz3HvsYt8ENIw9aC5c95woGhoZgZKP8sreJ52qxo41YtsqaUF0z9tfq
M19JuP1l8oJeG72s3qmbzCbZUya2TjKOTcLNPznL7wH2UAiOqUPILOsPch8EyBD/7NEEQMyxVXZI
XiieuUsKb7f4U/6X6b8kKL/zw9qQ2ovSWzPlN7NEvmnUQASfD8SkPQdhBLOraxOG7xUDAzhQ1VJF
niuTZvmRD5Bq8y0rh/5JEQB/9Vv3Fz9RGfLqZ00F2SYZmKYQnJHUTu+o9j4r74GCnpztGVOFnbdo
DzoN4XbG0VlK0khVVsSNmyu+8YiaxvhDwSYlcTF4VRwT/zOeTmQlk/pedi2qYGxag574RVPIonZE
oshEwcXiKiMNAscVvLzqaThxSP6ewBIwJP6hFTQoWUK67WIF3hHfb6lVO9BFnGYgWF6RexWIp0i4
wjUKXUvSU2wtYI1HGdPuec3Lv5drMW6P6o49X4Y9JYheX8IQ54FHAWQi6zoOQ10ZBt4yq6ks5Y1m
AxxKMtNuaHE09WnurMEt/zALhxYLfpUgR2Hdy9LTf+jUDJmWHOcVLgn4SMQVQvHJ/ocIfzYuFk46
NptZuVlyBXZhu3ciy5iZdTPBXx2rCOObIg/a7uihVRO/7719idRL6SMOgyeh6I1mhrLVjzNbGiJl
KDaw73BWezzHFYaqNSIO6w+J8k/j+KDL9MeSOVSEaHdzKkDIWzAPBETiySvhXMBrP9xBHF33do8Z
gkHdZaUF5sLxIVjc6aBJ/zusqUMI2kiwm38xJPDHM0uDZ/yeVnoBNHffgQrl3cE8eR0BkprRCko9
wR505eNI76m0j5j/f/6wykR5LZDUHSQV5RPj3C5iBIJkAfxmRvx1LkBatnsPSmhBJHfVgv/oHlV7
8QZ2mKUvV6eQVabObe1ryGJEy/RJKndfHWZ9aZTOnVuKdSoT93oiF7OZACnPpi5wPMD2cdVrDZXV
biPjDHC4LGwQOUS+oPaHev+9Z+wlc/OQp1eNrH4b+aclLCg6n99WQsmjAG2tlUOJXAf7uzJsMPz4
l8O54Di1WXNdcnWZaXy8C90sWKu0PuJOObXzkGDFSrkslaicz8FWvS/JMz130G2AqH/hFd4aauIk
RZG/QOgU+9R5mkB2+af6/ws/DxFhijZrqrFDkOzC5+2C6kUgGtb6x/bkagoXUXgGUeqrv4VGkPXt
5yy/Am/t/NbCZp4bRstl5bWRwoRoVZGjsG0Pp2levMVCwG5tt0BxnPVVcTKu+cf0z3B8RUxSCeBJ
Zp+tqwmbjAV+uhiASarwkOoSI/47fEQMc1x3Trbp1V66+4AlOf4wmRjpvIJQ8D/3Pf1JO48MsNvN
LDqbdqc+cx86jNTKHPAj9+WJqzCNHz+ZR/iOE2zG+OlQYoZxQt/E7iDj/j5fZixKP3o7uJmcwsiI
dbss1Vtmh401olDvGMTxFCu6udMGAybi3VG/KYqs9CWIfD9eSDjqKC0X9UY6LXBzlDTL60LQ6EBz
LZY6tqJxQ/IOnRWD0ctZjvWwHC+iMFTK9HUEInjtC2Dnj2JnX4G8cR8DmRTOewopO8nwFRN8gG9h
p+l9wyxTg+SDRnD+A3UXCi930hOu+aVMNpR06dM7pkfxclDsyrBz9AOhUTpYpsARZDdC1bO/Z4O7
h9d4bV21ZD6veHC7xltmAspgS0eKyOPemxIXoFdJkuYNwQIUh/NWMIT8EWZSS5o+7dJZwXr+FKoO
+n8DZ5R7pb633pBUG+ebERcYxmO1tkdcizzNj2VCUg8a3p8NxVkG1ZHWFAWZzs3ec8NbFUMTGTY7
VH3VqXp+7cbYIETfYBpiViu0y6tWT5WkNveSLipwh+Ezdu4yn982a0mqf/m2nNtzT2MNo4OyVsX9
ZPsa+LF/ZFTDuu/yAiRvvV8UGeAey+US6S6mS2I+nCy8JUcFCRhblmwZJByqF6Skp5WMhNu6992k
IVn9W/XSlQPpXO6RRGvJ4N8rWZwS1LQI0IFujzQmUxTCXgn1NmlxSrT3fnN9b0WE+R5kZSSdptoy
75x7MD4s++NmgAQTZILhC9gxy1lu4qEVG2gJAFkF2Rgt3YOawtfAG26QG+eskvVvxqRGqvK9w5do
8d1cXtuTtYGBpAKLhAJaYfqLWDJPmVSm706HewRpx2A8R+7BhkZSx2p6sXk2OwmI5LZSXaVlnP4w
bBJhR5PXevMoerHaOMxJLGGG5BWPpdDz+xomMQOSqum1Z/Q/DsaSvDSvDKpeVQt3hEO0co8Tv7Eq
yDNQOzrjClPf9qEa+aUNBh/gQRNxLlq8WGvI+f+TCAuVBTTl9CFbqOJyIIiZ7SFnRbuuDREjJZG8
RqZvFtzWraQIhKx/eSrW/KektHZ2ZxrTFU6FZ5V8ET2axxc6Zg2CtGnqWDH3luXy60xGyFCJeV6U
UJursmP+U/jkPX98xv0t7ZId9XSnHqy4ExrO1HiKnYjBCIRlbBHdLHlymTCOKrlSR2DdIEhbpXf7
1H2mjJWiSZZJdYMVzKEPNk+ejQAHKs9eJvEkjBzvl5LUCpWIN90wt/Z0zMxi93YjgDAIjTi8bahm
emD7ByRWmKRKc/OFRN5P6oGxoIlE4Ytb7ZGP2c/CXZmP/0g1gl+HpItpXREsqwHZV1rsjRDcdStv
bcbZQi2SyzInF2ZO4uBuJ2kebUN8sN1ZsCbZE8PRI6FIItLfgDeZMR61ppUlcRx8mWuQBdL8CUGo
YuZ73aE4ZEkLldTOnlDGubG18r4AmI61wNDYJZ6tRkrla8x/LTxrTQPGTRPkXMVpp2K6H2oVjzM+
mX67eYUE+7sMPErXEESkVd5/tcxzzqNbIdLTsG2EeVqHMXLFizV+siH6UES9HovOK9C5xtdc2Ee+
G+pqiuzzzkw6AU9idrrMc3w8ELmC01cpvW6ax4GXis05zuGa1ndhmLTyvv/fXQHS9a0Ku1AN5Ubx
ZKNn9kbONb/EKZmJIcPwRhefQODnHScO/9yOqxhdEQALsZ3gpP7t1GuATxdCjl03wtlmUUs+IfLS
nV9Sgj4kqFJe3SGecpZJS+on1SkNbwO+efvyJwRFzqzSj/ljkLB68K5Wu8MxUCbNU/VL7nXRkPpn
F+x/DOpAppdxQfVb1+n0WzLbi8+i7H3zeIS7ZeUPcB0EDt8yb1PM8DtTXhWkVJ/b8OP7tgaV7pY6
2syL8LHPSMCBuJy7/2emAHo+pdWJDX+G4SIAMYjJBTkamW7q2Abr0ocv386fgl+SQr8g0MPHv/XV
zUewL1f9NNMmXex5pwTk5xHuRCbOVI0hgXLx8FzZGg8emJM0XGPnziWBxlPzdGuC2vP3v05Gbo7D
iYaVvmZU0QPn3lHCXifVEGHSXpL6+GajoBPYuVdSSUtJ6TsznMcZn7pLzdTXHNj/GZyc3KCqf1pH
e/YHtLwMzC9+uIXrmmMJTbxrQMZj5mkCG3qH3fvQ7D0fcVhRhc++PeajXiGjWJnscFCaEt7XbPYC
Zvp8DeiUSu55l3QIK7UKXfi7Uusu9AdYlAyUX0JqBRsCh3mnxIj8BAvVX7UtrC+RzyppfZiprQHp
VkxNbplyp248iN1mYdPnp0ZNwBFI0AEHK8YtgtV/VbdOktiAhzmgv3tr/MFy8tUGuW5w8Prve4od
ChSuJ//rcpuZsJIOxZv2pXlqjUuEw9Eg7sqJ/PZSSrdlDQ4IzbsHccQa8CcptNUXUT9DO7ojkkb4
Miv55PxAyJcjXBFg5MvEYB7lRMMkGheOsswyspc29SbA9FfqMcQsfc8w9K1MO7J6lYX44KIavIBg
rqNduG23OaXnQO4RgbRqKeq1jBosh3DmAiZ4CR8eWzIbloSaV3eCFG/+B1g/hykmJd8KM1jWt6bN
qtFhekZPv5oMetLgjHSTjhLRe3vvtIsd9Y2/vKGsRSQhDCns+xH3hZZju1feGgZMEhMjUR/hVpqb
v2cKqCKTEaF/ZMHbramBiSy8tz620xFlEy0wIFI990OK5HuCU5ilUwrrNx2SuRQ1KzKjUtD37FZo
IYxQHblforateuWA3c2ZY28XT7yLyI57F9wBoxj7sdrgTZcr6aE31mWo6xHfhHbIaENZJmMAOJEn
LDCa1oZJE7IEwRljdZWvQmEKzxkO56K7OFXB4Vn3EUjI7XLEkm11yB7j+e9xCy5oMbVkANb+G2Vo
bglphrp+U5y2d+EudA9SzmMCwCsesmmHPOeWND6R892e1fbARl9EagC7ng+8K3vHfRrNa0+Xbqvt
NjiEhMlAid/bv5VcZP+oxAmsNo+yr5Qi13COXWah/aHbvUvf4vKmHo52ZrJxLVgduuGECUS62A/b
cPxzy6PhoY5xjXhChIWVP2W6u7rsy60I7rhHd2LbFBl3EtxSNcSWkLOEwGx+jWkCILHhPPxkcp7C
2DNbjTBYMS4dNa4ZGtIK3y0HPlHhkC9KMtqNX7hlXc19JcUchcBCwiIHAfQdjTA5uvILID0BCS3q
nhkLR3jmiwEtuWFkM6CBMLef+naYijH3iwt48T1/YTBjb6T48bRqYVCgDgEMZHys2GY4jiut6Ao0
sfghE9K25RHKQpyApy3Sun/2k+/9EP9f0arunocKIdQqSSDR+60Nz6Se97O8baFbgpBAGtwzQ7SR
W8x8Af1/6ESZ+XZffsjISTnLtlZK8eKu0wi6tvA5DiBxjPLFVoDE9UPGGkBYVL2LikNSJErfFow/
tiO6yS4v1i0KGORLgO1PBflovGWYcepREhejXPy7IRC2W0m2yOvskb5qDlmcvjzspZAhge4rGWmQ
mOFCyWZ6zdPuhBiBxeWKGDln1cByGvfw2xZJ5Kx6FsfyG4dAArpgCs63q7LarI6Qu2sLUdGpjy1U
aDgjXxNoscduVLiRbpiGAiWiYigqxcRL6X6s+kTFWFxxt3lEK7d+Tx4ZTm+D6aAkOAhQefilgh5w
wBzghOS0dezqOEHfmerw/xS9le33JvcE7TBfx0wVkjnp0DKrh1BDHZT8El6bsS/qnNTV1HwTSPeU
oRFpRQ+XxKlL4ZSuBJgjlsWahs7n86hplq69wUalU0tiT3noE82t0XHtTjl/6f8PnVJqLEXGeh4d
q34+TitqklNO6aSEciav6Z8X2FPvPcWbBkasTiQylx86tYECvcXVBQLEdAbg8+ugunnoW77/OtK9
jBgO1s2Qtsv4q9wuIQwegACI+AR/8e9fhzpe3rWcNt9fT9g0Mf0OgnZDirZM+ZSRBpdwpElCf4zl
afBaGhz7pMNyRsh/Q5vP4pFuWx0VrqZpgn4IpvwkE5e18vBAIU5ev0jbwt42/Da+4OULAqqzwhvD
bnz+7kYd+PYNoS0mHsj0vnVQ4yRQKUVOkDMQY6bmn3PIgWJ0wYIIXN78EFh2QcAE1C8b6wkgZwJO
fGOu+0CnL7lryanWZco1FeKxd98PKPB9EdVUER/xNljZ7PQkVv/VB5qJChAsmpf3XN4sjZetH0t/
8qdV91OXsMCKRB46oxZ/k5TjYOqmBMDY1lCoVxPk9Te0nVxuXAO4BgaD8HCEIxnCu1zMFw+cQJQj
loCtneAOW7THEGSR8tUXoIKqy7zyQLo5DHVnt/iwDyx1nRNKUjr3V/uLHrNFpAZTkCT14KDlujI8
A/fgpVTik1GRyQvItx1rscDTsOH9P04lNtuizOECqUPZgDiB0vYszPGtiMQayxAVpgZGThn5D55I
Mg5u+VFridJJRRmGKKLN9AcVHtCEth0iKcD92ZvAD5UbWgSbbPK7CILBl2WQ0JyLoWF0Y5sVt1np
5kyud2IjYP6eMPRvjofQ8O/WMpi/h+c1ojk2ZKRkb32v9gw9f/H5S4qznw+z6FGKyuIB2ToyjvPd
XoMFvMC8E3zPcyt/b5IegUqTse6dzBcvSn/GP742Ox7/IGbsn9yVbqfFJnZsUlWGDhQrJd2aQawx
pGiCaiJsyh9dcuLuHVNmg0xMXAeiAFEw8cTqtFMdg/ET0esHCMcorKkwavLkj6TH2gkLBdHxfVl+
dCGhvlIOjjg3sv0fovErdVeMQjl7mrPBoAl7LYmsWKgqzUjWx5Xnk5HBwsGJvcUvV0ob51lB8CI6
FPebY2Ud6GsnftsHAyi6nUj2XUghZ35Cj0xnL69EsrBY9AlzBIc2VXJQ1vsl5f+tEgwAB7xgMxch
inHNrYA75DntRcztHV64PpNBz7X+0l5oPjfXWMB7vFKqvfRk76/UBRySdtVZjij/LyI5QQTcSjzX
7BlNr2oFv0EYhV2OvI5Y7NWcNzxTvXE0l4g/G/2w6GQ0yIE8HXPNkpUAuBmzbn11JzZJaPbuMS22
mYxhGOVDVvvkcBJLSiXi99VGqJUwcC/nr/IurumHu7tKcUpvYhNt3/8429b/pittS8KZlQzzoxKF
FFo/yFdE/3hbofCx4L22KAercP+XGa6Z6QPqTG7zLS9uZXnwIzhCcHUOX3jR3gGeul10TtBsJ+tA
GJyqoeahYFoG6p/XK+uJsGZxpKwztg+vI50GyvqGmTZ4Etp54vhXYxZSiv0YP3ImTPhMizEBKZFl
nZRjh2EjLVS+EAUXW3kDoxHXMzsv/h8TOukpUGyd5PlfHPDt0UnlK2qmdbcVjekyL4qyiyPud+Ns
PkfktuvlhrCbFk26ylTxJOPHCJRtMJdo9Y1ljmUPotkBUGhNvY5GTb8O0eCt3x769ppNSMEkI0n0
OwS504yN19JnSe+W6O0XDc06jfRUweEQY/i3vnJATBqMas4p7mL5PPioQKxrpg5hoS1RjIWPZe1T
mC3jeGxlttpEzUKqhMoUmkb1tkwQ7h8CD40XozX4Fadx+kaud6GKDfrz7UYDXlo0nqnVth7vv15M
9EzQDSQep4l/4MDQTgexIfUzgrNrJDx0F4WS8go3JH6scbnpB4wPWcfy5q8DzFKoUq+qMNzDjG8v
dnyqQ5KZlT3mnahpKjyxOrx7O/Mthab7u800xlGChTwbQ2Y1vplCRPzGrLl/3m6OJlphoTe6DVMS
wWXXLwDhXTpig64Z4g5aS/LKZTAesuNrt3lcyjz0ahJVqYrIhq3AKAei1F24W6uTXPwY4O3NqbGz
k0vrHO5dIXnzTamcp7iobbB6XttzppHzN7zNt9e5vEYt2fTvp8/CbVxIpvrHx9i/b1RQg/YxHSJT
K7NQuiVVz00RgYSpU0GK5H5dv3y/Fjxkfx6K3YTbwEKhKQl0i6KKDV5hUFmAdSyzGwrgYGIqKF/G
v3yhkrV+xHVMbpWfE01WVmF7LkzeqqqlSsNEn85TRrAZo4zkwxpI79EW9emncekb+oOHSqEG8dtz
h/nFD3tKiPODIdSFRw2K7M1Go/FpvJA/+H0Ci5W+okycWv69VbcqTq3F8g5L1JzYfceaKuH1TAl0
atJKa1haDBR8SWJ+FhYhtBRBAKydLiX3Sz/rpQyY7VnxWJ50i3ZX6h0EbfMPjHCLf4HkJsry9uNu
qo11KVP3FnNhKm+0wvfwbXWUryGax596p3n2WNfieAAU3va7H5OK5V9foxW8VBUU+xRijf/HSoJ7
lBTBvX55Kra8ooLrY1310ztIWbekb5Zj0tED9gn4ROz064GhiDLHk6yk1+4XZzqaPgxo9ax4Nzpu
9a1ilYxCpK3sfZgKxXsE1psUUpnZ38LzerI7sQU3LNPdlD067QC0tpSmwBPM1EifKT5PK9KLlqY2
iapPH8ybATZtCuL7CbpQxYyKJ35vps/KHvapHb67krVo+eFsjcdx6wLjlqs6ZuCHBns/bBK0VI5Q
c9kMkh0cXkhQkn8krSG/5HKB7q7U+OmSEa1D++vZNfzB2v21AU6yZr3Pwcse+FLR9pdn7X0HkPrp
mnS1E9lvn0dfHQZrooi8qVFG4CqO5Pxd2dXi7SNUiF0zDHmefbvobSw/AyedkgH5YQgXyhaHgi3E
zkbOjqBRkTxOEX/IkTYHjgFp28GI87rZ2+b/ZJGNGPb0ywJ8VV4BTWBwpTLA9dCBA0JJCs4tsUX7
GMX/j/zkql1JLP1lM4J9vvIn1+1Nh1gxUH5GpK4Em7udmB4x/1zySQFk4dgVZztVw9/UwSIlp+7j
QzY8NhqKKa7xy4bNBnDPHSftfdzAYoTU4PMrhOrlPVf4fm1eN/Uhm5F2CqWuRahk8lm/LRz8wHTc
nq1PA2Kjp5Ptms2Fky0hH809WGMqDx8ZpN1I04HUgbL5zAAp98Jxd1cdxdp5R8i2VRIPtHQtshuC
2szRMxcKf3tresZYOnwZIuMyojSiZFMbyUj7qXgRIFWigWnbcM+YSVliEqXLTLfK1xvmOfGXJ7LZ
rF4BvFxlzMGSGXPj8EkdeRs4iW/UjjX7NjmWd9s+FqbpMvy4TptLOBzoF4uJHs0ImSr2akbS+Pec
2R5MRJujP0KuWVta4D2MUJbX9elo2HnmrC2mkKOfyTZxuRi/WQbKrZheNo3z43h9AvcwoImjtwnB
rU8s1X3/fcY2EM/ZqSc6Mpi8JSrzj1ed2SjXj+toguLE9DE7OQHKHho5XcD1NDUWzYe19SGQKvho
i3FrOYIDiRbK/ileNLIsjenWLMeBUmxywTBgRWpSj8akvm9gTb9uDX05gKLV8dG2VRv/eciAd0Jn
b1t19eHMtWR5B2xzDT1jYzrHC56ccv6WCDzKRUC/BZ1nk/TH3ZIZsXF3ukJVup0Th7tKvxZFvwBA
R115smbYzwrSywUcZEcm3wlyfBmv1JKvaYnEkhbmedLV7oxdjATrOHYOBFpSGwhqjPvTiUmhmgt4
0rtH3+oZado+ZZsQuOYdjaHynPfMTHNjQjG9yMCTTNPJg/jdJGy1B2jwhmVyUCX/KcQeWQ0yp3X2
M0J3L8JLFN6G0sxkZIEZ5f40RYku0vmyoxMcNrI3uqo+qvlA/yDQb8VAhW/ITtuxNcVxOEqzUPC7
9SdQqb2IPe/Yya7P5LHSw2y95HvfkUCigRQEqcg3NZFLj69Y5RLYtX1KhadX3VW1zRT1l5o65Cnt
8zTDpATD/l4haobRZMJnHkzqrTewhY/HTrHgjNCvk2a8vrtKg+xKTx+LNaWi72YlhVdWxWLSkGiy
npoLpGtWgS0FR4vnhOO4/mnAZ22DPS3a5NYyWMks/ss19yG6bKeEb80QJ4z0A9iGclputVZSAvcj
g5CHfdaSpChNyPhkwF2bIR3aB8kDWS8bXxE8lDcY4aUeBy949vOTixEjLy9ygF87IZ3/khi98pqP
SyGgZSgaAV3gpS99fPbVO3QqeYLqGBeu50vtBMH+Ws992pQjnN9V3WT0Pd7rZZU46mBywmEphKWa
midC3iZm3KlRf1j+IBisbx1Guq+++y+DOSJ1iRqL45rl5hCH6FY1Zg0RMl2w+DC3+TenPCWbaxOB
/1ikplHGYUCUdPXI3LGprcXBPGiyy+8ssRyMCI/uRnfV/iWz2Xqvbv+6HI4ULbgDcJLq0OqU3wOi
3y92rTR+6fsHhI8MIFltEF6SGBpzrPtSrnDdsHNzpbyDI53jU/SjsmrilwclWk7qCAuxi7eTqL2D
CiTlMIZHY9VWkOW1+U1In/bWwmaDcZLAm1SdBOTO8c3J04ujFn/jLt8Qx8vE8PwM0tbaJptCd9ig
666doB+w6Uz1FjwmceZuzq5BUCl9xHnzPg3JupX0TtpmrF8KW7+5cyKv/yk6Y4ieJghQTa6cD+fT
YivKBpdro5bFMOhJFMDZpvxwIUDL1aXgZyyRoDCrOVC1gXMYu33R+fMqX+gAoqFnaGwGikmEoogA
IU7jil35tY825Xp1IhxFOhpOTClPZvsedVHL8eB3MStL5/n73N24sj2padjTI7Hv1ZXPjqa8jMP3
XJqMaipPSmsn3ZLwW/gEjBV9zD+uIyXndwVKADKDzXhK2j68P1QZG5vNt/fUq+XYQDZjFwFhWHuy
hos/1T4/oGjE/yx32ltRQDRwGrV36KzkZ5O+PkLlR63iTMrXHBUWfKVZub7jbBHNtaT7m7j1XJST
Rm+B1gQRwDw4fga3ZXvCvR0jw0/Ee3GNrpSc2oqnXAqbHkSnTasZK4ac2S1naG735G/Fcg7Cq/0r
oVG2PDY/yL9T+wr9/25vCv6giCeqEgSQ5Jp6GgUGgRIx7JGPN58opEE5ipLlsLNOy+m4w84eZx8h
bbRgfvbpQt6VeOS+cJYlZpNhcPqfrBYt4y58t7e5Xh5TshyPIAq8oPed0nceoteIe7cGq/BWBR3z
g5vblO6XcZ3+yxGt3b4GnC8qjwpckM1TKXfKr3cJb4CQdHFc/lRkpEpdXyELRSH/1kBBoXHSsfxa
RiVOtpmBJEjK4vwIRY9PoUWAdXSyICnN0CVLJLZa/sl/erbjwRgG3pBKn0K2N6L1mvCcecBVTWAy
7IgUelkktEOpHWPhKhyMsLVbEV3UhwjlgcogGAZfNykHenJCvvKd3SGDthU1Z4Jtv3TAzgDdM5vO
cj/Tq0ipAdS8IFMBFMGM8jrrQBUgvL0i8ZJE4BGy5gSRX4wwx/wxGnxtFyv5WbSKDf8UHgVsCzS6
AHgEXg2qpew/xOmAhnvY0rmzToG9c+dD3kwrEmdfRu4HBLDEDxn9uZtvHVr6En1r8j8iEgm0jtrb
Fh/yTnf4BouQVVxJuwrV6rL7SPKE8zL+kGa7sA7UvT5m3xdOncO4/dgOOonfZP1XyKCzLIAgB5yX
7IMD/zR/4DTd3H+8klVL8yUuCK3dhmK2pbRa6ALaRt+OfEZ/d3Z7EQOZoiyohvYnmM1nvZywUFDy
ZfGifacYdTIESYWNZA6HYq1heZH/T1pH/0srgFgplLTncg8iVJgyr5fQzjgCghg5dMYe8fTDFj03
jaaIazEEqGvcPuWZK9y3XI99MAESeABusLzo1ZmWd6PYkTtnheVVTupHk9L8Z1STsDfRZyVRdn0l
TH12Lnwl29pRCUmxDP/10Q9s6eyowyVujGnsBI09c+Hs0TnwB00WEBY3yemyR3A3DqKy55gJrr80
OpxU7TnaElV0H+zDzeapAAXDjE/ytPMeurZ1Q8REvGHBEbz96ov39YFMw/flEUfrUmlD7lmhSrO5
CJ6+82h8Eysjgpk5veDC3halPR0bH6oPmcBdb42bgvib2LpolWyYwjPymlbY5o9uEuhYox6s7xIm
F0+NO9DDKHRV7dFHq1lpk3edWmEi7/y8qGoAlkYqxLvazHxxc7OJY4gOxsV/udugIHMFWJikbZKw
bmeQ6sRSjuamapCxu7/ERktordqE+5wxHf3Ur16S1MY1D0x7lejJguIZ+3C6wdJz7IW8lCbvIKk2
J9liAZLGHab9xwJ9Lqsf79nM8Vwxcvo7F/qLA+Hqm+Uym2CXnL1B6RYvUi4SpydvhDAMnkJ2hAkL
PJxforiQBVFovXtr5d+8S8e3zgkp3SLEZaH+m0gf9/6OzS81aiGFvbPSU1vtBoyWvZ+Gl2Hy0qUA
IJJvqRFSQBZGrsDvxxRnx2AcyvQNexhtcevmS5cBb5DIH18/Nxo8i4CHUUdY+3spXXTMSDc/Dfc6
UUjMc/rcmFFgkpjp69aqemNkh1bmiDkCUCoJHeU6p+uf0WHGo0qtGDdAanDOeIoDuVqxZ/vqQEer
BIwaNrWVFgvtnol5chIpcgRj418G36gS6vyoTDPtF6YLxdS6+5FowyJ8A8JAezFf9LvUYDyR+qUn
3jq5/8TMOuLn1MWqWW1YOFbRMSLEqLYTESVEZEoghGAPNWwnWWRNkwiIJcbNG++F0trqsFQW4myR
Wpm01W7Y5boHK0UqDyNyGumHq8/lkbAURpvyyzCk2LUT4oE8Vi/pRyZaX1WV2StpnhdQZMjuFvoT
xXckgjXKCN5TElk+yjuqKWkJVhdX3ogMfKEo6Wq7jZF2stXgJhYYviTdKljSh+kWTPV8fm4YFlnQ
JIeKLpKQAOGxIWOigKuJSxTQgIVLFU7NxN24w7HfTBGoOP2z/E0t1UKwP71z0Jf8HRkBVVC688e8
QNq0Wg0aVRp4dh9PfJU45TuGy/FYfE9lgCburF/B++U4H9ULBHfMjPoQntNiDOMgjqedEPDrsq2W
EhxluKYSn1TbTgX7l0To8OCOTdQxxDOEmn2n49fdhG5gau6LRuukW8HPfUh5KmHdlJt4K7sZGX8n
dgw6zzGiGZb6MW1lFNYGKjgKn7o2lb/K8k+29tv4gT3/cP1d6EvuO56tqTxgMIhTodKJP1s3yqoG
CPqmRKY0QTrAr3niKiuzEl1qFPrRY/HrCbvo565dvDnrdRih/Es1QlwB0ESiQUzbxYasZNMOIdb7
0FlUweUfpdAlSZ6EBhaFo8ZPJgVhUmh2vGfTbQ5okJUttUJAEczaSfO9jylOWp6lWPjgQH2nCu2v
Vg4g+OE63ZhWkXWH3US6i6FEHYKyNEVScGuZpi76AjpI9II58YEtUwBnLrM6LjgFa2NfBXvtokME
oPkwIhD/4PAdq/HN2BLjUrcacIvkOCL5aJQfwE6R0C8JpUxLKWq+J5960MUJXkqDvbMiJDzgE1WT
Iih2tmL6++DxoLqtZg+tvekGuvEuKwTCkYecES5jImIvViHBp/pMpGH3rmfQdcjjwvxkjTMV/NON
mSlNdNUqfcRfpQw607pDjw/Sa27x2CMIG9FMB15q3SReU0Pppka0YZyhBKbo2DpmXXcbcE9h2g1g
E9pAOBdZ5SY6fT8+aKrrW90Z6RdR0JFpHNonKL37ZNYbsSvYtxsfMiusgbi/CUcqlAkNd+q2DTDC
fl6XflniBYH+mda+jOkXxZTiELl/Pj/4+P08AFKI4OtZ5IZ8nNdw45bJqyFfWBk68RkqbWjIZEc+
eQ39/TNEmxZo35ft/mue1Eu1ZRvvyJhMG3xF2opDwK0eeKwPUPBeulelXFFEtmcu6qc80bmOxl2r
dJPyRKtB/1s9pIJSbafAWTz60ulswcN7lmMeMu0Fq3Bc/M8Af0ahTB55DyX3MfF9zHRsYlRSlgjE
w48frAUWsG+Kl7e4jxjBD73wWL0ednpQLpMCLJDdaPkNVT6sjLdHTsy+gKAZalTc5CHhnihM2ewe
FGUpAQVpTQHU+94ogZngQRLi+mgCAM69fw7PPWR+KJRLNLfqL0hNxRqAEVwRRrYSA3wdoE/oUz9H
ofaPZt4NMo9RcCt7FxUziVRgxFkk/xV1XqG61ouDO3QcJl5IIzWwbvu5ctOaOgKwOaqM6avZ5X3e
KwJFKv17q8cndMTHGzoGn61jp1lHO00g8HeYvOECVFG0cdH5qNmnbHvhHXo8TSvRFo9E6U/vm6U+
oaxaJKRa+jLPwvnb+VyHec59gziBUZ4T6uok+FpZh8Njjzeg351CnKBib4bKcHYPdPrjE9V89Can
8iBMDRWYb3aTl3B+1a8l2c7hpQxD0KOWBZBlQGH4q3/7vJpOIjmB02D7MLn2WESAFw+iBURHcet8
m7ASsvqT6vsAs0K86Tns84D7PqSXTT6odnAA4zoBUQ6Az8E5LawiCWYP68W0T+KcAcHx9mDJ2V6A
fEps30clablnuy34TCgho4j/UrRmnLWZ/7v6bqAdSCUcC6eJU9J2uov6vCTg9mzbxG66ocQzkwm9
NBlDayoFk1dIlQ7OGYDJURx6nz3HHMWwqlmWLxvZ1YBbb68kYP0gt3Jfs0EZ/YRcD6/A3fq/Gfam
JM9arILpDLSqPCDNpKJg2vcvFt8YitcNdPX6cCWTIhG/zM1b9cAx80tq05Ctee/aw+q8uV/HNQrp
jgSBpDdfPfAyUpgdwMaaGXZBo9WipNt0joVOs/VyBdAaay1Y/jfaEr6/1Sd+t2GJq2pOai0A8E62
FcW7SvDoS1ZGuJX0K1sqI4zKHDAVPFBHQPBVI7vv8Wjna9G9Jy66UAhWT1TyO8ygoiQBz/j86EL4
GRQHE8ORD84G8WKBMaBD12ybqnSB4vNm9+c4ZwCv1S2dJ6lm4AcAm+2LvJJcEZ0KKjQ68hv37aa+
3Nu7eaRtc0oLi42XvRzCPkQjT+PsgG/6Ej5GfF1quskjgbjOrvLrZ1t+zV1rEnYqJ5D7uCy3m3DR
DtLfYZFNqeh3sSNdBDrgSqoBY0DOFDUegETWBw/R4T3T+vFXJwjXZlywgfCpQJTItGrSkW9ZYBpd
CuXfX4KR544dwz0uw7xDt93XGQviso2PYgY6OoOpyG1RCgvfDuFsaYKuhVkwqgvHBT9u8FEb1T2+
JoUWBoBLY+54EdP7pVeHR9DTpbZQSNo7DWRxYV5H0QWwsTwRlhYiq0XpoPmBOfKod9Qyt+bJZKj4
XDolZVNyzAlgk3rsz5xGm4yIHDrxdZ3ZKPfMN0hhk7WYEwDy9PLhX4uJUFEkiM0M6iP2Sub5mFdj
i1XdbyMwzx5AB2dxBD4BJaM6m/9S2wQGhpd4jI+v79ekgRs67L5yCxKKwrpQme4q0XdNA75sq3UF
8uhMAWPNoE4B9z31QGeix0Dx1tnvWJ+RnWADP9Fqe4XzLpDhs1wW4RIO/sX8rHjdAlob043951QG
vaGeTGuP4bqWLxXWf3T/B4tJ/FdP63QpgfQ2c8bdg+ncH/2vIigwy874pXDZ6BwHgK1ZHkEc9PMw
dCj5UGolPZsxIfa1jtu0j6jpJr86mRznuIm3/elLNkjxb78vDEtQnLoh174x804AxtAMPKuGodYY
rqANnrmXDJ/VzOf97xfDmvCXGIYAsaW1m7f4RSZPoROQ0QU1Rxa9xFxvx2Fh78crftQ4oDBkGVQx
rou6S7yuLfeRBSFpCa4TWW2WWvPO2ytG77nf8HSrh/VffPEP9dPLlQmLBpIlCZMnds3bz0vU8hvc
vCR9SxRBHQLq5K2VhcP+TUh4y9Ikx6sQaq6kmA+34sFrby3lQrJHDOu6EPeLRPEzkxbg6zqYPrH2
efTO1lXWWyVhh+bLULBa0twNfSr+hPDiHAeQH7cjOBauRM42nRp3n0URLXIAKknY3mSg3InnaOj4
zqqb0ifaHRDEzjPtpMLjfmVv0LhJ916orPWZs8nEqyx5Qv75/wnaM/HXLt25VN+RGj+YwEAM671P
GcQG+SKmOQCcjKN8WaL90KlV+wkb6A6hZPUtKSbfedFc+RtpTXJqp1X+uqYB3GUqUonnQGF39NJ9
/MHfDiB5IADfb7mGfW6MQUuxRRPyqFnrJkzpcS/i7cFAENU9GRj39eDsTtgyG40weG73BjMBW3La
1c/a1eE26z5t5g0+uPYmroFu/aVloZ5akOa1skc8Y8+YBZ4L5X0OsGN0FfiCs1h6XAE68auZd4d1
yJtIq6ZLx5TXl34exEoTDC/oQhydqzhSE/h9wJWWWyZ4GuuVq97Sj28tZLR9hXvdelabNbVAzMQW
zfXN9wke6+5Xfb+9qkXrSc0KxYLk14X+vIoo9/BXD+TPajM2SgUxleu3N07kgWru/8BO6w65FrYS
S0GT3pJGigK3YixBkHw/afYq040omX7GvR0xejt7iR/0c9gehd7e2Gvic+vEI4q3zk0nOX0c0oo9
Nnl7oadLRiwNQAblcZk8gzEmIkpgrQgcn/F9+LtfV3sAOl3/FuV0MWhLojcNbivB1Lyzy3YzNkq4
YHYu5/2gmUt3WPeMxynIjDxrQe+H+235+KrRo0qXzNIvgITqClLHtay1B1rne/bhdRXZCh7tCZwO
K9FTnvGobZG9A3znmDY7PUbLyG8YjJldRmGx58J/+UHKbsGABm01+RNYI7aW76HcOwGi2k4GIJnn
/PrYYJGjLd+3sGeKdDs/uSX9HhWsH3Uga40d0lo4NWL32+kVzEz8DEK8Wff+7K0/skHSko4qqd+r
Ue9nr0mBFRi4iYvGhgkFvyddHzgReNU31iKosFrUvBmw0ucBPv7Vp4+jeqAoUqtb/DkVIHi07IhG
C4JUW7ISlg+hjSiwCLt59BuwFlRdX9MLeNR2Zf5yOfs0X34uZM5vjYCMEVHfwPX9NgnAD2U8Q6wX
VvDIV1EbRMk5N4Cq8Kcd2gE6YlEMrSh0dOqJTBUGhlu4I3NttvwyJd1dDWMMEJuBoyJFHAOm4i2E
AM3ccztsAXWCjUukgk4OYZLV6CSvyL9F4ZHgtf5HBE/jTnMfVv2sPcpjjSymLNXNBkgMxIfxtLMq
AbB9W27wYl4lK4LVmTOzh37KlMZmPQ1GDbsytDz7Nxoktcs9jk4/yZyF0Kfr/3yWXwWaPbA4y/mm
7PCVfPgm566YqdD8docPoMIopkx/3ovV4KDzi2UV8S5kchOMJcMfYnyAhTtX61YwZsxv2AE4/yMU
2y0mEq5HDNb0UKKKOlobp4THsa/k0pKUBYZf5qAt+pmW2zQfgy/fSgkrLS3dGTEyf3ZTVv0K8qTM
aIMc3aHwC1+4x1wYxVs5mYLY3yFblQy3R4rRYKWMyXD2WH0s6DNv2BbipLpwSNNnJe0saVexUAbK
N9VxhEtxh4WT5iVj65eba1BvXbvoJOc2GT7JtSFCM0Wg7YMqIY1M5q742XRC89nqHI1T54gKnfLX
6aVU8jm4Ceh0m/1YYMbA0GiUIIOExZrnLAP0wL2a/y2S/9MJDtaDd31Q/Rztn0TE0aFA5o4+cRbR
WLmM+JspL2NAVrxxKeGo303Wx5XV0DEPhCIb5Lc5yUJ6I2DWX48o3bTzHubHW2yuDtKJ/fSqPc9v
rgOVFJLpy3hrdg/DOE/F++d19wHn838E1S4jxmQ+3RPt7CLGd+D85WhFF75Zp8cBuq1n6WxRBaTf
AA7nm1ZzlfKrb1WON9TeflPUIWfMUcH1jbTJd6kPCDsRgYLY27rH1rgYPCkiMt9wP9CT6VNeElBy
gTAUvX84l9vvaj+zxgbs1K73EomRhHtiLzQl4gPz4g5R10QE+EkDvP+NJ1YJKvGqktBwqg+yhmO0
XMUj6XaMfmZ2UhRbDmn1g7GYt5C4RiA1m/S0VlVOtZTkO+lG4MsdVS8UpMOjDFBFHwvCLUYszeG5
SOTO/uRHbTa+kzkrLdPLFbift2n4zaBkTa3HFj/BBjxpV8q0cBSxLRmX8x5ehQQCeN6vCo05XQ88
HRMvTsm9ekQkbGsbXRB4K5wS5pxfD9NIC776bhAswHSck/PV6nsoK/OF2R6pfX9Ndc+9RJ9cVyW2
A9GCpkCgIBDR6iffUHIBWvY7xHqYe0SrnxP9dqtT84xBCqtlG/6HpbqakF8aXRLLqHN9voCNkA4W
UoMGr+OTrb8u5Rg5WJOXcBUsQYa/QUAZYarBiQREeUI66W/t+mhqLdib9MtlDZuTnWaKZ6NbaLAm
BcMUZTgyjpwMcPxuv3UbXK4K6jwLFs1a6K/JaJ8P/t79zLySoRY+chXogssBnGlcARqfcgV6S/Jr
8L1hRNQd3zNAesKFqJT74lFSJxwW/77o6Qe79H4LfuGM3wM8r2Yyku7RdEw7hcqk+6TCONfKOQVp
M/S3WBVDyx6veqPArXKMhHg2Rt0k7NGx0nbCbjUk0SPuMM7YYvqGu1Z1HRxm6iNYswopgxgDU7tN
XpbTmZSjlPCsakiMkBJ+/Lb7wJpJ9UboPtyohgVithYUuDcUqxTpmZ42lxUT7fSw1AzD6iUkOXvy
3lLbhPA1veVkfWCUQzQdJJOuyytha6h2B3Cn0fADXRtOvA77sOVwxLglshCGKiIdn7lpTg8jTNo3
twrS/+IgcbWbDGM6+1bg1u0NdovXGeMRhyhtMt2UnHq2qRsHGDuOrWxQ4ZKsmpixKHDZLHRL9p60
sgBzFyT7XUayJqCk8LZ8oKYmr2dFdkxkq+zHiqALaY0J/wBDiB53aBu3HJG8Uct6tVSJ7Uy4Pwvk
kUTc/y1txPJIcHv5U264bgwmWFIfLhWFFDLPk4BJGHgQfscyujtyiClqWSnWXjuUZiJQm81DiEpp
9+0dF7jp2pib5UPx3MBlSeMjQE0OdFf239lp8672MGTrmnEk36MeY68StXZI71H0xtZYzGFL77KV
e/pT7x/Emp5ZlsKPbkSjOJAxgKnpfwRWg7yM80o86uBTmMSzd8LjlOjgpCd0gcF8aGgYMQSiOF9q
8jFGlj8pS7HMjFq2ocKhVfntsha5l0Lbonwa17Bfw11QiCKnRyPkfQFqgUJHYqSlQ3EDJtxdbSRL
Rz3uyqixNQdpCWJrZ6j8WiDd3O9W3VHnwB/rf5+kQ2zsrR5nWM5CcF5fx4ujVmnMygfbtIbTuJT6
ySFM0dv4YNpxUS2O4NUOxcGpqwO1FqaPZP2icV7NGdd6N3pWM9Ve7+0EoPoX/VRRDUnKcntp3o3h
2jgX3jFpJQNPromrQgperaKePHnbStjUPA3rn96Ne5vq8kbQ5U3+d661vSX55MpImfgcD05nA5ez
+cfsYnjRHvypH7qH8JVhF7xY9jZE2ALyrH0mJVSOORKeDcBw+CBwPTTGCaFjhA0yJ8oSTxJTnJNP
FP/74Bq7te6Mh7nVMqAcTKDTEuR51gusVPptwjyofQvbxvjbbjivXLIEM4N4XFN84Ex9COvDEBGi
AkEEe8COafJYM39HOQXp73FSxbBHikY5VO6twOOO5haB+J2MQ6tpLJ1rYG3JJSiTGBK7EJmr57Er
/Wcb2udyVBe1XZ3brhkiTw3yxj1TLNBJLQkuMOSI5Anf5yaczHrESyzLDUBHP50bB8NrTlbk0+FS
kM3AFaCQbrKuYJxYMH86/i6dlXU3E8eYvTZC4L2nnL4FnZxtLWBDPjaCSU8jJ/rEzUvhuMtqeLxF
Q0s0b2DVMebSW9lj93rW8GWVKL7hQOEGBpsATt3fiVOYd6Itb08O9tQ/aKQwpN06zhEsO85TTHZD
GRlfF++LCYr7HhG7hVKLPy/dB//MjDy9rup4pw8tjgp5fHFgFj8f0ALVkGgGQPv09fmfXci41f2h
Hws1PBlxxHclhGLlw6u3jLeHD2uRH0N92zyLT7fARCpbVqLcvGvJBt/5qkAl8ozFvDPEYrky+7G1
v5hprSnSZrLcA1MX3jcASvHuEZUcMTbo5j2mu8joyNGO4gvr4bY2hJ9+ryBzj78Fe54Y76zzcUuM
rSAST7bEkHA7/HvDvPh1PnsurFjIqxTVSK+fTP+IRnxCTSdAmiFRHCL69SugY65ACPQ7Ump41sTT
5VGFzguvKsr7N5Z1L7NYUtN9j/4jOdCtWyfoQ9LwyCOkmx8sqLT6CAI7DcmHxccqrBf+94KZ2LKh
kM0JVZFxOa1uYE5YtHmUvjTQkGVmZOPdnGTVV186SSVqrCJYs6N7TBvU3rI4g9ek2SuRkgseCwcH
9FRlZnTwlTiOuJyArTfY/irpo/TWgFxTNfQU0tPiqkigAKtRn6lMEIFPzT5xIUEwLyKsZZ/teuw/
LimOC8vLt/j6ehMe2dh5Eqd4+NyWUzB9b7knD9iUXcQn9BIJfaGURxI2vWeQPjHTRC38H6aC8jbH
UQfQYLscNgdr/7pHw56ZQMXjYQAkkbEkzXaHed6A4LTX2sZwxhW5HQDWDGD1gFBCBltVwl4Zmirg
Y1KcWzIf8vkmr9aQuTIUpAabf2jqsOWgFFE91IYYmrbz3A15Vygl8VaH54bOZj4BdhuYH6v64txm
j4pROqpHYOW0SIN4gjWYl3pFpoS9xPiAenv90f2dXY4OED9n5tq8vawKNGpxJcmH5iz95z+si5k+
mzsTiAa+5C7OzjOAHjwYgnFPnUhNXM/jNVXhjO5fJ8HorIhilCJuJQ18VLTYm+abO2WqtP57zQna
4cNgTQ6MQJh1z7a7YGcs7MqbkdIaNuI677h1NtVaXx592As8Vtd7nfkZKUW+lZij159IARLXqhgh
bt42da+20VgNUfm7HgqtJytcBFsZ/lTEDiVOryL5SUBQMcIOdc+uioErxpWZZtpuW3QSRQCZREWR
esbSv8BN8mykzwz5qVIPAUGWaMLy3YXlVNczV+H/Vys4g6qVy+qpWnpv1PRXfzI+MBsnfbBnF9Iv
0FhjQC8JQKk3b5jPVTjyI23oSmWwtxxb7H6l6m3XK5oizeBWuNSRC4P/oZwkn3nMSR4xBync3j4S
9QVwu0fZhUoBLUXVWzszzfx30kWiLbpH5TvpfRUtQD7jxc3DLlKwU8OlfLfjcWr+8qSCHWS2IBB/
wSd0he+/lmNGY4Awy/e1bDRkZgp+9YTMvtaJInv9z47umIcEH0oHfUohun2nfVfJs4haIpuh3h4w
Z/iMAyTDMyDXOGxS2eEFYhdPevpsgsZlgavw+H2ZbXSlxUv9Oog17wU0L44xCWtVfhVzEHDoE0Xu
W55Eum2X7HtduRKrb1RCFm6OQgX1I3gwo4UuhrwTLrZogfrKLLbU6dGYEPU71GjhB5lpetDbvReg
auPS4VTEuzAf2XNGYdmxGDXBf/T2jejxfQTVyHImPel2Tgm20t+Sz5bxYlikoFhUakNR1WWJC/55
LaBuhJTezmu1QjDNKqgciziwA8D08cBz88L8n7yXcMMMFP7EApQUac0AxVqZtFb3hFmLN4w7fOAQ
ZvBQ+PXz0lJuU37wmGKwiMWw+7gJGBlqtC4jA7Ix5eWroYb64cotN2b/kKRFCuCb1Fv9PQFJe4CN
lWMMJBjE2dmdW47OkwjDltKadhIj7VOyW3vK40sAN2DsD2thbYllIIKPGGiA1y6pRPG+OF19ROMJ
Oh877bunSL6TOXX1u1xTSj6gS6W8r0Ezk5XiLPfA8c93OEUcqLlKEl1mz1P3C6ZKsGlZ+xLkEnFu
p99UCnJd5fexIQiGvRy7PBD3IEGCkFt7xO2yoDe9qLo+/I1QW6gM7ZxEO9+ZdfL4Qzb44MndJx+i
zmv9861WPs5scI9BfLX5ajUArovaqA2KXFokl1BTzbfDoZpbOruGFtyPWh38Ys67X1b/fjflX2Yd
gapt6OErX8opoqpBtRmOhkEfyyEp5pJ420284oq0t4D10veGE8tY+CtAlgtFYryflfymQ0KmH7Ac
VVpqlCA16ChKEDjDW6HACDB1aqqHeLVXruH/qv9pT3LdN5jx//L8lPn4QNGa8VLLJT/J9hFURbF5
9WC7/1qRIyRNxDg/PXirlfZDkQqnxGip4pguMAL/W7BX4M8NQlvnB9n23Jg/PEo9ndyrDL3ATUAm
v5pb+VTBw+uBBMEmBDVIQov+DmfV/BfUBN8TmZ7THW1fcP5Rxse783pMNy+t+MtWXjo0fnhw8bch
06g+fJvfOEnL2hlufZdtICrg+61KbRfwOy4FnkC8zd05IW/bYCkGEV8vE84Rnzf2wZKJaI/5Kioo
THM1EwKEORAcpI0VeBcrEVH0wdzdXhlVsovvAjpFSbV+Ut8GtxVgG3xtV4HUaAvDj1+vmkT/9kYG
5hTAG5Hgm8Am9dBcFUv/1qEMToMTY9kCV/kTfzxopz7WDbJW+ZrUj+So8hZq8724nCqSad0SmM3F
bJD9jY+kiGPXImsHZZG0zg1kdbMYzOMnFimE/QAD+KlmOSOAXWzKZDQxcrGi2n0QYH2RIRLuDX8f
8KRi4Uf4rbOnreLrDuNmjjsirdVW02SHlwtSq8btIbJA7Vj+qzdsoZQdFEyhVbfxrJyQvtn/cdmY
AN+6VY7lT4rR2toQBU/2HhMtesS5fVtZGzkwWSxe3arwGqKTPW3qaGszobqvmDF5rHG7kjlB1W9G
2CAto3I+7Pb/dO1yJBXRKxh2284xvY7hlThkAGQIijpuHhufRbiX5k3ThoznEqScnwBTCo+aFHX1
lF6Lue6GX5VvJkh1GC0ifJeEFr7ix3WjphepyJSI+utuB7Idr0KdbhVE8JDaYB+uSNeA9RoHPyXZ
6KM5/NMn+aTCafYkwMfmZ+wk5kKIGQuPC0UxH3IHVOkSCtTn1XGgH3k1G6FT6QISodhqylySu1Gi
l8R1V+u+n0hzIbW3hRT3c2BgUXvMrJxh5XEOMwWU9eG+PhKG+s5B0269FzqQNk/0PPsQjJqJKAw8
PAsnya1wZbY+2fHN4u5LBE+89VIcJacMMwWXfecgYCPeejYVrrygbIVbOJkU9Gs8VyvC7SpGxvdy
uDVqnVPjarA9eW/aD6LJFiQHaKDcDhc+fMwZLkyGWb2/EH+S8+vG13VqaLmZl9UvGOjDk1UBFMxW
IHN2+tmg97ADhKb2IhSuZZG8M3QTNx8j3+Ex/oJQz/I01jgyR/HyPstLS0Ngk/5faH3RSIjHk73q
VLDqt55wxpBTrPGpCvLpl732gO7cgxMOoWG+ztFhCaJScJCSAvDic6nqfyAoptWDtwYX/b42wNIb
03SBToxL6cC+2nrWDQISt81EDuRKAUIVP+YNba5lqhQtKhB8H11qqFvEf0Jjq4SDk3rMamB6VXdn
A6RDmThS9wCpIqVfmzkj62SpaaPPFmfKix+51zqiUlupjT7j/ITofFibP5oxD+x1PhNbPt3RiEA3
N0bU//ELQtPFUSQUjX/eRZz9J17y5awqWjl/ybtxW6yREc3DusYkHLJBCl+qi45uAfJEm+TEv2I5
qryKW6BoPLlgPsXe4IK0A9kS6quLy4Dk12NLKIH65Kn3IDr+gil4ZL7LZIbOH3ne9T9gK3wnlgh4
WwJgwbOvPj634RJpr6IMHYz/zZWrnT5iTX54BNY/8TG/Psd8NqNs2h7RfK0b2qRxNeBnUugvINiY
1q+jijMyVm7r/jel4ddII9DNrp9hdpXGYjaVrdequsGlMuxZqUz/egC915ACA7TtLdDAX0k6kS4a
sY4taG1rNFCBkCTAWnp6hioeq05WDWYypaSKRExsGgub0zTSi0lnjYq15njYawZolXb/4ipS3jKO
0u+5TNIrU/9qgLNwBaAF2m4aqRTcKEKVvGhNyJf8BXXUidErJ29UVQqyY/EoEaF+OTRVOQvu9Js5
Cn5FVBivB+U20zk4rfil7BNY38xnj9zv5SIwVJaOij8D/9GCSu6ajzdsJqI1ewis0QG9iZnMnky4
zI4KUmeSB0sbt7weuu1joHIuKIh8VdFyDSTEMJEBKvd5Bfp0lT1/rw8xoZxlTi4oxoM6k/jdwKa2
FWuTB8vo5CwXrsJ6cf6kUmCPQ/8HROzHRioJizVBasd9SI7vttqFDagTSuZFobs7KXGY8uXynqml
CeNUcpCz8gid7vl+SfifMh34pW31XpkfF8gJgcoqk4WK0HUIan25uahKNjsb6AeIShD+ZuGcnG3f
FjevsHSsyjRxlFIwn6vqV/EewI+6NIlSuzBMctxHy+U1U8jqp7nNbD/2oYtBulM9TSpDZSg1WAjt
3fVwGpxQ5ce6nTEjrvZj+xoVVyN8/x4skcVB5AgjO3rKtrxZng9J4JkcqsQqvy/dj3iswpp+JvEy
lVCCy36mMbxKRoQxfrMrwYtyBbcqH5EQkmnqrOu6TVm4/L+LwxC3KZKihZfjattzDAeeEzHhoV33
FTXqWU5nXGdL8aDQPuj6eObCjohPF2DYAhLEQV17VOej53Xb3Ir1i12faARD/zf6kTjO2IFDBdur
MS8qKq2+E7A60v6t9kl0Cn+k00UM5uxjKYTvAdoyk4XLCBdH1O8FlMaRfcFMfhDPee1zGUJeKaMT
jOJfnbZ8eG++mn86PiF/X5z01RZx3BYU3jkPDe+GbdKXC1C/a5PUllPDdO+JdLfFeSEf9gqeF2h5
JDVloM13HE6xuOaW0oznFB25qkYO65zcxkKv/w2l+bGVdDVXF0tbzz3nB+E7HL8KxoLpszbOsdSH
jvQe43oL8rIymI50HD+lvtlcqgEtBNMFl81dHJ3AZkD5W/ALBeLa+TpEb6zySccZx/hY0bHDvqQT
3sqV9YTGBAcBg56l4hebsHj7SJ8mR9Sp1eJ+2F8MVu8AEE8KOEMrdxPL3OkzwcbE+OgMeudKQnjR
Ug75BLQ605lIiEi2tjBSRAlCEGRaYLE9bsDbH60uRzCY7WQYK0WA7S8Gi972XxFc6YukWDvFObgr
JSuNRTPQJvCHXelJpQuUBaa/7y7aOq9bwoFrIQfGLmBM6W85X+NmiENBfnEF72v3W5Xfxrrr4VMH
UXyYwJppurNVIbB/0NXGCksuUTYz3LyjTFubjXCDDA1jLqoNGi/P08bZM+rluw+tNukMw3F3p8cF
kdaAa8goakicVb2sJM9su/hmvhx0mnXmNSLTNF0Go0OpWUpvH61HxHLx4n6+JlogeqAXZhX3qUqP
A+hMhxLosulLLfyds6N9tyz84I7qAMSQG/KGb96IfnDrGYD7JeknXnppGMeyqUtwyz793Bx9t1Yy
kkPBcKLar869wqaldUlXQqmIYRDEN2SDSCLoyggySipZOUtd16BViIKwXp/df5eGaZeZcIg+8+Vg
jXrXsNSDQQxNCkz7yi7P4Ye48+qlR/o4FmeA7NuPsYoP1jwfWrmD5HHOw+EzJkqR0jfB9KWWBan2
7IHHn3gi2ly7RJuu6uGUZN06JPxtO6reKvt2kzySXiHt2pgh3PAczJfILbpkVkXsQU6YtDmGQHgq
LeubNBezdwlhJkU0kcFY3vHSq30UEq6XGgvLtfnmuLZNLPmWcIgM6fN/espBYaESDBWx9PMWVg2s
mXdfQiDFhezxmVvyhdJyivE3oDEsd8T9az+Heuz0vBm9VGYCSoolG1BQL4RuQXaTP5MCtwUsKFsi
6G0v/u0hBoAS6kYMwLoFBj87G5d1X3KvxDbwSkfEdFn/WHj/4uCxxG8YMASkk0yxEb+JTTqNZFW+
5aHwp3xPu07UgH5pmftzorNZZCTWAlSAfJ3qhiPEavor+GydNvXE7laTX0jpwY1LhiS9aFSIdyd4
oHdc3ulr14OkwJbBogGOjBl5DFJjKUrA3UjdIlq0EM/32bTp99Z7u8QkGAaMKm4SL+3TJxDO1f+7
fWoze648aMZn+PAQtVHBJtO+Xns2nbF4V671gUg2Cog+IVwtmqQBU2QXZD6Kwi1SnrAqLHGnznKK
u/KJ06/8HcXm7RP/sb2+ut0VkiFr7RRGzehzFsNiOgQ0HkWk9v9JQpBZHRHXuNZ0xmnBCELPVlIa
g81kc7zjrBg3CB7lh5RTN/kGRBGoD6YuOJKk5iBIMoLeekJalcsCVLt3Tbs7yvpVJaE9FSmfVxiz
wRZ5n0ZIFupELqRFLIQit+SlfoyjoSuaII+KInS1Pj9cEzcs0myr5XgavpbojTA/SAbqeMIRYmwM
Ok5+5Im3CM9yQhYIlu52Qwux6iKDa7jNwfR7d4OrAnkPCBkNJRqfq21dsqYSJbAkepm89IOxJqlQ
aW8JY/q52T4PsjMPWCNDwVNsE+7GfY8qCfLOZSv++CMmkR25OdrmdI4kZJJFAdp51Pok9KY9l/LN
bqEyRn3S9KfBLKsv438kG6XKQKfGRT1M0fCRlLdVhgBRgHkHK07sBpchS0iWeKrTgro60QQlCVSb
MPj1QTVtQpQ9qHP8aSBcxO6lN20z4W4XtYpBm0ipADO5/aXaktyW0TOH8hNVY+8qhpWvt7yvYXgJ
zjFVllbDYxDwcIE//Ldu5xJBIX1rLQL/S23W9GE8gQDo3U7K/QEAlKb/snB6a7YPkicJLdBP2ANG
gM7166T6an5KVdVSmnpyL1edBR7NzO+OPVeEkUc5TbrQVFyXO0S2Umod8zQJrFC4SjUpuy8UZCZw
Q2sofDk+HcF+sJVNP+SiyJ0QxZ7HRQpaMzgAcniJ+XXE83IVc68SWWESodN5OKxghn8vgiN68XPD
MIYVZFAJxXORaOFmDbKqrIqO7vYpmh4+EL+5C7pGcn/RxVmKICl3EnkIv7RVNvh/NDmQXgnNC0FT
4lydEuN370161gZT+e0C6HdIkTQcLklCX++NzM/NXWZF9h1wWmlOQeKDl17Sc+akHAL06AR9v9Rn
Iwihg5OcBW0MWeBGNdfsppd7z8PDWaG6vZ1RbZUPGVVkFo6VgHsH0ZB1iFN8TtGl9vyBPt9G+jas
GgmOHX5Q+b9CU6bw4ZaCJEwjvePovy52Vd4Q1VKYgqA9dFDsh0oYKDKrXmB8Pga1iG+Xq4pnnkGC
NIV2GASZqapWecUi4//x7GJPiy5kps2KfxLbJBrrXH1baxzVBl7AVT+udPvGEc3r0LdZUhYAawJt
XPw/5nIAgM60hmlzeysd4QjiGAL3tGCvMFogO7nbAgB16OSxOviq4wj9sRQlVVoXMfYqZq39wNEB
2IZ2snY+HCvScBp2SjBacfLa/jy9oprJYyFrTa69t/fzUkc77O65ud9pBIsZpkXNdJhyeuVqYlwL
nQBRfyHzItsODPntF3qFYIvpIDOXak5Zr0uyT14tZxga3f45u5fFs8lXiWpfD12itd12LyU3Vo+L
JOAR1mUB8D5Sdi/TnN8z+kPp2l1RfLD7uywFHqpYSv4v7DaDjnWdJ1jwN5jMkECEG4dJK1Yh7Z0+
DDA6C2x9kBpbDrrwZyRmarDZmXy2sWkxrGWrm4Osk5Y1357p+xKpkBI7+A2ngshxu/qiUtfYKw0j
RhhlbEBtvDKwvDKmH04OrERJBO0Kyo0sjaYUa9027X1rWc0vTNfic34isfxrgXJbGspkfC8YbfbC
0OqKsCysvFJqnb49TBTtp1HWBK8yhGF729SPDKsJPiQJaMLUjbc2KY7jEmjH3aAlhCLc+GgFrqaE
WvBeHXj1eOInJ89+u4R76jtZRb8l8Q5uejpsv3mA/xIQ7ZysFM3ylfKUHXx7OU+ecQ5UTE/828yl
0kb+vMCYx7xly759mwvXqwvm3y22r+qxRVaegf+U/bk/VQseP5cJKCebcTj7D4yLjlthEOaF/fLB
/ydk2M7G4tpSn/UACPCHuXevrlZGdRbb0Qf5QhXV7VI9t1rRNC+szI6BP/N50AKU40E+8LPE5xIc
rsS61Tx2TlTaRogNETU7zOmBBFlB/Y3sPI8bAEAZJOHhV9xZSU5eANAT6E9Gb+yhBbZTbNIpOhls
0xGze0k92YwukcypnBEbceCk8p/8RKfaTYZF9Hn4py9cImzQ1G7Kp9tvTRwZneKX/K7UT1Gvn2ax
EmRxOQVIROidkARYBx0ELEjP40DieNjfTP6qHIoLn44+IOTt/jUqzDwNvB0Z7QaJS35BZOjh4gj0
ZIghywNSBKrwE8DXAwKU/WsHeMkt0qSBPyo30MG2Gc7SnSnpxPQ2p1asMEdJdJhX6EOMQEEHaiB3
i0F63aWgOCUG++KkMjsxLO2rqTHc3nVqIbn2w5eAh2chDSoufLCIZAlhEyBjTYyFZ9nwmZyUqYhB
8inh8jml9UZUkMlfCeJqFyeQD0ChAlBvHbGT9hyqFC9aG1Oza8aKlAb7wcKjtUHH6i38QORts7z8
oyRpOajshBPUmcVGNMma3v78VrfvxBKqpUhteirGzBAZ/NbZUxxJjBW+V1I1MEbgFjYeY31H6wfF
EVODbP9ptVxeF+fGgdVfmI02ZuBNUCGxW2cGMy0Nfs2oi3N1Azhsvxcnr4t+D2sVEfx9xTy/7xpL
9x0YT+T7I8+v9XK7nteOSfLIjV/qRcK5zV3Q1syKWt/94WOXiwjhZI9Jxz+NjVJdroTvYc8GCwi5
lwintyxgjWhAgXhosFGadzIqi3rKGdZAkzuDN8z2tktvuIkBYgP+mzs9rqnCR3bWGpgHFyQpIsr2
zchJI/9LukaXmBGvcIQN8Iy6/d3iZ8bJ1vFadajolatTSo4KTVJMKx6Ip7yrCYw2Z/XnXebV/Jap
F5qSSGD7lTdDPhC6vUay3Dr89cf2IHAnGvVI4HHIL3tb3FZ+p1ncXkKN8hrA6xmirOIJckEj4j7T
BOiYzA/ba4dcHp5ImnSO4LTI9vTbKpF5ghuuDFRgFl4WuFvRrLK5FN9D+GfBeTVNdw7EUD+5Ba6q
a8pAezSAp1CD+rL8EOqZNB23/v21atJGF21In3QBZwwWIQLilGT7hHAbuAFeoM3MBcFkgxTJ/srG
F6Z/SPv3oP2um9DTSIfFpP1OCLQk+RobaLHRqt4hfG66N8As/Wqq7mUXJ7z9RFQfyCIxiBJUyk+U
RMjp9YNkBGnNAi/kWXLNjc+exeN8lZWyRbZ5RAl6rrct/cAILjJegKRpb8LqXpu32cenAFaeqhPS
s+QKI/hh8KaKQGMl/KKMYEhf3RUZV6IBJs/q1cJW5lR2ixyTQvT/2bVR9B37DnuDXe8cqEO4dZA8
R93PLwC5vJDbfU+nerFJfHYI664xaX/uzh4DO8BZFAvUQxLUUT1U6qE4QA5GJk84ds9IKpnAIoKa
JDPTLsJy/aA54hk7DxxGD9D8Xv6uOOnPhF005CXRjOsleT/Q+NppAX8RLLSTuYvZzhpyQBJF61fu
K9KIYjz1oFRcDTbfY3fDAwVTuvuS7HTN2OSXhR9wA7MJvKprQMKLbJRaPoVvIgesK+bmEniv+wTQ
+iGpM+vK4sAnfCqI00G0F6vSx5bkCuLuA5eqrdtj5FRUUjXyP0jpf3X3IzcWAonzBU1H325yRA8U
UrHZC8fRQYSgyaGuEBfjcEo0S+9hi4Gi7OWafU6SAudfGCifkSJXSr2RgHo3j8IrZBZPV8VKJ6QX
PhaTGVhg+wpzW8ozBvh0SQLqBRh3Qv3IF7L9TN9Wbzy+qMJmxAoDwSmviVKgM93vOnOoYblHYZwi
fX+0e/DqG7sJM3VZYyDEvCsh2PjrW8DJHeAoOLO2p6yj5SPG8Vi/Sogk2zjkOCHQoKqFD8q6HQm1
PChI060t7TtqfGGgdlsj0r82Yy3dNCcaVD4LaPSk/eIxbcluR/GknQ6yYlw0dkwyYjBoHWJKikwW
Jsu1KQA3Erxm3uHFooLfesgxaAmyKMiu/8kgHEQyzQ4kcd0NXeKrhNqL6FpRbwcF0iXbDUJ2iyQ+
HDUKVTr4TVw521o0Z2hMI+SeBhYTQr3HO/e3sPa7ue94U0a7iK2Hl6AnfDPXkuxxaShG77w8o9WO
p0yRNh2bnid4M44jarMdyV6p/yLYcqZl2yMgvUuZ91HiLoDYJmknTArBwE+F61lbmkchH1fOK7O2
nZrkZwn43K3MmlN7HH9DuOq/4zzk5/D5wm25Nmb/yGq+QcjmJ0NzSmcioRsjB2Ht9hX0NeiVFa3S
FsaZYn9ENHYEHQHVclzRUXkS5os4QUlh93pv3BZqoRmjTe5ZjBhgfW3V2JB5/vBSz2U8Soy5Axa+
kXjm0WWbXSxvtqqVx4MKnGDQwfPR4epkoAxT1f7g8muF1rhDkSX5b8zUqy9E3pu8xrmKICS7iueU
/qHAZu2hukU3HAS3eleVKOYR33wUjTmZT/2LLAGv7eFDgnQdgaNXyRBkDFQbUzaxoM1nkDwSVmuQ
0oQqAXhyhF2vNNJrw15WZcK/4bxa01iDC93Ri2eLeWtwbNFnOTJ/s6VPausbnrCiwsFZVpCcyQ2J
rRx+Y8uzg5f4YyOcrttXXKTGPWCTuI1LsIK00XjNZ7u6W+qIzWhXSe7R2OviIUAm7yAgzzP+JNkb
W2fr3bEVuNYiS7sIm9nPAOMNL3RY6BatUOupsBPVoeQ8TMxUCJkNSQRVC4PL3GzpywNS7/h4sS0F
x/hgpcwktfsMcIRBxEQDq29DAimybwvyibp/r9cdD2PvydK8ygHgMfojpEdtgqG5CZjXft8CMPjN
aa6JqaXBJ4W7OgMw6kgrpEw8kj6CFekQIB356n2szcXkE+LiXqqD5qdzjP4F/ufNZO7wLsXPQww8
Oe1/rLshgLqv1k2rRqRsh7fKg2hLJ2aCjLjO/7OZbXhJq34G+MB9sknLq4qE1zv7ZSi0gssMIAFk
wSY5wU2HESVwf91ZG6M2MxncxnIvFxLDq6EJwSng7ilQTONKv9+udJSfxYgQ85Q8zanmDES47b/O
pp1OVGlgiK1H/B46JHO9BXtcKWOrdU+bYmxZapSu/cDLKnNGQbfmKcLOuEFQ8xRAdWo+lg8swXLY
O7xvE+AJ8JAda0c0W11h42lsB7JtQA1K7uwaaWvY0owDjXIgo0QTwaYIt80zPmIKiv5CCxRMkgXv
eL779pXlKEgHhkiGpbljfVPIKPQQL3UTJZzZtNAPcP3NkD+YtohtzKKtzYsQfX82JXQ+G12LyLn/
s4DN1iQfMNaXmqGXhdYMrQnRMHQn4DpfTsqrR2fzq5F1e/gBP49Mbt/n+MCyMMo7ywuTbDtZF1R/
TI4Emdqsf7Cidnld0fgfkb7F4DVOAkbUTFWWv9qBKbtFl4kemPfVtyyfK4Cgh69qzMmcpZwgDbNo
mSGKn4daFYeqZ5aR9cB4oraqsIys82a2zBydF8la2sIaobVHfR1qxt/SSK2StgYB9utFI9auY/QR
JmMUEKyNjxHvjgYXOqEolbC3od2r+hGHXT6XQOJRAqVyJDr0HcueouvAgb/xAmJHnioIHhzfKr4u
ith4SiUnsGO9wCCea63nDcIP4NjRQoITeuO+RADteyhjSn+DY7mJjjlpNJOLaPFlcV78G+NBP41t
P0snuSbxhRedkOtTmTiX4TWZ3uZ3kFawGYKGBPWib0RDyXOHWNGzAWfLbKt+Bo9FApQ0X7c5d1O4
0qmA11+OKcMjfoAtW34mF83sJ6jVLxaEi0uEv7e51hMslIwCQ7dTJuPLlSG6BGfhNUED1rLIdWK3
OLXDkNGS4wDuE3AyVaxttpejQvwymYlmatw7QqQDY3eDoTmKmqUC3g4i62djx25dq+jrQ0oWW6pm
rLYB9qbm+1tNXa+aabT7/ncWyYfsQzopN9Bv1zQ6CCtwg4Cqohmn/bjy9NgXHfQTXlbALVxzEfY6
EdtQwul8aXtPQCJSyUEytbo+vhGwHCfsM6zJA6qFJm8YmfF/UGHRuWFYzIszyOyh2BzDFcKhmmBe
WNwftX9n10m4zViBHu9st8tkHwukwDozR10Zl4uQVj4euAtka1N81Z5mn3XAwuRVZfgETukapMbI
Szf+z3BoF9bEd0tNYZ8LeDVSYKU5hvSWYhA3e8c6zeSV5uwIi4BGdDsZq849qLwDO+38sO9044oz
IQ+EEXTcUsTGLm1Pe8JxDPxBV+rHaU6vuVVs2M1qVI7GC5+9z6BicvuK5dydIYlJKOKYyvwTdmqv
1tqq4PeWnK4p44PcVnp7mUqeBEoiTPwBazKxbhU/qYpkvlSrRe7PAGwOBrX4fD/GhpaoD1LkD2MU
98jcbeIP/FgeDNGcyaS7mZtb908hVq7heiBRvB+gmrI4sonFeNlnBDXEEFVKbWp+xIDQHjQAHpgW
u22JyVHTeyZG8e1xq6ceBmBzM+ISjH5USguPJAeyGPrCMbF7/DPaNSsp80Dz8smQhMvkqMAJH3zj
kj56W/w2jw3f6Zkfx73dqy9OMeZS8N8lyt+Fn9vbcBjGvF7MxCsjTjXQ3N0pH8ZN8WhP6rR62NnC
nB74Q3Tz0gE+J4JNT6jdkz3ORf+mOX4Wkm/F2hcPQJNzay4zp0bdYyP7E/LIbJ2e7iwmDFeOJx+9
NMIjs9DRIW5IHk+H2CQ+FDrJ2HnTJddZ0CUFPRMYb1t303k2SQlzCbfVZw30lN9RhiDdZz8f3SFU
aKvpaQCa3Tc6KQH1kdO6hXzJFRJC5ADD9OyVRWklZscczNcIz4K+twkZHDYODM2oOYmQNUt+JhHV
gir++7sO2hSC0DXvMkuDO8obEM83/YL+NdAM84mxPvPDYPIGsq6c7GPCxgsf+nymonOSCtzQ2j6o
8U5LVp1QJa1qGPaNN8jFi4nyfiHaWPuD/2dwKvwIBOc5GUIwaCt38Qgqj8bB6gunvJ+UHRWoTvYc
rdKT94rolcN4iqxGv7pWFUPPQ8brn0w+QUoZGuaKA/vHHFB3vmtb+iCUjy0q+kGGqPkqt0SPe6uH
VaMbk4s2aKwIUZVK5KV23/AOeMCeyO+HfkI+pzVaXeRONlcgypFqiaQRC4PR+lqFc9d7Z4TDUUkM
zOtkNHG3wcZFPyd17dM6kXF4OKtEj3CgkyoPXohyg6qiob74C1HUX9aD1Y4wuz//VgYWfDrQGPmn
PryiuaH94e/syWMpAXTEUZVs8hROOqjzU1mBdf6GVDy1awEeysp0BfX62kmzOVbqml8gi2ziWW19
2Cr7zJa9aSNClCzDUeqZAlnjy5Ww2mp0PkSATrEvAq3d/XJDvmrT7eUFRqsn2W4/BFlgW0TYrDTW
V92AEFHUYe1CL26EsSsGGLGGG94HTNFogAIGpoTbhu0xlNsJjEVmKMeRpM78KK1TG45DqhIrruoN
rlsslrOSgDK8oDH93CXhBiYjXC0ZMgZ7YS9XRvN1ivD9aD7ujcIpt164LijdQ8rYFumpqT/l02eR
qkuEdrec2takjtXNQ3K0hsxzkgGtMbJeEZkCSS9KMNAFnwJlltm62iK/ijxOdeuCFXmZ5ZHcXlCT
4Cg8JNcM6bvCKga1rgmMAZNQRCMpFItzZ18ovkhrQCmJ+pZ+FAHW/uecuGsLk2ndHifGTwJgbZNB
jJMygZlC/a8ErljlLyVpYVDP9ha8v19FavKyDUslnyjjanKahfRzO9t7U+vwHTNMJoltCZGLEGPj
tGzMiMMts6ycxjX2ncFDl3Cih32p4QrBxBrFG0OnUwamwxx4jHRjF0lMQiLrnDPb6U4Td8KqrRV4
CeOAh+nclZYkhDpN42BMRwc3VgYajOFYYqNGyb/VEc76kD0PoT0SBcHWeVJwreNE6AzlpVVzrDOS
WogXJaivPXR8QGunmeGWkNc0HY2WKtLhGyYDXnbrYX0za2h4s/x+cBQlrpk4A03ZdV0YLK0sTXjz
pJTc8VG/ZneMCLU5aI1NvVCdETFm6rsdqERKLfooN0zr+MenJKqaD7fHOy+EfZ9r0aIUFsXL7LgT
hcG3+eHQAVSW6LilCMXlZedKy0CNPP3Gtsi4UZylftpH1D2YjR1X34Fs/Z75/vBYH5LPe7uAP75h
PUbEca37Gk8NEqkUJbZM4A/asb2Zz1WBm6Da4kl7Nu+JOru66w4mhkCqa8/PyblHzfVX+Y6xPoqG
BOZfbq30UmBmwKPyG97pgpzcVBXvM1AD/j56hfXKB4SzcO6SFmdAf9360lW6CJrV6Fp6y17YIH4C
RGuS27cOAhSf7IZkSArmn35siGiSTw8EylZJ+7TxA96iGiJdkyYKveLIlkTBHaRi2fOvmMQ7cmcq
AsjovL7DZBl+M9z1sGwZjrLghQPGWJKJj5kzK7Ephspe7rhEBtiE+KcHx+qqR5IKhuPfup3P4wU3
U1ouPn64Bs740/7LAKfcZ1UQBIm8E9hz28CryXetiGLu2yqdHOpB0L6/j1r8vUI6blIL0ObUDQAB
EtorihBGKVeoutdOszljvYO4Upkv4RGpePTkb01HMfzjdeFfiwaVArSPo4oCqr3kWlEfabianOC1
zB7AK6pW9xMcg+duDLkCZscyknytq9RFUXFAcWiE40myMLnkVNRxm9uFeg9isoksdLOykO94V4h7
kg82LPv5rG6oCv+QrLyHWPturg7j1NxrCZRZLeV7aG70c5+qy5OdAJh2bZdBXQXPMdIZanv1HS8m
3QhNHpBBgMuit/ukDG7GqUpWUwnIOUWM66bhkhZzhIo8rj7uOWVS3SIzjHobCyj0KBOZsbZo5Gau
aWDtTtG+dCxP2JGOXJEUOCyt0ZOFq0BsonPXt/exzH8RCugp6OkGIBaFBM8hkuzvgTY5pV5Ol5z5
cfdHInAPKkQbxlKqcxq85Ao1J2ZmtBupofMUpOo/llywmbCIQDz+UggoGkdut6GAHBBkt/h8G0Kr
LMWFXs/YJddScAzocwTTRBxcZuysliUbp91b668cU+GRhbvCE/07nKDECr0qE0eIb1q3N9ohM0NN
WoDechkkbaUwuR66lO86OsVXwdAc3w5RkUlqvQPs2KIBMuGLzu8b/4RvVcWvgZIRFjZX+tctKI/L
BguRsfgJsl3g4U1xWCitahD5XNCu3SUS12oFHVgbrHC/wJTPCFM9NewlqdwK6OzLQDOuwlHTqqUu
nMRxbPpFmy5rstX+hySDG+5N1jOx29ZynJw/MyiHPWPPpT9w00GUqnCv3jwpQXDjm9zbPFGZGJSl
gRPjFm98DDc7ZGMXqBe5y6o7e+8ziiG3FvGHV2FxFY6hd0rHJLYEqjiB+wR+a+0M3EcMT7MVH+wH
OuZnzbCVcyY4aDqwErUDTHFr/jHDP+wty2R8Tu60nq8Z0SJkX7ryKkJ9aFlyoQDzsYVjFrRXL5jK
TGv2JvLE1f2rePMkxCuZGdrU8f05whCI2n9r/gduIahE80GcoNQjA/vtx9+yPTUwi768kXDq8wPP
CfWmhrcSN+JLLY8BuiIl5LCTCoaC8KBfed8n08XLIaLWD2/E27hf7D5F6JphPXUIDnwOTNQxJLMl
X9nP/CqMSiNIRR9sbzUKkHgd1ue5TAFGs1K9QV6vbowbpu0qWnT311ZYa/28ibLoVgT85V6Ixa5O
+muEbT4znnKyUaVy2R2MtomkuhZYN889KpWv7/c8OnBPjOy3ZoSKlRgqLNoFWna787glnVmxKOJ0
jzDBdBJmKTbbYWRNps6dNXm2Jg1G5Q6CoaLBJc+5eWbC2wCsLWURyX/yaEg0DVbaAUbsVXoootZE
IdhKWW1FqJUaE/2BEU6YfxWWAAyDf29ddprxudoKdS2fNA76i0RrYyxFcWrEXcLDS4fTdDa6X2JV
SVIfuXqUUJOAf0+XYHiiQPn6fBG3VIDrX2D/+4a0llAcoRruMlO22jCvFDkmNVcHu5AAXh+6B3kp
SZ7vQlzLjaRhTRMJsf+6L+FRL85xohoQjbbtl6TmoQ/cD0lWvkgHzk0wFbqynljpSpCA6yzNKA0M
Ykx6tUqPSEYWGHK+bGrZxWw/cKaoKN+wp6NcuuwMeevvsJQIJKfg0wIrj619oKXqkMaLRp8iw9Yo
UAO5urR6pIHyNdHzxhGqQMOBmOsFk6OLmJZ+rWufHOworR5V4xROvMN0q9NnStDopV43Lz2LQXEA
voaUu0ejdxU7cDRFcfyuD5eF+7+8eYEehWUzvt1/Urn9aBjE4FRNyzeu9BZOLnwzG84y7qLsZwxO
+IyufLH/p6rmQvEQp+6mmMTw3L2pMjDDioInAtxtcpX5VbLBvE50V+OUacCJJMdfi+lKI5ycj0gO
eqiNEqQgqBaD/twdf8EqA8X5ZN7TZg3rD2M7npEBCmpz3wYdjnivc6eTK/J091Y60YtEOn1Udom3
FRbZ0A9RekN8qOFscvekq9sIX6XMbauvcqg1rENGoRTWjTZUb4vEGfo2S7abkPDCHwUOzhafPCYp
LdXGieEJ6kMYdHwOudxhi87E5S+Exfb7k9JZVO7X2gk4xTAWT84sFrY2jaqOCL8kM0gboQWXtPk5
lpy8CckNeqLzVK33Z3zQLwN6311qA8NWjxI/Ger50h1Z2Oi0u4IPm8KaIV4r4EEtnsArQ5OTwyjG
tq7Tl0d5STF+TDWQyibp8kufA1C5I0WmHcI0otQvneWNLVPS1lr66lC+7Mm1B5g9JNCllGDjZ30Y
2c9x91l+zWf1gBUS7+vy9PPHnMNbbZGeqJbSGFhBsgtP7MGdvYo47K3DsVB+3XAiFLE8lKTCbfdU
iso4YpKVWKA3O27QZ/ZU3cPR+nDX9fLjQWBD+kEdH3LElXdRcteLa5hQbDWCRvJHHgBWt4tMn2/A
NpC4Z2nu8mzonwmgBXAT2JdZlquhYfwxz7c2WAA+pbb2/ZvqWDCahY9YhMIjFSfcZs9YFzWqc8RW
znzsgJbzg1bgyXjayv46VkyE/hYUnSkQq1TUIYXA3uii8R8i+Efoxtfdv/BMF5g3tSQRQP+xZJFo
PUIfksz4KHdZpsfNXOYP356ZwHffDjUT6Gmei3rjFSxJd68h0QVk3pHHMotvBO+sNqvQEmnXpYSR
omAnJVDg+MWIZJu6OZsqYHsQN1j3ttat+vcSs/koUVMZ9Bhhpx0GX5qS3pfpT0GZ8sT6YJysv+ZW
gVMcyTt9iDbOaDkV68GRhU5ALqY9uYsM63m1X5UAu4rYd7FCi7VjJlJQOUUS/Xgs0noL7NsWnCAK
1RPv0iTRIckWy74D4gnIgc/yKPrVn0bTHAEqPc9EFm2A+8pe0VynDMIXh3b5uFKLFTa3Nn5+U90j
j0od0BmBicSKmjl3LJ414IFf5wxxUCjJwUHLvGlH+VHYSspvhVb1lcZQ/IInqbKevhvxf/LS04pL
csZz6Nkp3FYBuH3hH55nhgP2auwaYnzbH0+K9TKTkLVONgS7G8YpC1NWDk65/9I/AZlwlLcTH1fc
StFbOvSATinlRruOsawYL3TLYCq7osSzrSyMwWUHwvwMdrjV4Vqz0AkG+C2erd7d2HWFils0o9jd
mEhIqhnPVsDbiTpQOrt9Y7LS6MpZhHgAo0K7ivq6sEriilLB1telYGEtyqe/3qrFjvJoDWQtiEyr
H6BgcIqaOoYus/kHjFn8JpitBMPb5rlQyqJAQseHNtdRMDIOfHqFtlqvMphlhuQ8b3v+1TcyNuxN
A4rj/a3k5ypn2TU/5dFZjlMQun2QuJe0p8BSLqnqHkggcvh6RBVGH8Ub1Za9FtNI22Uu+L+O86Xm
qTrM58uhf4hUDHqiffBX5mG3Y/j+ItFJKyfBfvR+TECCelnG618F19uvfwBA9CeVPVCO4CID2Avc
Ve49DoHWUI86eeZOi1ROWpexiamMzwubYjqPcYyFiBFKesV7mBosZFoFAlRel1U/KEz3Qn507k74
LdhA2vslHxlkNJhw4gvJS+MpWghcIYlhlE6auJBhR6hdeJnFXZIzNt01ueO6zItH3mfDGS/oTw4y
q02XnoEJu0zyC67x3J9HTmwv064P7sdQD+6g8rMYLoSkilwKOFt2orWcaMK8azSc/9PjlbtTSXAv
a5gyfnl23bKEIlIHj5G7cPODiYidPHc6Pp1c9SrC4d9V3zEx4uRNyw6BPAcyYLFXz3YqzmpgEEiH
TCpDpB4SHvFthOjPRa9lsrQn4g6Zj8oIZe9EeygWUpAOffXUTjT6gHucQ2kYjb+U9ZZ1EGFRtcCy
mI+4rU8tFCFm1DoLWlL5TnCiMg1EWGnGx+J/5pRm/fi0Zw4ELlDhpvGYrEY0Vq48HxynckgTtzr5
RagiQcteBeXXeu2p8TqOXHn2O/4v5Ij5C5/uuDxRsmbJrWTKGLa2mqPC8E1M9NJgpRuRJZqpddGA
XPManpxnPZsVglwux3ePyvHHXgPgRy/RH4UeklyFiSLWT7wRNj3NeIv9tPCrGdTVAoS4UTVo+s2/
2BVFYcLpEDMfGedtRij09BOqScUaQbIOz167Bs1dIHE2nsHcDGrQFXPTNm4LaicixVaL+It3Rn2D
wnPqgJpsNagtlv1IsIY5nos+LQd+3z+0RyM1vCrqEnBx1bSn6V0UseTUYTzJFJaaAnoO2+OCBVJx
6uYa3jA5X3Bj2msX7JnGfGNCeL71GwBUiyBN5DCWOMH92w/QA/qNkExPue3HqvzfPf3QCZRm+/p9
uYphoKWXbTaLSL+K4XkzLgGPvX6mNKbMWH5qQDsGByfZHMSr9DuyZWNCZDWy3A0K1Ram3hc3B/eJ
iI/hkbEIK1soMogSqJHKMo7USN5iGFGXF/INq/3rZtoVkOirSBGCEXlvJ75bi2Jrp0wc0rj+tR4e
RTewMJP/WLiSVgvSf990EXhF3RdyT6oGGYa9YaLjPcOQ43sneaf0zPXr1BFKwSIdxt3Hv3BGKVho
NO+7Bfp//bML8l4ElSWSB21PID598vgRyXOE5bdIa8WGylsZxRK3YiLXbz2xpGuYITpMZMsX7h2F
iFIYkyX0uEzEWFRCRImkL3mju+b0V5PgaV3WW5VHXOWSohQ0xv2G8V/wNMtdH3AAfQBi3LmeE/qx
5eWTqX2bx0iMAq5cUr9HvHY+7D+vqW6TYivd7ieI4OqE0hWydpVDBZItzQYxWKqhN3il49Up+/eD
Je1cFAYTx+t41r9Mi63mM9e2xe6CrC/tZ95hnUPQcO/5ppQ9Bdb9N6IjQ4f+WtFeNHRX4fBCgLfE
C0DymrkcJaQSrSRNN71rIJuFOKOIlRLodoPQLp+J7/QuZ+NHUjlkjG2tlXLz+Y0AC8dO9oxX60EK
R+yqCUHf+4snUQdVDAzqGqb0VgqpdVGjY5yl7LkHoSmNwpFCpHssGOxSdEJuE8eR2wjlCmpEmMkY
DG6dSuFLOvBLtgZJOfG3Jzo8/qIoD6QZQ7JLSYFpKK5BV5j0jnxDFmrStvM50kT//1scWlfoBkNe
roNqgZoLjIxMiDJjipbqdbijTzBHiOYOdxnmn2HF4noYbwUQ5+2abjjKyjOZUdI+RQMPsagrcCS3
zuwAVQOkljTAz3anq0QwsRXtZNFoV8YfmoimqOO71QS9bmdOpb8LgtQRgy++sy8cJNwx9/OT7lu3
f6qVjTZZFek+csx8LIhRsouZuaIlwIDJSkdt9LJLLH+pnJQaf2ObJY+O1F6lOEuvk7cjf5Od/c3z
zg5Apdd/3qeXOGWw3sY3x4bdUzq7Jx0SYuACsBuuMsYCh5EYRmMdvxeNpmwvfxgP/Pmg/meh4H9l
tDtnk/Mr5gG49bJED641R4E1wM7hqLGxvmRyQoEIrf4DrEvJHivUGlca5+QyqMu3KFe7kmNSgpjb
s2XGRGKVNE7EiIs/krzP92cPlsTi6LDi9liUkxCRulB9CF282b+SSXUhQ5olXT0Cxe0dU2Tl/X5D
CARrrsOJhsvPvxBwefgPnjXi5lpGCNN8n1xKqtFGeJjILlf2fljIm0VRTS2uwMtT+hpI1+oIUIxh
P1ZE2ZWT71eJez2MueZQwI2emeiNeTg6E69QT0O7SMSr1GlU9Nbem0esnrOe/8TMFDKx4TwS+wCw
muYuhiGZLDjF9uzpOqsBWXJvPVNi7DehZM7jLeGg197mtw8xIa3x1FSF83g57YAuV5SU8uUwHghg
prgV5Lpo9WkoyzmCY0orQ1yVKnZMtWlRp6waIUfYUWzg/HwfSm/vHPyQj5Fkcmydl4EU5hQtSjSN
72B4F4c1fV3CBmPt29M09zaP60gthgPshPU4iHqLPam9aH42xBR4WpL6NreOJx8+AzQKR4Y8NmRO
LAEZGWIlXaLhODOrfKs9yuIg4y6DhMMduXhuXROLJB5Dg6VLDrTrJdmqq+zwB8vLlHeoXL4YbeEJ
wKf2hkcFgnQKOJ3bMmr1/rvfTrxArW9vTd17dFrdnDllUZTxgau1o+WYzrvhEEzxP4GKG+dzZqto
pLtaoD60V1lgXqTCLD4kYxZGY+Xx7HH86NezBzQ0sin4iCvW7q0JcnSMzISm1duvz97s9ApgCDsT
uuKXKDfGLwn/CuEJLjp6eB1C9a5KwvK6KcClMlMlIdDHDPVxD5Xy3vvqhZSQYxnJyhLhgqaa0wvL
sPieFRBBfPyOW8vlwG8RjuKdeh/Dxf/AnLEzJS2wftX5sFbm7P33NZzSu0a19lSycntsQWKFDKnu
V9zQABshtrWqCU2lQ7O7JflndUB40pklUT0G1cgx+CS2vtiW8ZpBvl/NU4W/UcKwAS1lndiY3qBz
m38hFtXhzOeuHmMquy1L5m0a6WPsqfQTwLl1W5TlUmb8fa4/VV9EjkfsP+oI08+eE9AHcbXzoEds
oPOoKxa2GRWe5gfybm6ZrDKH7Ehg0KG+qwu/ol2WzBZ3Z7lEkrY5wXaShjUWN8TvlcdP+98OcUTn
9P0nHGAX2Udh1SwXzcw9Sw88d6diQQ1d8XXXlFSuh+tIqGmd3QefZxz8iwMxf5s+5p8Kc+LWsAJo
4cQJKAaI5O/XWgQcMliun6SSiiaTLHjN7aVAzHtmP0st0u8wlLOVhOwJtoRSBihKzoBFtnWhSAwI
Gik4UMkw+cKQPymzRNhXrKE6vIIqknF/8xTRcRSodqaw9QGZRnbPQG5S2NsppkVEeVaiUP5LlFAZ
Rnfd1w/Pf+Wt1bSMZKXRo7UBQFif20XORc43N4cjdMtxb1GfzUYH1mQzDl+6yCMEJrMtCZj0UmpT
Rrwt63U1WS87tKZFVVIRcncvV4+JA9YVNXHfYlykb9xyvXRkYG7HUypOHEyC2ERL5LmW8hXdGrBo
HmWRCw0MicC7ym/YYyw0lPcG2OvozOpiw7RGoxtrbI8ZUkrMVBSN+lkA94o94uTBpHkHOJRYR2yo
heNtUljYX8Jyg1upp1mlnFZSV0V8Dm7DKnhxOoP7g6BG56F7imx0ggs/daAS0jSW02rPfDw8uiX8
QA5AuW/IfiX6RgkaWEUKddJqFVnbkzmYkmzprvIQU+z5qWJKiGDlr0K8mmqLXP0hWVh8f9li/snq
QJNVx3T7y3Cy2zEjU3Z5gVrqzqIV/8mRw+tFIpESG0+bhKfFR9E3GpuIgdCgH8Y16lu7b4eXwqXf
eEJitXz57OTVdEDlhReyXGuU0Tj3pv5DNG78navIZhbruDABJpsMu8DWSR617qCl5ZKbPes3Cir+
/mjtH2OtnBaGacDvdWMDy8qhEhYG8YBSgKNGAsmQm+hIxFpaaXRkQtPgSi8sZHEbUCn+brAPjdZF
aktcpUCZocdyzp3oPVac58HcnKp6S8tkPR3+guijXttt3L9FxVIehVitDM69bzljtEiV9AkIuF1x
ikE/JzEpvL1X6DZKZryTaSiKDF1dPAdYrCc4piIbNK1i735X0kp0eEK5DZ2fAyE1KkPGF1QExeHS
+1zCKq4dBh62xSc0i2H1B7BNwgWo9BESdIVfiObOxdf7Y1aNzf41MgoPqZXYSA5iwHWFJhppoSzc
a75iaRP01Jqt27ssRkfLl3F489SsqGofqUH88IajOuPZxiKBxMZbJMaDBBqpPVWL9EveEkDO7QKe
0U7fuZYZoWlPpBr9JOdmNyT/1au2t01ysc70ztd9zfYACh3NznGBS6CXHrLb4e/IbHQJOlwkNNZU
0QeUtW7bziFvgCtAM2ivXatfLP3AoL3IHg8dmZY5XTK8OcWYe8xxxfTvqOZ8/aiGkYCUuvbfov6b
D7MpSjL82JS4fdfwuhXbLxtOEZ9r6AUn0xjnBb5Hw0uj+TVmpS5ES28+1g0RQcGAEmZrgJzS+BiT
JwlOsEZfA7qddzy/dcwGRirN1adzs3L7D5488jfZP1IXYhp8uTQaDBy+DbQLTv2OTmGseKIjVZTC
+diIiNh1ickJGw+Ql8y5KHOVQWlCt8pcxogA8S6a0B3XLYZxmJ2t/im+i2sUDuVzs6URmTE2JhYt
NaMSIjztz4b46S0jNDFQDKGSUzaB9Dqqsfq9lav3M99rPKFHXi3Li7FszHQRHbH5G4QWtgMZHLa0
pSMXZsjMI+LxbnnReecVW7SQtuAnnhnFSEmP+VVzxy1nNW3yr4Y7rtoyn78DLWaHvvcQzta0+6Tu
5vBUQ6QFMQdHIzWYiOePDg6Xxrr6Q/y2/sqhrQb8SsNtC4D2m38j32pX8MLDfDjSDKN7nlAmCbN9
Ry5CGVFoc2RUhlBLtRKsDukTHAk4xgyBV6SsmkuxA+bhTcMGP996PvZJ9hGtx+hKT+UJPze1W9LJ
k5vWxMZtzrCZlVgAHhE5jEABzZR0GIwgylUT+6bhFuwtIfY8IkBWZEjTBbhwaiuccO90wlRSxPv4
x8aVcwI+NqoMrwLbKdTKdX8Pfr/ogdKrr+zfFr3xjCcYniVljL4Xt6jPA5D+3DMOHoxnRLgdIXFA
zb8q6hVmb3DKeAaCAEtipshoazH3qhotLSxJ5VGulBNTGbZNTgEfgvOP6pEMtHU39NUL3Ron0Usb
vwdYivGECfz4yxSM2su978FX611T9hjiI8IXNP/rRxWElZ19tBusLBUSD8ki3YMq3YxwzPZKjbcd
4ROrFFeQyMbuUqp8bmH0DhrbToUu9bqZgUxeHFke2MCMLkOrnlAlr7BAWwH/6Sl+YMXabc7RA9sO
pQRC8MFYZexhngUQPoF0P6D8d8n2A8xVFnhTJxwrtoba6tN+aP8VOTtexFiC41sJqj1M/FL2T7as
eKTZhpHhJjfbe3evmj6iCYftb57hvHQfb+9KeH1hzxgy9ZGj33+fsm3J7rDimnAezK1ICQ/OYE95
GPmv4udQ2uy2RTO0Nf70+droI0K5DpzqTqTvif6raN6R8LcrGBmXEUc6m/iNCZ6WCn6iLys2YBsM
F7RzVQYE5fyU113Uc2rqQ6RjY4dI0GsdUiZ0ZXn679+GebErheYXkFB7kydH7dux/lSrAkF/Ek+M
8DIfpS0C0w39bs+7qcHzex9sv7tU97+tG3ymfqPNZoC/q2BJfLAlN40XqY34hGHJwyZA+ZJDH8qc
p0eiZMfu7DNgPIWYGwvWLKfbFbQnEWaDy4tj4F/3CpQwu/W6ER3apw6NpdwCpGpWtmpUgemce7bq
S5TCT928azEL0KuC9NjniP4h7Uwb66dzn56V7cNxS9Mki2yTDmKCrw4g+cIMIAw4/SPK926v8djc
ngHcAQJVg3iOnEsS7SFgPrm7V8E+F4+sz5ttVoLypLBg/g3D9BF2p5j59B52GNCqIVMSjNF4cC0r
0igBn+mWJptCj9Jv56Vkiv58ZUsxokcIphMzhWZguQziqhcLuhDRsAvG8zYSLAEUcLZx5OqSdJ+K
8/JAhtWUUQVCHFxLD3plSQibDPSqu62ijv/0iIxxVPpzfXHKQ90/gIDI8WT/nulbY97yjyQY5vRJ
Ei5vVWLDJ3vUPMGVa1tVTRQcm6TWboXBq8wy3ytY0gS4gVucXRJaZ9GHcay3/VSsb+Yv9MBNl2Ys
WfxZa3NZ9PFl/coY449ccG0NK35kUzm58TVgSPdKiD7x2wzpKGL412UZDJLC5OKpkbuREpdPqxm3
Qw8zApfRs0y3D/zT68axsAJy4lb6+c/2r16kIeZGeoKRURsd5sPQTNkEs2oMCYaD3UrNbk9To/QR
+qkyzaNx01U76lPWjHxVtldaSFSw8uNUwspLR3XlpT2+yKvWyscVdW4eCwUhpVE2xjKhVsh7C7kE
x5cHYI9TSeie/itNbgo0VlWI4l4nl2HYhiNLGuXpXmHRKSiRimH/uOU0gMKs94sz77ZurcmlHAeg
hlFq+aDkm1Cu4kAxkVy59hBWQN48pnejtdAxSbtGPcrqEMc7ehJkMT7TYd3dt7p0lRaHCjswuO+B
ad7ZZ6rcdH5hRtv4JqIeoxIzAHDnN0iXOonuIlkeRkYHB1+XAP9uh5TIu0DdVU5nKMUGx9O+saC6
ZbfObsCqPfNvLtSI/XekYX8MGF0dUG1pRcPSHiWGSQk/OFmG47XC+sA7cOVu6u+qAS4wU3aNJSeH
B+9ftp3sztDZOdcMo7B4m52rMzujuJlMdAcf+SGeoc2WeBlYaZTvCedAwq8lPmPOIUBw0xiOiiE3
lawiXn79JASobR/wQeLEzJ/hHNoSXMMvM0a1ERjimhUBXqEyKHED92eEVFnu0enR/2T5X/zSVxml
DhsEjGS+KwRBXYjqwC8R43kwsREYA/qOA5Z1+yGEFf+W3J33qp9zhvUUbtmES3IhlP0KW6AtGPOi
jF1njXBopfHSsfQ//2HQZ2ml9Ti070k58AclGWli2Ps4w1AXF6RnYPuCfrfxUvU/VFg++Vc1CDcv
MhStlD/50bvucnozvoUDohivrwF84lUXcyzbJDMLq1hpGeqrr1dmGQZwn7tU0K8oew1qn+LKUL4t
/MHfNa9fDZHT/rTjzr2Hv8CpRzFZURJf3c2zeBOEtqhPsFYg49WpubSBe/Y21h+C+EZwC9U+vFdQ
YgBpoIwQ2Ihu3sgu1kYp9ASFs/z2nPXnpGlgpgTI4xPulVj8KsCjgH3lOan+tS7zvFzbKWQTPKu3
k5KFtGwkp61Pi/FCAAOKwg+mUlvfLidw+CuEHkulXCtq0WLpWsLRzVptXAPcvTxaZ12fUiiTVcE1
fBwDDXSIfeowg3VlJ8qQiGc9wmk+LRP3HO9Bsg5nrxjdp4ypnP1RCW4bStVpVpqEbvLF4lY6iPF1
lgq6cy6YcqYoIsuR/TIH1pq3QVRTPg+q8un7le7s/c/jgEg/zR3g4YzdjqoI5eVcTJ7PqOLNxVJm
lQ0VPKkiCdDZvK//bToWzN2DwUJbpSKroIQ5DE0gWa1ZC4oxIgKUHNt9iEbz1vOiDMB+EbxCll73
AicDsLlGP3wAA4TK6b7uUO02nOPqTJGNRuDXepBNPeltHrcYuStPQirZPsP1b3yBKDKAcqkSdP6k
QpXERewxuOhHjYolZ5SXkVltLHc4Xe8eKLX8F/Sz+7T2p9f/FEw/DhO9hgMMAVLSQJLSZY2o84Lf
ERgp9vYEfs1nns5ojQ0a9dUZd7lJcWX/Affdr5IoFM+YLGXn9Cm1YtSroMRAx/E6H4h5bAq087p8
45rSeIKnAiZVYaImN7LqSz7jwhL1I1kqwnqAVoiOLbAoG3bt/QjSanmF5BcrJN2rfUGjekk3RLT0
5F9kkOL7cQNtDmGtiFgFthIVa7cHWp757HEvTa6jt1J63xOF3KHy6Ng53S6HPlT2ODuzw/AHsuMY
t3AyaQpDpr4neKgCk7y1m2j/WIjw4/IzGKMGZHkDCGkp8pCCi85GVb8gJN/3qwZvVPdb2/Gv6Smd
CcJ7evjj5omJOOa+vzma7Xi6lesYgCz5n+WpV0tgb7NtBpFcKEooo9VOm5Obz5RVsb9tPU0z/8te
Yfvm+f+LsHoe/3o3MgT81cv5PD1FjWq6yC6pC8LsP3Ml5zQTDZkBBgefvP1j8IMrA272nkuG1ea8
tXGdzZC8OXRP0XVAGrO/EsPnU8EQV64Thyl/1kBLR2yVY9hTrHjzNIWn/z1EfiMfVUUKGXFn4cSq
ozvLgSZB04boVMAxGeffhx1KFhb6T45QX625hHRUZ7IflPbKOSKROjXg614Dn0mXw3Q3YFanZ+a+
VGFOGUrnxo5jsGJGDCnTSQoFqm0TbGAZQCWb8yk3hCRdDZAwrUWOtk4TPexiRewWOc0r06UEGNSs
EOUQENpR2tP2hNy4nHkn1gYjc5GpuVJbQirowLHopMJsOPXLbi6cR+DWFILo18pOdinG3qKFHoet
HvSVihzZUtyDFnLgsrPHj2yuNeNt24oYJeBao8ES55HuipH4mQIE90WIZiGnapXoj5tDQXeGuAP6
95XBHPtOl4SWS//ASS+Lyh29K6FqYu0v/njWRod6QLGZyPS5rgHfKd+LhRmcv98qoqLQGdNwPbsZ
bGkW7FGl7A0+cncLuNCzcd3xir+MCUY6hfuGJjBv9XlYSrQsPFMkfjTe76zzeJmF0JLkewc9HqRx
wxj+SRihUFEfl/XQW/qNwk9zP8f8WiQD+/ZBi2KzQlgJsWeP94q2QOiBgd5YnR8nO1mtK2BOqgr8
yT5wTMauptnBKGMKM+fb/7SsBAHJZpUYmBrbThi+/7rDfZdr+bmEf2ObGkivERVj+lSE6BevVPUq
yNC3q5h2ir8CVE0xg+bDXbSrjAMGPKdqFlePCdSnJ2CC5Saiut3xn2zBfFYfMLerRlafZmwGnDGa
uZHM6D6JYRUZPzLW3+OE4QolOnR0ZcgOZxkLlxMmtlmPNgynPk7DOAeKWDe39v3Chj12WG2Q7yCo
8EPMg/iZ8puldpP3I27lDqDH1Q0REvHdcVtxED5el+AIQZHMXfWHgQq4B5eHwoinyQQtAC0X8suV
rSJJ2YIWN3YEl5SSfS341u3GjYh4RPJOpBa83NZgDMaxdk+CkoMSTBQxV63ltjwjpbNVUMMve2rb
9BXXiL3dlCMQkK1QED9sJFyr0gopG98xLzBeKrekYVDziPk5S2g9ua4EiEI1SbY25DUSjxh4ZHnm
sPHEIsr81qX3pK5oN6vWs2eKfo6Ley6c5mqSARdxvCAiOFUgFPEF2v/7gICor1lkNvjQEAiKry6g
V2wg7H7cMX33tC+R70YKfnjb7y0r0jwO1uhq+Ng+ApTm8q0+51UaErK6BfCrlxhfUWgyGNlZMqoE
jH6aByl6fA1BlDiJOU/KNOG9vDpbhPDbS8FjymDDFvCU7pydLdTPM2VV7n1rIkgVGmHorsp5q3P6
2NhhYPbMsZ4Bb1dwyhOqCz14cuNPzwKxZY6h+QWUkbTwk8WI15yH+Gn4WNBaVX6Ww7r39tpES2Ez
xhgpAJpxvmT6ndXKSqqqUm+igDy6geDbkEWq/UJynTCnN+8yVga39xQFDiDwYP4t2zbAOLci+9pt
RxkK4KswJuchpTtyGjRUxiDHcL8VgbZVztuuagYJnbhhJsGHjKxkWba0lGoA8OfMm5H/L05rwBOF
8QPXPXGg+5yIatrYgXx2mYQmOIkkMqIj4HsxfMQh76fsXBEEkmNH+nlTDV7UP4CAg8Q0HPYHXEiM
zI1wW9JPrZZC65HedO0awLw/6HIAbJDl30yOGfN2EuP8ZLpQvB/uxXg10/oXFqEcvuvIl/6ekNCZ
RkFFQEhBU85DB2Lztz0jdf8YUwN94e2mo74CEEC8GFHeC5Iuz7bSFgv44gN9gbgZ1+zzzzGymEtz
53pHFn+oFC8RDX/yajQz3hcDUXG/iq1XiPbXuzzWNrMDqNE9FSznizp3tMv22miiZ8TK6o/UjsxS
1+/84GQFQ9GwfirJAo5q+TIsOVwnLQF/Hwjj8aYdcChLEkTDysv6xkdXdM0vgoo9zP9btM9Lx++a
CIQ0yPlZeJUyFyIIbWNjwVRvTMWJvArBdAtzmEUmNUMa1sbLTZQpEtwcoBnGIP6fepYuLlJCouWf
tyI8qPhm1dOldKmt9FZcSCSk5J5Uw6b5+orPyiEHNGtp5de8L0wbJuvIivd83I21OIyIubMi0qXn
0589S+TfHDL5K3YVPTQWNMl9d2zU7PeESx+Q9Y8eO+/YaQJjY0KQ7V7PpcoR6R6mcXWhgM2ONNoG
a9K7r3srkcLz6KZE/GjJbZqS7P2lDwMbvngcyaLGzWqZH+F/gj6xDTA96xxk3H30FG7i6QpiYr83
FcxhtDShxportcBf/aorMYa64zgFnJKs0FGlqXakVExkl+DN48gRCXx4JAOYRABUYUMtw2CV3R41
u6/vsRZq2GkiT0Sggt+QnOSw0LP8CSgEf2ZWo2c8wJduG1Q5mvIi358vf5XnA2BtGQEUatEbvu2D
HuersUtNkXqUmHcoNFrYEhwVh5mqdPRnVW+MNkPfEdvJWBCb3XQLItCwrnkAMbpPLEALHKbqbWVL
WAGYPs0vdY810MbCMc0ATBYcz8z27hrc1Jz/0WbQJJ0jQgXZjNwE5DKDZI4SDrihWesk3Z9LARbi
7enyZ5aCyVTY+T41kyO8EOtAlKcFCSCWc6/wePl5CtcFRws1rWU2xXqAwRcqvUBU6xUtFITpIizG
XX9FEWnHDIbOneaQulr3nWE3rPz1R7U6D2D+XT533oXCHI8blYftmf03o0oYnTLM/Yk8f13Q82PY
XvSOzQUtQLLc9xKBBBfpZbdHv5tuMjNmF2iMM513qPXigqeoikoQgMzxaTr2UAgfHwPwNq8SMlq7
B/bHfMG3du/GfO21bXeqzvZmX7WpFkhNLPaQMb/bp0yaiR11YQ7ZkzLBkGAijBZaZkl+xGDk3ite
nsPjCOxlOmCgF7YM+moyYvC43Zp25aM0CW9sH3kHcAZ6bGvwkAPKCUlU719v//5/4RGy/YKfugo8
l4ixR/Ss25pGhSzx+sMfJugDTWwdXr/v4rRHzSf4k/2ZhQPLp1W9+YoPR8XSGryDFUDG/+Wx2ABS
EFYA6Z9rOgYYDAD2l+3uvs6vDnmHIrvSN7A/WMeFYEYlRmNkL2Z07JBLX2zcOlgnHs2OEq0jjgmT
sYjDkzb+SOMBR6MKl0ArsYYp5iNJAFn+OURe34PFop1mejhQS+Ajwwxf6IrGaHFtMLAv9hNcfJ3D
6tE++u76h5Al3/OzR+3dpQhS3tBaANqzOqjXdWrqbxLVGUJxlKjOV+o7b27bB+PoUVuWY1tj/7je
MaXXmSot/QWQzsPs++Ehl9eZ3YxKzKWiRvzQZ0eltOStG3CuqSzIjYs3LAbjKhygHJ2jP7AhEeOY
3icnu0CNgYV/rlqQzRgkJ7BEOYvbYBPTclAWldm5a+7rQClpqjvguDYQDeDCTKlOQlKCiWfug22L
BhPS7AuvvPCekshAjqOVaGUf9YApBKsV2Y+4D1ANL6nHArtH9D/u+8XldBhs/1uMPdnvhb5qjhcT
V2s32859Y4HMcO4MSvYngnEmbXJqZo4S7Fw6c+YUkE4k0Y7/2pv9eqbHOi9oIXOElEkkU7tiCqxk
I/sqqQcxkQ5IZ6SibmHPT4P0zBy2vkynZ3JDfBEmpe9YKAJz280I9OVaEjhU0XPkwMmY+UDiP36M
B//CcUWvg7bwgdaHUkZbdy4XmYDhjtFpCbVJ/glTLypX2FyEXuFzWRuhFGU8kKD1BDOL0HJIDRMi
RFjlO0paWoAtBUoScMfaeQdjDf8YVbSjir8roRpzoFUIO011oFSiT2R0D+Qo5K5DoJ4siLjc0a8t
6b+qOxUJbPYTs6hCt6l7XvF4SudFo3cvVQ0CQ13IRKGoJ4zzF27vGcYBRgkz/8nVGviw/wk7X3Ah
DkJxAAy5xftKBO1/1l6Mk9FJULGU6gWywt2GDF99B/t8n8QHaBtQUS8tJtWw3cOz3bDqf0q1/ALC
++RZqy1vkM9Ko61Bd8hgbTlhbDO/7pF4CSWoubwNyxV5NW/xOaI4eL6145Oh0a0sDoKLrc0pGGaR
LWAe/5b7KbbRmOM9mxlskZCX6aDILGqsX3PTWpxrUW0l8bH+GDHbs9rQxdmwFAfRRtm8xh++4GsY
Uh4UV/ny5QjEMbwN2pxU4y8e8ffvv8O+zg24t6Kj3SCtHKRGRgt384DTVgDQ2Hn5zyktlPOjlhZJ
6g4/CbMnRj1QrVti8yJSeyJ0m1f/V2EX9Nq1XqBA9PgRCYlHNtpx0hCVozhsvgGZuTSqX/7TSRzR
oHCheL0raxuCplcvqqv/zeZwjUrcFqTr9HfU5tB+k9jPnnr721X7mmuGfwJsRUstLwIDh62XBWQe
H0S7E7JeYBHDUl9M6Gu9hTHuWHGeqPDUte3DyA0DLTc2Tt32AAdsa7fbGPwuttGVWdP9RoKgXl3z
+X6B5suSprrzfvvWtlXeifQvrwXGITkBo1eNvWuTGdymAEGO90JTLmAIp/PgHg8W962xZbh4XmcE
a6fq+vBu782bHUfhToCAXu87veGQIioGPndRaSBaJH0X677IziKvOiOIkmi1mh/X+B+mZgxzFgJt
CIW+VXHaXXk5f4OVFH5PtIBlCocK9Yw/uTA9O0w70LYxNr4q7zK9jT51enfDErpw9uVqdCJ2L6lG
pBjxfbbAGg51DYexwoq731ui36qm2Ue4ZDxqwfWVOXI42O7Sj7xl8qWNZu+ygG4a9Y802CG3m+B/
+pUdGzkbuACp56T8KxHdUbMbBvuLda+f/N8zO0ce+u2KoaGUgpuz9mewNPJsRfGP2bs4nlkrti6+
RC3HWZijWTdoi0j0YzEj5cBkjYNZe0CV+bykCoG8SRgL10kMICZ+htptgV62mDli0+27g0YUtbFk
K9J+azwDWI8eaIuwFjRaBDdmUBEH1/hu9cKJd9YB66uiPOhkjoDU4jhhR9LGNHpsJtSQ9Jm+xJPG
sWR2mqIUtZOLYhT2QH+x4Wdytdw+VymzwVmvbk1MGzjxMBMgHCwFvYAXftUtDq03RIyrTrfMl54F
/+GfSPdSpCiywKf+nnKqCnP9mp2RWlF4IY6HJ5obznR0/ZLfBxnH/2110e7c1ddqRotCtZblKQCT
OqUzXoeMPmBHv5R/Erp0CTHaaIyxx84d9QrpumdbV18Wqy9/z2sI+Xt+sWU5phsza1Y1ApiHBk9q
fwbWnTdX7bslKXwH3EdAG4p4QVMP/2mODhvv0jHeYm89deiAavtdbGfJlbj6oivgSzkJRJ8ohnbP
j+HfCkibXm0E59ToyHs74znjZTKGDMbHh64JLuqesoe83oK8aWi3mIxjeH5ykE8tEAFYBouFDOqT
d6JVaxlpxfuDeLzmBrvbgzhmnhyoMJVc0zU1rNxIeQVNGfQCz1xk2qSzMlggM7FmP7REOfZIgEJn
4Bmb+Y34YF+YNBLl2sDQU5hTjT4ByM2GXjiXho7YT8mH0MREtATzBQRmvGOCbO4SBoeeZw/DDCTc
VUjW1RFPTUxTs+/3wIEzyttASXVQap7Ya3jfDQ6SrsSKxRDRI42WePH1gsxDfr7Yc7DJOiXzXFUI
+CoeGN2IhaOrzE7sW226PZt53UzoGzWMYsQACoaAoRMnQuRtn7vudhgDhZRDgWgIP5fBPw28cBdK
bLU0+k7W206Ysd6THyNFLrVyol6LLqxTWZTKsyM+EtdFQeKQjPeOddU9rZ3h3zbf6o+4FQiKIV7/
fCoI9Q9O0oVjAx45nzHNh7F71y0c/mfjJ6HxZxKObq3vPNRD6EnyIAeTivowoUkgNy2A/GEYvdve
ey92gYzWyf16cLmtjd4aIa5ZYyMO4Wnal1LHk9CzDe+oswDGd+doNd+1c52JjjkJ1nivVwNPR9R8
k5ykgLQYvGkwhOtpeqsa8A8hjfclcCzZ+v8bOEDTwZw+I1AHKfprJ+aw3LgLID2a8jZktxwR8jHp
SbOFbyZkLKTpZt2Ow8ZPMyvDN3IUmCUeLOOJRag4mfaq0bZ19YDLdkpvojdmWUeMp1W0Jy6sc/th
GpaqOqQhRpr7Td1N741pppskFrMxLRP/GPaI5qgllDHRF+DJYkRoekSLwao6eqS7QQDmcpR1qj8V
GpbYJcoPOL1om36XjeS8YT33jPw+ufnWGpL7WSgWHM6Uf3+sCEnBZEfAUcGREABSs2Avy39FHO4s
lnwE3kaj/E5H2HrJWCm6aPnJP1a89GOD1mw7T86H0q2xh4YYGgmldcfjcxquN8Z+I+pTElI3lS63
ES599VoFueXL4cXKfHFvnjWBsfpRIsYms1HTbgbeQ9ajsMbrlAfKKQy6Po8Uq+uAbjfUOzbe2WA4
X2YqEowPfYytK4P8inlY2I81NF5/Db3NPRjnebCmoH1lX++a4YShhokjcSkmz+rbGqXH0vFZ8XA4
qADqX9JhWKEf+kHRUOf/9QmR9281AfCyeIB84sp1TLFFcYm8gTsKSDLwTBW78BlO9Ymd9Pn8hucW
VXA6aIAHmxPUnViG3iGnQgDTVvyDuR3ETB9p2lDN/AZgZMr957A44uHYPHdebJwo7XKvYYZO9anE
C5zCzkAegyVbfOxQz1Rh5f/vCPTDaOMnm87NjLAKEy1TRJ+0mBgXsRDfSOe2YuDCxBVKs8qf0FVC
prcqNhqNoALtLbpcjgDbbCqyZYveJ57yWQbb9y2Yeo2ba6LB5dvQ3Bg3W3AtQENhQwQ9cYLslAP3
V1NRiS0ft6RPvVK/TPBVGCpkeoMlevCZnYNVWNfqlH/nfcYMsW7+oHCmsmPqKN4FyDiiZ/Yexmxt
bRU4NZXchnj9S9rYZyYS/L2l/+Ie6EmJoQREbe1MIJZHQXjwmeDzOSKGNOFju0DgXnWKop88Hco1
8AnMqdLeEsk5NjMOXq9K8zBBy4lzlJDqJeTQDpGkTFV1Xhv1OfOxpbo3elB8UoNxeOpD1O5bdfN8
eTjF5VRwG8Khc4ESXjNOwm6iHVrQZyKRCbKhRqPakUxmdgvxR1DcE4SqWOt0FjeLmXYzWRTK6PEp
yYgiGGw44QTEhe5Z7pm2R6ExYh1ChixtWfSQtVIWTcuCkn8zCOZ2/ZbdVAdXW3LMo2DmwKi4w4mc
0rc0InRmuwv3+wQ8hptaJK6nr58sjzj5Ez5r2G+JJhhjoWdPNq2DJ16BE7xGQx0Cuk4ICdJQPwqJ
xLQ35FDqSFYutRNFoqqrYTDgB8RE2UVtFNZiJqbtPnsexipjE1SXAHyI16aPErg2OB+YKkCfOfHQ
RO+imHEKTtoqi7t9RTtzLHBcRkK5C3cKxudPlZlTph4Z/Hk8cnzHztNUIrn1/c81LvbqbbBxwisu
xPYs2dwTTq2expKgABEHPZc/SIjlDPsrW3aV3vPFjobKOtM7N0l2+vV9W9lxiKOJlwNXyZokmPQc
7cPvC/l0G2MM7Rl6QZZzoyyiHS+K4ceLp3RKnx7FeMHtdxY8Ieump4kRIpv0isld2nhEsQ9YfGh8
p66u5B5uFS2mFSUnu1DpgHS6vBvjKVZGk5Odyh2a7WOj46TXxqdlG2NjKDrkE3q4VRSRlzfwuXep
zwk+K3FM2/8LtjRyydoJvxv6qyTN0dbru5/Ldvutb7MM4gc0IRDjyIC48TbBwJdirIwfun+CJrHg
xPTD0YhoI4D6U5fxRvnmmEC3T32u8TNhaDiPUlZa/wtyYRWjC6RhyOQqaNINfxqDQ4ReuBoAlo/x
3A/NNtSCqQwGe6H48acIwCYaw3+h0CGOPLjFbnLkU42ULcXg5hPEDDNBLmujvDwjrnFAkWtCS0w5
3NXMxEmSREIgOik5wixFOyHcc9cDquD51bnhTEJ/zW1tKFq6Jc8DSt/NeyOBbKejbEF+zrz2MOBC
IsgQmGgDXxg1LvYbA2WvgAvHmd+kXIPa5OYAZtTcbFcMNRwEfUyfLwo+nDs/gwn0PszUKFF7z0VM
iCBRb1Y7/5Z9HZLPFX585BF19i0JrkOsvy5ftOfz44e13dtaOuXxNt40uuZz9euDtiPCBqMJBkcS
u2W97DlPfq6DGt5rqvyFiw4i3HomG+Oc2LPyf4IUhpLUHLvUllJILPRZG3PIjD3xg++sYx1Txxw6
Yi9lV+6iG1G/DN2r4W4gb7lhofHAZzzfCuG7DJBPbn4FPwQvByPJ3MLk+1yn1dvRDY9Brcgz/eW8
AEWsV884zkHMb9xvz6Apt9rewS5oLKeXKBmv9yrZFThX8FvW/jNihFlwoacvH6IRSVEATbM4VYpi
iZK8hthcQqp/LHq8kS9XmPgZjVuKxRxqLndxj3AYnv9Cll99nBcIOpHDhZdAlcWCqQPAjeIEDTmK
vgjhWVTwKPw53sU+RaPgEk+76wh7pAMfa0eiR8LKwuuPFO/Pl7qDu1T3DS8uezFzbmJhfUGhVyc9
juH+Kmu5f8qUogYknPLQ0+1hIZ0Wpt/yBysGTQR7Ekc1yRxSo6l4PxrrWC2ocoNfOwfXktWu/Rln
8gHV8Qe4dvhE7VLPGHVoq2NmmX5h1wlVG5FnRxyK0M1UgpD4QTaJIZS1T7pMFfy6l20m6cYRsPvC
rhjd2lxkAs3+8F5hXtuPuEOI+382xU68e/8YB0/1CqjDS/18WxJWotNgoCOB5XH1J8RNUvJbgfW+
Rmxxegzlm7eOYUU703v0Yy3ZHmENf/eI25KMDJucf7VI3gTjwPQG4jLJd5ycFDYvW/iBwh+ZAI81
KdjRXFyCpQbywRZryoA00LX7Er8AF1AunEUqbfyiQq+buZo1UbW8vJp9OA1cJ7n8gedbGu/HY+V3
eMXsPiK+jxiAw1Dd+A1cn/euKScyHwKmRiORPBO8oVhNi6yxKkhjanJ/yX1LDezVOQZyqV1TgKAy
i70R1/WzwwtCUF08bCnPkQb+cjcKOj5YAxqLWSxVlBkSzVcJHsQ0BXNEHbSQPUdZo9b/sHSQlxqN
LwxUfUuum+bCb0hDiCCATA6VmlM2Jh8WroFTNEA3A6s8lxdWhB9HwyOURx8O6Pb2nmiggylitN/K
HYVCiB14Ysdpo+IUhjk4y+dHd9xipvhZpFP7MEhHPuHA4FYGAHO3oMnd6s+tedlB1Q7nbW+infZd
1ABxvN4ydHlmEq/wzvwpwcpZUHC9Kj01uQULD5gbp8vU5kBQqF7BaH2XAM1r+/5H6+vEsRrCktdP
JMWlCXBaQVSTD7uoCJPGA8b7sc0/6UqN0Dn60d1lZvisk8ysTTqQJ+mTPVYDp95HX33hPl0L97uz
oun3aZ1JnuCX8XwrD3LelAO3Gsk4Z7OxCIsyn7MoYdI27nUAKHw3QXtZVq+l1LvUU8S2UztR1gc0
OhB69EQxHzfvxyfbyddU1oZA2mGIZF7QiT2v2HX4OX6HDmUglYn1wmVtIFf12CIN138OaVJByDsZ
fmkiD1xzopsI+9VPV198afaufIVESmUcFXxhusJSN+i7gENcnmjuDwX1Kxvx/k96OCWBFOb2OpqU
t+EsZ2OEIIFFS5NKtdtCe9f3QN1CGZhSrabt6e2G/hz6VvxNRE1HnkQtzHvSgsPU8LxNqxc/7kGZ
gKd2w4jk90qAgD2dN8nwAuxBHXzuVSq2byGgduMaF1XfRcn9NNuB2IxNGIkh7lJh9ITcmLIeGSYV
6CxfaksLa/hrEY1j5VJzOT4/O5O/hWe9qm5oEBPXK55jdOhgNrn4Q6RIquW9d1WmEMDA6rOlmZ6u
9PJ1gCX6OHU2c1gYPKzj1z0PdEJrlCcyCfOo1kqKXYk8YPLyLKfNyMkxfBuAWHqCtNeJNCI2XFja
BisCgseRu9l98QWYJSwxjfJyepiUeSzlA6aQtomPf6ZtIktnEe09gZ8qwsJE7yk2gwby9VThZ6/z
GXvQNIO+8sSh7v5A873COOZ8rWheZXellpn7sgtoh7pGcwzMVlcaNnqWVVMSfnvdlO4XXxEvqMY1
NhxW0Y0XA4lM4r4+l+9pZS8oJyngtnJOll8r2A8LlYn6oPsaUfmI2gh4S+VluFywWM9zIt+mA1Ar
y0mVT6c9qFDWBLCSTmLzBpVAFOEi8d0tMyujTXSxvpgOJdwWuuy5ziCfAwbk+cCQvcb6fPjVcdmq
IaGnT+BGLy//Cg9Gphkteb43KG8nWNb3QWmYWy4s2gWrqe9gNMkpZJoOjW7MNscQx1q6ou7APW/6
9Q1HmC/rK1JIaXt36S8u6p7OHHf4yMx9V6OjvxvIdWFH+Wn2lzdV+XhOFgLWSHCSes6ADI15t9Oo
a9460H8N9osy9fjhUZZXicTOdQED/P+3MI+nxDURa7D3NKaNZlVYhE+J4BPS8w6mIhr+3NjrnckN
lCYWn7Ja19BMJ6t6neujONHurpwcLLLFsgv6XiUv865eYcxMJ0RTCXV5yrbneuEuXjcPsvRTc9Hu
ecLrCME8c1vwhi+ScTo0tUdU7CDrVomykh6Y9qu0S+oD+XZMYwzIsFnfMP/l0JMe+bN9eazZmsjG
hEWH91oH6gkOwAyXB2mr74VxyFo9evDV6Z5+I9cG2NJfC7SHhkti3PxEvNk2PlydalbdlL1slIZ9
YdQUhV9IbLGAGpVlBOQyq+B4LMDlDGtmkW9/uB/xZNB4HKadctV5FIWD3/uu7ZlqTQsioOr1kCRQ
P3IwvyF/vX8sBjI6MlR5+7wPVUooirIrO+3+598UdQtHehQpefOVdyze8iUTi6dhY7z7w3v0KrE3
Vzwh/E2nTZDTrs3ru2sRVDESLY1TUJ61zN/cB84cu0MQbt/eZA4bk8Mk1F/xONvvRbieT0IWotys
zByyEVDTuFqVpqvRs9zpDUUck9m8tJXld6shA0QpEScrRm3s3fGgDIPEd3UCwPH78xdomv6z2O/Q
hkW3CT/FjC3jt3N8SDr9QGcYPUaeFaC323Hsfxhjk1aSpde7S+QYMUcgc1dTSSfDsR47rJVa08Av
sxKLuPuLDzy2uB9H1pQprzpZg7ZtJx03or4GJybFst+0IdZWGEyfxnYHNbbkNGWZ8h+sjJz51psI
mIUTUcbN6caymOSAfsFy5ajddtioLLjSBwwXWPPHdUH3/poIUIwl5xZJjXjyQrLC7eBbDeop3yDR
Ju4CabqhlKghc6wRvbkMX7Nw8pY8oUv1LWHvLvcq4xFXJa7UEpEMad5sy0faUCkUBjBBzOizEMAu
u8HK+uTd3evwflrc8mnXbXUhIleh2+OT3E7JiO1rTXwAn2tWsPrHPKND0kxTK2OkbgteXjqnOn8d
SL53LH7oUqjcB5PP8pQ2bzaCx7W4RfXgp8f2jH6wCNNC+xiwSTy5thM06grXBS013OMWwqmzwkgw
Ig78mO3GSrJgfNwmPzkr9HswZC7XKBBg/9mTAieF62gZPOGiZY8akHs1lKAaXHg8/54ZgqNmVCy3
ZTFPPAhTaDCXXt2IZpr6S0b2Hm1RhyVgP2O/6W50caayeeNpxPJ1v+t+UjoQQuet7KppYsUTYEUq
eKd6DlkRBh7HNWzCTqq1zRE9VYeVHwWms4uKdAgrC0OioyW2DQH76wSsDLziQSu/gPLGsUuvYZeK
63jSiha9sTbmCwYMsFifBrMHyeFrwnotVcm5avD72Usdki+vxDP8bJ7x9gCg5Wthfvc8QnsC1WH9
GT0Q3sByzgHybGX+SN1HUdIzIFwKDazfJqXdZJnp4TLuv3OXPk0U9d8e9wPWZ4tOTJaf0E4JZeau
h4FzFluGMGIyld65KmAixcKH+WWvb0yM+z63Ew3y2ga0m+G1DiXHYX1ZLEQMukn8V0k7KlvniTwS
r/Mt/QnGdfatnZTYuel6A2EAtBvOx+IB7DnLzOXyctXErM9Z23b4eqMxSBHb6GLN2HF2s6WjB43V
C3fm9MgcBdRrUU09ra/wLwR3Teku+F35x4QvIlJqqZpna1UYaTdPdcJvc2wUnc73IWMg+l2B8RRd
PhjbJ+aHMXHTcbvCUG0Mrz56iultL9TojuM7eWfnkeVD8zpvojvU/2YHMkBjBYP5fHgMxp9t/xqZ
4YEj5jv90bXkZVh8b4aB+uxphEpmFBVZr04Jzltkuc8VMBNOd/aWpPWkUIUvtTzR3xfcAEkXxtAp
XUs1obdqaxWcwC1pPM5k5RdoGnoiXtLnd425IXx2nkAEmKU1SLh2KthHQ4hkXuxZf3JpUuH5HXrL
scZL2xVPFBpw8ctqzEv7gYCEodJUMJVMvCQ9vo05+oH9DBx0se5NTj5PNt0rUZcLp07GiRA9LiPV
A67+BM2vqr91swxCnPjLUMOTU4osFCrP6zlGOZ5c7KmBZPvvG9WD/SFH9z8u819BTl23ZPMWG90G
1EqtXu868EODjoMVmqgnNsSPWjvj+K9Qaxge3cB1RXXeajsuTRlqFjuOTmKYcOhS1+++p2nba36s
hqhyeeomlp/17K6b7E2cNYb2rijzccptRP3bZMnF47UMTBNcchfTuiskg0hOXVTqMW+sWdfBzt86
/bSkDnQajNOyn5uTj4ObfhM7HylH3TsUcJBS+PUMui6ws7ysnaYJaZZ+L7sG633RkrkifZ3ghMHX
xZD00DkIniBmWhun9jAMou4Xy2zz2aXor1YPrSFxfepHuWHkUPNsqO814ahZyXUsbhT0Fx4YmSds
gmLLvXUDTkgaQaGAPZrx1IuMioF98WGJTUOnQKrP62bZOYgWIe+qTcQicuJz8qJMX3zBVC0IzP1g
x3eojIGE6UJ45folQnbNVetF2YKf4eAnrYuHrtOBtQ0kK+E2kZ6r38E0sVkfEAfJTEdRdrBx/W0M
WM7Rb4jboYtSonXajNxR2X4ApTniEWmbXJlMyvz2X5x5mCVlFdeC904XMKJHMsk78s3Q48pEFcgH
PuvRto3XSCLav9x3VnQr5pT2tq0G+HlAnnhQk1qCWA2qcPDPTdAb5aCqn6GZKXezwiAMEYiT2hlO
i4t6qWm6i4WFpwl28ArBhHvL2A9lrWwn2kpxkORIKduWA8/irpvQbGyZ7hUbQIZju+Z+iS9X6PSw
i+AIJgYH5zt9LY4jH89mGMKTjfDkFv+lkdrOCNZD3XbeecoR2rpmYImniOJLqAg2rE1+jpySn4Iw
o6MnahbSXCLZ9G4cJfW/1SAvtiR7ILoeIqPw2m3IU5NDGCBfXXL8pzMox8KJ0O3NVaLnfRsU6cfz
aSHsoCCXyjydODN2ILXP6AIpYr1bdpenGl92V5V2KBiP8VXXzcgC2R6JbCMGpkxQfEvBM/6DZCjr
3DUuI5GBQDiT62bk+RLP0Y5fsF6RgR9TTfZmvB7Q5kL3XhWl44n/ohAzz2Dv9L/l85teL/dR6cXl
36J6qRgLkjI4vXRCcKOSrZPAUR6M2Oe1Fsuq2yflBSDmocXISDowU2pSPmjipwvUfvEIOEc7GYzx
7cYcViQXQ3dKqRZJdAx4YCp1EC6ykNwsP3v5RFsYyy01Q4x1AyIlz8m3N04zerXKx46C2M+UG5ZI
gx6EsRreu6uj8ha4efwKB1KBnFYEXU8LpvLt+qBsz6PpSGowqOojuH7OOfq4KfRlp94vnHxUSCB/
8itQv8dj/sNNjqGKLCiDFMPWylMeO9pv9YMFcDuiBWfSiBu6nqO6qx8Vl7bgt2WnaUBKvIJlY3SF
7m2QGwnQgLwTqUsH6l2hlH91l5eAZfH4fbxmfwBFhpH0Bbdhjfk3Xt4EHl3fViBCNQZKb5+cHHfR
frJ1N9QKXJTU5Jd2SOxSskc1TMlAFGEJPgxwKvhVZok3D2hxq82Moj8xao4deixt2wPphaB/a3yE
GjcQiOA19Qblm8j+Uk2OHI5CVS5FmWXhx6I/Slic9bxMzcvHrDoWqU9MzdP4pUQ4+WppqpIHUF1N
BbIbKVnSns6xwt2pSgYhzyghbGINe9iZszjfQsG1M6X40eIbNhLcQd54/w6CQJdrNffiNOVd0w3Y
GwLumwYAJQ7HQkrNVgl6cAzSv6A6ieZ0mZ9jj0GsBWfPW4EgVXiTd8zcVkLhIOV8Iwpw55Qka5QV
pbypnUHnuWzk4QedbvZYiUrCaxooYZ2KxCdTyM/4Ymt7r10Bd15plVK+YyFX2ZH1eBNpv0z27NQq
gbqihSaD9JGDSZXqPgdkNdL1HsF0FEqDDraQpjYfcA+tzLVD2IpvUqvnvovkW8x1JfRn6/7mHIgg
bUPb3hb/MT3lz1YrXf7m/MkAmd37poZ8O08y9I6Le90lQ0kYv84+fLrKs48wMPMrtB47xwnu8eYb
mjtAV6ONiXIZyZ+lMnYXYRgmGg6kNmZ8h/p5F7NU5ddIjG6GhXgz9qTVgUzRX8YQRXOHUQTJjMf5
hTr8r43wzt1b5go2IOtatJCqXblbAobjpTlTZpSEihi61ZsPsoFosm8NI2utPwDUQD3YWpMk7mjv
vQYhY3G74D2nBcYs1s/E1AtpWC01msBv9PtRKu2vuhcaTwROiPv2jADKYYYRKGD4Qe+mMNnzAlvN
WXX1LUcsM7N5ktOYVGdqyb0mUFchAMbN2EgLKOqVfmobQCtNkbCK01FJq1dSHCvGKUKU/zwJtQIk
/Id6lNMgpD9GhyuVujRQAKJoyph0styHXIc31xIS2bQS+tN0+ztUAfBPfSVnaraswfOJQ6bbCBZw
hdOY77xZRsQCyxVlzuctLrIwSYS6STJRwsyau4nBYjag4wtvm/nfENvGhIRp0NUV2s0Fd3t98qjM
BXrlWjplhrdV8k1NMS8hlXp5L/tPeC+FWoD31agqZCivGGHCj5OVxdvUt/QdM+khJMmN8NbTnLKW
zfBlmd+SntdW6mRlNGhQ2zKMiU8iE0zBvyzHSWQFJ7mVjF7PR4FHZuU2QM0kdBdLUADZTZCGDu9u
cg7aCd7CBSskUpXyYeV4d0sYkQs1bnTIYIvNvZTV6mfD/ituu/5E5XhmbyCIfrpWsQ6iXjovNYMc
+4iOXBR2OnID4ZTOf83wJ8sZCl5IjEw8ATarmqnuLih17oKhSkN2znAUqI2VNlAnEuz20eH53dxu
3F2sslB30aOkbe2RS2BM4mbUQPjSde0Bsh4sJfKd/FVX7HiCATZ4Ct6cdT50q17W614L/QPWieMi
yeBBv2doG2/vbFefmR3/XEIoTzi0U3Iq9SSRSxmxFCFnlNBPgFlBjo7QdkQZC2VpRFBPTApYkQnq
KBpPD7kG9K43R+qLQGpzCrS2HjSV0vi7zT7OEVHDxhB30oBJpj2NQRj5oTcwvvd08oUkQTGZpmlR
sO/pnJD4GFuFdMZnJO0ewkcmeLryydPtiwT+b8qCcn58OFV9n1ykFFpfDBYYLyU70P6ZnQ1xmi2I
EC7o7+IKBtWHZksU6qMNOO1e5xnBh2Zt6zgYKfDS0f1nXXyiO8KcgI/q7s4a5EUWRYN/ingxBH0l
+eWgxa9Eg6lN0pQ0dxOjX/e+poTXxdmBpbjtkNg+5nmlT6klxNBx0QQ/cG2bEHkjgFnBsqdGD2Po
ZdiV3elqb7V/tx/2nPyONczZmoh5wUmFJz/UY5Il7LhOcY2SWAHVH7HIVSsbx2kAkfZSIPRtaZ2x
Wl0isxfEA4QD5Zv1lWlqMeYcVdrIfv5I479S9cIS/cmhbQMD2bu1N0kX7APkUVmUgY4bQdYp/xYf
pqxbJRi6gt9PNthHtnzfYD2MD3nsEI9VhLTRmSQkVCSjPzjvXTGW8JwEfTCYBDYlEldAldJ4rMMg
Zux/pss8dGfBPq/Jg42PD7ihQ1+VxoDRIiPNKxNv3R8AvF2GeujFccmAnKmHzuVjEiyQ2j1bFCLn
jvKdyOKoXzla2j4CrmlJge8hrKsle2Uq1056LWpII7hUqE80wXLEE6MWRsW6RN6USOD+66SG1k1b
+tPx4gSGmx7PTTf3q4ututUUcR/FQObE+2U31exRF1ebqv/8v7KrZE5nCVuCMODqBvtoQDaR6Dy4
MKwq6wA0rUhwR05kuVRVhMuthQJxe2wTpFocJHHP/ufd/yQQyfmWJRu01VuPNulDJMWw4eVGg87S
oW8XjEs3gQFFpTAnWhACAWcqG2tRMVR/9mMLnbXlrMHLFs5ZXdxtNzA6q+pcsWbAL9VEGNm1uu44
pQKhcwgfdmENdlgncDt+mbDHt3odLrC4UArqFMSVhKF8b6F53+nSigqxn/J6txTp2ERqh6eG/S+R
OU/k/AxZgfBVDIsST7Y/Jlc9LqvrzhWrDxyXsCPvqytUtNt2qjnnBDqESpumgHCa20TyCUqqJChO
+OYl1qH6Au2melAgVBgSolSje6ffwn/PQjtsHsIkXCSE4QqKFCXFTIDI66bWaDt/VFLCMWVWdWrV
fkd62doaZB+6gCU0wGA3rgjTNnALpTzDqsC6KJXU3OCFzgL9n0ladLBsYtpNQaOjs6MFXvXgpmHn
IpeNeQ1XNLe0ZqX6lxtb129QjkftSwxXBu0gEHTx66aZHO5WZUr7YGYQUsdrsQRhj1urJTz+6lwR
l8D1TL1BO6dF1m/2MLOZvLxxfoEunAVcOyU78GHqZyp7bxwc/JVv83BYuO2vuPGvPxKb5HEpZILU
qE+XPEHGf0JuwLZT9byA1T8xvgv1lwZZ7v5yiq8FIJu/sd5CxlxWWRDq53THiwO5yO2wlO+ZhrMV
fllB3sXA8YA7osgy8+InyxXTBE0ZwG2RzAgBg/UYPsCmxVNC5g7H7Qt042d6SrsEYR+wr4bW3Fdf
MYWQxLdGLQgmD05qTryYdH2N1ZIp/RGyJvk1J/qVi53qwJvChvCWC5I2YsSXxh2H1L2dYCWgZdOq
F54JuVxhx4lrNtj61sJAt5t+f0ImszF1eCru7IxSJy2NbULwOxQeY73H4orA4yAoIIGpykn3pRu6
PMJWVBz526M14VMy+NrmYIn1pdKmh98scsPWgHpNrR9x/sLJB5qHnca5EWbgH/WC1cXB8gAOfz0M
Nbol0gnx/Nz8q08g8y5EPxOY++3e0LJn8gCTOA1Ni8LqbAtwHJ57kDJade3deXEoFNJ5RPFUDaFk
pe5T6JFbmodOSZZ8K+VGsqQnVxfd/J48H9/h4LS5ryHr0Ui/QbEsCBvC0Bi34bh41+NS6x3fQ87a
aW1zOAKkSemzx9eyUdYo+bCsVqOsTRv7JoQVd7DEL7sqITX+4lh0e8hCWu8eSLTZBpSihP4pDdlY
GcFcQThh0tGQ6Hl5x9ijTxqSUzQEddxqdw5eC1GiTLCc+cqRQbTZAaBi4sWcpqWnqpPSkTMv1i4+
f1Uv6tohcE/U/zQFpD9Lk8UF9sBAqcLt3wkeNc46v3pHo3chrRBo9GEpVyvyv8TE0Fhxv8wRCFOn
ubyKFVjgqRyOvuaoyUfvTnNT40ITp0bJvey66T9CHea/2ZgI92qRnvhcSYuTqhyKUJ3hmJW+SW8M
m30DeUAv5oYoNEykkmeZGqYPgt9ZCyKwRDWYUtmX8uikga/2MTXQSKfUCADkbsejYA+T6RJjTf+C
giUPTzkMjm374kalQAwi+fh60vRa/r25iexOYQlXHrmjoZLibwpkk9C3fRWQSNhPlV1PVz0gz8CX
rKy+4Mmpp9uRX+C3GMB+ZcTcMMERM9OChUSPlTvQBxUM+QV4OhE7JEzba0MeExiqJWS3SJoBSBNK
5+uo3KvbZqfT0OwaJCtI+T5vo/U5prPViYFVPCSPPXApM8zmPV9MVD4ESjOBKTJfYLWCh8ooFzrX
M47RqlxiBwTsrHONyayyU85YSRNzTRxZV7lddwGqdiGuuma1iReZyGAR5HnQp//tG1pmWi5A0B7Q
SAK2XEGD2an51HJud4qEHzdaJEUGjdO8xGkrJ6iRbuUAFYd+PIJuJaWVMfH+MOgsOPX/xZVXHxZc
JNDv5Hk0e2QIazZitUFMPmaCUw4xrp9Z0rsBw44eTHRNA+rOkvnB03OwIMhxzdv2odZpyB75ojvs
HEh6ogvfvTDiYWJtGlUPq7jYEs31yat7pQErV4GW52EooJQVrYgv5NtoBFQQTqBgti40BknZ0F2l
p5jJk2cNqvnMuQ3dnD6q7RLBVB5CX6/iBxH5l3Q038e+CQShR1/DFm0sD5cVcoK8CW5cPiuTsclo
yxtRD0WTyoVdNX6EAIl8++ZDnLpl2/LJqjwT200p2LzHh9fv2yGOfowlU4yTs4NmGYjR4xY0OwR2
tnO5FvgdJKM08MOgOf4cRBsuPmfSRP4zkBBRBi229FlBFOrI4mXwcm+Z7NQXNwJwpRRm+zi1er8r
jv4gnm80SBG16/ijFevhx4cdItErvmyTpBej8npEACqfTXnSxI/4jIqX0bmYM3L0+KOrJZgZw+SM
QEpCm3RafAEOfPna+VCCBQLYk1tijT/KOGDCW7CDWqaGp3YA9cbnfDNOl9r+yUn12kWJXrGfqNlh
85+hIFAwTWFdld6JnRKl6Kh0wmJut1QCb1+GYz730qU7l024jlRIrpxSTMLluH0PlwL4rq3p7iUh
ZEed4RzzuX2Ytpbvqpq11O/pSnNvl/sFOUdspnldKMqzNiVZdUw1Jlz79XuNmoYEILM0fMfW04Bb
w1AMBspmf1dMwnHwbuG6tPiscPTs0I3RhhXYVHAiQ4Ydlzcb/fZzpMCmxlAC2IYqZAIVujMwYpNq
SgU2F1c0ijDZ6oMuxS3FF1emod3nhtqf3H+jDAtIgyEiCkRZD+i1OGd9Nvv9bI0I/QVitKWFD1sC
Ddk9C7CyAFWbbJVecWGctRBsI2we4K4Kg2Q3KBMy5TfYb3BIVaAWD8eurP25O2yTbkN6Yaqp6kHi
Y+6mzyat/WwL7MLRY7QTK4M6f6wSnhgOsqHSHwofai3fEYTTrRdbFOStAQQnUpafWuR7i23mUkDe
eayQQ+9HehfKt4gufKFe3GjoOTHZSYGSVuq7WfomPufARfukSBHvFB1MfggmIpWnVqKKXOkQ1xBI
ldRarUUquQrHNka9Vv7XawKxI3DRNpZjTwtWuCblOWTtizVyR5J2vSnaoog8uImNUbnfnA1UY1Gb
QAElPSlO8KbFH894R/lHoOMxBZAHzcq86pBsblKoPsL3cc+DMReBCP6/XaPFqmBbmmxMlaS1T9oy
y8aGySO/xzcsHDm2HA0+4jOVO/pQLOU2B2tcws4cGzYMjBZ8cQdbCQzVsClCK1fduIeNbnSsq6hx
yg+037ciSe3ThwQWK9AOONGd/sQrAvbp9I/8VmkfC1MvPYzwPOLvELUyDr5IRA73Kx5hdhvAxz4r
5lMKe4Hr5+RdaCuISDtZcc9L2uenhxO7p1gFJfT8HfamvGTU1ogcYc6DS2XiaYWLGHKizv5Hwrns
Her/WQarXCJn0JOlCOQqVghg3UQCU3Vvstf8IQ+4muFAP/UZLipEo7vK/lEzhETr/KlNMfXzS79K
chNRckSMCAOFtTgO/SQW1sd/RJhC6FSmRipjgZ/61TPSn8it2+zpaK4wsukxmcN9zaXkfie+IfYs
XX1iKLSZ+NGUozT1nYWSyhan80dJiVFpLYUKfoBvie6vVc/7ulMOdamOTZAAl0vNrlE2TQofczc2
7yg3f7DZMCXK0pz0320AmGMSdkMwOZFcyeYNrMPAwPUB1ltrN1iVm5kmv0PZg5kE2shE1uEyoLp6
LsekOpC41t0UOKQZJZhgrZvFpIa1r2383jJPR/T+yWNiocTjkRWotYgn+iHITqW5O1yDUOG01GJO
dQ2GqES+xhZZbCUtd39DfrygLjrCKZAlaeOGI6sj992alkYkorTfFgFLleBvwrv15/hBTUzWfFEv
3ivEjXIP9kEtM1dzhswT1nNBB4nwsHquGX0eks2tBDGjwf5Xmefn6vazWK114e6M+iy+lEnL8tiQ
tKSqUDYZ10ppQKXgAeiEKjeolzfXhc/aivVIXZ+tK4aBuhHh8BrAJsof5DsoOkIINLLj25NSv1U+
HFnVRxcQz7dhd5WLJcMMjJP+jl+hFQ8mB+HFYWw6AJUWQ+x7Khek1PfpsG/TUFMmkeL+IOSqlhix
4j9E2cVSD8CXDQdjyiK3qRfdgKHfNUKVdCvf99mShVqYu9PEeQV+uHaKN5ND74gKgefxdJFQmEiu
a5P1acIBgnamk6XKzvMh6YZ0KrjwAQcuoPknsRoHGTXC32+EopHNr5+G7AjCDbNEZZ9TsYEfi2QO
EWxXZg6s7AsNk3gkeD/t7skFensbQRvZOPkjWda6lbNNMiLD6IZu2Qb77QJ0zCcH3WK+Q0q0LIk4
8ylaPRjzT74BjKHZ6pDXVp0dH1nUi8SuICNP/xB6FDP+luZv3E5JSWk0OhCxrcjmb78eKcWusV9s
2+PBE+vqHF7YH7gzdHvttCD5NBKKLIjIfJeRmPiRiq+ScjW4Q/rxBXRN3/hYxBuN1e5m7kjyMOAj
WYY+3wenC7q5jTFJfSibzF+RhDoluSFklIB4Asf1Cva5cyt59LM/JVy0SJl9kWllTvbPkOql9mmh
0nUMQEFVXhzXjPeTsIfRInJFdJrtGOq+cUnH+j1drYihTyl6xom47z7kvxCuFxiluunCpfe1W8oh
2TX88dv3tpKrxSXgQ1Fjp4QQhiSycIJ39if+vNtkvjVxTV1rSgdUZ/ZluvBk71jnY3N+B3HeDMdi
3W6hJTPcPblO56nZUcosLcilcyX6zXES4soFRZHASgET4m2E63gAjQOsmEnrvIywgw6vgkHjdl4F
oPQiXAaErx12HV2Eyoku1zGVwjyPCwaZSvz+SM7zThBtWPJr3yDSMeV2Eehzn7pkQuE9rgAIEVxI
+WePdq+dT3/qVqih7yQHrcMiJ1txU1OIXMYA9l8d6lawwR/g9oa7ZkFQPRPFflIYrhZqYEB+Zl4X
FjD7gp2Q/2VsWEGcGOQbhyDR7f3MdLZ5MkPeo7ndhov7pSH2z7p9Y2rFjnX//7GLMA599ORLaWQp
lXiIgMwEQ0UfuGWgirQA1QDutstqYeVd7I+CZemtLqZ9/aV1xGwxQK4b+u8SRvH8JQLKGb6VAkSH
ACPzG73K6jS2d2Qft6zG9TLdTH491y6cBS+23VZgpmWYlDlxvepcgmBBNtrxkFq8YyuvlZtBmmGh
g7tMtLHJrnfIwMl28Z4ZfyTUgO+JH7WaoQ3MOLJLMW9BXssetdTDG2o4IETAEjKZkPRGbCmqhciA
H2jV0sZcwVswsFJHw/0RaZ8LqwWWQdv1PbJ83IApnW+G1950dQycAtx9dpOlAQoDX49ueuxX0CQx
hBqxtgaF0/YTtumKpEr43Ua5wYMEfX4J3juWiRE3ma0YVqirY9FKuHolbmL++Hddc2DasDEPXXGw
8YBcPgPz0zGMvcGFx30MsH2wF1P/iTFkgKGlov85+A5+cSdCHOxXCQJ6SYNH/EsYDyDvO71yFX2t
IsYp3HzxPOHYGP+6UGQ4g+z3EBxQuHNqrJ0vE656fsjpB7QM7Lw/GSv/NPp3hlBjlvQT/sH8jJpN
9GUb/UoJTfu3eAJMONm/TkRSo4U2k65XtXvU+8aX0/y+A68p0EqT/4zvlyWkebUqkLXP/n022BeL
sb+fVp9NRvFi3psQbi1V/7vr6HY8fKd/8GauzGjdcVUccAp2KkrlV2zSJlb5/G4wa/wsyMDllq+7
cDzwV46dEfAar7gEmWs8XbeOtdrHe/AOruCrzDB+etEFzXImRSeM7O7EiQy3xLcp2cTX/Hm0ljNr
oWfKH6PuzJowQNwKzAZswh5Au3HOblOObtjvO/cG3+mcg7M3b5/ShDwGWlbkL4bSLTpxOXKJ/pIG
a50PPAD03DDJrrd6hvjkqoPmfLybqTS+9PQCMhcLbbiAlD8hpBvIP024/Qj5OcEMxQflmKx3VVxL
By4M6oy3Yho+m1B8e/wlVP0PDpTT0cMqOHWSAVBdiEnZvecUgrICBxoyb2w+3hHp5l/T9XqZLuas
QRRERmLiKPu638/vh+UXNR0t9kjZt5Ts1KtM5j8rfWVF/pUjmuoarP7WfhxIcu0GfEZx/vbM3v+o
P+AvkOy1d5ui2U/j2g7Pych4rKOWVt8o4YWTE6fMTorjYZwitx09QraYI0gxtrbxF7ZgtNV/eUFm
oon3s4PRej8OHY3JovOBsvEbXoOXynzxHHvakRIuXb2kO+IvZhT3QBmw15t+EFAe+IJ34wgC8JsI
0vAB49i2g//X+LqwkDpgAhJ/oy+8ZNSpBSKlBy/Fv93nkN2QaE7SW7uBtoDNaCvE0J7uvTQbip7x
80dmWX0uwTWpFsXoGEuLX1PN13dU4i7GQaj3ii9Qk1l1ZaosaCdYWgdPVreiFgMdX5GDQPlY1bSq
AjeQTOMPzuTsriVewv4htdIgY/ttzW5q50GcSV1VrIE82edI9o2lofdUI4o0gnPTuj5LeIBWtZa5
6smAkFUyf5n64jq9UpqOFy9liWVomjxxK9mFJ4Gl3l6iiuW22WDL7UKg0gY3BSHsGtWZ/nPVBvJl
qJa6pS6R7O9VZ9YJ89QvWE4hQuYq0qoePUD3N8IRECluoxfR4ZOWoBhGgd4vnr4WLBrFrSOTtpC3
AG9jNaacN4ibCXvvrolfmz9okD6KyVHydWE1i8qAi1YWX140YJuBkZEFPwYimjYw+bTUfPH0l5zR
0Z2WRvpcoP0FpyAIhtnVBM3Pj6ABxofZUplHFMRj2+P+RokBF5u/LWeKThZN4F7IoN+l2BSN0qDz
sYt61Vpa8g6LKkYBkaNqC+ywq7JwaTkOB/PpUUrVh8rfOROFr23dC5x1YQmoAfSkBNS0Nb7SuI9k
KXXG0e62ifaYMiSL0kDXYnM9oAu1FcHfliBIw8lvrMI7+7UNlNMSv43frbcbHpUxGfDgzs5Iml0Y
nFxZ0WvbbYxudflK/6KIvuJrYxFZ+Z/FfB2gQWZNkfYvB2CI5cYHX93+s7CXDNTFQf0d6nO6T/j1
Mau6mU7Kw29SuZuxWfmiVR20tBZ7K3Lfz6MXyBZxQFzzA1SLu5Fq3XXTwjOV2fw6jzmFWZRLCFEC
gL7gUr4fqlREawePPnnhelIlCthWjUTpVrENTf8KlOL40AWr3/Uk2h4OqBu3QCAmlkzUrOIb3Hvi
toQu1BDn2ZeyDLYhq76jqfk1WDhOGiWgUND1okibHKDmFySN5o3kfvfSNgXEZfZvdHKoofDP1Jfi
/lMjKHOvlvwZ6ZfNshjvUopSCBxQCBRAM6nm4/D2psaxh+qqpd6mLADJ/BFJ8M/+c03RrHDFhMQ2
qP4qsQqQoZ2o3aJ8MxCFujF46jeBOmQX3tTaHF4IHGSpG4SAA0/Td6bWOYswNY8auDj0A7UfioM2
I30N2tX3QfMawrWYDY034AxoUkdOKyaBSaB05ppq6bGjErzEZD9+8F0zJ+jcjTeZMWzgcmLXPFZK
yGv+fA1weXbnuXe9cQCcXalYBWXjv+7XoGMehBuKkvEP9UsBZf38/oIg3KpDh9yRV22TZql7z+Og
WxUSNh6vc0bpZ6xj2a1VJP9sD7yNN8wHWQve2uhjzmxMppM9LyLGEZpv0fHRpzb9AR2G3YqKsRvN
qAx1zkfvhofNutmJth5UrR/9QFC1S7ST+FMLGZCKokyNeLRLGlEvAKNiTklsqBhpRIYGyfay+2gs
xH22CRpRzLWl0OOmpHjBxZwuZdTp/aRuzZksZwbAGskGBXBDJ+DCVgd1uKRXpHNf4q3dM+MtEn5S
uxjF396JiyLrcI+PSf8MAUldjQ5P60LY3vQuEcH5LlGtOJwwu8WPDJTrdmnG6gkZhl6EGxgZohTF
Y8cR7J+3Jj8Y6tfX/Acm2kHnwEsyFGQqa80NDspwi+ov7pwgwMiOHQobxKr9C2qS6ETDeRrlBd9T
XsokSR2Ah9dFjHkPVLhRN993OeprjEjxp0gRKD6k9keYPte9hemoE0VyZ3SJmhCPmL00crdN0Ybk
oFH/ZugIaYdIhrKhG4oABbCwEKwwiHuIPa19Ddj9kerJFftQZMTGjKVxie9qhWIKuknkW1dsNT1E
GVkM7QTEXLTivV4XKRWqkxLGsE97PFdSOoFeYTAaX9Xj436kCDfrWPYjX1kKYc/2l0ZCBj81OSLx
p6kRlukHMl0b1J97TkcBcA8Q/btmTVjRmg+27t/IHyHQp2sli4P4wHSXJmkY+WdD8kyZYlceHaLv
v+bt+Sd+cEhq4GUKH/WHlDBfAoPQPLq3Q32qGS/sHI80sQnINZlTpkE6lvTHqePHL2sqCj2gO/ss
Kffu3JqlrCGFgt7IKxO9P/8WNMFcUiTSTbVXVOZ8OO+iX9F52x0UtHbuAZvswl6Lcw0fA8AH0Ctk
cbT60h+wPquFbPhu5phEP5Kdr8OxqeEh3nrPa9IXHpHWDc2K6t/5H/FW1EMeFgMcugRchMBfZofc
t/+zJqz/KJ+36+NxEGsBaJREj58PkZazZf8mOsH/4gisAL0dAL3LIwBGju7TqpqNhyS4bguQLFOA
/Ocz8Q60Ce3BVxDjU0cHRFXVvqHwXWtHgsOJE8QjNNvW8HwUpZZQjTwvHdbNj6FL3BKL4e5+6cE4
3BMCtNiByUXFPql52fHL1tfJfrYHALfTUj/I94TRrA0zxBL/HtJr4PaqJcFLhSVk+h8KpONIBkA+
6nM9BjtBing3GeiPi85WYh+u3Ckk6VsB4cfkF9S6+i2l1Sv4T87NBUAgxzuASQ5ISSRTDvI2chiD
BDJHmSYNLtJPuRXlS8ywT/VF4XqVpelLjvCbC45V/K3TcHzHQZuh2/Na6f7wSUVpvTx4HmP+nSo8
fzMa8uyvJrkvR9NRjv+R5AYegMC77bAE1WexfQrjjlaWt3XbnWGsCuBpsD391DBNTeDm85KaTuDf
F1dLwKFgkN6EZiFxRW7LH80clVj5VKZH2bYDOwajgHm5qraeC8aQBoanFwPSpNaKB1rXIreKEvI6
wLqmzf38mwmmLe+cvtYCEjc8LBfGdskl731X7LQrQMzdlpwA2ohXWgEAmo1l58raruOuhojmZ+qp
ylAKLi+5WAvw50hRPHQvgYFMvOgtmP6CKy4biby5A6fArncWY8q4K4pLHudz9gAJLZxlEITBVXnq
V45dAjm/l5qPSBQpp5mFrEdJKs8IMiGlSc1WS3BVCU611ZB+PqZb3RLNWF+BHAgImoWf4PIxzUit
o8pQBRrG5n3kNrvfOevewEB9aMBXp2Jg6DuDL89U34zbyptXq6PjbTv9bl6GLcF08AcZ0j6KNUq2
hXtGDNrkNexaxNDDoi3V7a+kBpC5cY9VopzGC1TCihHtFh5ljVAiE/qkv6vNNP9muJ4zEIHzQRh/
kIhcHNe8sAeVAtwCsqTzDdO2wnakktfLzPu7jYabadpTEMO2grztmctssXI62qvLQ2na710rB3gs
nNGggWjZ/5nkoeIZThmfU6X6TvW9t6P/fklTiA65BGp8qPZdC0ris5p5gLGte3VAGVSRFi2eI3Ve
9Ab9MO5gjNERcy0+2sLXdbKpa37vXe4wQ8jcEA+eMPLIwyb8Vps6OckikJdp0mCXeFX1KETWimRU
HlsZmvPRi+HTXYMsoz3PJdOQYc1v+1X0oF6rKyy6alipFSnTVgybh/WzjEnvl/tWbTSadXDoc1A1
Ake3T9RiZ8sAp9p/kupmwnkdFXW5EuQWOaDb4Y7v1G807HIZ9nvRvdyAH9cSYFu7pa5QSxutoHoY
fpo/sktNZITk4cgS0DHa0rLQZtN7PcO7WF0iflqFjisg8BE4LZ+8g87bDx9HxJD1O6WvO8iqXFF4
wSkAD/pLy/KeyC+YHC2F9dv4g0XahgWDDYu42UrUi+zoiREUjduULOVb/zqUIrDb2jEH5uXRo4hF
SIUXz1hRUUNQXBEZPls29pX/CdCKyHv/AsWn0ADiCZUXAJcCaJQpjWY76ViT9HKOtalcG0H27GN6
SopWUjRKve2rxOmK1JnK7B22MgdCvL7OP4e5Ssb9CALG7QgvltxeSA8bes4WuarxvZJiOJhg5n0Y
FMy+UZ6iKPsp9Rf0iXdTBzwufSjEJwnNOUxOqIO96hebb5qGbKI/1hDnv/Dp869qqL68vK9GWffi
QKSLX9C5DViX4VJzda7qTTbRg9q/WPWLOj5Y57VO3Z529TIm1JvvXxzh1Ub1DDDKQRnEcegdSpFE
+DMwGruLZ8+BhluG03OQGOPVii+iLXNHlokxz2YLSOM6B+f8o6e2Q6T+GLmR42nyhBDfOzEZtzoM
dhXGK/P46QWwwdQ8ZyMKAYqFV5Klv9sKIAcs7p9W5nJYjc/H8lBubsVYKG7cA+gHCPqkweIEthPf
cAtz0I07mnIDX0yVZOSuRj3kD2Lhz7SX/Fqqxe9H6PTFnJJRiNbp/FxH/4wMD83FwLflxqMApmrp
sfcm5eYufv359zCV5TF7BZC0EhXsxyoGXs6ITnEYIGYXlRVYD03WaMR4tz2i14csUyQvQuCu6FKP
qYZaCz9fLNSHDhLlhrwVYZ0zwzL7Ko0CIy1kzFPleJgtDr/WRFuruu5PwEzkQ71jVs/HANhQcdov
i0mNBmWqC2Mlq/HpccljHNmDOKPlTgudzYepuTYp4cxopCubzvqTPTpGOLrUuWJ7rD40Gs37elWC
ff92auR1+0gThldJyD2vCjrJr4FdIXLhqN2+wKOtZVMA3pjVSGKB6aC/ooSdIylybb6pN3vC9/SL
qXick0hqi94fWb+kWo/HqAEGZejwXCddoq1XRIqcosQrcIvAX8AfJ78kCRlckfyBZBszTtvEM/HO
RslQCz0cLufs7Vkzsij4FOJJNkakmC/V2JKMT2d/l/9QuXoq9A4SNsEf8iPWxpd4tyotB9bAATB2
rg4MmkNLOsU3uGUaNQUlMEkkh6RRiM+opWsmC34I+WvBNaK9xjdOhBA6lgManaQ7gywYp/8K5kPE
gxeGLyxNmzZUolIIhRclzVRQ6Cz30LYEghW8qiepDIgqv2tfyad8BrJTcHREfgcf5KNL6i7XEDMY
ytg3ZSBtfAuog0owYqQlxQ3Ow8lTZzuJIt4xSlBOuUfM65QYKGpoo+YlTesJTZHvjKnOlgVfI9IX
0J9LISrlWpk5l9pBtQhVrzj0Kf8HDFFUHtoMBY7phzWSctplBGuPhivRhY5BRjbz9muhS1RloMfP
zG9BBZnaI2T1+S9c2H+h9CqL2q5MrXH1dyTsKoPAlCc548G24V5XMZjjUinh/bMZsvQDcDEo9GY/
0zluNtmYPOeI5xD5ByVbUKg3XpY0omJ9ew4Eh9B89DsU9zVQlOpLlOP/VV7gOLQmaXjEMd27AxYA
lsttVGK1jNbmgyh3cELGxzFRh0s41qcaGcI4v+X/eVpyVgztSgaJb9yVnOBd222A2MLx2QXWtad8
qWu7KmfkBP9kEzkhZg6Shs/EhxLonW6cuIxZikXmq7eXP6r/YgSLRIfXr7Dka80HHILnrLIaL+tw
gwYJtKgvur5mAfEf04GV2tNQLYvP/lKN688Bgu7EcHkBBMGnTpWVPqvTb1tjtJguSiIeK3QR2V/s
RErt0yKjGvAbr4pUPvzPx79QS0ybed8uxBKdhEL/nYC3aDhyl/b33P21w1L2YB2eMJ8VOlmoj4Rn
Nv75S68yOCfmclySW1gS6NVsrra4gCaCsLJ0btJL0iKLZfPrWXHZyt1iRIts+HLF9nC5CqsGGhW0
61k/wFoNY8XF8fVmiA8mrgQpRdTxB5ZpFZOR8i0Z+AuwvR7g0jCtXjG6AsD/pbnjatgzpOK4a5iz
s4fV/y3TNTx+aYgN1qNca+Pi4BuW0UQRRH01hH9KKuar75igRGeR49zRi1UOClEvQF+PYkJJzfRl
mrq6/Jvut+dRotcyqRK9S/6hOmucYj4kZ6pLiQcUCNOxfzKlkfsaNs1IugMP5mGEB58FgdvJCV2J
2WU2FZiTW8KCijAgO4FFKtxkhlOda37jsTZCTHM1Dzqnu3FfwY7zeNMw16/jV0AvUz4VuMFgL6et
osO5fVhREcacagHsrGYpdkcQoTad2wLnEh/LSYWZ8gnGl2j2rCvYPFqWaX8XnNyyGoQRuGk00xPN
fwQDqQCeOURwxNzWQSqpJl5nxy5Ke6J0eIfme7iMOua4Bq1cXImHIOtFUymJxMouMaYP30KQld0w
/oOKtZ53CuwwAtjDuW+NLsPaZPuaxHoDHBGh0Bk2qoG0fxZ2jyFurN9uqEY1L5OiDwjbfAuT7E7u
Q+o8j+spHG3Dj5IU9AEO74joRtne5Gs2HAiyNIqzJ4U0DckxQKwa0CcvV6JmEJRm7ePd/1GTp/DI
H62xgx13ij9s3NUAgOLkpYqLE+VD+RkxqL5LflBB+SI+Xwv0UfgzsINYMgSS4pqu1mNOdq1Tc2eE
Vjo7+UIWvio4sPAjpcag9xXng4YaQyWJPMdmgpy2O93Wqo4mSmmFSKVCLRLef44Z3SQTUOwFvIRI
bng3/t8JuZzwio/TvKVV6Cx7WsqUWn4X4OYPqlCLorIuRLiHeJyainJsO/lvRe7jk54ACjyYIX4u
m6gcJLoCc3u9KWcb8FRWv40uOW1F55eAPurQSbUmb7edn7Ott6cQAZ6wcTYEWUcmkrcIy9RT1Wnp
XxNgKCVzIOFmroveKiu7LtaWu8BskvuiHAdCveKYwVS3Ys6Uoxj+YTjBGpNMj0GlPhBhy5ReMNqU
U2oFi4kucGAg/lffbg2gRJpBdbooYSIs9fOy1nS0jPgUyfeTwQ76e9Py/RDs7oUvQN0zbPOc7cOR
5qmQehDikC6dgNRg+2K6wEkDqKE2mtl15YyRPEC4aPiODexi/uVKBIuwGFjLJuZS8uO2/KcjIQak
1IUamV7Mki0RBbetg2bci5S7WQzXnUsthlUxF3PXmqQd9aoBj/Z4h9pjqZHlswLUScG8lk6g2lbn
0FiyMkQ5eaBKh+hOVFUtxDvIX92BFpchdHnWZ0/1B1yTaLMXeKTwcs38tPdqAaVWbn+YQGTfXjHT
8XlQ+8XqefsqaDixhjFm7FPP8r1dZAg7/+LRvKYw7qY7uz1612JCbuNr3ojwIMRS28S1eKz27RT0
Vb98Q3Y9VbUYqYvC+BriFRxdSFf0DMGbVfiK+bufcX0i7ypIstUlsRI6jrXs600pag+5LIL/4aVH
JeDL69AUgoUWEX0FqnS3A87yBfvuknYBKSIuGIoMmpRnCwaxRIObPxd56e9URqvdfLf5WWeSlZTG
E6WzA0A9T0ZXocxCpJ1PwJZk4sXD8z6POTnQkGi7JpSq/RNpBVVVxvxiDOuL1mfivbzSS30GdEBu
JCmwUqoEyr9xzdzJSA/oWD/0qK0Hif+SQRJQDE9VCDH9Xd7re8cweZhUq668J3MEyhuNAo7sxoLU
gzMsw7T3sBQpse1B99vxLwjf0LrYxyWRkMJOb9m73lJxLrdT7D08OaS4LygmNstfGcJVfJBKzJeF
Pu7rSk9BWKqWomd/ASZgqLHSqPTOkQJMQicpdU2btwp153jWMhIZIVYQyr7kqN9urYfCUBmGIUDD
Bzo7ZX+wrEzIqvIH1Hikk727NRxSrs+SAktLCYhP0qI2Wl4I6VATEs+MLE+a+yHi4SOZQ0iQikfP
j+jS4/jj5DqMWgwVc/AFm5Mi8nWADK5lgf+xtvTycF0DhTprrt2sv5+p/ZlX2N9lBNVnS04CNvcO
KsrYoprtWLCmo9M27ZVbpvDtDHhksiM565G3BzR2apnKlVG36Mer9+Qi4NvGjQ2DFDoKHatL2EYY
7wJ2D9A+07ovjrCpafQygrv3pQj4YdsH0P/RNAqqMWvKv+paekYH3DEUUf4mK5h2MkXPyIgZjq9F
um+UBBwAcTrK1WpPjmseZvIOpzLU/pxK30isCySmppCNyPTlzAnvQRcFWoAOVeH9QARIJ8hqj0kS
7bDX1Hymx/0VlNHOuDidIeSWcG2GTbtFseN4ATp/c7cXfS72ScGxW2TESr2dvPnGImgSFevS4e78
bI+AnTMYT97Lr8OgFkFnLPuDLqkz2eAUeHRqNrR8wQjz2ScrrjH619znxL/rgIN24G0B7Zn2bsRy
vysWYoajPqKOHzsrZm1/9y6uRfcC/Tg7ehQ2+WeqAsPQxWRjg1f1DQbiocCK5PJqkE53z/kI2yOG
YVKAqarfk5sSOl5Ly9pN2vjcotIY2YkVLUV0419uh0iZMlxkyAhZKWlVLXggLzUsCL2+c+WsKYnK
fTYUVN96MALGGmDm0pQ2P2Lb5zvsGETW0RxbWWUjNKjPztpziHcZ493p+kWax7K3GXll+DDANzqc
2GTRZjQzk0lHaXHGNMyyZ6MqJXUjPmNbDVca7Yjy9vD3ZILAJDcFMBe4r12/+csMl6xrgSoTd+/d
NR9rcqPpUAqgDJjOe1K+lLq19mPXVVthZxdTzoryZdNyz0xMaDwmYN4rGMoM1XArqoF/xgKxaTha
jT7RqgCmbrEWnRhLY+bJ49rYwRNiLx5+3yP62Z0cAoIJ2VRQlG2f2IC3Ng7IwbYZXZd0IN1wRAlI
KLqA3o7SC1+alcMMDOSY+94i1l4YmkW9FyrU/y+oaj5Jhkp6eP6sfnukufbQ52vnbgNyA8ePUeGc
TLk9YX6L8Zy38ZVV2B5T31CNfep5suyueoK8QImZlkX5LqVXapXCgYnuEaYRvOEoJhlx3+3XBIOx
RxstxxqMcBrPSRj4B4EH8EyrYf4L4+ZmVAgEsvBTjycj16anx05LP/H+KeakolYF2qkkx3hymuzG
wlgbbnvat2yWurSnk/w3KPKivVna6+x8DZ2WKEM06Ftbw2hexfh8BoFrlyqHDPHJOBuKJqKn7tQn
tRExZS6PNjqKwW+31KDZt5bKqmgEgNSnVDQ/dEVj8dItEQyMyZB8wCLbQ2fuVClbu0C4MfvRr5S/
v0DRQsBKQVYNE+sWhZqrbPa7qRg0cxL4ln69pz3qz3iWeoxEtT0AZyPqZiM0/g0Vb7Jyu/QT4S6P
ZGAywzhU/QHSZ3PgwfEretDr2tvtsxN+WYJsd0f4KgEsITLVREoCTbRWPHUh4DhS6CY/W1jBm0L/
Yhy4s90SDHgL5xFE42HeQGPA6PY+aUaBOofaqa06IbiJ6AHGxMedUZPOTajsnIpsjYTsrYZvtUuj
KexMJ3o1nud0rhy4vtHGkX8j330EFxx8AWBCvGw0Vc8CkJQ9Iz7PSxZP/9qB73LqhIh5yP0qYsB5
4m4SWDTyA0FeGbdgHVhMZhIr0tJt3VZyYleAwghDOBOksWIypV0fO8hLfA91OkUQb33taRpm2KH0
LsNWE+/7o/GtM8V5rjjrc8LUqNovq8Hm9VYv5xKkU6MZ68CG8OivdE9tZriqX8YDkkrAzHVkmrxP
vKR9eWFIoQIHe8C2G9LiA80dJcOliQhQw4vmhfrVGHSPqDC72ZhNUC2IS3xNjdvAQ4ytB8Q6aKe7
Okdjupa0vaK9s6hq7Gtl8VwzHk8dd872SBkJ+smL72eAVnkpCrIgvBpoIIW2/yuG2LoLapgxGD4e
q1gWoWPmjQV8pr2oGxGtmqHgD2uDOYuYxrMrA1YDqFvMZAvhQj1J5MRfvESODr5EqByvkLls2KmN
g+IPEKeTucpD33F5jLGY+/B429HlbL6KxNwmVJTNwTlaH6eu4F/oiLT2LimqHzD3FLTcOeSGebDq
p9z5Mi9j7J3r3hVErOTY7lMoQfrCNfnZC+46JEZ9/UbGWmMLoWu4ursBB33btAlNbtiin1KbhBCe
CqRkBVAQ8uyi7uXivpIjcSZC0OXqqLuKv+Z6Xh18/I/PqG2pZiRAFOwKSwwDhL+4dZMO63vD6e/I
iikyhRuOncqcGhK14DuOuSA9Zs0oR7bAcVvgIj0C15O6lg1z2bykQUic0xRh71XdIsGNEaYN4R6e
Eb7Jp8lg0tvit7g8xh5bEN6cEtSG5rud7aip2kuJK+9VvqtMr5IjjDhr0SednF1DiyfKo0VZZYDP
tHiQFzhhaRyPmkl48vVUfP05NF9gI1IJo5+l7K/703qFxHrYJWXaGkE3YGSPXixrFf9DHHmB6LEW
jqGD549EzlPVCBzciCSWgditgG8zR0QXOydBf+H4cC22Fc1MXpBUAZjxPDLZT2kewzBMWHAePcZa
YjFPJ2H88kpGCRCmtXbumegxIxk9QDxgc8DvGdX8iVM+TvaPw1tizeLZILhLwjHrDLFIaZCkE0TD
CQtATCCKHX5SPN5i6S41nI640q3aSnbiMFIrHOOTaBQMQZRYqvYL1JWkY3z+/mALP8/VNOi3QBZE
n/WiJ9Zd4mnGpi2RAaYarAYyi1vav+EwwN6nwJddG8KXaj6C6qS7DvJVehfjGiK0TQb/wzJCDy2K
80hTrzFdbXYsdMobO1noCVYJt5xTg/RTmcaHJmWpR4GDYca2rBpunZh9QM5tORD2b8OHvqqGp8nq
Yj/t9mUXQORHG+I98So39zpSID0jly/6dw9yupCLJPanqDgwdMaA9OfodJKgZi4w6ECSjmOycw53
WUfBeGBs1uEcJ+uGp7kUpSBWZr/ItYqJhNvsYc+OXPDmKd5B1kR3he2JbnWnvMwMQhmE39pCQqC0
XHSadY1GuWrQopqWl7rB3StMsxzhb7738/UoadzYUdpINIYdr2/Bu+oUBrxmb61sspKRv31DV41H
O0dNkeHs6wSKWi5EBG8TZUUhb4xUnac88jIRGG2KnfX3eEKoXVGKwpmlMYeD81l6fEw1o0e/i0C0
2lFqpasgF1teJBWDmiQic2EeXibhbwYhlNtF9+H5RZRGBUdJRLjykHj6a5xm+GYjRtXoe2MiZ5oh
ynM3mbDLrCpWpR5c3ZhhVXA4f5WuCcyFM7SZqE1c3imPTm3ojQ1hel8hrIX/bp9EKrbwkDt3v3Sn
6WgY6fOYjKtCceIUBOny0ca15BRSlUthfFuGw9t6P4Xnn4ryadqCj7MISp2Nekewf8Skbs1+yhJZ
v9R5VMvuduQb+QuN8q6JJ0tvsrFbB7QsBOGqYjctSMMI5X0aIbYuW/6ClDfpAlsQYZvd6kXGhcOe
LfW19/0uylGdW+wG5wfIGJ4hAijrVJcbS73CvzXg16mDSURuXucF6JoPXsobmxdFKQRYofYBdqbj
V9ICcqXf2stnUdcHD1mlzprfuOl+Or78FksVPWFhRznKP51r209YdPH6G/DvXLcfdvx/srCPevcl
qGc9qVyGCakpq93PjFpZCI25Nchfucn3nkzh6tivG+13j5Ry53R2hIaUM8ncCftkmzdj3HA2k4Un
pAy4prKygn8dYO3wUSurKVVHQI2A1VDPd8M+CHq24LtIXWxNuuJ5l2UzwqZfrDNJYj2isnJ2vfun
brjOziFhpMOmASa7+1/n2M8fOmH19kqOd7hu2iufzX2BPq9edjCurVPJGL7y6EWCPcwD46YuzZdu
Tl2aJ4rqeMkmAT7F3zplilq6E2nFA5m50ll5oQbVDGNvBlSnqUcUczEpa5L/oS4ltX3jHRQ6KA+x
oWPQoucwnvQIbSMJL4C/ATXQQMUHFm0Gq84D8if0F1nDIurg/fuDAfvyJuqmk6BRp1yio/F7XMXG
JEQQubNwgMzckZreR6skrTemX0zv0bmLzb59Yo+jzqFxwb7ye9ekxtT+PJ0CM9Clzp1FAKVXUrTV
kMyE05AowaxECPnFOCoVoUV/WYrKTxV6LvYfaS9mXfBKe4gr/lcsDxTJl8Q03SpvIx6ROdAOPa8v
HVC/XXGsRu5m4vo1smtHUJoqLgVfSsCRUq95QM4m8DE1h0PYCoP97BGyzTvFPcGGQY+cZ5XG5CzB
yfnT5tBc9ioXGipALN9u55Oo3n/hXROKS4vlX5auFQnNfdMYLys3QDzDwgY1lw8JAan7FPW+ncif
OKrdkUIEVtsqc6gCYlvhvUGmKrgfxfsiVFtYxPJVjLBO7QcBIHnlgrNfizFBPsvwVmextlFev+3t
57dW0eRi34Rj//uO7s08q406G8EdGHLiHGfPgcpi5KgmMeSWpX5HMDnvo1QnVJMh6zCna7o/iE0N
Zkgau7mCLTReKaSLN5TBiTRWqdMazLR2dEvjEDE5vtfMsWU4IVyAR1SobPuPcPEVSPXcpxRoXiqg
+9hrbED1BmVy6DS/MxZOpbOTPunfwU+F3bIIDRqxGeZGdPF37IFooPXr8B903BuahBVt2PmUsF5K
aUcXZnEyJ30+Nqr3YZbdgVtRZX98B/A+8QeGyWf1GKDuoBhRsUPBpoAiH+gQAWNE/Gh9BwlsFkt7
xZ2OB8YFRtuLBa06Cfs6li16LfTmi0XXE+BdDyBF8liyvLArWNy2k/QyaVI/6YUxjmU8ow3MqVvL
yG1cY20MUMPnKmIZFzW5mBtAWyweZw6tQHL8rCeIcL+ZubE+AVXlTCQJX4YQ5YUs1ayJK+0axeOg
HLf0pk26kXdEAqBQ66axAcyx5wr9BX+lrrtghGwsCQbduF32Au5IW8UgAONu5X4nu9kvBFuq/1OP
81gbtEtVvzz8Q3QSXOcuZzFKdFzgn6XLW+K/jiKsmP0JaA6w4+g1t/xLI6qPYNbTTu2gtjRpWBck
+hEN1vhHk0cycPdmzritYWWe5gdz5UhgXB3oTY7KcTIHWAVfkdOeA8euehVK+W3BB98qEtWGwXil
93ULJpDL8pKzn3/WLqTeI39Qxl4CCDTXvKmr/Yoe0zSEC+m1AhQV1wl6B8woSC/Hfd39GYXzDZ6K
l0MmHFI1B8mWouDG5dNe7KHLWQ2lPnfYPxXK2n5cM6Y4JM5SYCy1a7LwNYSo6QQ7yWqiL0ARJOAl
aEfoB2wCYB0qvxecqij2xIN3pPHT3otM+1/cydJMwuWv/bSyC4AlajXT6tEarTL5Cqd5t/S+oGGd
U0fhbacyWmDzTMeJHYDRx2S5rn8rALWjesXV2Q+DBndd9/MJc3cptYGe+K7vTraW3dVQzhqsEL3w
8z1ZY1c+02IldrnfXl4BQr1gkdl+UjZ4p3QC0u71b2OlOfppqcfAMuasTWuMiCtdAgDO204JQNEt
otoWHA/nnzOMTsEbj2q6ssYtngzoYgHcBM6SqTm7ISKKVv6T92dziMjrwn5ZdH0Ph7p0M4g7N87Q
s6aAwEv/Xi/zO1ax6RwXRXtisI2LGP5KqwfQkqYjRMWoKK4SGMQmtYKyUvLz1M6SU7twMuKH30kP
sXqPF5T6PMDEweOEUXHOLCMsSP56mh2AahZFMuL8wSJi73bKbL3ASiscmp4R0bJazljvc3QqI22p
ttt3KinelISLX/pEmPotP6RUcSuHJOAOvWE3Ufqy0X9kMrtT3yNWOgZGXDeCQMFCIlh8WMDBr/rF
7XormNXx9T7uTs7hrsWWOPW6JwDxN+ZcX3kyfyHgJDtUq5HAaLBvHXYlt93vfPZLvWLAONku6/rr
Tx8Si34rMC/m/dnXGaahVaNLBkVKYbY6XdY7bbNx7zQHuW21mpF2tGsXar1EtqZHFjAC+bg1ZXbo
xGhZKJiAR5IlSHIjaLlKKr4dQqeiFlupq9XCuRxdK6XOfVmwo9s1xvxV8EaOxXOEcuFs5ttswmb/
9hcq7Hlzw8yB7g/RNimdHqhw+KyrcH+BVQUq4d0o8Svj3Ygk6LNE+7gqtAanfn129zxvRn2opE3P
lCmgpyZ8cXcgmC9pGenusRyBr4HD/yJhtLBn8INcjGKcnO6EzkZVAfzzkA8jI4aPKDukoNKcV5ge
u/xdAebVHOhB6UCaDOGTVHj2vqS6Sb6omR8rmWopa1AX7DQDuXXvbqsUZpi86D05/4whSMA9idyI
RpEgdhhJy7sMnk+TX7tEWSjaX2z27iJPKgivKyBvE67m+Y72/diX5HyHZTPezFrD8nXruTSM56pL
jXqGII0Ry/VMDzQs70eRKOr24SL8K54C16oD6VakOa668gjSR56QQIPVX4T0gX1IybLWn1SL4k+2
bmgJLTTk2rqJu9/0Z98k+H3FoYknKpvlX2bNI3x+NXsfoOHDjNHNHAqDa7Kwy5IXk85c1Mp5jJsn
KZU5U20g9oUZ+fI/7Teh0FgbjzY2obsa6z2YcGjhKlnqlKWpR0X/faMYltwwpQAbjNJf5MkMGMkQ
Mb2iUftXP1czlH6nX1zMDwZ3U2QRh/xNEja18OBOCieek8YmOSFMG/i3zNWxs1CFCrvTzaM/3X0c
VzuaFPCAYOku8n/AmgkvVVTgGyUC8ZE0ZGjwXg7/t92amxeAREOqmLlfMD3PueDbVoUTCXBbYxic
s67JxaD1LQsHl79pwuYKqUv3SyUA3ILOEUt3P///z5QeX79h7xY/7MyjOcejKYmVKf7YZMXpU1V1
llxuVJy9D5yE2/FNUEH7snHwkM6RZ0wAb2z90+rBUBlxkQzMZ1gNgDifXBMxahtmKdHwYBqU3mo7
q3Wfw83epQjDHgwLMuGXdp7BCjJo55/KibWpfCSe3FnygdKtcFpqRYVmA5QeOOdD4Rp1h7SJDqZM
vtOn4/sRAHJRsrDe5h0GT4DMiDsw3GEKxxvYze9fF41go1dftAGhFW2a8aZIF2Zp/k7wIUJYy3bl
4V20kk4svegCPOGQMkpTF3sG8c6ps7wC6Hncg0FBJe43NIDOpP1LddVgDAH1iwYMQ2CKW2nkvIm2
J25nkNzDTywQ4USdTUBUy5b4P2IiecAyrGoB28Vm2RjLFKwvrL+MhBAqDBZjWQbZZfTiDvK6gzM7
EzZQ/rLiqX6nwXaK6tSbamQi/Qi9MQ9Nx9vccAu1P73suXY4csn17T7JKQwqArP9cpRhs5EhnO3W
XVkTwD1tsMH9DcISVLfAQpE9X82GPHEWSA1iJF7Qtwl7s+RsPcePnMOrkqS9YW+skAkAdNSAwHq/
iYDSmXmSDeYQYyfuGWQWcLruZyQe4r+w/pTPLDtFH0jH80VueWBCA+nbjIACXEMulcVGpSaCs3xj
E06mW3IRqhHO2kT+2KbJeVD+hYlfFtRPYlplqzIdAyDiRlste/vu5GfqVWchJUuzF/XB6iR9NysI
POYNQ42zueFfvFQhz6/eW/HmtBuO0SJyhiKWnn4XcXxH8J4Z3FjOa+4Y8bum0ntce1CYpluWjG0x
cnf+B0aIiQqMR1SSR8CThXQ9y8hBcdFK/rKdlYXxzk84rWmn86B3D3UwTiIxh2JkUk6IWRVFqu2i
Nqx59D2FXdJ6OFbjH1g1iP+TDc9QsORGNVgQBTCDOljS5I+20CNfTAviEvMmSLvgTGZqNxYvNKef
QwQd7uOHGsRnGeBqB1UICEuY0YUywLcIPfbPCP2Gzk7uI3c25N3gSXnyc0n3xjsihQf28odh66WB
xhgAwpzQBgJmzJ2w5jD5GIYaW4t90mdqFvFmZ8SNU1Puy/vhKr7Cmn1v0+zo7ds0HejlMer5KRCw
YzlPwPdrHZqdicZoLobq1aUEiwl/sDGwcOboB66q9SsScj5DrJJz2LeM+WjNvBeHpeKxsoJBKQq1
2ZU2eqtSQcuXrxIy5l/sHlrlQx5rui0bPySpKJ33I3tJBXGb69/QIvEQOE0viXADDAuo1KPF5b1j
3eAFRxyUTiDzM46uRb8aaZBcDhYYisdE65i3q0XzfoilFeIPKmu6dbCpyDMO0VFALNtqedwsGHB2
YUWULuztcUCGFUfdFzfBT8d9/Iah6an+3vmu4voYicp2oWzh7rBxxJQal/+t+DJGHm/7kHoj9aIL
3rWaFICpOz11wZ1i3Raa7OCa2IPGhfC96P4y1iCs1f7OIWihhs7lnhcYFmdIo3RFQsj5wMOwX9xi
66MJpDVsiJxPMcTrPRfYM0396lM5JHHidNM3V0k2/G7DR6299Xy0S+JWaxR5tO6vluMwDP9LnINx
da8UjL459EbTO9h+S1uoMZ2qyVXDCbzacSapusPGycG0M+VIpSUI/AS58Ho4EvNNA7Xaz6XmEmdI
bz/IRv7iTN6U+BKtLi7QNYl9nlucbU9WFX2RbjBau/ICWqyqRAZqDBH5vBlH9CVn3NtaQboURrf+
qRri8B498qnJY6nJmG2j+Wfkl4A66GqjfEYSj6Gvv90bk2BVALrnRtzyv05CcG+CkItju4xP9w2T
VMKh1qPgviofYnbt3vyxQRobCt9YpZNj6fGQ+LyW1mc/4l4BD+xpl4ejndQQ71qB8jljA+AX+n+e
EGWsl7eJC67g6HkmG2tyRXw5s82AWlqAB4Pn1Wee4YNppoB0KRWl9IZA7Kg8UJ3VT1HHg/QZC4fH
U2IV4fBsHU3/2vWpMiwBPZ70pYvTRm2FNfHqMiXZ2vFzTOJGyo0oCfcjm1ClKWKUBrMBwCqiTdbc
sTFaa46Flr1O+6JbCR1DoVlILqTfrIzY+YhONS9p2DyqpwV7aShesds9Z52925zK6v4IkpuG5Vsg
PHXaFXyUjYCEE0V2aSJU7ml02qzGqePXIq13XxoS0rRi9l9vtsfsyCinhReFajZY36XYau8tXVzn
d1Fpf0M7k1wnyV48Yp5RgyXDa+zOKl3JAQhnnEPt6E8bBjdqGZ/GXFBpZyDhbUsS1o/kUNJs8X7R
a0CktC+6GMztgc/fdCpvxpc0dCvZgT0AJo/pxtOrRNECdB3Ur2n0fD/GvW3m7HfWYkjxSJEyWPvd
43LUX0UziIfEKNaP0cXxYQAPzAVJhrnAhYwI5Oh5+MeXm67B4ehhboTCGoomOrDvE1m3DzWyJ6WU
PdLxabAh1MOqaBPAFD60wJ7BsWfrBMRg2fvlBB8kUxMaNRhXxam/fqxKsrSuM7+LKL+oEZMOYem/
bpdDYRio533ibDwncKJu6mzTjo3KDZOCt+3Mn2J71N3Ary+zRTH2Ki7PF/d8D4Uv7HjWDF+sY0l4
BuWYTEwlS3yMMCFf9o32IyzFph33u12TIIK35+cgEjncekaJzPutFS0iH4SdnqcGS6IEc/yOzvGF
lkQEBe7Rr9GigePT75wDNINIrD3ZJmQT7qkZ8i1b2kkA5j+1dkD4hvUiRqUJYTi7Kt9exaIUEqJ5
xxEXStRgW9mARj1FNnmjDbPAp/zmY22A18kZoL07AffyzevROBgUZBM5360+EVsmrqLQC1dg3BBz
Wo3PM8Gcxsm60h+Fg4LzFET0B/0qiuyyMTTm2HyGYBJH/pbrV9TkWf0w/WTj1mRkxFRVdUi5o2V9
FooNnbr+5cYYke6ytzHKMak2rEp1BC/PG7SaTq679BMdIjXaS3P+ZiORPiPXniyKIewUWmY/tuSM
x4/3wJ7bcGMp5FjXdDCvz148appx9badqP5SfBf4peR2yJyl2Kz38e0AVAPGccBJxEL4tNOb7DLv
PQMmdZWIu+ZeFUr6i2Qyza7h7TMQVNoGI+uszhuL8lnVnyZreCsVX9VRFEcHBShL0hTXy+DTtoCA
Qp/SauglD68k3M0YsQ3HgZjxubsbyx9stLO7tyvt6wOs2QK69TYUUMy7G2rZOyeOx+g9asaEjluY
hS6Bt5pPFhYZXJ/Yt6xbfI77gOJL+xLmwlaT9zz2FYCqG97KEn17AIkDJHy2YH28l1Knhf1CJqaF
JAyF+akS2BeuEXRUjFsw9VQGk1hnY3tb3L53OXJMlQwAeLhBSmRwxOgxzcdg6UNwwgwQYEhKMZxn
anHP0EO5zvO2CvQ0Iy4Sf+hGaX2e/rTyIfoGJHK5huC4P89XyQAb7dqF9eAv1FgDNlVX/HdbdS6v
NrtPK+c11DjVBgCya94Myzz6zKANvxsniNvmhuek1+ywb1b7Hx47BD4qo1tY5UFRbJHqTgK33s69
adlVcXE55p1lEn+BLnjgNppzl/DcxxyDUD2s9u3RItQKt/4dkGMqY2P2CF+m+Juf87TybM02Wy8q
4/LunXwI7jlEDagNjP1mD0c1u8kNJwODtgrrBcOf0mpWHru08c1AbT6yorvJaGpLfSsXq1A1y495
/8hzJRSJjY3xQfrpL04NxHao/7942VCqhkUpalSEC0y/QmzDF7HUPewyzwBz8/PvrSmBi86QqW7V
0ADPlcjo86fUNX50+GkZXOAVJZ1y5quX5vSmLq5HmDfH0uMq4OBzZrARwYqUHYWXUIShNHKedGN6
fnK7czhzbmE30Y7ItDia4vjEKS2KxmmYTdhCQinOEaNkN8BHal99YkzvJTXUHKQ3G1X6/Ql7x+cE
VGCUGgwgM4YtNpCNGaj6f6xtX0XjJkZMav9INW4j6nRm+SHe7V5y77GwOHJ81KOvMAYdD/J7VIve
mcdjb2N0cIEqmFPmNbVi1Dcm40dDpYFASnPhbdfNMU1IdHFZkBajl8dYwg6+WbiA8jR5nVOyFdQX
3y8LMGM+DCgTUqUZWj4jzbDkLPIBfKgGGJ7luUwvXdCrWlT12vFn+yonHQRMA7PR9iPb2e1E8GOr
h60D129/fQAtUdgzqvxz8qdUP8v+ewBNTs5jZElEeEVZ+GlBmVDaP2vkht7ncN49lB306v53qh+N
WRmTL3gFsm1jBqkDociM61FzTLRWkZUSVzc+Hp2cu4HkiT1vIUq9Z6PttxF34HXLnu3v6nu6uSAK
c7it03JjzwDKP37tjCG8jW40Bukw+q7+bCWKTGC/9PKgZQ+z/sjyCZI0jz75hqPdz91YaqHf8hxk
mEXEau3VUSQH0KnbTiFeWUNWcLy3Xcjvg5HXvZmdNz61NtO6FJyJZIJE1pDV7M9qp+hc2dyYNxXo
zo5t9fSjjiFjOYpS8MnYSGzEorD3Mj575jHba1PpCXSAu2T4A5luHXrOhMt3q2pcht25XclNe4Sp
NK141X+/4Irns08dTrhc3035XzsPGFajRTjxPl+rTLV8FoqE2Nn3SHhfeF4uoIo1fy7SmHlHu+8N
C0u6a2nnMciz5pBZwsuaOazgmkSQtHEHxDtFLG3NEi2Qd1oFsspssY1sTdGKKqz7sT7Q6dCidPRT
NcQhBEpb/3hTZpTvtvHPevrTM34j9Uakiddj1GOli8jg/VtbmVjiW1lNcwYRs4pa4I/CCazQo6VH
QHVbokLwotSufaF/iAb77G8IdQ6dR7aucSLOW4CgEu5pVM4doN+RBEAqgwuU8Sy71h2xL8QIil4q
FJQdYxOXYSp65+tqR5qOxKvnpbf1e+ncFAXK4LA2nMz9RRhgPpVvqXG0jGmD/Xzj8rjdWZ+vYVLj
X7+1M4CRnqOLE1abx5CrIT72rSH7nYBr7z4++KMZj7XyP3OqJwl26t2VKW5gdqiANmiTPkdg97Ll
BPBrCXYrnRc2aZ6RpW3QXZdPjGkfAjviHT1P90KAKVpkNGxpm3+eOcZNYFE07vAx3PaGjCIctY/b
ilswTpLHX3XhDOHoWltfM6rUNpORQktaATI4a+G12l0k6AvVxoC1/RWkr7RbUeCpI5NElHKWbZPy
xh/my23e/WyYJdhxbecfbe9JaX2Ue/gJivP2DrjjeoXqBCoO7MWToi39mw2od/yH90XEyYDkzOIa
5feXP41TPC+rNQL21hJSOoesNq/ns4bQbDbnhb/qgUU6ynS8ef/sybjs1qLE+P5IvQZd+26UEgwC
95+du0fd0gCUeW4V0TLBLabWhLIJ2iFlXQeHzvftflMjPH6DPcmaYE+LsNCQ5Tka6WsVjuGUyLkU
oQvKW+jTCBzVmIYAtvoEoK/7wH4CJkAzNaGx8ZqUAtjmtPew+TAGL8VdnZa8z64ejauY70z/Og1x
1HlJo+dkz1vsXKa41IKsNzlvB81mv45zBG6uL1Xi8qjjNT9o/+gBQ4mGyf5LQ3hM+Vh+p5F9HOrN
SsGo00/IoeULHMa7yVpd6lNK9ZmgFWO+XDg5TMNAh3hHKwiSNbluymT10K9pW6t6a1/81zbhsWoI
EoPDttuYXrNPpsY81/MRTyUL3ivTk2bF2UOtUgSIR49p2loKucko1oT2u7J/IYNVJ8fdEG0ugmIM
x8xMtyRbtw6MfcTjHnFEMLNjev9s+BhyabJVcMnuP5JeKj9zjABSF96kHXi33v3dnkX1+EjdJ4Po
gXsdZ5AOUgxppwjmNURI97JTgDkc2i2ZPFv5rqOO+gZpY1eencAl17CJT33Skavk4OmDcGyXHdwy
Z7skRsHmoElM4vzlOu+pm7ggl5aZaERsCOYJHxfzNK/5fG9aSDmvhiosr+NH/yzmJ3WXc3bEWQPX
EoewTacMR8OCD+S+G/p05noAqpGS3eCSzs2GG0KluLILL/zH8JUcrfts4AgAgGA/XsQ9EK9Twl6K
RU0URRGaQqehgR2YhXhp6oR6eEmRiEwe7/UE/95eQcxGDqQqG7GAZTcW2L5bPFig92qWt4RTa13S
so89NPqPO6dCZVFaVWNs6xEJ043iPgKTO63y6lFU88G+trnszNhISL+JA8P9jSPNcwg2uz5KF90I
h1tQJlTPjNs1CEb80+OZH9VJiNX4lxzmXscsUn8XcAEpmvx0DVzh1dRaJ0vyqR+abtwpP/wSQEe1
b9I4lHXhu/mUqJ4TheJTd+hzFCGe8c4RRydSqqM/gVMFKbciWfwQ5l4eY7nSG6m/yN+W847d+XH9
Sclj3nZfu5d6tAexZ5qTxA0KrfLFhgxHuPGEG8IRoiSHvNmhzmhl1r2WkyMyIoodkUWZj2buMyZa
l8JHBvY2uBKbn4qRRcSAS26jhJLNgez/fXwd9LtiyBEkp9lxeojS/9as2pU/pHdffbzK1hIMas7P
XBNP1aJV5aeK6pBpogfTlPPLbeL5CC9t5Bt3ORRw9kY79ldTw8teDbEpQinpEy8NESRtJg7c+eZe
mpq6CXAWR+h5JeVgEWBv46V5C+D4CwyUmOqniIdf2DoFsubkqCtH+JAB1qO4YRms0wDjRj4THUmZ
9AI1Jn1OpONG5TqujOSSVlw0Y6DlNrWoU6YJtlOTPC4GFvxvgl5kRixkPUppIeAxyMZgmCUYtjVm
BX7/O/uUY8qoWuX3kaWmP30wwcRULC9Oidv8duO4rU2lC8S04u8+wr+7FqgpDmrA8AHyB5pZEF6n
Zj4+CZ0zKPF2ebitT5xNFZdmPh+Ol67OSnZfrrEJ//sjNkCh+Zuk74wujxgV+yzuH3/4q4BTE4pn
1zD7TeXUtQN3+0RB+gd3BbgrL5qdiHtr92Dze/0v6Wj3JtRPrhs5UlNuzsf8GH90CTN9yDQ+SqyE
nTorHwb/tPFy98X/Nofa0ZfkY505Jwzp9XGcw+aXsHnoAT5o8AjcsQ2OpEsV2NpEelCznT42kFEd
hK9N0O7ga9RN9HdDWGJ69kwb3q9VC2cLQP9JRWLpMQbun1ZiaUl20Ekge/WuSbYxx2TnciDd1j7C
ZILwdlOfz1P/8WWKVoClj1Zusm5hItmYFo9W+qU9zgrrx7YtGiVPCnof6w7CBozbEMdqSUvgclrA
4O/eTajFRfHNpGVGszND9xn4Kx7EiFFvX+Ht1WBkjFzKjdc0b0M9V2Au7BGjudMpWy9rKbqSaafP
Rj2EKqvahU/kED9cSVKUqJlqZeS4QT3xbLZowjbrNOWLS0MNBUBdXWrlQzwLIPSp1pbNdPfO1Z1/
lJxtFZSj24uIoazB1wZWzz//MikjMkvmBQ9BQ+cR6HTI2DAQN0N12otAr+UUM7bQIGbORDQJgqYs
2p1wC5F5+x+JV/JrHceny1/KmYQJyUJgc4aRU8cu1WTtrakvQ9ZUa34+iFqCnGVkCogL/DfIVs1a
G5g2LMRMG7mWIj7Vegdzlg44mQ8x33M2+sxKGDHZh24YQwXY21KXmey+DdSi/bD6+3Gbj5R1Xekb
Wdb5UDV75nvKfXyTVAbXCZnTOWm2lNw5xYwN1d0pLXdMn9FyHZrWOdX3kf3p/q39gyAo+aat8JvP
T6j5z98S5oYx6Y5TcFh7T63rdNgZBS2kZNQA89LHtc/hgBqFDaIxeXR+xll4jVzlEjywAeIc+hEP
7TeQYqfiErLllFv1cnK0PUJQ2Xxudbx2PNV61KQUzjT9E+F7RGp1jN0Z91CoJa8xs3lE0U4LklsF
Nyzjxj43iGv4nJ7SySVEzX65GYABtyOQaZUydxLuXt9LKypyvn+hvrzmJqeQalECZpYNNXKwEmDd
llmgk/EsPe8YYHLTIa6J7GAxPHdfr9Tq6vJCxLFE0XvwTSU+FGMSLvJ0I06+avgb1bkHWRiu+fzm
r0IfEiGgeZa22Embhq9tIhP8QPK3O5F0EZHuaD61qbZq/jTo/YOPCW2kaWF73YFsYpBOsm74TAh7
unYeXdCfAi/iQjZKdDljFhneCvVLsu7dqZWE1hUoRRtwMPOKjxcdClxYj6/1rCvSRCC+jKDgOJV9
v1NqWBrV91OEx0B42/GeA1uq4UC8mzMOG2bDAQhM7MwA6TQDjn4x4U/N50LQ+zV5vM9Mop0z7C7X
jzk5AAhqeS8ZIDS15D+TGI9gP+MGoYrb5XVuk+pYZQfP4Op8kKBVxpS4GCepfUli2Cbfz1KcEk84
5dd96N+9vUckde0QdKYr9SjwZJXoTnz4HMSGVvkN4/4iL4PtDUeRWKiDO1r3x7SZPbsSmNfPtqet
KXeu171PMT8EX2dj775OjMb3eKo07g3RHnuyljqZo4RW89yfFk2FamVm+pl4XIM+Q/IYHfZBaQFX
IUfRw4dyDOfZO7N5lkzr4LB8n2R5rccTM04Nz/q05PjbHgRMhx7UIAHdGVboVoI1keU92EL7+gnw
42s/yLyvh7vCfmggwwkmwrOF65Xg4Io4w0SsmNoVCATtM4uIoCQciLdY+vjARhL16lF4D/8XnlTl
jWKZRikgAh+gCGq14tVXfMzOlko/P6aQgX+wtypS5J81zPM18ihlZ0kCrxSYjU4i8sLnIQeg93Ld
QTHCM6gswIRg36CwrUNLoNAWOMvr5M4KOdnY+lA+GRcB9/uU5p806b8m5j2bmLdMYO/T9CUoG+Ur
AJVjf67HLFcrnn2/fs1sxaSYKLgXImblRKV/3GEBwebpJOP0SBCJHVAvqu3yxFnlihFVCUTAqznU
PkOjdLJtT8iUt5UssRJrT67EyRZDIVNpahNZkcVN7SJCRaogv8V7ermZoUq2h57h1+XKXnEFbBzI
ENKLzBYjpJHYZPvtGn/9qfpUBQ3PBG94Px/IYl1jjJ4M8T3wKT7GzMdmhfQnGH1qsgnHu41moHgm
nGWVT+sDqbcuOkgg7RSmKEG/SJD73nlPEYor1AMuAPVQ6MJb7L3XFB3NctUmk9XqDimrvDxHZWPe
kszO50GSjZcSd9FsYbNuCMP/oLwZKEa/GX+ycbxIBMZdO+QirJV/sBuDTxAr3mN+5MeYeAMX80jZ
WuT7+ERwENsfjxk+FOaPieIYGQRQEcOaDNHBowpY1Ji98i+x0rNRhpVMsx5pAd5itUyA/0Pr96tW
/1793qcfB7vwqZaoTzMFzxD4aC1fV1z9BhyTONY2tsWqZjJsMAjAsvCexPslRF+E3haubEqQMqAF
FLmS3d+4x/H18ZT3ZuDl0QthueAyln61+cKN0z3IAn7JsQxQ96mvAuULb6Dy64rlcoqfm4DJrfT8
xTEDBTqIMht59dgLKqiHR4Cjp+i1qpieNFVyQfOBTJo91re1TJ6p8jY5gY942zXF5XgVNM0gnvxm
rnOdw34Z0sDrKOm/X93k7L0xcOgE8hE1G52k8SQhwAtI5FmSidWYpQXDIN+KvrCOMGGiXnb0uObf
iLqzlebFQuO2/bo8B9vEnSWMYyRWM8ZManiqyXF+yIdKa0pZZDS7mdI7IR+DS+3jOOCLgMdHa0hO
m+QBb2qLYhClrGVBOoIeFgBwC4E5dYrVvIXJMZSXD73oeWci6G0tZDF5yd7YAGpCvzXZaujgzakt
7RIkfKQ0v1LLxgF/hxSU7Crhk6OF6GwP8VugTaJAqTwXTAMyHTagcf+qTI1obwewDfCkiOZHodUd
htwA2Ot4Lv88WjLsLYJy8+/HOwFNk3W82LmbhpY2pYg0WbNKSlPjGG6O5eXGhVEzG+DWg34KxMOy
8s1l8xIler49/PHIvMvedFCwRowXiDz3suo37v0f+n7Scrba0PhSqS3gvjs8L8vJfEIWX3ABSJaH
SZwAPtV6zHCl/d4eU8O0TnglIgPO5TIjQL9XCagyOa3F9AerktQDYU6SVmjZXy0PPiel5hNpV5q+
zvoCOVEOsMkqXL+M0bXr0FKrWZnzJX4JF9ImAFoHhVFF2IkHkRdE2oLAPTdxxrWl1ad8ivWxQBhP
PVvNliWXQ5asmnbHU6XWiw1tn3SZQ8Bt5vCj85SRiaBRrq4HBiL2sVo8ZnpWKiLmxgi+paPUcKM4
E320MArqU3RQt9VVlpNn2+7zyNSWOSHbYT4/zg4WY0/Oj2bE7dF6Jr7meDT6v7koPZf5oRVidLF/
FqvjvYj8+ZlDzBlpsXD7yhi/Y8NckuLZzE2h+dGs+A1lKzHbcxgE3DS/6AezpoiF1TWL0eQ0nn4w
yzxMTBEwZU8ehwLh8DAZLbYuKxBXhpmiE0fhICpmETUrJt82qdIpy24z4eFLylasnIqVk/r097dz
ztB1cq4nY9bkNlq44HZJTFwHuWFQ1RlU2nF5AZG0gBU5YO5zoUqhqALNo1uCxR7BPg9XVM1k1w4Y
G2qiq36n9RCfBTsn+pbwHYfCynyfrwa4fRLlsipDhD7/S+300zZDDtDif8Qb/iIszbjK7Ca3RLeZ
9alrDavNbhNPwdROmhzgCvVmNcnLDfwU1t/btREJJcotQJglMielpqVRpN8QSF1CbX5LESPbteDd
TtnPIYNAcbFP+CL+84yqKlmC/mWy2JyXarzz7RmBHYPcfgp9pZyoZIJsV88i2Bu3QmwIHrj4GEMO
IklJSk3oT6eNPHex2nKmc3wf4gYf0s6c9hRL7Hb2tKao5rU5IR1xW3+JU9zxdfP9SkASBEnQpijV
Bu+eIN5REVe2kIAsxeYWFXVrcL/M9Vj2iXFQEIVGIyNP/+dEeBO1ART4waudUHAzxlKC11vMF9WH
VXaARNotI/zc+4NFRAXyHvSmW3k9ScWDaUi3Gt9r1ccAEtBg3VjMiPiaEssBJRCmctGXSLTccshP
mda0kJCLLqbhIbwMWzyfy4F61TGVfYj0QaA7cmAzUkEkf5bXYrld+lVLWRzjDo7bpaZgCeJoRm/w
XZP1LkmH+T5fcAuj9LCbC2E4QT9OUsK9TwNnffm90mixkiPURrxQ9FyuXy7x78orRs4D1qgTWqpr
le7NFiCpJXGd/XTgAyI7HFrdrYfTVxFDupr00ZVo3iwUnCTudlKsvp9jqKz43VJf/boh3oycfjpq
y6zvc0BlvcfbW6encPElrd0M9+fP20oF/3xC5G0WcuwFRA/0mzLeFbtdisr8pjuaDhyUU0lCDMsS
I5s1XykTgaQYIgNzHq0xjsVs72JxxZboTwmK2vzPe1YbFXPOoMqfUWUc41NfI46gnl3jATldxUSd
hfqqTwQl/0moHrYtpUnF4SDE3f1ZTQtYz5H7WGxLaruV+OYoLoHD0Y/TwrZEvCmlTrRn/YPjb2W/
ry6j8waAc4ycVhF4oG1DVuH41aYls+9P8Mwq9CIidniAjeg/aQH2au5eJ44MbbJC2bnXxvYAU6rT
nj/VkBH1JpFhETXLw5eixNDkiGjeBiUSgYD8m9w2Ao/8afglI/T8stSm9p9lxF8m26Md4kOfJXCb
XhiOlYnR9npsa2IGJrg7t3TPGgxKD5B4CBW0/fjXCqdZBmV+H3nloIxIfxCL8va1Phdc9ECEQqNF
HDfgp/goj6YzduS8C7qQJtFdeZ/LFo8SRV962WATovBg+CV9Zkoc7tS5NsCCuRgNnruMPccOVK/h
9x/gzyyr2cyIS+CkHBgTf5irMK9LpwHinmiDcnK2WTgjoTkvgzyA5SM+KqGjGRGmJlzQu+tRsjAR
gcW4eREMfvViKSx5xup+MfLKZ61U4WbBP3pD9uVzsrIU3iShb93ENYADF5i54DrY2/zA8EpqaxBV
MhKOjrcuXhmOvg9tt5AWUuwoiLqpBVEFi+6S8GFZZjKcYjj7BIOxv7GrTtTFamrnEF8V3IminJ/D
/aveRFAlsw+kkj6zz9Xfeyu0nN8QLPgHbH2AWPsYgEtqMoZMf/0qFd8xfFH67z9q7eQYq7xQRVZN
UUzfMPRTc3CdTTu6iY+FcjNuBOccr8R/6J0gqxXTiLAl1DV4iENo2JL5jl0aaMlHojBEXp2m4thH
vtPrpIK/NnRuUsYclznOmvRzsqrrqlCmUM2ql80NAp5lqh59FQCVLjheatt0kEMxJkmtqjDQA8L3
fyCkg+jV3snG6sFv0+3/Say1p4Rl3kasCEULDMNtGRo9fiqv7ewlwDkHJa1gbOAKigQRGQJToUZx
0ii4LP6WAXY4tyIEEH81nHqrpe5tg8y7erUIKcOIQeAPwlY1J1euSJNOe8y/2/Pnq+uB9TOmEoL5
2xGVbceJl6orMapper2o3S3JAPNODxMmI7VxcClZFGCQudzYr7bA+xh8XXtRnhml7RmvS1uSZQ+S
rCrzd0rMNr89BYIcVuoIZTg3lWxAvkzHu/a9wqepPc8stZxCwc7u1a/LzUT5ffBrQPCYxE8pJ+L+
cmTKRaDY7OpBFdBZaRdE3dnCvPa+6EwnAX1m55OqTHeJl0QYOazwu8tRgVliC9tTJUit+Zw5gb8I
A631awyLNoZul+bDW6x1a+CousSMN7A3UBVlP7EvCn2u4PjxH0WM/NafeKH/llZB8Rz8IeSsfAtK
Mk3jswS6f6yDdJAm09tEiVA06BUal6uCoXOHUeji9wfeh5ktq9ekmfmkO5dfKj/rerJGnkteyeaA
88m0L/+JkUiLQlh3DjGRa980uXALUAP4qOn5TjDM/6CxRXUYzGyjBvgiel1gDWuILsCH4oSmYX+6
/C9V1/0bXkrsJD7cNVkl6ZOsxmYrZRXzB8e5M00FjiHkPN27T7uEDXYXIlCPlJsIw36ERZbenHOw
AxO3xqdIQJgzeB187Qijohl9gkVgxRL17Z4c8TmalAGU8LOGv00JviNcAmJv32Y2WKUUAnNmrHDs
B3yBrXUbcEHDskEAw7mkjjnVyc5InLZ2Z6x6LF9kRRmNUNpRYTKpuNDo2aigEHCooDEzdAam1rGn
wL9hGcrIfjBmZVENkPpmizlCKvQ9NM1jjZ7SH2k0vmCSEDRe3VXScoK9UhDNbpEjypzT7NoHLpdw
mag1SHQo9+JeGVYkpI6KsOOAC65xZd3deuQIOMMo0oiyct+ylWGvRi5yiOHy+FkGOo1ZaItygPqy
yf3NzV9iStLvILJB5ahuUBgyY94uuzrPx2SLXeOkG2QbFqIyJu53fUdN6D/VA/ebPlDOL0snRmGB
beqxolysJZDsS3DDwp9pmjoQXyYCosV0JmTq5RT4SAd/L4ZdNl28IKUB/5gpgA7vabeCQxU1WqP1
73gerQEaihptohcqeMlpraVp6rZQq0a5jhvBzoa6PvoZ8vokRVubb1TX4iXHWXHRaUJTVaDrvCbp
gBOIJZHyBls0QFKabLp66Cpsy4BkzlcrV2E3GOug5Ug6QvyD5OKv5AaIDNupK9BJWyVqe6ToXhY0
D4fKRWo9cEZdjYqDwuLqxzxos0h0kA/0FsTO64oBk0LqxdMkLOU9KSzfTGc5cNaUhhIqV9bvsHWW
huQaQoAEJuCVwdHULZgJrz2vCPWt1zDEjUKF/rDsyuJiyBoAXwbwoDTOaWrL/t/qtGBluuOMJ26M
9JLavf8nttwVTOsaTKlik8iZ2hUEgP1PDVmOOaZvlTcFwzNN7xF/L3/ArnzJKrHoLYZ8b3vCRIr3
ktWxAwqCivb5Wjhp+qRfmUDkVAMtvZfB/mkl7/BP0wAX7Chz8u6WYxH1R1BnyAk+KlNDCPGefOuc
NcF4ayO1gDfwSHyl7DFk6Hj65l/u+tk/jrbynC6MzT41RDvnZssaZNuN2zlnF745p2bRGPklGPXf
ADrfR+sfrPpdSPELuAdqHUJESpU07SUU6VGKMSG+hIR/a1fPVTSaMw1UqvCB9h+HEPq5gDpHCCIq
mxWkJX1bcgiNJqNbWRUQ8DjuNpmB7DFpvtep7Vkyrf3hIhzeeX7B8R7WyNHS8TGpnvmLMJwMbGE1
QUpDKoFvKcn17+/6u2CubaPCU8oW3P2pfU5+BTURJxGW9IWDtlvGx4hzrb7XpUvWJb4xBS/stelS
aLZ7vij3LA5uAR+WBFxaATjhRD/N/+t0DYqmhZf5W19Aq0RsgnmwmWkYTxmjv3SFfIJuWZa17svi
XsvN4nWjZvHTvvgl9PjJJC1KTuK/8NqH1dW7UPGkZYpRhWtA2vu7oNa4jbH1tPp1ut7PwepvVpzN
JXt08OuE8dpLjIbjLUM9g13MGoivRbxxRDGSlAYnfIMV5VfHa1a8H72pYQIlgLFiYcv0NqH5J4Zq
jQce88cFMVAXPxmCAXbBxqxOek8JfjzAUmaLgByLH4lfsNlKYviZ5oh9UmlnZtwfHt6oOrIbk9uF
K9Dui2Y+kWFpdHc3QfxGJwWRN8NNY+5an1pEpaWIB+7E7izsmw28VScigkyUZsbPqOGTZPwG4mS8
g+BO4nN8kx92UCA+/0vlIRguVQImTf4G8omBroT+1qZaqx+Knd4FAlJaMoBsudRD6Y2OwlgTdgnl
wEa7kfQFMcCGF8g4Fh/5V8cRumGoH4OJflz1l5fmAwtCEbUuHwA4qBuFtdmg8bCiv6hbN3YB6h+X
NpC1BLqQ9RQJQ0TBLlwACU9YRY/XfzfxzzFxzYIlpeyFCLIiKahOnoOA4LkaGjSeXZzs3MVHI2OW
6OguX+pWBjsqW1vQE50leL9NrYuGCfwkPeLrl7cXLvYBbXb9+dP8tv1d1mXtEhie4l6IIWlZigyi
fhZ/Z3lB7Dj1vYud1GUA9rUhGqBoFSLXHsfUpSrqAZryxjlJdUH/jD65ZF/o9Ni9sZnpnv7Iz62e
t4aYL40KiVJYXVTLA/FRVAzFUcT42nu+c3ZROzmeWfEFVMQFoLEvlJ1PjP+qniKuGOxEsk2OAJfL
JsTtj7EQ03GNzlLXJaGAzyqlaiNVwasOtyFjb/ejMkALBeY3VuMIGEMxgeZt9Rx38UwXGVWwMfNB
3wpgDa87vAEdsH0F9z/IXfTlvcIwKvLT88CqoXElw56S1MbhjoGDHELXIwbAoPJC6/W3OpDntv7W
f7SJVUsyZyYRgMeXedCN+DxIM633DerEfWB6NLmYrmLT5kr8WsYa67LBy3ZCVl1JDIUSLE3bgFHh
gWUFf3AQnTjpYM/DfVSnVgrqGQeMLWvUsU0Tg5yLjOCGbWwMG4/jTGbXQsMkA6Z2MKqNJcLIlpTt
0LPRcjlCQPgDpt1TPU8v+k5Jh08ZMuwyyTZ6CLOMzYamdpozdS3GahvgeLmUZgOiMnM8TD190iJu
BQrDBMoOhDah8moMSFtJC4qak9MfXNjqUftcsgI4b9cwFEyaaOWGYe9TFI/OHe5Itbcs3EHGjMES
LM3BrbF2cKMmnhFsTB/zm9HkRB+NbbXNtP3R6tfdn5Z3dX7fKfloLdaYTiKmC1pOIeEqSyf2IMkB
7P+rIjXfVFqA+YiKPrXio/ddLq7hy0gQUzox8tdX1GFEsU6Zwm62ixk/bdjcNsU9vfFfx7Fj7uUW
pl/mhLl/2KGJOwo/NfsrwGQuxYwWwhVxnkGr+tJoAUsaDZ/wZVvWD3E3Tz9DxaISman4cLzMcy3u
jZT9DO3XFrL3HIG18oDxxqBi4Gu0ePPzgqH+qQvBiFjQq5D0vJN9D6g2iwzP+p49ks5MoJ75vxjI
MBZeV2YEQn3uO/arkxaz2ifivBc5r5H0zth+ip+1zBAj+T+sDSbACukoQ7FIdSz7etDTkvS0Z7JF
h/MYBW/BjvBX74b9Yz6XNvkCdu33LrVXJCWoGVRVESYc/bsm7T/WG1g0XDoilGvCSeX+B3fbiV1i
3y3005BAkBK9QHcrc+HTct5U2+MzuzVWXdmYjvafEYRpLsit4dr+YLdfvO5TkX9prZz6X7gHidd+
2v2QHyP9OBfSN6EyA7AQ6FGWV1FLbX+jQgWlTgh/Ruj+ti9ESffda5yBu6a23WBLPELu61SwEb6a
DrVfxV+GIeMdne9iOtJlax7vkS4FFXi5HWWxmKCofrWj3gc7+5HIrWSYHTx67k3qVdBMrMwgYChb
TzgIP7C4O8Ifm1JXay6ocYQP1OVPd1xv6dTNUfBexkyhI9J8F4BkSKuZ4cLHvkRyjyRplx7FL0JV
KBvAZpNMxKUgxT7nRVfiRfLimjm484zonwjsPbQFoOdFps7aQIA76NVpcaI0pYT2AxQ6n/VD9e32
VR/XmAKk5vs80DvwfAnPd/PsKlObHzKGi7Oacwyv3D0Y/6sEuI6t3l36+8X9Avibxt30yAD5dlXP
o7r1hEpqtd597XhOyNhpBKhxV8SzhxxMIl24AKGJCxN0ff6KHszkQ92Jg+PVtp7eFsV0IvflAE6A
UgrAdYvhRDnZJPPdDDdU+HJ8sAcig0iE8n55wRGGMD0KWSdLduj479HBS9IgrzZsVR1BTWUnnG6I
HCXVT4D3+PjYUpQ/KnEQ/VRgSGtEt9Uwh/fGKO/n9maekS/vH3dNWYSxYUV9YOdFGO+MjeWu49AZ
qylZxgxdVfljQ67o9MDPShGdOX201J1wHtgAlJ82obwI/EzpSNwbFekbX2ziFHFREgxaVL177F/a
VYUd2sDznRbLI5U5yGxj4NcpcK1vJTBP0XfM05q5qlObHRzR4B9ocM96l78YVbG9oEO56QIOfac9
Svl0SS3Hmq9YCdAVPxJuvrSQiD+dkYLbsdcrfaXTDdEpi9s3rDOkhUZazPm+tf7teG4snpSE4WLE
dlumWIYbHBi9paZtFTFPh+iaxks/NuWPiVTgVdpdADsW0sIWmnS4IoIBNNOCqE1sO0pPsXvY0BeS
wEccU9Wt5JjRCXXaRXcOF0YsJl/yM2W/dQoxSLptMPTbAGexCise6rfH1rZAM0n2UmaH6/kzs/IZ
qcO749TYs4UaFJ5sfO1ZTZ1K4//uB+Ow1yc668g0zyZ+mhQDckf2r95u6s4uBrq0R/pz5PRyPGNE
t7I2ipXz1i1eApcruMo9/jKC/bUBwqMfw+q41He44CzhWT55kE5TgAMDaTJZbA8+vJQhuni/VeNg
HLaBnbTDYxhM0AdMmEPOHFPMk/bUnQ5r3u3ej7Cp+zfGqJJ27jQE0j/qvM6QyU79ET2bIIxYdOIO
iKtIr5BBgOb2cW0yoaE+rX3a7XcdReZsEROMeQTgZW5h917G1eB4xiLmI1buGAra9CjK0a1zNSDN
EiW9y4w2QuwmRQRFEKQuFsI0vw7Q9a2h1nTKD7BjeV5hcLoHmVsX4hp+BTjrtzsvJ0AQ1OR6xf+I
eE6CC5/UQSMOnBHpeAeZBDqzAj/3ZdM2wYyayqQ12GbogFBWEyMis7oyC7zq+OvRfNsogQKXKpCm
BriQDMnYDUeMyTQwL7K0kWKLbY4D4fEts1azcZvo2K19fZDJcj5vdSyGgUt0PI9N8dMZxi6IHi7K
dsXKIrlYO87zhB29mTyVO+El24LoMBj86q1NKHCT53ebukOV0KdFBiB+9M3Gh6zmDwZe+A6Usbrv
UFajhUUEKCQ+jQowudYaHzC6HFxYZ8rvprMFUOv8nER621O6OXt2LZTjORA//OEeycdhsGBC8six
uj3zzWKsD9KLld3Ghk/KlbwG+XD0da94SKrhxcdVM69HgoGMXhlhV+ojcZ3vKLfxtSpW0fYerKGL
ePgym3JeCmhbAzXAP0UlnCm1C5EnvI05z6JJd0EAy6RBw5Qj1uL6ew3IFm/c3ncCT4ZEyZHtgdnG
FI3kHDyb3g7PEclF4BoyqfWwURJMaW5H5mdV3iSzSKxbnaoXyOWXJyeE66Dklcbw+oTMxqdZ4fJ8
02zbXTVssAiAUK3EUhYVCoMZ5DSHNnJdsOtoN0TeLTRMfsoSO2vDgXFrWT37zLFFyU7LQrrUJFpE
Dig9o0CkT5HX1pMXUandmOIEqdofPA0xWhe0AQhce5gTtCwhuBRPZbGV+WT6hQFcL8Ng8sT8xVjR
NGp39TlzuG8jOD56cu4jvAPe29YyY4HSJrwE2sD17cKI9VOgBbOKdrMv4rtJ2y0zGzZ4D72L4kfb
ZkBsjYF2XrpVWgUM72J2dVMVgW7l3onqORHzK7qjd/lrkTg2uaPXf+SrHnFNmvtGCcfvsxFT+Dwe
WFbTduZj3n+pQTWQ3GMyLqvczJoq3iZJWbXNNgZMclNz7J53rygUHlsINsqgcEzkEValWJzRI27M
t/jM9LJruKgFzUGxQBwXf1rh4oXp37x5ecKUgZaI3RL2wqbd/pWTQb8YK+SyxHXa7okcUv1bACTW
VQh5YTSF/kRyatfRiyLnOFLPDiDylD33rDn3sHWi5HfeavOjYnJ5iEa7GOSAbu5vqFOB9mfddINe
Befx153McJMHZLH6wAmI3+bBW11OzfQEQvnNjoh50FDn1fAspqFVyi13UQqb3t9W5MfoWcjMYN4G
UmFfAiZ8qOpbj3MBOT0WNntU3xhA8qsgvdqzyUm9lQ3hrUDsfG8Q/qc8Q091kco1ksnemPDId/Sv
YdQCTzd/uttBu1/m/WwgfqP1XEAqP3bPQMIEeZwl+FTPym4HfCOUiNtQiOsE1W+Fiy7AeA2V4iva
BrPUZXVIJMYrL49uhUbZ23iYRFaK6OZH4CXAN+BLYLZKv8KbdWy0orJLI5WWMbyguodiy5AmLdJz
/pKnwoX+MjAL8mPNeA2WbCqdOfp6T+lgORC7+w+Zv8GKOpq3R5L+NRySz4ExeGTOspQ0YiqPy+0k
IK+V6qVWFcveIgDFMUnr2e25IzXxctqS+V3vuhcCGrakTU/UjmhnLfwsgdFJhDVkIBp1vuHgKJ81
gApFy/lDKZoDxsV89IchGW2tg9Qbqrb2yQ1R38bu6Lk/XVVOO6jmayAxbQCxa1hYOdOYO4XspEoD
Hkx5p6yuL4EWt27DXl56Ea+RdpT2gtqejGa/DdFNYOBtC14/wgynf6S5ZvZKBPys0OBlkqsz19rv
K04Xybispo8V6Gi8HTxA1GxIz2mVgH/torT3Xu9GrUY28HKSlmt39kkDDG3FJzQ/rlupWg/eTEan
k2Yf173sWCE6Gi4/uK3qEMxJYf/W7v9vwjszIAJI+bJwyljUf5J6alxHwsn+r6aZJ7Gi5OJZpALv
XOVO7u96QLFDQWV3TxGE15tIH526e+cmawtzugbOpssnF5dtTdRx2M0ECkpPYhDKbgD/3s9ipmbn
D7zWs6bf2nmKTqjD2A7odm4Lbjc3j8i935rJB8pv19SqSteprgAOpWoyhMNqQHTIwKhojuOm2Zxw
DFsIg1FiSJT61D7rBRS/fxxsHk/sJfew1+3DTq8AyRGbEUsqJL8BJjPXJGRIxZ/QjhfCDARJrVde
lONHVC9SXcE+Ng0iKNhHb8xGfQRFN2vLieg9fKzoMT2S4mTgK3SIdP05ssYF4RvmI0sr6OAQTs9t
vWhmn5LaGmuEPTHjvbAOjYWe4DzJaA/TfpQ5g8wkm3lP5kebr9WqMs3IUmcXbv6DpTbYwpS3+P+B
j45I3buTiLUsbomkRIDPBcr0uJv8WB4qhLpGrjAFftvdsrbdCXaRyrpr2aEtiGGXIOLPbZ6I53H/
4NYM+cvVNuWz5aM/1feVjN1WkUeeajcDLFNcFY+PDe22mMmSN846xWJrziCo/7HyM96LJaCOq5rE
u4nBP+O83TRNCRgELw+UwDF7X/rEYYpR9mi00392OZieianNerPLdKN4if4vpkghm0DeZpR2k6kG
FdOi1KAcaasUQkXdQiu9K4wSFbGX7u/W5ch513s2EpR20Q+GoiLdE8XJFfv/R6jKAOHMe0IE3cVI
z7e/A0XQ0rtZmC296/CQ0vrXr5+DSpkK8n+eK9a97KjztGzaojAlls+/7qln/7GCAZH+Rb2MrgUa
ptoL19DrPBQWo+o4mEULlZRDqFI841n/tq0dryte1YgtwJUkdIrTN68qOFwOU/ODI5asE5BjMVoB
e4Ej7HJXmPynp9eucn0CpmU4AvTiHDPxS4kxSd9uuIRT3W6B+zl1HpWdji5Aqsniad7C42dDo521
NEPOKE1plTjWb+fr2d/87WtW+gCzw1gE9ffknI5dz4H6ZrlYPajCgSTpUE2FT2GGXxaVV85Ffqz+
6+Wc5kzp/9lKNHwK1Roxkabu4AQxzRCJA9I49PAwtnuChDMFaySWsCOx5tTC0drreJPjhoq3LP8e
ezU3Ki6m0ZUM2FtpxfwQdMOzcvK9GsQTbdztqx0mX3dO8jVJMldshN+eYrUeizy2XjjK4fQNWtls
5ifuCslGReaHMuxBk1Bw2DtYlOulX/3qWsAMs/BtHsy5XYZVHG+J8GOq/mHP0Uk0i635OKhlN1Ol
iU5a8OWbuCT7fuLsifose0XShbIOwRq+YYbwUL4V2a3rLK6BiTeWt5BuSzkW9N//bMfb7Z8TvZt1
Gv2hb0Zqj0tdzHl6ux1cJztti8pPiu7uPG5is3AgJO1xrDqEpd5FAQE8J2wtlTKgy5pCBmtmTZCp
Xa98r5rnzc3m8VYlk78iLYXSpQfVJ6eY6bOpEvdrZ3qEjbkwb8/CJJ5YaeBMA/cmtVjupQnLuSsD
EYWxBPIG63AMC/CWrPIjUS9R6VAo8JTzJ6j+DFr7QHECAbcafsf74KFJrGqUJM2ofx5o/8trgSA5
tjG7quDcPVeBspHm7Hnl9iuf8jiJMtKRYft4Y+pvhJNiZAJen2VUQHi8Jw8fD7hvpZaZ73X55tsi
aw0aVP48uX7i1kJdatBY2h33o3XxWaVjiZRyMocXjlvVXUkrm2y9V6qW0uYJnAVCCJYqtl9BfXIo
9IXStR+Cza7m2mXfFXNLUVAzEHeb8DjkfE6fn2ySBDpuzfIdcdrL27KpxS19AydCAVQuqSPCTSAc
s1h9vnVaGQjGp4BQPKJ+Xgb2eyYug7/jJ2RF24Ykp6vAhkyUb/i06SpA378JB2ob7zcsUfUZDjk1
PWQKi0A/0xIYw9LfRX6iXEP653XPU3PGXWLc28dNUF2sTDnOx948L89afm7qLG8Wd9tXgNxdMfPO
dCCL5R5C8Y+eUfy737cCQ3GiXIVoxzMfvAfDQ4YRJJvt4SnDQqsDyAhEkVzzgkSkRMcLnXGNk1Nh
rH/v5GLCKmizQiPCD22JxizCR6MgWqKaX2CVDTENqz16RJhlaXIcbyBnkT703oWr8JC01QHQdsq0
LuTucnDVerOScn4mqvk+zkBtgW5tfj/bKg9HkR71GLxpiXlQ4eWLLEAglAraTJZyyyo4fD4bC6oX
SFWoHlEyudTJuoRt9SZFuKlY288zpEXySB/Y9t+cpumR+C+u0L+6Bz6BnBtLRQuolryekBxvHOlf
AUzpTlhoULEQG+nik8J2pNTdkB5m0omciOeT5PJpi/X+iyh0iS9nRxi1imsQjGrFSASs1D0DChOn
RGxQJC4zqG93HHxnoJ7KgvZMsPy9gxRXuPu+i7gHgaVZW/hXL4Jw0Y0R9dsRttvRFgyT4OzjPW9V
r4E01KdEDRlno34tSzKyrJrSqHTHKRSv7jnqs+A/5JJjCptCOkbwSMQKOwrveX7+puiJgbVXtj3f
oiOb1SZo1i3G+vfqqII9nI1rFe2ozK6gztK81BMvcFmzC6Q4FjxRYZbJMutHjQj7WV2OyC39FRyf
Opz/E83a0yLEz77eH/RlZUcQ6hoclyTauHvDt8IdXbr5ElGLP76UJr9H8HFq2gOUvHWsJbxhlBPx
Zhg2j2uGDf3oF2IXexvOGAhcCUfPVA9CPt2dICUggDqx4R8tqN9gOF/jyTeH3OamPxhz5CVCm9c/
QBHaKDCCwFE2goYkzkMCdWpGRCkmyH3lxmzV0rYM3YK2cs8g5visW6zdbG8mgjcrhdvZdXR9FrYs
GCyBWpwruxY710+Egy3FoL9RnCfF8IfvBG1zPyjkE9rppZfyjwdwWb2Y5wl6ZvwqmtlPx+2Gn9ub
N3ay4nZWn+w91LgH9MMpARMX3EFzp3KG3389wJX0xYgAHRp68okY1nxLPkFTzSHJQTmxp9DW1Alj
dv8n66zFRiQGGUZUVHRPBoccvvslvxR5MmkM//LemEn4uSYBnsQD0AdjnEAPVIX6irnk8g+P0pzi
aFcHGxDb4TnWvbHZFmxAK0R+8V5TZBmEUopfhv3pG2J+c1Ox9vIlEpipN74mCYhmbfwAuvPRSbky
dao1KN7nqjAKPdiqndqxE+Rkxr1WD5ELC/H5w5Jvb7xhOe4ZDgh3CVsIa0i4gfYv+fqMyk0OWBmb
Dovpnp3U2BcuLgyk1e4IedaCRgTMofqnYn8ZIk3cmKN9tuM5GXQDDTaiGw4rHUPrFNsFptm+Kwlf
tyLTHpgtMyhsq61KSvVKvTn5xVRX/TwNdsvUfAjECelsIMO0Fn6q80GWuQQ03b9/Y0NbUOd/I7ky
9+f5JUoUzDIdQzGWQvJH+Np75VL8rR5o23E4aCP16BTx99z/LeVFd48rtzbxWIyz/6LznHO3l5SF
9buzpC2vJwB/1oUWgw0+/VjQIqfTHrO5gw58xQt4H8vbqdSgCwMa7rk5W1lAsqxMVXnoIMVD6nQm
ZPlbswJgPjiJv2my4Ta6+i4Fu6Mj1Jr8TEkWtl2MOQ5WoC4+a+mVwAxqO+e2AD24YklhUbnLy/Iy
kyrf9XacqZRJ2hXpKYwtJZ7kPkN/SQAiVEhm7c6ytJd3wdvkR2Xctt5DdXPnEDeITQgekaW0njzm
TiJvSXFVNJYhWpphBf0xAErjKgKaHbxVtNH8gLsuv9MpxrbAzdJNWO/Mk1NgSfcQgD5wymYi0n9Q
d09sx9LhM7rjDnDRnBxYvmuIn6CefCCu5o+Eis63mtApanI80aImj7bwxA0i9Zer1dF3c0gN4xdF
v48l1o40BLyP3sVzSaM9QDOi3fL9w4UqPHlIu5myYP9v1L6ov/UF5ecunbf57SfxYBgUFWA6n9wR
tp0A55+KftGZTOXcv2s7yT6OpLKtoU0zRt2pFFb+mnHUDdzn1DlHoA7s+OePKKHkdvs9ZpelMvfi
sjzZkXUkC6/MgeKibmlSK2cHdh2GVPa7sowCq6X5T+VVm9oofU8ylH5stcIpY7yU6CtG1loxljSB
WAFBtgqQTlvFK37xvJiFZWKTiE3NCUVVyLTf1Syh3DpCdWZndTyVvCADXui/85uOX68a1BB+N7V+
gNIBeIH/W0CP9f4RimLdERRO4udXb+Mtqib6QkjGOEz1QOxRmpek1wdZsk1FgOIRAThGDtq5iCo0
hlit/zq3zRmTTvER+9HTFMl8pZJU4PWb5G5QW67UtKgmQ0bF7HnyYj1mwFHuIkiLsgQi1PqMEIg5
M+e039ANGfODVOX02DqWWCcNG750DT9tMv71KHA2PpvsVmayzKSjRi7J7iJhkYiG3NtATMgPCMEy
AAvmdYa60ahKSzR4GmnB7M/Ri4Coyrcgk++QKMIcKazmJsxuO6uie4nBF8QUOxLZ5PH72AwOqPag
45mIkxYyPzBxNfYr0LiEjJPJHxdKDZPmloMdgwRseCb5NYbfobj0Q5Fsr8j3sgFFMsnI3zHPkAUB
1BimZVjlMw1Kjo5d7TLEPTYioVQP5WBhZxJWnYOAgCVCGayjkDQf2N5bmRszZWPak3VDJoYFJaPC
pJNX7IJd/fM/GqkDNR24jci+ESIKflFZ5Q0URWI6ABqZssJSKpsfzcNLFdLRTxPv1G6v+ZzF2B7p
qtWujI9nBC0CGgQyH0xmwZJsTh0ljteS1i6v/mB+ujz/IJmpOOoH1qfChQ1wl84MiGN8y5XX/h/q
gYMKuUORDc7QgyAZL48huAeGaoaxwwLvayfWQ9Ca1QJO4eDtw6VLRLmwdWvg7DnULP0osvHWWHvR
2W714DAK2JY5QnokSmfP51ElgM4uhdgwJlcd/AuZq9KxJtLCm7ZK3clYCfiQAe2c1LPgCuLKhavl
x48wH7sVrsZYhQVQ525wiRxZ6BDLwtPqafdoPi3wcI47iUjCG6YXbkzQzUMAG5yMlyuHk6tMwVuf
DVUPZbpszYj18Uhm6/nXCz2iNobgQ1rZ5lnanWfTCG4c4hGEaIg/jlr4tmjGOyYCQQBuR0ua46ND
mqfmkRF69ynbIM2NR9OtEXdFsJrAc3+EksobH8ESIH+i0MzbRKcUV1n7roryW4N5Nwyxl1ED70+M
b0YYXTPGbDX1tG2fC0nyiTMeyHiMdW3zbKPSA4NPGfDlSzOlz5/NVLTS3KaoB+T+vdSlfNtSlYco
S76UmImHNB5tzW9vIhESCJ/XTdy6RWC74uCcJhlqsWTGTOZwCB5IpiMrqfksKrf8J21Kx7QOPRa0
OkdrI50b31z7AcaHFTWiciBKMPm6t2DeudghfgdfJmzuG/u0skBB6rwW0Ucme6Vgb+iPTgKRXKKL
+CtCafIXyBTnlJOKD/w9PVFbmKfpZ7AfVmqXxlOm6GiH/nfGXYn1GnOllDGaq5nmwZ13qxJuckOf
pE6fj35Hr0PoVZPldpFDmoDrRjyNY3VAPEtDW60q0SYIpzCn3R1UIg/+Wg8sHMuMWBfIZWtXfQ5z
9Oznj2HQcB0uy6rA4XnacMSyAR+E9Jh7660ez3+wx9/+fo1kHiTil23ow9J4qFgWm6+6A9tpwMrS
6JziKDVoN7pKemVs/R8rE5SMcgJCfOj/CPsOyu1yE2b79alxIpjN6ceft4kFLlWJvG8pM/h0fR5S
7wnqe/YrHB/AYA1dZLIW7dcuvnGmyaU+3ITqE828hbICD+bc8yy5mkgHn9i7hlmhW8xJE3Acrlel
9E5BaXKxMjCPvvVp4NtTYxh+aQV8wplVlRSv7G+YTDKegjI7nBUJp68a994TR8f4qnIInAVNpMWf
vyK8+6u/YLK9Sjcv6zqFjK49rceN7zlb3EzWZ2tR4GFDjCGxSLqNkib9FwBeAB6BwdF2DCcUJOoa
SxFRv0rMLqD+S66JN6PDbi82eP2Ftd6b3D4I4hZvP+JrcMDCzAKqegbfcbKdK5Fs4bpbpkXGtGZQ
Ln/Kj7FvIlwymTgVNJ0CHmkQhCUnA1H6cGJp9NfO/v4OkmTTxiXlTvQJpfWTs6jduUGxov9uPdMZ
eFAnTmjvmaZf8n748VitOJNrzu41xblsWV/H2QyjSlSS76DSb/PbFpY4IDtOqi0RBKLo+K9winBO
Sekneo+7b2UEu1BNE63hmOZtnvj6duhvnuiZZU728kavUF5Xm9w4cT5qSbAyWWSo/fyFWLIH9lGQ
nXCT5eR5FpXPbgPU3dFQjMFZpKf8/PSwh8uneI/gToEZxpZ4JQAFyDCS4/sDW83VbfxxCgM3ock8
JcqZeDgKcWp9/lCo8mnXuYyTQqnaT4jFmwaDkPIQWP9ISSHgW2yQi5mCPJvai4RJeUHxgUcs7dvW
43hxN1frbcWz5MlhJQGEoIgqidh33yX1gZf0g5Uiw/2TspZE9QRiecUgQu4cHdANDR5Ybbl1Uqal
gg4tGyXJyr5fxmkBUf30hXM6i8DFIQIaL2lVEk1zERlGFl2RKsHxZtAnnjaD5IQiDI3VuyTDzT/9
tOjhOItTfBkhdkZSdHySHjyJB1LCnEGFYSW/bu7UgIhV4LGikcFeBqC1zW8HL4RIzddRNa6fjgJZ
t4jp0kQo00jEcVZkuugeXKyqnOppOlmrm6GDpsUc0d8jMN1WFy6aSTWfAzBUamSXeeMvm3Aas1kZ
x5MPBPvGEfvaXVO6ACXQlUXMX2PVhs/GOTOWaFKHWxc8VCSzYHb6FEi8wwWwB14kfak/4hmDq3UL
8OrKPs6Qj416VLIJWFq0qRo2I9UKEzPufnMrJOhEAv9D3mNPGzH5huiiKQ41X6UMVO8xgJjwV9Wr
GV7IexcFLz/meHd0mQJQUYDViJGU1nM44D+IwXBW2yQ3+Y7h3bLcgLuKEve4uj0QJnXJPMHftoyw
sbmKW4wes8ovfHryqzZh66Jto5uGLDG2wNmu68Ql0/ESafka8553vPJEcBEL+GCFl4Im2nu7RAvG
9KmAzwmE9FrQ/6ZkwRaBgjSB9v6O7+XFKkVq1tsGOWaV+DRyyfZX8KrhRcWxMzkNIyEtdaS0DL0L
LzM2EJ/QXuwZqso5WkOmdWjxsEqrKtiAWOlNv5n8Yvee1gs9hr9V9/hb3A98fmSB9UKxwVF7gTG7
YQDscv8sepi8Zo3QAZG0MtxzknhaFF9vuFhqUwphDtYJ/doKKo2aBI66MYXmGa4Fib2VGFZ/YfOl
HuSvEg7L/0nTKlbxHYDl6Y5PVnL67eqhitFzFn2icuqeHf2n9Szk3DJk6Lg6VPOtiKUsaZj3zp0E
fWzaAiTY0pVz89plVayDg8fmNoGBfBFBbncqFZ8pbF3PC3RHgIFWgUtHtse4UiXSlk8BmBIBmAKx
lZan5KQIsENtFF7vOEN+wVzZL347Ug0S4kM3k6W/6V13ukXtM2TP7OCRSBpn9BVGJ56deP8F3LD9
jRknjpaz+DnHgLXVPrwHxYZ2iZ53RhWY5E5Y7ub1xo4Dl0zLLThJ30ihC2jv2foErpWlXfzDoO8P
QuekxAlnMXL6MrL0Rz1lvmyimNmSBTdnukIIijG/VVrDj60rqptASVPUrdo8aaIi7yXe2uRDI10u
ECkjv/M7HZMNJTvLtCLchbrIexOtK+AegsKdeSEKHiBkeTCLwMB+GBXJY3pXgXTYSIxSNDWNUE5Z
S5of8u/cPtC27LkMyQyOiW8leFIscj/SKABwTJ87rVgsULY6qBa9aNz4caBBNcASQG+7AQMYxc8Q
6Xj786yE58nIweEjInDbxUIOlSV1B6IyJx1E4fn/nMBndGGGkEI7kP8pHIV3yp2ctMc+dokyso94
s7/8SIp0Ymq4iAWrfBIkJcP+SGK3iKfounsgcW2Rh+ThCNUOzOfEeYKlQQJ5EBHE85ZqI2hh1tDE
doLS2dgFf0APgCe5VNunEy8QUYjEKhbVbqyBYErG/CHPK2QeinjOXQaiqv6CRftSsex4ZLjj2QOO
Zhxds2b3uZ+pEZ8AUm6SA/4vWcERp5nQzI7jl09AgdBxsVokSUz3jUXDKbYHqacFrArUQolOReg4
fjUYQBb0uHmZK+hYaM53Cd5sAWlUqbHtRfWcPET4/ToRwaKscWwoiYe4e3+vzJnI61hPRpReE2YL
LpxCv+msCdJ4D4UXDrCxQ5GNTKT9JNn8fKZ31tnXVDhVj3jIueswVz6XPu/3O7hA7hV5EZct3dl2
YmD0bmIDAtRFIKEIkB/R0JyqsU31dauEAUqJCOsr950/op5SBFpWieI+Ww8qrJHU740LJFOJjVte
8+wwAxSuooTduW+rdnsMriG+KlQsHYSZtOi7hITSIjbyvmkyxToDbsUPtYcvFvKvq/0n2Ma4T8tg
i6ELb3m+F7e1pAHWZf/FdfXwIKT/Mv3hGP0WTPXzgecwHKOPBTzas7cIY9zWsvjnz2I5uUdC3RLr
4BooHCcMwZl929ecdFFmuw1ZD5dvI4odB7dRypTHxXodwFgYAC7FIHH8VhbZBseTbFr9lHGCn2uQ
On2GQlF0wJe7jMapStut6/9mSTgP0q1o5fzQSA/KC3oEsIT5+VvRoE3kHK8vtnufl3IuLfukLHGc
ldA+AFdYj/fmpcMeDQmw4AfiFwfdMoOfsMmdDDVVDaHtIL5a34DAueAUAedi1jfIW5/CmzxfZtF4
/9ewoAd08xpSejIJ/N18UId8mxWsdS9onydASVQJAaBhWImsQha1sS8XxfD75gY4gAPvHyKx+ywy
7tbTs2WVWlMl1xha5BGsT0VYpfCCFCuMH6/H3Vpk0Qgq3Zk62WiWRjM7UmOA7Sa1qXmdvOwkbEMG
/6nH+9nG6Mc8F76wDTAqgWLFbFX+trz6OXQmOs2j++I9uh8Lq7ayqzo+4pIUifrixhfMCIB09q0K
hnDndxAp8r1XWxQ/ZT+jdanrgzaOTdd0t6Fh2QcZv13fPQXo+Ddzjlt8eQBQ5HLCFVyyQvATm81A
Rm6CiR1kZoFSZsQ1vGYtPSlcPrxHjPe+aNV3JerTiN1wjs09XvPGoveOx8ahfiUiAzP7iapbmnM0
/zDhtm1//qSkf/VtR++4TAiibYZB3kEqVbx6E8uDeeXLay9jbHG/5bRjfjE16D7p81sSU6JzfD29
xbQORFuwbqdT3yUKZL0TtWmonJzee115RNiEgE7/+YZfW7I8YXezM1Noj3u27lrD/5euLYWH/WbO
p5fGTt+9tekYjpplWyxdl38QbbmfYdjhDKuDKdKDInTipG5sjOeWodBnQ6yIpJXLA8qqQcG0eUiM
P+xpen5gtFWrdcWtqdvtimH41NinqEZ9KovC8ry3pjdT2FbrweB22rhEfz2Qif5YkfK1rEaX/uoW
kRzCcJ9iD6YjzDnq6dVbLEb956vc44KPWY2jvFTic2NNNVZBsjaNnqh/Q16ly/brVDCq8KPyKVdO
ZD0QXnKzdH9q1mjnLvj/NUdHVHx+ZAvrDDyFfojs6TETtFvMLY6kgJwMSePcuAkcZv3axQGDs5lk
2r2YsMkKsgVOiKoKE4PTc/lD9VRWL6kYP3LWbh/O3dVJ0EjWP1Vj+BfOJEPxTo6x5jaRPo+bpf6N
1iMQKiMzVMhxc39LKGEqiwxFGtoqcpt0kB+6ljrhgSEKxDIF6T9/+36SfziIC/X5jfOsBtqWMGHC
bXIqDXaJI16c/hYw37kUcO8zCYdLHUmUcvsJibh+ErXZ+QqVLOXiJHrKaYoIihPmKGyDlRPQuWS0
o4vPhKZaRHcjj+tqpiw4Sgn18PAxwcUW0/Z3GPJAI5Z7v9iSHrpSAg8qbwz1JCu/oFIEVdWoDlPw
yl6+Gvsjzp9P+NarYByAoYvrUVqlObRp/kj54Vsl4PVQZ1KLoXCFgLGxwJvSid46FK4VfnwQcVS2
y4OTiboSlRytDM/FKMHJpw1JTWHthYMNz4eMXtn0/tN4HT+auvQe0kiFpo15NM+56JkaTBYZKCfl
yUbASX/s89sAUrUnMqhYA6chSXMVv95nsNOq34M1gptxMbo5uhSvVCjlOaN6HjyGGbk+1VQik7M1
k+VCnRES3S5FMs1G0bwEZZPng7x2PG88BP4NlxkdhknUGF3KccvBPkho4AqBNm9h53o3859Y0oLJ
g5bERjpoIpQN1E3kaNjSRsEOmew7CbHO/DWMc5ER1Uidiuh7UjbOFG2bJEUodpgC6Bzkpau2U4Qx
V2PsOPQxlFEFFr2xac7Dcf7EMIPh81twfHz5cWkIcIAkCFd9rs65SY3xpjjzNo2Ztr2awBii2K/o
SX4I0oRlTkb0NipUHAKdGycwZdGi6iVixxOnHsMA213QHj8mjOzkf69riqVlwBvtx1dKMhtD1THR
uy8y6bvNz2GWZNjKi9+njqOPHIStYit51LiC1jMQ5FSIFm3itYIWhVV3burNZHB6LmOHtEX1vpxD
5Y34N/ZfsWrcXvGoEbkpWAXJHBnPoxWKbsfhxcIor+xW7Q4KYBnKpKq+6Wk7bEbT+5DnXWTMGXck
oa2pGYvbRhqeLAJFnNbiYZN8sAYiuLN+0Mnb7GOCF6qRjSMER1Tc/9+W9eb8wxf7lAv+TAuGx1HC
j9mh21HadwKM33Z44LRkEmKWidW98vPyHcvf8pGC0dIdP/AxFlN6OWZsksmjP3ojTxOByfrPx27G
/LYcPRFlMTndNDs5R7Dlpm0vrccQC067eYewsFqbH7E1+/hXCPmIWFmxSO4E4TZ7PmhhHoZxnWDb
9whKjalYX6GEHMTxdCUBRMHRszhyhxaRd/Gu+eyne2FKSle90QPW88TXYmxYAb1Wg/C/ezArWgAT
GoPOQ0SEl+7X6BRO7PQLkxJ9hKqU7kvRcC6rgsPu9zwJEgfQs5gfxhhxwr+waCK9Yb+v+aVATI3R
Evyj7k1AdnlNj4ebMk8UnY8tckxaLiQxQRncdGrlLizly1ph++EpVWpGeFrNq3lXCoXX0hp61Xy+
+g7ogp5H1aLwZqx1We0exBEqjNM9WF2qG4qymbRkVl7IcLpLmlfKdglnCU31DeZXURGXWbwHxBNG
XzkyNkuApR2tzEyzXTbP41oqN1CBRnMl/deTfHn3FJh6pjT0C9uNULBz7sOdA3TgEEH3i81Rn+GF
TnWPjk4SNLNWvjQSKeo7buj99KcN5ob8GUa40jTMbq+Go1udcX/s6jLKoOgd45y/rv8COgQNwVWJ
RMDz/G85aMryDX1SbphRiFqBrcy+/ExbS6OHgYVueRN+WKTiCUfZFIGWsyiHgD/HGA09gq79+OYT
8K+t/ieuBdqdpOhC/x/1L2rsknU0cd8iQHeNJr3aWWz003Nj9YVgBqtUWumJMXK96hhCDe7A/SO+
83PtuAYkuTB0Owlptb8zdHdmiu8mQ1+k4zaY5i0zTf/od6X92ttl1pm7KCNe+myxImU6CKYPl6to
TOIS/SrcwvTEfEHpQzmoRgsdO1658le/B3IBF7K1iECosuOP8XKPaqKYneR0ydcdrKRXrFFaT+qZ
sHe8VDy15f5F8teRtaj5liAxtgWp7IojNf1wJPdj+l1CdLeJ66JOhurHRMQfZaqorEI3UPT7VFyA
QBaS8yukJDiKQm5T90VB89J8m1popKqp6VeIgIRHI8keha6GzI4X9BhFhs0qeIbOP2XcWlWfazij
KDzW5b4N8F6MUdsIjZ7qLvKYPv2JavjzDzfMCTQZi+AWA+0CctpLe9gOn3he9VyXDtNyxiCFnC8E
x8S87gJ/eSPO5/8J+6AI7+8AqoPghq+jIHvfLprBtcS9kHK3e/5BUPGsNlNCjVe8ZRr0ptPaXkKp
ZDmn6rp5HjuTn+Zvs2tY1/8l/hU0QKC33aBjCKUFSVgRtX0+oGd6fRmVWFNccfGbLN/qAoKtxuxL
tHtctJY5l/6qNlwPqlwj+321RvqFBib8ofwLzHInWfz8xWmw9cFY1Cy7MzagwtGvncJOCB2WbRio
ihtDb5QGVZZgkmKJFlaltesBxLbXl0NaHKFq/uGjcUAoBoq5nY9H4Ciz35iCt/m3RNqtPt/dErqd
YfSvNjtKJzgvQ2/2JhJlHpDqUzr+ZYuEr79nBPVZfz3i4JWE6S9Nxf+a7Ou8H4awv3rlw3PpFBZ/
ymzl5kJLXXK8NaU0mVi58cb83xmg3niUeQYXQI9A4TUC4l9i6ll6uJFI2tW7dsw2wprCQRoyc2bi
1TEQgMEnfBXuomMOPWQIOO+vDq8662Qr2U3HdB4rgmu96H4bXXPfSzMmVpJl2CpRIbh6VhoiJHKf
f1JEVbWg573jcG9/SKsGDx0IZJy/+r+73Cc/2ieU8QEEvjAsSKFhCMehLOswhYPG5YOZCpJMmcfF
D4D/mRv74tE69yuJenm6amZDATIMivSIfR2ubFvoCq8i3YhPzuTMLkkjm8yuCvi61+k0hOVswnNZ
ZJurPYwq70/GXVKANaJV88SD6cGz3M1cCEu/sdENRzOzr45J4GATcHIlibJGRXRjvcpYhyyiGs3S
yPXvRzD9HjiprrAfEzve8IebPky/2bBuod4MtFcEvOO8gRRr6ZqEJSyTaZ53wgHglSCIYCLdbW5y
BrsKb/mXEhQaJwAY1IbGHpyq3cCtblySD4vHT6hhJgjiNGD7g58lOyylnO3XGvx/F3HBshfvjD5c
gHsSBtNt7MHaThFiDqU8AaLYqNaUsPZkbvPsiRHx8WaUhsKykinRuGtRP6qkzhga/eDKDEpwZIzA
RzY838gVe/KdYfnUyWfdao37YHhcebuUqQhHc/do9W4DKRAPlDtRadKyV8z8GQuUyK3VwFu2fuYe
z9hGcf+JswvHiarl9l5kNS3OO7lu7Iep54cZfef9odQUzdG5rBhrUn7c/5QPVOBdfVtuLAoH6yxs
0HMlvM1alxWhx+TXwO5fcV/0Aunz/gUJFwKcaEKeHiep8freCzlK9AJ5RKpgy8wYukJaODOVjQr7
3t3/FvdwYvoRmLlNWu0gDPjvz+yKt1KmOBXK+6lNu1dtjVQgd6ITVZYNlasFyCl4QgKVB2f/Uzmd
/ZQTK+hxUeTPZlSp9JnMzZm9n5cbD+UTFvUjAlXQUlNcfrW4f4IOHTIT4UGOcDpoh0bf9o9inuMk
MByXgrGERefTBTIDs98YgmXw0mkZGfo5gG9BYXNqT8Gjj9pvlFiTku8/otOXnJRSgZCuDUO34nFP
ka9nT7PzU8D/ybppJFmH7ynm6i+YQYIVV+AgCzRy6YeQM8Iqh9SQKlT1Uth2oGCm6/hwsvryruTa
LXn6oEJ/+CdrQSnKQoNXOg1z8ZXFQrXjZoKzyKcn4XLamB+kDFAikNqxZ52j2lEvOxu23FiYlcRH
YhFcEkr1CIXWoINYQwzn/k0SHus2BE00d/qQKWk1d76fohQJOE2E0SVGx+NXRKPGPsPJxviw2/+e
KrWkCDjujdODqALEEUCEXs0AsA6sXyeSLG4v6sKzQtTXaUgQhiO3z266CZG03MWnR6rw9o/qpbwW
bcOSwu4eKc7UsUsKTvmtQ5aU3diLQeZje7vFAB9sXgXFfhEuQRwtdS/NA7PWiNM39uH0sH5stkyT
HKHnsLpv3HdPyQMU0hWXjWd907ZoYGSuNGye9M5lEw0W7gqUT0Pp0TKdaPY0j3wt6fHmyBqyjarQ
b5Kk2dMOLX3NeWsEE2GI1fcBrVB8uaU8Ukk3LDaJxHP8HmDw5hWjK/dXpdGZJGue93AAt8DB4ChW
tlVG9lbLa4EJ1Ukb3R/FauCubfXgkP/gIu5y9xMqesiGgZoCPViEKZjpS7UZqevgoYE8Ddew8nAl
rrZJ5HVTwCYbuUSQ3Jee2yS9/D3PFA9p6dYveDv/WrcZpaJ1CEcHuXpcQhgYZMi6V86ROYdEeM54
0ruuVsr8LysN/q7hmkcTvUlaKgNB8kfxW3OycurIyB0ConPNzK2Ey8u9AfYNjtywsn36WYPjlFJi
3vwUs0AJVAqOPjT9Ydo02uiFBHYagS3hc6LHk7FOurD4tXasDj/u+sbP48+OdCnrvfvvPm5NCMmV
ExxQpX3Y6C47BRg+jx+1STwQ0YbwHhNmwA8WXeLXu5y2zEPQUy2L3RW4tp5ByqNNVKmTl2NJCNMH
I0Jnw5cM6Tfx7ufGdDNAQ5lHL0IF2nPWXkn1Xeex+h4Ss3kvBS8ajdvEbeyWBBadEWwPRaS8eUr2
WYBSqnrhUC+4B+1ZhVkOGTHdI+JAZbPpDKhLqEVsKuGDhwa5gjaHJI76vxyYn5iGzZnUBsFw8Jm+
+w+fWxMe4DYY55QMV4GGh5+ULXSpuNMSgLXjkrUHQrcv8E3eCLjGiQVYcPIwbL4C2j//g1d8KVF2
AVaYugC+LOjb/fzrx/1zKPAMZgik6k0yE9uLH7fBLfT0Za6Pj0pcwkFjF+DEdFQsVJqMNE/9LxOI
EkownresBR8IkSLwugmLFwth/3/x8YaD32RNjecLzNUXPc74MyeaafIA6CUPpQPwCqFwvtgvNEhX
iddRpHwzsM9JkIKXngZyAOi/R/qj8NflOxv6MRxJ/HC1O0IoZGZBroO5Y+0r+zEfv8Z8cyK/Sse0
PoC4h/s/1mTbBEWgcLnBrzoADDwCA+uAMxxp49v8XPREiw6Y+gFho+a7nwtbmhHziRcaEKxNfZdQ
SSl1rIN6bvzuPQ+5LgDW+sgqbLe3z+jzJeLzIArpzv5wMAMphFHT+62cocNTtiOnLCua9ChtcCCh
jgwvqF5aewy6070p/x5Ax1OVC7+XfeXffZifMmDbNswmgEtDHcD9JyonX3L5pds53sGq4g/l4NhG
xrayYb/rdwTLguENekEX8+n9kTWQ2RiVPFF5COk/PsIenqEwKR34tRABVrdLS9H9L7hUrDAX/VKL
6IURD48QZmyauVTNhv6bh9IN5jRevhZJG9CQMtYg81jYynkxHt6U5IhpFMAFUcgfXBsAjYuQan2M
vFFK9ie0tQsL/eHVSfSOpGQD5LphLNABLxsuQgCknIT1rl3cRQEcQIIIeXDtHsODOZKTRcV4V58Z
qQzi0K2E922bUXFMQnZrW4wa7XyfwcP6U0TG4/pNP12H6nKkCUi951QUmYng6ktoPatOFqa/a1oh
N0R3pzXDww1wodGSLWv5iDwuQqkXgNuRNmPB7nuB2cgw8ooZS5WdUsQI4a/M0ksdPnQRZlCmPzIX
2bofg1x5AAU1FDyGscSxQpvsFqqIo95o/w47eoPFIBXrVLNmSbfEKBOYXkPPhkSwszrIrHOhScGS
dTeX9FdnyLoe9N3wT0kzn7z7yfIGuNxryywHtBnhWqAtdEClpkG0MFKxfbeSKjV9WmFF2Dh+14kX
68/f4wILHQhaB34ayy4qNzH3k6QqHz6ILTmJpZXmBaUPNl+abxhSvAoQTn0Ie8eZMbcad/KN6nl0
+zetAj2QDTHCa3ZMudjzFF1UVebVVFAI3o699M6QTiD7liHVVNHopjU78g8/Ijds8fJQIiHoX3Bw
DuYUiO6qa7N0lWAEkxGb6L3B8Zl+2Zy3IN8l06c+y0JgYYNpIfQvpNyOkav/JJwSG2uC1fPOiVQq
8kW/swYfRdE7S9L6VnNtKMGU6BghODC1N0sN499bW/G2B7Z59QJdwBsuY/3y1WckHqJvWAwCL65W
OyGHTxrMhUMTLfaaaQLaqf5heeLttIZQFeD3FjDoeDid6Qe9eWZJjgUyVJnWbu+pCSvjZVhCDyQ1
Vncl7v+Fif1AfmqF0Lr7mKdHO0h6mTFld3lHUGaIahPJhOkQnGujhckkrhSk9OgKPL3wfPblqYle
i6UvCY5gYVkUTlPUTpoNYQV/nVhE784HnKqcm+UnYhErr0+O6jVRL//1oPMPCDeEGrilkckBd9SL
uEHGbvYgArQPugE4Bu88JQpTUHfyQlul71NehAaGBqwY653kBdxIeb30BcVtJjBSSuXX9ahsrZk/
Y74PEOKOX3EFdTGDIML7yIasvz7sH8gnxdZnE9LbU5B0vghymB+ctJp2wy4ZLVOBHjs/82cANsxF
MvZGLoPU+NsVAZRXy/EhIEAiXPiGFZ/lrGpZgQ34QzOWLXHgjkECLKnskPh3bJw2+z3zagYJKvkI
qCQQmQ89DyQTYZHc3GtHLqFQ+x3roZaXJf9LIi5gt+d4HW9Aarc2i5pxYUHedNJgGVTAEvYTJJeY
W60hPGvCewNVQkGV5KN8TYYVLoR5MufNDB5IgLjHhI3caZPW1nIYBy488s9I0P77DVt+kxHwP5N4
6V/JYOv2ixp+P+Dlp0ESqu5cHTwySjhWaNrb587c7YYsdGBhvQI4c/z485/qK3Q/OO8cIKR8ALwt
lvfXABWJdGNp0TK0ezjldVE1ocsZrIySk63DbdFHPDAgVwSqm5Zl2poisCGZvPYNiVFxA0O5/5yr
Hshl9x6l2G48dvSCTjBaHTz7cxRm1y++ItpgfgIzSEJegXBcl6e+5vApt8VKJlM1CENhzVBQZpnx
Y+ceOdnNDS1gZMRIU2D88XmV1IMyAYUpcjmt3ICpp+d7KGe4wO4CSdRvKDQhPhilfJWPCFtNENK+
y845K5Jqd1FJ4dPOn3+bw1P7wB8bq8FvAYICv/IAnlQZaoEVda1s3STMHnGNip/kytxmNaG+T7ZS
KMxBZVYcm1U12aWs2Xx6QVeA9q3pGadRZf3gx9kY/A89jxwc+WQHrybF0HkhSP/suYdEAQFYqhLR
E0QH8MTS7XFae2sLwKXVUb9GLD0Y1bWLRgIWeB9oa/vE8iD4RsxsARn/vk5NIj95dxbEHZnYosO0
QBjgqdQUBbR+MEPaW8EMBvJMZ+m5BIO8/XobpggyYkpPbmyXyL+YEnql/y+JStGO7vLWwOBti9vz
WwijkxpkHg6N0UGVuyEWtmCnusP9SEXUqhhIfpApTtX9WgobC2OZNmcM6D0bcj4fkt36eFFgYvet
W8Qo4Ft76ICsp+eHp/6G7Gd5IrspoCS/vIyIPdUngAV5tH5zSsbCU+sClsYrcB/xibGSXkR9gLxS
eaYtQzKRZcWK/0QUNAx2wFPoJkDtAO8qNz+xGLpTsp9AkpVuWZV31LTHLCA1iBFmU2N0t/nI2LwX
HMbg8dLmE8LE1wvc0DaDpg59LQXsw95/dWhUfh5x6le4CddiIXWNt1G6tilRQm8hpTGznbfcryPO
yQW8hIY+4H6dLkYygUurFtJhHRbsK4Lras3PmLs43Zt5sn/VsbkwQzvWNtVneySjupkqPlYA68Jy
nRNpKzlh6Rws3iAhiwxlHq/4P+T/nyKZATa/5B1lo2Dc4/y8Q4+Zuu7MWAC/nkY6xJnhUEF1Mkmf
NFRhxPWADSEXVOYS4CrGiVtYBD0eYDfhO+in0182iHjr8s/WD8DYIlU6Zv1V0ZumZ+MXoO7Z0crF
tXmiWrIHrPQaw6wFMZUlsMlUCmLbHpFWTPzGqqyvC8gyYXmpuJubURHlElVzv3i9Ar2foaR7Yxs8
y0ynWHavFPUwLkX5UA2F417m+C/xePL5eUapzd1GPU7fK+kSQuI2iep7ZvzYr5y+w7IsEgB/S/6T
1EIAS53/3UQ8oqN/DcG/fxSMdX9DVRxMg+LtgdBUJjufI1ydXDuW6tSs0G9zZsZYHARAGoJGs/1Z
yg+Sv8KJe/gzzS5IfoQfl44AsACQIad+C40qBVtSoMdFs46sTvS+qXoUXXlLDP4o5B8HkUUOc7gC
+RgdeuZUh6GYbQHzv88ezz8Ki17KgBgH1IMnd+AamWbEOX2hhDRiGS13TW7uWVtqowIKoV3p3YZv
kw8SFYDmYeptbqKfW0Xi/EWuFZh5pv32YWYv1DwNxwkgEln/1czroS59yW8ykGOtMy/iwm+EwOEr
SXyFWpVYdoE4jcBHSoPVpMtHS1jJOMUa9U8Oi1BwKiDGX9xQQyAF5QQjsjWcu1BAdaPwhWKOKcgM
2pXDcBU4X1UDddxtEGswG9vRZtDOEwWifyRZs4PwWe+V+UJcITCsQ8VVUhN/5hjp//rQYRKrsHFV
c35weDapPJYLVQiDIUMsx0A506ou2Gb844Rh2g6k7DnYlEMFsg==
`protect end_protected
