`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ch9jB6bPy6KffkJSzr1VfMMETaEtgJJUKhSx5d3HoHZUA2srR6apVHHYwV9FAwpejQjVGsH5GfCf
D0xPNHQK3A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n3mIjCvvanIKVPl0SQoPFWXUAEVrLY7i2JQvYL2UNwU493BALA6tcSTs8YB8ghJKa7VJrXByj8pu
swoBmlOgI1VccAzF7IcQYGw62Fwtf0EbUg+kQ+QegYAYBtOUMBAMvNUWTVRsGDPJuLMZKKgTlSoQ
YyklVJ2hLF6uIgTJ7C8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H+7gVqZq66Cg9oDzE0RyFIJ/eNT6OeflAvkFT4v20qiry+Gw8quHQDuSh/QCeJsuYVvK30JrwPHK
e+QDzUSIPjLr9CsuSuKifzNZzJLm8elppD/UCZ0D1in9/bRB4Mb3wh1tBNQN4r1Y3CC0ZJG/jmHl
dv12l6m7KCCQgGBgdQXCYPo/1qRHg0bakGNbmRcYjpr1cVrXn8qw+3Dh/HjKHqcWeXyu8zzMxZ7U
w1uVM0S+HrBeZV96pxvBQzGzm8f8u0FIzAUkjoo/wpSSmlusRvf9xnyrgpdck+kMM97BBN5xhvGa
6vHtrFc3kOyk4pqKYiKvhrV+v+d76+Ula/IBGA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hc8zs9UarlZ5hATlg4MhVeBchT/DV1dIS0NF4yqD2QiphD08HMWhZBp8x3lFg+8s1z1Xwi5DOW0s
syjcbooWyA/eVrMzzc1DznTwpIXLejhCR4bKyfIWnBfOSxsA7/7k11h2apiw9eKaKpcOyIaE8t1f
0ao8Yqa/31w9IU6WDHo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AD5nada64DyjGv+zT1GzqzTaUxKcTnh2fmmdf1Cc9MNYWdveRG4vIIMXlpCxzZt5ZqPI7SPcebUg
2HYDqoL7oeWnwu9mjQLNB9TTCLIVeC/eO4vln7E8G3KrWhhT2OkPysk/dMGF1Y1GNrqfQoxIQ0M4
UlXIHvTuSn6tXX/ZFpbKXiLxjIrbWvz34TBQTi33eZ1o0343B42WTRFYSQUdG1zVQ9mQDD6gVeWH
rSW+eE/Ce+/t5oe/RXgFNLZ2iGgkmWrksz4MNhvBh/vYfTGdVwLlcxVkR4GIA+SDIvtGd+cdqgp1
XSXl+Q6ZDR7vBENFeqE7OoQmRqw8BJGKCf6Vpg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 82816)
`protect data_block
c3Ga7FVO4TphgtKbT7yld3cfDRwhpnA5xQAxgWMcy7hAYsau8j0QHelg39CTRLQY4hKW+pSWl88N
San59tmT8zTZkNWonU1lXSskXEzuLwg5rhX708Cv2pTmFyjDGWMBaTiq4TThjVMx5351CLgylohJ
kUnqjx0tnjupBpjkhJM8Kk5axNiyZ5oLKp1ZWLSz3CqeiRBt+HrvO96S+un+OVXuPdDpwm+omoS/
eTBNuPjXHM5FZ1jplcdzY0iD8zmZrzRurrg2KD1D54LscKp3iJCLoeQpofvnVivniLe+qJcRV0th
UQo+Na6UfCzege4UQHP7lnUZXLnWqDDploqZRlvhXTiP4FaYHIk5zGOL7vgvLe6MfbswatJPcEsF
30t2JvBMsaYAGXrchmz3tMcp2PfFN2KnWehYdc4S6lMQ8V34KWhhFfHAXbwIM3MDUTZ9mg2NxaMC
W0kRRw4vH1wT2IrPR9mIQANsu5nnojLQoeuZTGVNnk7TWOhjMQKfzAp7Onj1xRT1Opw2i+4PdxLg
U+7eQ6ncLFSZt2jeehjdm85xp6Ug4eJL+dC17KdHpIDDigu7YKJpGtNbPYGRQMasLU3wLWjOoH/p
JldnDfMPeV/wNciFwOvdkyh1KZJBaTCzzvAbrWXiwwPRJQXiOIW16lJWEE7f7Mu6kcZ5Fd05tUXC
j0CliuT49rs3qn6aJaK1//+5ruRPSJNhXnQx3Nk445UfE1MbmpzwQdCBAPYsBEyFDhv1BTm60LWs
XGi8RG8AAu5ywEM65kY9KL0xBMhMMVpcLbdxy2tIIvkRPtY6X5JbPbNEwVy2vTQWxzgyo26u/+UN
HHigc3odVShytZEupbdQ0lCHxCSVK1hlJ5SRl285qEqpZeYlrvyv9VgMtHhFedHqmxHw00N/NETk
fDaZe6FW5xLR3uxtR+wHV5ZFeOpj6O8Zvp20NSbFpmpXxM8JLuMYhatP7zv0XtK6oNs8B/SenvqM
K4d3sKq0HwTuB2yA8fngk0uhZHSGs0KIFeGRJC4PL0zFD3h2c2tBl3YkkGwg8/1meennf1IdCsAO
CWM1tMvLzA2b+La3NafY1kg/3Q3MKAhxlrCtiGExs1bwQEf9rURgK2pArzGcWBHECuIrQOUsNvWO
Uu6wvLMOxQ4kUNF+01xBOhC+uyH60FdKq/6sstyert3McuxDgXPgiDm0K33OFShSrryTi5k4wVB+
eTLOG9ePqB8qVJsqymifdE/6D+iWJeoths9cRJYSRT/AkrPohJqGi6A6Gy3MfHt+61YrTF8TDpKU
U1ILi4DkQ7oxmvG9BU0lhtKtUQ2huwoANd73/Rq9a7VGD0C+yduQmrServri9sYTwD2ZkUR2C+d2
7zLIJ39Hibp/8tM0VuuQ3X7obaT435+ENR4BTd/TGp8CA7VCoGeUUiqsTIp8ky2k/G/3ndW0Uj3b
LcGs2wIiNtUo+uZTzVMpnlpz79OE2Gp2+k5MjPFVh5zOf6XjlOBbHloBxGKM5PxYel4qA5u+khjq
n9V0AH5M4XOqkmMcMLZ3st2JqlfiVkOGc/2sSh8nOROOBDlGd7BXr4kppOF41sWkH3podVmg1EBd
Peus5/VMIBRrJF64nwvmFq+i/TxWc9EAxAgzDkrZ/vaGVf9NYAhcREYlhVDuYc2rWrP1Zairgxxu
Io7iSLeBQiR1ojR2j9enyhLgDsC8bDXknLqR69o77QhIvjOCdBgFmhGfPNNsTRO8JzTiILjS/05j
3QXRl/dGj0180JtT9lnLdmNuWCIvhr4Gc+rSFAO4rLwllnIXxgNjDAGKq4lZ7LX4QvHcrqgUuJMl
PUEsNPONf5kh/OrmjrfzufXo9H05I35RPuewtZl42dRz26BtxgDdkeEhK+toocBoZAn6ymjV2cFP
EYd+4ABSCf5C4wLIDvKgj4EtQ8jLkHwUg8x6DdKPDsB9VLV3YAbpVbR/+XDquUo4nSj5+aTGSWkr
joAXskWrTPOy3Sgd6gAq9jGF6HPTHrS520KTWlzwsB+8uNYa7punuYxqbuxHDPJayswYZ1sTNkxo
tViWrh0ZoV4rAQIe/NNL/ntZhX7IsjbrISHLgznFXRajvLL7AOM+4AqFgfg1vX522OnVTw+mUzF1
DfcP3ZmiQHDn/I3qtS76okW2Tw5Y7vsEkhGuqTqk69fVkOZTASSfOjVKIOIqYWNysdWeVIgkLAoV
gJLatzQi+YfDhzA4UCl7qgtu1Y76qwtaiMNn1PbLEyFzTNW9WmJ5lLtKUNwB+WvaHvMXjHA5P0Rm
ub2YYHWmdtQ2v08WeMmkja07Q9ReXsaxXFNWqsaRdR4KAUTGTyHSo/qyRge8k6JgaFNPAnADTU1K
v7YRhzgVBBiixbLT5SDk6wXj9pndEWpawxd8kH2vekdpauzJuvmZQhNzfEiOMxzZ5/237ahZ4z9K
y2nYEHxhc9mI7Ujb4NofMmqPLJIgfg+QOrT6GryC50StXWU34PMv8vnjh2gsHxNsCN9fRoHEGKqU
dZEx2Zbib6xn9JvRlQ8kdpQMiUETAS8/cSHlEE2p/2F2CpE8PE4V1LnRUvDCW2dDCb/YALUKGyFN
ymMzODIQiaZNy6WF50njZXS3KSr35lqA16xQIfjM6h14FddGLKpg1d2lVCmytbN0GzfeIvSD4T+x
FG0zXsPsGYWNZIkUbuXIQRvbi9SY/Inu65zlJfT1uj29kH6SDGBhNECLpwiqw7iQfy4K21eDKUns
Saw+3xyLrNmCToIS5j/p4fT/KzkwXBvJ93Kwvpm9Y4X73fMcOhk5Uw0Mdo2LxacrYfPGBXxQ8hpp
NeuZDWGExiHUkkj09s2/mGoHZKYNK+379GxSavVZHYwlGTCk82lXhQLfg92e+e2TshFHngBzSNFa
x0YBftEgv9IgZkp9RT7B5lRi3w2wWnldxxuN7sg75Sf6wNglXRHRkX82Z0DA0HMHDQMJ6N0HFEoR
DJitzCQyMQAT8esPvZGJPm2Mbcw1Yej2v3Z8WOVIX+yBi8B4EAUYT/bMkxHp+iSNgHTWTYIeke0n
JhLbNRSSgi6ji1Awu6I7q6SgzKdhZrTGsRkIp4hSbzfTx+XOsxv1sb7G8VVihEBWaxUBn7N4mSmY
Z4OeAiMJfro2FY7Sf3KByC0LrYdvvne48lEC0olYUnJOOw8TUG4CTK7sfIDItCZwzlE8wGAPcSN0
8/5g0g4YY0Mt5FopOm3U8/mtqVsbzUXhxtSnigoBY5ORp5QvfQNIjxuZ8PnC+6PR5PS1u333/reV
eKvkc8MAlOY7SJ5ph8htXP2QNejWPCA34HvdXn3hJ8YBof9OcgdCnPpeRzW7BBeVxTLBJr4DxpJh
TeLRQ8T0h/k/hRx1uV/R+QwbCPOdKaSUj7IUkcxS1c+IXGI77fCCArhw2CID9nv6KIi3bLYMcT8g
a5zJ2iirgMHBprf3CbTdanC831CAVdilqzdun6F1nSCCIH3mCgVBvSJrzr5KRHptY3sjI9Tw7tPy
kp14mA9sMYHCjh/5VXK1xpaaOh83/u4+AnM+BhzqHCyV0BjQP03T07naa8oY+z5151jXwNzF2lX4
uWqPAfwON/p1BhIuTxbfZ+2k3PNDmP2ZZwgeMYEjKVuP/hYXrRWMZ7xOuFT5QvN2WVm5lc5Q0WiX
RAMNXcgreIjYLv+rsdlDH1eCbzLUid5rklvTifci8kFkDPr6hYGmQ2gXg+OeZpz6bLyVWVjFnEYQ
xGiDNvtkEjA6G9EaXb8/QMY8aMRoveVwHMgjAKaV4miPFGcbm+UBx5o4Sq22OqoqicWVNV3SPmlb
KzPeg9JnOZWLhfvNoen9DEabAjJ8VPf+mdjOo1Di3tReyKBI57mTFPJehMhEVHBnxzUxv7UPKGlX
j9VwOmaMY14qGNKU7FzU2YnUn7yXMNeyNtHg2s+kCcnRFSqHsjthTM38/Z7whr2vUwQEattxDJuL
y7YjfZeSU2t/CNNUwwv7jxbre/a986bfqPvggDk5ALw2vneVoKerVRsJKDA3qJOkO5/a1uKU1IrV
8WEPtrvbd16g0JrRygakFT7o6BvM5uG3cpZVPwKK0BrKRvb5F761SObl7zyIX6sBfJxoje+ZdYyP
8mDU2wumMA/s8wFvIBQhgKrz6Gxt0hPaziRZZZsb2NRM5bqs9mipuqh8vuQ0KqmFDVq+H7Kcx4nl
xotGTculdaDx08/Ptl5zi3qyyPg4PzoLRpV/dscUGO9oLFuVBElBw5sUE9MlpC4YrziYsF4tH8JZ
8mCECLvlw1MfEUT3txtMrPudXocqVpS+HRF+gOhVT+pSR3f8tCUUNa/O63ruwapV8p4GMVOBKdQF
rwVQ8yrrjtKSYmlMqIdJ/GFKbLJDkLPi06mNdOPi56ZgtFMxb9xN5NsU2+MsESQ61M1A+jpmpN8w
cvNpqYmdUhF1XcdTOgDG//J4Dk95+Zjo5luY9PDxQcb8jxPqw0UFnhyrYXDeoVtnBL3nVh2xFD8q
suxzE5wkaXZEroRYOnlXTk0An3hrRJJJmgC0bGv+w2KlQ/iWB152fWeMzElD50CeTLJI9Jhomxp0
rT2WfaPImr1GEJxmEva5qCWprSX3F1J2NjxaYRjDc6FZDnDQzMRHxschzfoSPTBoWtEZidogTwof
f6vx3rKbsY79/Lkr3ozIFWztpcVynEKZX4N1wza3B6TZ6TrlIe4+95fkIKVU44RfHMy+PUpOhuKa
gpPaD50IGIdY+4nmtxrQGZ/ANK9wv1vWps18njvEG3Mg/k7zQNJFYLhEOcI4KSrZYkZ+8uxZQrwO
EsEBi5deXRyx51aEKkI5zubc351xi5aD5EiJDR1HVu0LJ1H5/6Ixq1Qtmo9GPyRP3IULa950AROy
gy+kgY+esV6rxUvmlpProbjqAeqI68lwTgIUvhkBt0SL167AxKtaz9XbFaOKESGfSIfELy4k1lYO
RB1GqVd7ZFLkc60Vnx7rOJk6eJBMhC4HgAwy9qZ8vI+OmQ8MIfVQ+hUIKPezR6OqNUWI8JKJVrcz
HcWdTfwS3FEzkxs/yFxH7H0k5vf47kDUwzf5xGX2ggm+zePB9KrKeEYuiEoe7JX3L3IfhoJu4guk
FnJ5aEQmibXG/ajEo9t76zZakTyL0Mj5kf6W4nyNJDgiqhI/BKWAbFCT2caNsu4DC4KPWqCgu/7W
yLJR1xX6rqPEqBKwPFSByIPQDD8uT+e4XguWbPd016FLbjoSD9YFxsOiAEM1FFNAxIGXe97M/DMX
qLV933CAzF2z5azp2wpwF+lnJKkyHKMSozUwHjJ7pLinMYZwv0bMtXCbCjl6ztcMsZKLwSNit4xF
4g3ao0jHDOP8ZzuuuF9JfKaAoOx1uXiRVdVgrRda56L7n3+k6sCstDs2dXSF9ov8+3y8dJo7FrnR
MmtoBjG/6IwjgA3BSWRnpElrLEMtzZP/U58SFam7q2WEAv/0H4GxywCpl0Gv1h6KQKKg8awhFf4u
2u1mE7rjpV8TLUscrctI7Gsr3ts+QlR495yhwioS6XEawZLvAkBfb4pSDWrtxTewXwym1DXeGFmM
e3FpzjMKz/jTMQFKkUQJUBsAHds0A6MYSuq4+rkJSxFMFzcrnWgqS2Ktz7C75bl2kddV8yT5/mcc
bSzyENKfxUFWTfizmY5qgYrtColfmkp/w9TnJrRG0EOgMJclT2T3lqE3bW+m0ovRF2pWvqVscRhF
wPJc911BxY6W7xg4I34ytL6hws03dpRLsdjxPd3VKJJZOJ+XH5tZUZjf74dI6vO3XZDXfPh/AzT5
ieVfMFKtxVGZ5e+WLOTeioHSC0BvymSprqD9f1RHrenc2NZ/gNtZ/C2wzjK2nG907E4xiId1sz5X
Bn9lHGA/5rBpnVwMdijWUj4Z7bzjXIlR5If4RuG9nhy3QvS8lkEqxrpY8VqFdXZYEFgQyu+c4c2j
BM5OHJtNdSkYoyWlppxQGV+1N26DFn3ep0t83nJJmZtIv2VdHkiChkKvxkEDFzR7dsAF+loJyTHE
4B19JKaGiZ/7aEZoY6h11dxKDq/EBVSoHOeQUHn9KzDMJDHb40KMff3lgXEaWOCUQSUvrrj4P+Yi
4wv3ICIaEE9k+Dsg7iP7uv0zAYCEXncEyL096xvXkcajENtGFtsmHt3W0xRmVZhlFXimuYdG6oRP
Pthx83LJnDXYs+CoRORC7jsU8k8VmYevge99gA+QlzeBfpNbTX8aR8BzJ4X10i7RRDQhthhpIiJ6
/SMmbrKyCk1QibbpDEuys/5lqkUjhMT53DbZCtj8+g37WP2KYKFJhrr/ZRKZ3uM5oSoM/uZ01dFR
/g53Ruda5o6TppssRdvj7SgKE9fhn1SQDwV2MuMQFUl7oPV9cLKm0vHnmtx1TBIJm9r1oRKGCHhr
Iq3dyHZUR9JM8TwwLUK7BNdZCVpQDvkJp9SF5sAO8l7RDc9xIRxqIypLVGChbddj+OY097XjpOm/
05qt1ApuQTi3roHVlayTm6qIA5IQ2FyrePkDlNMCBB73AlbHNbPJ/IhFGUJxW/5fxmmq61xQiD3y
0QdCyYhW3x0u2AHvQz77VqC6oBUbD3EKI3qZh66/+sTDYp24qA1/mCF9rCaCEeumbR/svx3hus3b
4q1W3VS0Rg2JQuYokeWK2JPglGRw2GhBCUzZk3UGFo5V9Vbg5YP410C+l8ZlrrwXMgCcb97ckfCm
uUj3CXnCYc2qfnLV/Ak2xJwKyJ5P+NgK7OPFgDAtJtBP4iij33cwoXwVsEanxUNboq5RD8ngi3+H
QAfxJ1RV6ln3bj9ZvjCKDPtofGZ7r6bVvgamEKfXqAS1Vp/anQ0DkE1m2tD+JxSo/DCzrVfZVARV
2MnvjdzCYe0nYtU2mFvl5xPiDD6Bdm/b+CZBz8HPTC71OYpmqU1rfoRfVtU7azMdYi32QA/Z1ytc
W9s21sn3jrqlBBHc3BrN/3Eeq9JlPGGBN6HR2OwGVoNZf1EwSLY+MPR4c8akRZGvhI7kUiihOrH9
vg7ZRofrGLVMS1FA/hnRfrmTEQP//SH9liOvdqyDFsSB93rug3i/HdD0UAcfV/LdEv8puQ0oB9Tr
JBKK3zsW1UTm8qkHUgDXblLdqD1bsJz3u7Vg0hKZ/wphSq5PBpf9wlyWDkM4gI0buNv0zAFJgbM1
6w3vi6W8rHBpMScuqQ0xRqU2JvBRsp+JGqI2MPv4Gkc8361dNSxDBHvlE4QRURGLqYbQKpd3NJI9
jj0AtBvyocdyrKXqL+rCwlIwvHqgRezGskeeNwtOWQZHXXv9ui9Qhexcj/NLspDVSo0Udp8TSAFp
+3xhD0gIWhVkLc9JcTelZJ9P1j9qsbXA3fXGTx8DALfXd79tYubih31frVdk4bxs0deeIWC8EEQN
v2UwDPPtdvKUQqFpNo7xe80xRgK0qw5YOldFFzFGkf0IEe3qAI8LN5Q1MOxKylrll5hyTjN8LXg3
kkP9RZnNIpZ0Mcf15cyzPkKr7cO5oe/ny/HcZ+cBVsoyZ5XHTyINIc4QrGzBQD2jE746ND5L4V22
dNzcFkS/koSv515X2x8Yrx8iWiq9qw2SV7dAVCBiNg0FkKavVIfzEa1LnRZWdC2egD6oyqYLUwmF
V80uVw5NjdnWInWvu3H5gRGbiOtmm90QRFe5JLQ7XNEPTgqOM53NAd+5fc2yUGBLcDMH8PEpk1ti
8cDHB0hm2dhVJLrOsF9IzP/vKrYIrUZ4p4JmCf3vidRNLz9W0dqRp6L0Hfeii20J+bxNb3Emc6n8
EgBu5Xal4tG++cOt6HGuVhZ6W+VDvuMYZKTdUnEdX0Gwx3ScgqErsU70QKVEl40B38v3nvtDLaws
CKzYx0OyCvcbvPu2lqTLVmtWtxAyk+bEEZFF0ugSzpfz+OI3TzzGWg23vJHmVFXHXBZv+m1A31Bi
WLBwuaqneD4EQDyJ9z6D3MPw+PJX8Qt6EryqKo2XzScu6uVCpcr77BnbSCHqCHb29dU9Jo8ICLHX
GNFlq84OVxLZBbLVB+81/AekIeSYPGIVRBcG2wuI7U0vKHBWw1VBmjKwS8Pfi84MUyQVagktLWeM
Ge7zjttvvMBxDfkQ2QeH7YQYjaR2cCiCJ8h0u0ZGlIrxB8FRgObmayjZQUb+JK8W9MN6UBvRRb3F
+7Q5Seiv/lfBb+J5uGxPpGLJoGxTV/ia6q90+t9eUXew5PjsHgGz6o7y9au+K6+BeeNCHJWq39Sh
aQpaW4xit8WfUup1SPd9fvBHMqpKHVOvzTAdmmYT9krAHzFKPLlha/BjQTQ/+J8f96NH8j8KU1iy
oXs9MIzenzULaf3+EPeTRRMHUXhBJKFXbhUgBhcVOlNGWD5ebwgstSgDywzYPqui0KFguB010Dxq
SpvYfhWTGAVj20cahhz1v1rbWlHbzV3/NJpQPnUJf87B+8lKVAUW0LmQjODloMkODQI2lsa13qaF
/Bya57wU88f6OEaz2TPHU2Lx2m6uztG4H0VImqC7snPnI0pPnQBl05vuJsnIUWIpno0WkosHl49p
gH/micTFGWY4FVG5XfBe5ziSvTm5iPI9HcVoX0E8/HjggpGQzzDK6BeW/5V83sUnkQSAiinRRKcb
DvU+2AtE7oppvlQRcGq+HQJDZ2uMrXhGZSTTvL2MSetBXnNphGvRY2ce/mHcnAv1VBXEeKhIruR3
Hqgaza7NrCzM+8VsNoW7f+M5Pa+9mG+15evVHlbLMN9yqhf5peX3kKIMLNgjAaEs8wnLgPZp/iP/
DdKFlEiSRasCDOCB785m824i8g8lEfGuWqFXrlzHdBi+t7h4/o7FWT9q5vpkA/5h1T1acHwtv3gD
/Cx2Q0spi79D1e4vvqEdsZxY4FVapQ+x7w9tWcWwIflz5KO2xXNWqxfhSqmoh6BWx7ybPoVyKEpv
by862ZRRklZuY862T+BblEbLVnhfXugTBgMHIjyjv2I3zd6H5jKSkJ/scOL3vSoYKuWnemlS4cGf
eNmD1a7Yu+qADG3YdFL+f2lw0hzDs2unRjKUvMnWbY+f6OAtxjGVmtP7VLk7QGf9wmzvJ3WacKAI
pS5orfywL607O2Ukl4CqxPJRNZ/cjzBFW/lGxKPL5h/CKXsUnjKt5l8QgQtb5U6PUGP6g6vvxjlx
8TktJr6tWqjFe3QFHRGc7+OENqSzbxZ5jcQz7SyzRMHhLlX/+aDmmakNPIQE6io2m91VS6ygLGyo
SciQc+bc23zP+nb77RPOklVBecXCi1104xRGVvrKwBzFbK1trJTR7QpRhegIEIUjOYyXW+LwJyYb
m060GQ3W7dWoFndTAJII+boNuUXaqcgJ/NCmkaHgRSkVGb9ycX1jlVfswkycrTS4uof9CiJVkdKf
9eFvmWF2F9ds8CmLe0pW9tZ/Lj8LKBG8pECBqeRouie0b5kmj/E6URjaXWR0Wxvknzr9pMwwM7Dm
4Aszt1bB8lfRAeup+uJWDGldWJ6oOGH3Nt+gyVuPjKbgx540uAN0CIVVrovJ+gsY2YXDgUpSwEMN
+CuQpo9YAhlE+G6cSKleHMbCNQc7UC13ll3n2Td5MfsxWi2YgHsCh0P2fjEwOB6AG33LvOD0quST
4ZV2C7NHVjfzCrVAc1uOioOs02OtLOKBFITLAWHOzqlnB7zn7h4Nk6DvwpMisehts3cQRe7RlkGh
0XNF2HhKwiXiqMX0ZK8bJDvtDqxoxA4j5iB+pIApycGJyVONblaAMxztEXm7Croq4j/BBUTIiBBM
dOay40+lgD+SBACGrpH6s/TZGItic7rMCnl1eTViwhYJ+InOvVfipz5NgInIioP6DzX97GS2OdYi
N76391lXSgIOj+r7HlJRUpMwXup/VJ1SUp+g9feAHkxsHQUPjJ0O4ICaZ0HnA0BuTYTz9TTjwNRt
gLalp5GkLSFZXrQsjk74crGAt/L7UDiiKCa6bZut3vuoYCVkF9ssvcnn/DhU0QDSymSRYdOY8mRE
cnbrKatUf2BSaasswt/wj9bMARD/LPV8DI4SrRaAS2CundD+zI5GonK1LJhQZMj/0cURvmVkAxpX
/hfyLWxI4vFyDRuZ1zDFX3/AEnyQPK+F/e3lWUCGoxO0ayfPErQxZTReOQuWi6gdksfFnP3gvkBF
E0Hq+fyE/hVuZMqXx/zeBUGuBLN+X8mvF6vXuv3+gz2niOR+xI7RMEFk1J+i4JtKwF90Ro3fbJ9C
/w7V/xt3fwGsMVs5pFSbbmXBsp5LYZKi3BUCsk/7vOnMS/w6NWQeMOJpuuV7uUhvt08ODbQLCgCr
UYh0UmAhctbbw5q1TKuN4C5ZNWczunHmznp9emwC33rrLn8oCzlN4bUaMAAvYBkaD8H+1A0CV8mA
fhtCRytJ3/hnhpKnECBCg1bmo1NQSb6zo7owrKnr0YxYh8MfFmhtDWD1liJQoGgR1P5x/eTQihck
12yP2q8Hiuf8k/yTbMdfOHEgZdp0HudXRBKU2+YVaL/E5oVegmv2FgaelU9VsUekqVtgeB++wO8L
R7LA836T/Qlo9mXmoMGUeo/22BEsXF6355LOgMQKYIzltrSKFertF8fehV3cdKjp2kHqHwsUqGs9
au1OmFHHfqMHqv1ITw9v3l9RMCZDZdFnPtVcO9CAsOCxku80AKO+J3cJN4RkKEbU7QAKeE7pNqYg
H4gBkyBU4QsHgUESloIseUmNo33hdTuWlXFdeV4aaX83T4O9wvLMIwKag267MkKXQT6KYsDdPNGd
U1G19lM7568xXO8xltK/GXo3NIcR7oeWswq/vp8qcXpYJFEtTD2nndD7hVclPhcziLrQXhzU6hrp
CxAWlvXmxY43g4DzZ2sUqTg03C1dwj4ddR5E0lTiZOzEYUiQKLLItmvKWlu3QYUVqsLm/GMmWYEg
XcaHUXwozdcIGawxmI/Ttl4gNgMqFLUb1bA2f954ijWDdIHJqRdU78JtRGV9ssVN7u0hrPDhV/N+
3DKZvKWSonLY8RMReHwyjFdI9+jyz4zsZJ4ik4H5szgmtcMmHn7SdiRC6lxopbAflqe1PeM8Za+H
NitJNrsejpNUhVN7Xw3WAXRU10uhUGHyJVq4SfIYqFULNbXrPYmzZlW8Flz0Az+P0vZgrjKatHEj
2Kl9segwG+NrXopG0jt54/XFJQiHUqVDf/H1ei/La1aK7p4vp9b+4NYrpDqvuf5TkB7r87MdsoUz
daR/wBMFvd0DlfD74EpnFslm+npJ2+xMoJVT09SC2sNAmG+8J/hjSGxTloMR8I22Weti31jmxE7U
A8IbfDMdcay9LgOgyt513cI51vtZgrqYVREBLROdCasyiCMv3iOHHzx2u/GHDo1QBM8gOpA8pDpj
1CmbfzguRKN80HGx1ECz2gnBwauWlGx2KwtJIBa7yuaZZcF1WwUetv+x09DHWRbbzI9Tfm6Go90Q
AdhaIN9QvLzKcTyIgC/0Mr3otTcaayrCQntEb2kIesgX/H0rkegupk/r5xyXHQcM0npJgi9+78mS
s8DaKqVmlrgkHWHgf8m9JAlHAyrTvsqLvjnLy61ycoVUtVpoZaFVAxKNyjqCA0T4li3n9xLQFNjj
nqu+TeZmL/hDKWTjjSInE8ncmr/hLjwaTyuZjUTIZDD0eu9+PLoEPIee2EaBXllDW+Yw6TbIYP9f
Za7vc5fcyPd0la0hg/SKF7OvXQY6GGkM/no9RHlBeDE4pxgS1JfOcmorDkzgG3ouMbjh9i0IVh7b
snpeHarvmShEyUd/079l9pGOh4SzGKp+av63wibvG6u6uDGUVqNx94tnfs4r/alSxtQ6igXgdi0H
Dd6Jygx9Yc81LgMBedWwLHwhqZk+rXfZCvC5R+zqnGg36X8tuGoP3J685MA4EOkqlX9Uzgmhp/2O
W6AFjVuADCyvP5j/urdhdJ3pMrzlQAfJP3VkAW5/PgMHiskkO4c3I5J5h1qnmShc1IEd5uc/7yFt
kkqF88b5jVrJJjcN/7eYJJyaLn54FbX745ZDrwKP20V2nwcxiO4VoxC/7S6StxkKw6QGMcfiVjj8
V0vpYmor7h2aHuHlKyi48qtzB794ecHHEEMR9vaScIG3brWymtqgNbjY4N+lwJI08LRg5seKY4Yr
QtCiUOxxXT/ZUV0nk1yKO2dL/VphJeyEvD5XdQgyMNW6ze6vI/ckwYOQm3PZ+ALYdel52Ux82kL8
kb5WsQHq0qiTGe8xYKdGPsmpUnMPG1Sq8OS7MKsEA6cBAJy04O0DDJzZIp8CPiWLS6xuj/wACf1L
cuVhe+gjn48mFVSLeUWAPY6LbVoxusq/oF3hGdn/UNHE3ou6vPiPGgGW+kp8q3iTHL6U/Gt9Jt1r
I9lFzkQqDT34WTx0NAuQnu2wAvnKfGnk4Vyul0D/+4o1IQ8RhHiZ4uAcywBP9Wq+8DP+RvwoOOD5
lbUDrMpGcjcVZTtfKXLLfIRvw+RbYyweeL/TjEviuyAIJ42TFCBZAjvz2KjBmWc64iBA5U8V4M6X
vpJ9eUtW9yz5PUNyt3JgnhMBfmBjfDvx+8EGlau05/4ILGlsLeFOU2HV1W6sjsaVgnvIStgIKPgK
fVoN9vyg2Kfldx2gZRVEh/NdCUrOUYPdOngAk3EC5qT12iItnxI4MiyhGfc7AvbhbXLtVdti9Hxu
rk/CmQ9fC6CY9UPJwKKtMF2iLjPX4kZp5f78kQe9GaJlnIHaLiq6x/LMiNdiOCz9vMYEXhNwG61q
h0ulyjGqzS/eRfI8riRKy7h8z7jCZCdp2bh7/XSgzLX6p3nPGC+N+dLji3vZ60jB53UjaX55ZMEX
zyv7lwwhl7/GUR0YfDzv78H8v1DvFRRbzkj90IN/cubMSYptXg7M9eneAKsRBfzPpTdueyQfapVI
rkrosq1P4QchiIsEU4RYW4lrj05VsQOQT5qiQHJyx4wCbNq3G64zCxrHYmf73mfBSjbcz1JR/rvi
Af1yyPDjqcyAdt3M2Vu4Sne/cGW+kKoJSpaf3+V5y247O3fvBg/u3Ms7g7ZAa/3O3yHHv16DaBBY
98aGXP/f4u0kzgYE2TE4HAMEONpqASDhfxUMfmKbP/3hJdkxMU9cv5LBQwwOfm7xyu1wn1ieDroc
ib4GQz8h0EQkrlBviSN8RIwT3mG1x7/n/nwC0btrhAG0GU50ce9EMbQOxaX7X4DjikVjmwwIoHu9
R0SqOvkIvHxMdLKEQPu0ZlOA9gKcEtBS3YJ5GnIwgagwgg27Q9GKRqakkw//sTfQBGtbUP/h6ZUW
/tBRh38NP25hx4X+jWmiraksMGqUzxvDp8ThAQilM3ebCXWSWJcus3UK1Kf1yUpkLNPEJVemEEcE
GrKWNJU7jKyAbWtEvQaqrVa/ZrCjnIGvsCT1OIcO/8dkJodNXEAg8EYAzJp7PTUZoAZRxTv8CfIc
gjrLwwmsr/ZMmHZvm1XBIEKV4K0kGhm4zgqRWT7p9N6wWr8Cf42nRcZsAl8XqQ6YFtJeHG5gwz1g
JDEiTAxY0LUGMMDKCErLPHGGvZSnfgfxWB4ela/eUOLeecj6zIt/8uVFJT+wolSQXVK/4XkxA0WO
pzWGCnm/0F+00pVrZkQkkemQUKaApiFpN99jh/7BDYyOu4vl33wDsXPhR+RoLMrItYwIEnShbE08
0twzYnzIYGR/vQpS4BeKiYvknNOJdsHQ2dsi29RTea3NpvkjN8qiKebWnIdwIFcnStq1D8av8aA0
zQ7lSsyNUaSJ1VMAkLeCh5RWzXrF2Ies8LIaNshoEWOhU90SatXLmIKUlCdf7NXXuQh5HVSe1nX9
ajmSW5tTuT+mFQNUgI/wE+GO13LQc+2sxmvgJ+4J2AJVUUJ9tHQ+LpTgl6e8fjKly5KAHhmGZmmu
PJ4ik6lWOua6u9nFRTz5/CAJ/qqsWUF1BWlgG4ZgwduD0Jkv3lmHfbA8jz/iGapwBdtUFduQU1CC
GhXya1oigYquB593Q14VlLmAj+SfurEXrzspxkVUKCPV+SzKVZEIK7snSZBIi7CKwAH00WQIkFV5
YxWXgmNmKc2krW9z5FCj5zDfwpJVjXcAqYtmeCvapDui3gK8NW73qGuoavBxF9a+Hj85I5u+C7F3
8nQ7k7IbFI3IruZyCA1SkRGcR2aLqtzPZ1DUXyOT34oYWfe75o3HmY4Tn5bCCk7TLU9NnaFKqogS
pYml5m/iiwdANL5kK80wRFEdsBe+WWvNosRO9cbndQGO/z9yGv0Y4BzrA8hLgYVNDtzmZ6Xp4Rlh
knhMTkSiYuPUpnsYWX92ZSOK6bXAXKYaI5DMFcw72va5xWZbULiyuXh07IV+jgdyl2/HQFnRtnx8
99XJY0qCK5S9oxXI5bw/i1Ed6WiyTO0K+JOHt19RjyVH7KtxdabyhnNVUptqLnGfTdVZ7pYx9rtO
TTT0LMg3pV4MkKraF1RSj0J/CJmlBEadmFAP1o/z2Fv10Z3Fpu3KmOh6N6RfTRcNP1o7YaSs7YSG
gW11XN7YwyTpymYBiE2NMMqdRKBrU5SgH5BORtNCN6tkQCnpJr1I+YjIYsSm7TwceIDiW6rrWQKu
8yBHYBUNAT/M6/Vs467SKGUhszkOPCRZF0wjjJy3poartng/qZquXn8PMK3U8U2MmkDyuMD+5izG
dhVxTmZrW/D7mXcP/RdXzC9dLmQov1cH66uw7rXvkwZOkLpP0cIfKnP1/6adU1VU3V++brBBUfZR
cX3Kv17Ef5Z6NbMCVFl+4DTjvgAj+Qd+6mEl9TU1eOnxJKYAyexp2Uv0A5YI4XuJaSYqI50stBJW
DHktQKkuVmvUAfLxTgibEolqsGw5kyb3KC+qX/xd6QZ8938z/P271Ih6MTqZ7a9VhCE+Fw4DGMHa
1ChSlRZeyQOJuvdyQGmg3vdvgUBZMFhuyf9jVU/5uNbqojQyoUw3oKmaz6uuN8cV2CGNK1QW9Tua
ikpasDlyLKjdYZLzDyLrPuL8p+QL2OcQ5AzzmPmM/EKhobG1BorDsWTsTC1c2uvKAI/TEpuvO1Tv
o2fEGDm+rlfsYQKZMt4NYLbzzP657oKG0LBqx1/wvJlPyzGk95yVJbIJo3UoYN+s2C6r3HDbaTK8
apmJw0ChU0YanjnfXmQym7rwN+Qvbmquhk9nz2HksLkaGPISyHADn/jC8wW2rwufk2R+SzWtFDJE
n2FgjL23/c7skrGfiUJBNDipvd2okbTsXo4FVxpY/aYzMQziF2JICQDNnib8hJEnIQHwPFhrEZNK
uHAIkOrG/pWquORpgBQOSW94oz/c966iMky/TlwZ+bkoY6JiZFDA7wTH424RdPoxnkmZ8QvEhZqd
93mxceXsIqmqb/2x5o7DWJj0/YVz5x93LY+EfVNf3mi7GzXj7mUlugLpsafTh/NfBwu6xLM+Puso
Tes3RqnZ4umdHHC/ND6BQ00QA3lWEm0al2A+FX9oWSaLbrVNkLNzJWtm/WPhG/v+SmuwLf/jUzAd
LJxEKqiOcErnc1SQKunJFw9wnyCiKzdkl/hZUyIRWwkjsPCGEIwVBf4fSJ+JU3NljBIj7J0iwDeu
ceRGEx9O+tSx3MadoZ9lVRJJLrLwn9TECUq7EDz/r0SScRxAFUHjrcw7+wzEM9wUMk7JrR8VZXsP
65OYzMsIT25pkgduYQiboh4GqZF1AHjCxv1SCGyWjMaYKDiNEH+Rh7mN+7tQ2LXnGswj6077+/bZ
oj4Y9Xm0GDDAnL2YsG554uhWW6K+7prv9q9/zvD/PPOQW08SRVqYkGJIrhQp1unf+ldXMtXTs6sI
XKEKa9OnUWFSFGkxU3SGDVAflrlcVeNfQUolJ8w8pWx2FvaPy0+28IFAFOmwYchY4shOXdqzWHmF
pIZGRsoZk/6aHE1PUNA8n63Jc1ovUgI+XndGrUU2S55CN2Na9kyxwxrf1L/mT1tjrTmvZjSySejp
zRCnc2c+hl498OWs/mkdUUN7ef8BY9PE4J+4iSaCBmGIoz37cGbtfJy4OYEDrNaw+HyVdNBy7UHf
be2JCGuzoSrAVNBAVua3WPWdqvhPFJMeE+JIa7aUWRrNu6VjDdAcwPWTFzBTzh7bE79dHq6YDfYJ
+o/iOkdrEd6z3Qq1b67lsFhwAvAOEeAuMFVy4PTFFGedUEL6NjHjgdqHxxL+QAlgsuyogpa2T25P
CSfKU5mjBw9vByPLP5slUm95ZNnc0ztSEhipWRwOXRriYIAsjO+insfhfrESi7zYiwVNhsNzZH3A
Q9LNX49rzj1sCzUgJlil+HXc6ldqeFHwcxdaOIZEK7Q92Koz4eB9SsR4zlh5pouUH6Jeab1HB21D
DEZhGVIJzMYf60VEQgM2O8W3gpGZtaBiQMHH8vm+cHhlgJ+MCH7C+sp3LLz5o0hmuukL7J1/P/qS
cvy+JwSqijeWONmKYQTwcK0T7YtwhGa5jxhz8gi7cBl5asqsUuDsAM4GpChQ1t5pBfBKT8i7A5D9
xOK+LoAA9jWWXtHHFQuYU0M3ESBfc9zdMEQQwRbrL5kauwZ/XZmYReGiuFxqjCWSpzJGM8iLHfaF
DGlZBkG3TEly2FzUBqJ4sbje+6CrMWodJ/5KwSTGgLTjyeJ4XXpbXGNK47+ldjgXr5k9x5l0wZ4t
wSIYNN3sEc/mopnIy0z6+YOCWKUC7R/immpdr46DaapsThrRaM1yIWD66347WcoarVlxbbTYoWrc
wIMCqfzngSfYhzvAq33vkqbuY1M+ZvJNv2R+M5GpTRYwooVao2cuK1huNOPdsbQwu9YPZcUAjeFc
+TDFchgtvLJr61UXbPjp8sFg2dMlusz0Cdo8Lmt+ipjbxS8h1zbpKsp03upP/efS4QfDdlV8a9wG
7wEaz+YERIsLBiJEbwtvftx2eq6bWoXOqUryvHljeFSpY5p+pHwW8oz+fU3iIwQWJhnrdPfFLdI4
QiNLU02c49hOfJndvh46N2sysv1vRKS9UHI3Nh8Z9Z1uZ0O/yceGaO1sj1RMq8vf/OT2fEyj9OdR
6i80FgE8jCkUNrzR9W4ggS27A1OQ8bxpLb72TMnh+25LphkoB3UhbIp5C32Dt8hDrV+73Pfk1Vsw
lZdrwsgCcY11NqEQmQ5BYJ7P/ZFWuNKZb+HG4PDRXTuH0CNDUQ2+OB41mkRRR0zfGmOdLpSUH04S
wiqy3yhZSdZ8vz3w9RpaplGNa3P6tYr8pb6zGIQArclOqetZqW1zyS9E0v5LCXAR0Be8mta7zc9K
xRcx4bNy0miwOF/xCjZhqNl1JVXuQTlVfUijOfcB0nkbpgy3rzshG7reUDlWrLwwW65VCwbc2mTl
nOpoXffqf7v6l3gPAnZSYLnSl6p6no+uaXCyh5n8aX5Z/SXLmz6FsSt8EpMrKbiwvEK61hUNRlpe
R+S0mljcyj7zq82wsmAHCJb5n7oQgMTJsCUlXo4UMYDV+Auq7W2B2joulkdyOBowb8T97eYSBeCR
Trul6w+vBYn+oW0jcSvNJDI3322KCQP6QXP26wk1KXhjeGqLDFcqy7KkCAuFmI/Woa9ExG+L7ekg
Xq7v3PS6Cr1a8EJ4ZBUAwMJTYZMwkSfETjRujfl6kMwKmLGtTYEAi/MWTOj3xAAq++atqee/qXyB
UF3Klr4JlYNc7ORQDnivppuuQfmXpqi3aJ7yKuNdCItt3RI880q9rodO5pxD99j/2r1EH9VgDPWE
98QIIU7L24aIJJ0nqu0s1KZK5M0doTYW/CPd+TbcvkSNLvfV4aVeAawuMZ0z22kxE/YOH3kOcVb+
1gIenSZLqZ8cNacxIAvoEJz8NUYTjIs8NXZlFKXpO4blv6DSlCaSrhTzpp2qMvdeuPzgLVkq6KUr
v3r1r7/Z0RIABlqfDb/AwukLYGqw5iz8ELNH9F+AbhMhgkWu03QYvIGp5Ouqbs1ld7vQbfvAhQ7D
fzFRQkjprf2ryxtDcVchY/PqFfrSF5co0/a6imoHFOCtiXoZHDBWno0gCIuLxHk3WThMhNwYSHTG
ZlRKLve7BAe/LcnmSeTBTKx+wsLNazfLGHrH52icuyEv/gcQksYYxqkVOS//AL2eb1jumvvNEo9f
0oIRQfS37AQhBQXW2FVff81TCsd5OsUrkM8gEy+sL0MBxc3LIk7/aUgb4LqsRpZyDQKZQ1VxhwiM
7pJb9L9A6D2bdpvNzeMgINbI7tkBBNPbrG3ZXSkUsZHV7FaGXdHzwwnzsrTB5ZZcihY7v0mJGyMd
aWoC7icF8gZxAQ79TMRPc4EDVxP3/eHRaEHMIfmtdmZ3RG8CSzHsbunDqJV2Aec01ybnq4qf0C3f
7Vftjzc0SyawCNFmH7ctpKaqyyovGl3LQ3DEvp9o5L1hswLWrGLVVCE4eVYFKP2x/YUxvUSjUF9d
hSIUMaQ2ZysCo0ooNfNTvGIM910QV9RTIDENZoUvb22pDBd5DaYN6eTz1oll3OTHi+J/vvg7EFjp
q1kiiUREFKkaRB2Vq61wvkg52sBM2dgzhLR4fgv5neYbi7046LN0w75UAuDqyg4Q7/jtWqF9B/VY
CTOnWdrzeoG6r/MLjrD0aSP706aKTYTmDBfNDV7E2+4qWOj2839J5XnVL+E8yGulhzVe6Wp6X3kJ
Rn3aEDl6O+Cht+le3+xD7VL3TCeYdUhlhBezPZHp927QRleuNZ57StrwRMoBV6Wi51OlTKDa7X9v
L+k0UY7Q3R7+5mEKaVZKqUU+FieuXYrKG35IYCPVtZOLGvqAQBuc7u1eU9q07IzBi5pq5u83kGhl
UwwdgjmNqLNuxY5C8LNxRHjtEDuuczdxAlHb+fkBkJEe1B5xdTE3XWyENnfNdVngL72X76CfzIVv
vuZEuovPBNgtzdcMJDA1BrL0mANvByQB6/CKcx49hb58010BEoKoX1wIdk07sb1CaV+23H/3wSzy
lV4Qoz9XzkO/MeJpFSOQituO2QuHyvvPjXdanAvaQIsAkrQQXmsdnFkgS3G1bct1TtcfctpoIgKF
ht9Kj4BkLqY1Y1wRxRrz/Yu0WzUE0NaPlgL8LIoHoojC47KsFVVVH7zmwGVOFOhND36hOYdvu5eq
RiiFSHgMwKgM0bPBpkK738aPW2qPDcf6R/LBFgFdCq5H31ZuGcI9OWsQpD5xix+Ah7Q6HCSA5YBZ
5ZP9Xf0ovoW16pm72Ehpypm2L8TqGRdTZkoFAWEEhoCnSPulENTb1WXePiDjSXP/XB055x+5DSBL
n///kvWC1r9PeNrBgh3sqEoiOBek8zNOi3EJr5p7My8/00a8+OfQrQRW6jWOkn/fzyaACXOczdAt
fvsd5uTJdOZGa066/zIOt7piKgMI3cG9/A6t3q4y2DGQgMdCgjAlE3AAcxGdzvB91h2BJjjFIDz7
lKWS2cOWygvcnjVow924+3GFLyVj2WVm0XM+PLOM/+sc4DTxJ/uA0hEpzSz6JYr1jC2DrHIuRoKI
OCtBtCIYKFoTW5GyXrlLmKWGFsIRdhCIHc08yo+afP6irvYRU1AFlVDIsk5w2hR0hXLmh8HCS/cq
QIpQReB9sWJZzzrcNrLFV+VcCWWyz64s+b9QW5ZqCsPBrIM2JBdeQseHhK8z8s6WwYD5+YaeFGDi
lwOfH/OqgRkKOLAP27IHouSK+2V3j10tq5iWgQFE1JUsz2ZPZ/Rplm+NyVV4CYfi5I3WHse+Q9bg
xb+O6dU4MsrG3HFQ5NwMaGsmrxxd+q+du+4TtpDAmSIUt5OP1N4zyiC14Kbo2cWCLOzmq9i6IozU
Onha0t8CosqsgQMdNiwBnDHT/bi/knFCzV1KT3nYKlcESyUDj7y6JjKUEx9dfm68uxXkApj/I8Zf
PVIJjdSH+djeCpxx8u9g295BH64gn5LyO41A8RjC/xTMAvAjaYtCbaQVurz6jZo/artdLRREsar7
k+LFkxZWmnRRGOKkWZLe3m0F2WaoemkKRVmUXbiQoFmBf6vTJV5p7PaJjsNPJHRps4blnM5F3Nrr
gmwX1hTc7ym9s+Zwj7F02AO9jLsebEVwSdTyRCkjMKQKJ6qaN1avOKdXuvhjCHVAyi3L85pIZ/rt
93NHbxzXGq4g7QWl9QStbHJcrVqVDmHYAvaqM8wvNE5GjOScRQvSqa02RXrLrZTRMEsdBFvKfD9d
dVyjUBM9WmRx92tcjr8bLfzPTUu49tg/7XtEg4BsDhHD8NVYvXcwD6CIngHp6XBIGtM5wIGgzF4a
ePKscG/wIgLCJB3qnk2Vpf62eWJnvsKvu7otRXY+PTXuHq6+MfO5QNQF8I5sYy1j1I/oWxd7OlUw
3GWRDNZZ0ammiE7d3Xs2/dxiUh7Ibzx5miEe0wAxxNpnMC5ZTo1Q7gHF+2IVbxgqpen9YBQlMgW5
r07YsYNRukoFeGm3Nnz1WNN6IMipDX51nDNBDYDv9s8dLUfUzuTfqB65k8KO+GioPT7ZCn88orLs
2j6t1egbWCZLXzDb6bRmH6k0BzWjweCPnc8Zyi4HfV8bQAOBZymI5JvjudcRzW492EYitNWFP7x0
qtn1YghP2thA2tm0SlkRwT7Z0bLq9q/u8JgUNxudIl1516D2l08vF98O3WVkIuDt9kxepW1opYcD
C+pXDjmypLhAKLmL8wF9RBXpGSjza5yAAh9HNc+PmMUVRttYoVBEsUnN4lec5MsV9kH/FMUezlAf
coLc5RlVawfj8RNgien9hpmrSa60hE4hZXLfZWFB2IxV2aBU9DE584JI88Ze5scLqQnxHT0rrH+m
MJ16t0sbikITaL6vaKPxXSpZxT2kfQ5tlae9kt//s62KPXLGgCqBhhiMtEQ2na85cY08YxOgMkpb
DnMfN/nKqh07DNBqnxSnZYbt9hQCMZXH/ctq3UImnDlLUojEFdJqPC6/rBOaZhWsEjTe7xXSXC0+
zl1sigyjss7DRbIXbCA/V9i1i3i5QLBX+Y5dpkYzNQn5kKc9+hKPqXhwGwORlKW+qYrMAjJ5K18l
9w0owqBNU5xWpjAzRich4SjqUu3w+hs3EuOKSBgqjvqxrvRvhNCHprcZiJgXIUitj2OC1RS1HLm2
oFMpmyC5W5T0moCYykWUwA6qelOBRU4cGE4TJh0bBQGvBrcfB5wuDoS6JftlgByYmYDpOhtZDjkL
1md8A2u2RNuxn+k9CPjbuz7CVeDXzt550qMJbWK7gobXFV7zxHK95tl4h98VMot/aoXmFd913/sG
h0b6n2+oyJi3DRlPIzxRte6c6wT6IThvRStKzEwPaBRt+A6zyXdYIUU551RacPhVgAGzpdvWDfmB
FVvfO80gbrZ4MBjwRKo4pN4IwV2PhuN+KNorCvzRsTUTaDrmtd2/v39PGEFIZUTajHrTDFEeYKN1
DEz6npfwCOl+NUwdG8fudjV2qZfMo2owGlg0SenMOFrDglEvydm777PbZnd3U/sh9+/U0Gb7SerV
GV3Dw0bIAdMw50rVcK430SHo/nic1cW7VG3c5iv2gXhv0G+sl3Rg4AXkuba8Gfmya3nS0YTPDbGG
yUsJOXNnyDVJfg6T2Y+dZMEqe5kqUZK1Nud7DBdlvSz3RZfoaQDmCuEg1rwAo1gLta2VHEjsFVSD
DuaUTi9ECSwb7HXXk+y8Vtlv+U0OFkvNmf730YT2+9xwq3i/jg3FYPPvKkSLrE1I3ZzDjrPd8C1U
h2sXvojjZHLZrTCSR//7Abe34pztvZ95Yk2GCLy8scxbckOqeXn/jPzSbWFtYrO0KQm2EGGWIuxp
ZsGzHdEfCrna9u8HC8Xf5GFmf5oVeVfmw8suNfbgz+IEjT3U5Zy6mdf96a39Jz3m9nqBLkIK69Yr
cs1UNhCFWGFDtd4kUVjNl41lVqUXLQ+9pO+77wIHKSPTTcB6AYkhmtlTMwc5CMuvNenMTwawUpTY
ONIB9ssXXQs0Gx/4enE6Ttuqr5airy12OftUB9r3syFkrCwEmL4B4Wbr+VPwpdWPq9Ud+vPOxCnZ
yimrmaj3XwB7FLuFtEG3i1iITRFPn6udZIU+iI5HNYX227yUi7akL+LKopNYSW+f0kv2HyqF5dsk
15YtAeKca5gTsq625HKB5ViRp1XvKHFuIQ1FUz1/Ep9GM9jZi/fYzXt8h8b5itLacgPZ+58QsR67
aUsnxi7hgJTVskoRqEIs6HIfk292CzTKZYLAoQntTPHEl80LB/U/z9gFGXtDIsnqnf2Ke1obyXad
byBqBxe8G+OdNN4MIERtur2bRyyqh+X8GnmxRioLn98c91473hLd1gW7kkmdavtaqGRkq/Pt1sv5
VR3uyV7SQN5bc+V46vc//lbIDKcrnafy3sc92DwaKxmvglpYZdngofL7Gvp6U4Xz4FLEyqvPmDUC
uqD3Y/ucnxuMXg/196Hq1JiEu6DvdrwE8VDIMJ5xL5/XjsHyMZzZ0zUjfjVVlLXbmsPyGL/zO2rq
f8bXe4DqwRv1tSR6evQrUY0KNrNGNfpIEJtTnfSbCLfmUqbAl9ECGoFDpZuExXDzA18EomN2VQn6
3IY8Bpu6oTETjoCrxdWEwGnZfrY2kBtCcre0H1ErP3OBqRfiJaWNULcJ4oPgp3VItDO8pwzWTzxH
bAScdfg22ne4+ipptN7Uuxz3Q01lK+giiC9bwraE5ZiFfLU6GurPe8XP4rSatSADF7qne58X6ZOf
RVttTuaQ1s184uMQO/7M958z7Aa8Zr7zRjUe9jOr9VSXlQFWyFL7/W93MbxTu0vAZwabS5/DPH//
sit+ufsMs9q5vMfkSNQKYkpq7tln7/OFo2gmCR0us4Vq/D+t1nvJ443m5aQumYKnbMrqSwSwoI2l
OHyOrteb1kzroFIMyzRZrhXmiWIGH9frHZYbZjqp7P7EOzMXsKs6xX6HW6Ol0YNxNQM2lrVpfn9B
mAVPc055p1s9TXH/Dz/lcunX5f5W/yJXncVA2P869d7KVIeT/7R8gZLzKcbN6diXZCloSI3FWHJK
0vBFGsO4piYmL1yEaZImHyrOyW9U2o0FHlW5wKmLsl9SjctOKeFzhvEwSCKpsO/rnVBwQiIsWjI7
LiuhLO+Kbq51ENcTvZNifm/qRcklhc/kY7Fp6GbggyyYb38i0gr3np4ERx8ZkPyQuqIxgfhMQd2C
/Hi3Pku1vr13vmTLgztXjgoQRkZHEo5hcuRxmbPceJXSqtVGcaCg/mKw1x6CWwWsgTgf237phkGz
szFZcpDJ8qzlvwkuEThXXeZbclOu8pc7AvKW2vfZydglYZJVmaGtZVsC3H3eVfadJr1D7yBjbfZA
r5/7oeLdINi5jxdje7itDcvFY63dl6Qi4JzeCN7MACf+gMQkeT0Y5gJtaWANMqsQdNLA4jAdzKPI
/yD0t7KkgSQHAwt8ZwCARiyxYcMnaA3o8fJJo4YVVUA3Q6in0x2SkuHoY0btnCXUJZ8YgjlyMayL
5Ie33r7AMid6hznX8FVhS19jruKSO1j46B820fpoF1VMYJTQdjws6pyhygb/U1wakyjtx62SfaZU
5IhxxypxRilwHClgPqS+bO4HytHmTyXe8T1dJfRZAuh3eKkbWvSKAqRhso3dN1zgnmSkDgzNVcIb
PPRWcUksJ2HBoJ4YBzVxqqkG9SQ7o8Ce5qkG9qhtjYLbCJd8rmPQqjTBhe1qw2ef9j8wUWqqolCV
P+KCJpcBz3qIGMhQn0b98WbTDbss/0z0xaG11EOZUTkqCCnHfHu7SFUoqsVoiIGTxx3um7s+RKoX
LqOVUFrYslcJn21kFjRuzndwJkxIQ3Fp7kxnQv78GCQENZr7uTVc6iA+K6hIjo/9dc8p4ezbrNUb
VA7yMerVSSUIidDRfrlbb0/CKPgR7JRNCwSKeF4EOtQ1znELfamRSQFMK8xxcsPhf2wmYStxqPy3
tXWDAqe7nZ+FSCt6XUJt8SkIV4CdivJCkCV22ULXtsKffTvKeRSaClBSC0DmRrYWygIiYG8fpehb
glFteCA3vnXJQyjYnbv+whjhzUaQ3qkhBe1bmcyj9J0hDFANEOJpC9vx9xn0oc/sC2X9gNH3538N
xX1RigIpUek06Vlp2wjma3cnS41XiMgGGxsTxR4PTW29ac9vDp5aDOiHtlZCt6aq/L3YPMIWEdhW
/xgXXgK8BqykkTa8Bb2uydg+V2OIuBSLJ15uyMnAkHSZ13XyPq12Uha4EsDT//OOcmFBNSWGkd6c
MAK4wv7sI8HNiLA7YcmM6G7YZyVIgPK67kNX69fuRKDwe2jRZJO/7ke9j/N2gu+3oGPy63zN52y9
9fu+gAJhPqkXHoNqaWEvBulEB9xm39HBrJXNo8Dqv5FxfHvuvEpEIpaL/GIwLdVlfFkRybdH8cWw
hhlNRYYZcdbzhyxnWpVCk2YHsg68Zgzs9n2IoorNaVJaDBkc+nA5IZ1qDd4pl8D9/gOi1hJkQHPx
lNbOq2VedDd4zvfn3nVe4U5Q6fmsRmJG9WkWpiNYrNkn7Bq4NGJOvyt5FRm0LJmXfF24umyQXitf
qF2WOncj2wEwHSL5mVill322yew//pxY/m0xEnuNW4eT5WaymvwJR29iaMFu6n6M2VwdUetmHGsO
ZmmGLh8gm4Xxo1vn1oQHI8l6y/ah3A6P72Wtkg5Ho6ktwMiuqibcxQhAy+Nd9lniyhTK3joRusgA
SlvYPnvzif/5gXPTu4KE+KtMMYiJZ1pGqbPBJ4omaEjDsrVUMWP5D5LCvwwE8q+cd9T0pQ/zD9a2
+dKWn6FWZ46gLNe7KjrsbQaZAEPjHFxpkfsFZ880XJlxrEDzGvkTE2DXkkBQREFS1HVQV6OBl8bj
BS4TJc7H/I2t4wUW29OEzoZPvl7TAm4SoPDXtNjxsUUMzZO8Zny1p8SGVPpzIjPvNyqCNzDz9AtS
sWrWwbKIGvyW41Uh5T0Jf1McCccM6iO/3Dx/+ncxQf+EJQujxbajREYj9guzIXxtySbntBsgdMgD
qdUWH+3SfE91MO7t6huW/f4I28rKidS1i1uEFEI6RF7T/avoom89ORxirEdvTzRM0DlcIna49I6Y
5mkGPlxxZONdnRJ4EgBf6SrCskjQZudgu5aZTrTp55gpL2ZiKQpclKWfLci+BCOJG3jJ3pRaubGh
i3yrD0Pt0RgJCbq1T4ipSbTGLeJYYa10QudpbK0kJRnaUD7DXqIum3XiGgzRnuTHPNlmB1/NFc2r
Rm4lxqsFI/kbyl/iQoIcqjrNDAciSNlPFuEKwfljMFhaXyhY2QqhrE+/NtN7EbY0CtcZ/ZXqPPhF
TKV5+MDim+UbU7NIS/wuyWgaTswesB0HbtcDsSWWhEKOEj+zYhYxJLXHWj72Te98RPxH68SnQrUQ
VvE3LLQ4VJjY9E3rnzK6bn+TuP2mYj9QOhkGTBfZmmvXDPATHf5kWQX/PHSR1dC7v24Yi925ZGUJ
GprJ/cDbOlSLoPlBsB5GF9SzVmbtICd2iNsDXgMBeREXsTTlYfD0edbPlVVykaYaEzO032Pk0As3
/Z07PcgmLRAFTH38/dVNO8oBVDdCb6sBTdgdCNUiK74KBeughfaGgC4OC0Kxp2fKsQ78xYzlrrbx
Xdqw9H6l+Vq46R02Sd39ueP4BWrMU9jarC67WYQIevh10VA7HoS6XF7thAnfDKFBSwkK/+y7hXqd
gvq+jPfeiYRVlmh7yU52PcfYeeJWelOw2Ox+GDPgbYI569yPT8cWF3ncAN87rTyU+zSwZayLCNES
UMHHK+edu7FKwkMDJrLsppjQEwkp4yAOYGCf0TymhWQiRiJoYGV30RJFhhvh2G8DDnnn6DVL0wd1
D4JZAuk20wchgGcyh7hm7NLDhKEjsfTCJtwpnrKhRT447pmTEt4k++omTbIO8jflbHgRThJ+DidR
T3f689g6YwykAMbFhYxDY8iaJNB+VRY+EQwjxIHS5CXW/rWuDCP/peIyubVqOIk5SkARaJwd/Byl
XtgMmfifhbz5dm8qw0rbX5Cc4JGqPm2IMU2D1lAldAkD8TRdwru62xUWYqArAyHpI/560YWg10G0
WCwEyogA5DGIiTdqnqBgiE0adzXFkPrsgvOEmKh6POIfUq12Z6eW8wIYk4QH1TLDlvnbNwllyybJ
CoQe5AqgW1IYvEiaLU5HQ9v60ZgfvIu33LURvHL1xL3ws0Q/IFNMp4zqexXTB4lwYsWnlXEEyQCN
jxH7sehzZ9vDRIi609V0eEKUqwklYmInpiAn4KYk3tXEA+TCSvkCGooe8HkqMZSgF39dyfKFf/dk
pAvW2xrUWx5V5IN+Q0sTd+R/cV8nAcPncmyKjTcxaDd9L25rZfkNBCTTFfDAZ3HXoNDnVLlds51w
5UxeCE95ylrXj7ee8swkHNnrxm0axmWq5x6bK8XmXzHcAUbgrGpNogIzZN2hgSbNUQtUpxt7W3++
xCoQhtLF/pNUkAQ1OgxKd7vIez8wJQwuNnt1HK4UiQFsmNRdWWNDhh8Cmo+pnbIKhS1h92esQW5L
BUEIm26+Z/QX0DAtu/sdpMRK1yQzy6sjGXBK7FD/iknO1Ml3r+Zn2u292V7BnHO+xz6++G0TuLXe
y89lFQ44/puzka/PMJwGUM3CSVzaMfARqkV36rxJOt5WXwtyTI8+1hukF8CS8FmrvYcZQq7yp1RJ
kErFzBVwGlviMBHeMl3p7sc9QAQlY9TX1IPIVkgCRcmebCjGpKiFd6j9Bm1yHOOq3ucGxQ3nyNxl
io0LHNCxHHx3KXeyeuarlbJ0zaIOdsqlpFvrHgv/KqhSb+hwK6Mmq4j9x9v2XTYpYSWNL9qdbdcX
xl5TsHddWzCfOwmN6gBLjUQG4OUEe3Y693qbIRA1YUR1h8Go3N6EdA4b/an1cc3a125Bmx4RgMy9
pYftcRULMr569/eQuVaqnkUilgHdcVGFsCra9HUVf6LAYxrKzS2MXHDQI598yi2XeYNqpULw9BUk
zcr117XQIDv7WSlbvWVbzyeHspSA+3SUuFe8q9WTuUqhi6SFMaJ95ti7qd/HdSPNB2++bjf69OxH
6d6/Qptz63tnLgGJaq+XSzCihULjg/xUJiA8MZbAkjFGd1tezP0aax/KB7YI/EHDOOiimNSqLmqE
mYo/w1YQFcHHYjU0VOI9wAuOrBSCkxc5JiY6zutjx9sZN+KwtIHCBor+uJgglaxwkmWowuSTPKfJ
v23Vv/wf+mqtvxa1e0n7bmEWE/TOGJSSh7sV7jwlMClWoq6CFjvboy0iKQ0Z0IVE3TLEF1bCMTd8
OUGt4MizXHoRVtv2m+0yaghhmEbeY/VGTJcBDXKzXqHKf11r+5yq7t/BmxEOPqOg9Gpa0K+Xbyeg
95WMR0ZMnCNIc4+g9sb+tzWXIRXmZrT2VfqGitSdvm990oMdzCrbzEA9W8zasMhWPiFiyoE+FtGE
20UYPkDcyGJQ5ergG4f4YSAUabQ+9ScKMj8yyIrauDgRYWVwRfbOKMyU1UbmhevIsUDt5ux3POhy
IikgwSYBqUD4zTZOoXv/ssnOiBjLNkoNb/znDkiBxhvYYI7PKOcMUAj4aMN6I4KUU8OlOCzJT45q
0F+7QwiDaqjrqp4FFfRAWq4T9lb+FUChZD2LHGy6KFhY6E1pf0P9KaXdaF1+Sph4SJbjG8KCtEVa
OS2XgoE/zKV9LO1oMYMzdmpReQeIa7ZJGYHc75ziN9n5HvFuLPw17NgDPINw6pGMEsR3teaIOtb4
cXiKpjKOOnYiNiAvO5Kqx2g/lEXtlwCnr7VS7C+rxhES6M9/JGXRhAa+z3vh8AC+lEhE1razakpt
3J3sUXspU3BWjSza1zN01+sF1kY6lXjuEMrcw5Mg0zeEtT3bmlwV9vSb97QmZEtym3/9pOZVtX6H
xh4JgMwaS8i1rtM3fd7dl6zVvImv9SdqcJi4zld3gJ3iURRxrsABNFHH2DfUhf6n96+QcQi0RNDP
hq3HInad4bn/OOxxSpnepREKXlOF2EYTkcceItqGEPAZDGTxVSSuVVK8uo82HQqPOiOsd+HhZ8M+
aRqY2mcnv2Z5WGWcLgTReNSU6JB0rcJ/CP1iUxxBI/jGbZMCxn46oGzjJzg35wAO59/RCng58MyD
ShvGrMpOeDkBAWxZp8/r3B8q9IPLqtwNGWk15RL1/xaqcTJzTOhss5Tg4MJsQ2PfTlKcLIvq98IO
lQcYeBulcQgIy+UZBoaVQkMPQOoWn/f9z7v/WmtgVxfmYegELLNpkSGUZSIi4rIeNmZvkw971TBl
UDtNBx7BcEbB48iU9G+DVHFQSmFvklcIbaXfjUxoimHmZNxSPneRDY0zGDtPQuiF8xqqINUkEYS9
a7M0fEkjaZe8wks2pJj5w5sOXoq4GKvE0C6R/q3ttZqyLlCpFe5NPyTGYhO6ZgDTg1I76Da+YnZI
zmsescvU9TwhFGSs2N6UIHqWVShHB12vDm4xZpSzB1aM/yBx8w73EpCdcx0io6TNkuX17/fqzeIM
G3zz65jkJeRuNE+BdopfOjZ09g6TND8gDc36Cgdxwj3M+Q9A3macTRJ6NwBDPLovvO2a42aWmyv1
CzopMPoo2gJiyfDwFTjAmLvubARAGn4S+6bFxU0OWmxdZeTkpb6cyz3FpYN7LUp5QlJzwX73cmDM
yaF+tBjFfhV0RrDJS1srkRknNl9/gHz4RH3xwDD8flbmQ0eDxAOXmE0EtlB84n8eczJs7W438XG2
SRsQVg7It6+pfEI6RFaxyYIAzVvgBhBlmjPgze0YcYNqx4/FZBR2ndJir1lCsm9/Rh3QhqIUcKKh
5WR96rjN+xheimCmSLWGEaJWDkIRHz6XthZk/Uzk2C3k1YOmuzLGBX3cf1s0+LBBk8r5vZEfhwy3
t2t3Q8wehOKempyXeeBfZtaUtPc2jeTH5sOmZh0NIPBuNfBPvRAFQQMiTLGdASbMakI96bFFz7mN
1S3oXbATMhOnkYG70r0vHJRz++GGyOfwpIo88krRAsCm/XXQ5Q75+a8ES7s03ou6oAVNQLrNO7v/
0N2L+MS/ZqKHRK0mmDhZxccMddB3hkrhH5kFGzz4CApa4aJjkasYMD29aw2LWclYxFlTNk+VXs+L
b5GZ53XKU1U0NSHuJMur2oev/KYn++klCqcrifHWoLVyMfraE808BfEcqFDRBvB1lZfNf7kJVPrp
t7j95eTyoNo0SaUmJSCf6np+t5nmRYT8ZuJ23aUpeFfUtxwCezyUN1hsl2t+FMKbdT/G56KPAfdX
QyqHHGncOop41Rx5Szdigi1oC4We0Ld9fDvKXcxy6Af+rNWcZ/cfE9mt41XSv/hlEpoxbYI8D3yQ
+IgqnioVJ7vsa8JNNL9sMi0gLOY/MXNTmOVrMSiU6aAm+fY2RW2PJDBCkxMZA+uweGxSVSe00dCW
3+l4BAUl4mCNNF9XtoQwXAiBmt9zHdt3t6WlHKLuco3bwSAJ83nzKudCtlDyPFGw1dVDQMZWdkOg
GmvXGX8LbVwgwjBqSboa3y6p3+rDzW3NXrQ3EW1N/0buWhj8aoqBGGm+S9G0UnuPCsjyhLW80PgF
0P2MHULmgriUBJdI/pPjgYwE9cJKdyV5ICtQXzm40aY2hr9fU7p2sj/nvQipMVTXa/SKsF4HHuN2
9VXPE4/zorOoADguHuvoLrwMfa9ODMXUnLEHnM8a9VKz8f6J2nTOh6f3AEDg3UHRMsXGttHMRfEe
Q1tjnbqU3h2LExdav8ZWRGU5LPy9fvIgYGAPBo913mX9tPkUoLF7UNJ8mNrElKwsoCtGY+214ciY
n79n6IW5phI2wPV9NBboLgfvrooYjZB1coLtyKtJrGmjS0499mDOH0VZwpiibSiPUxW0boNgP+9R
LOIxLebGCGW+zuE4pBLlQzDy0R3Rw39bOjcRDDm/HtCK2w9ith3WPn86NlnVvSinsrZaNzflC7Zu
YFXK75qaIXzrfsGGas9/6O2VaoJhHbohDTFmtEUcEIqy5ZpNx4nQuquc5Ov348VsElWgcbV0rnAR
vsW7285I/Y07S1qlK2+ujlyOnGLzaVeRlzKxRWk8XVLkNyQJDxAQqHYwUj1W8ndmBqblb7fwQU41
/hr5UfztBwD9TPP7bZ3Gv7ZtPDdA26MKF40OhK2b6z5krbyHYhMITlKlPDU6kczYy+jiEoZDUd6I
2NqAOUs747MIaJa3/ROPFeipu+omESQe7k9MOCBeW2OIW6hYjrouGEB5+6c3n9z8oVdYmQFhUMIh
cLnbFcQ1XdrAdLXsuvQwET7FJqKGtL7o8BAc4uLP0mPlxAXf2Cl0u5EzDI549mwSw//VozAqMxG5
sTrU2T+E3dQ3Hligmvq3heGjJf0Didex9bsmc1G7g9bJobg2HpxPf5cD3hJUM3xFDROcvUYZNO+e
xuxSMLqdi3HX5gezt8QNumqCsbBWZXRBjmbnyH7XgGO7EZoekVfPX2CxooyCovXzPFnHRTLJWP7U
RFFTsaO+crHuyXZI0mdbcXYvpd2DzIFlWQVjFk11RWQQyRqT+svL/QmoFDkxAYkQp14WuJNsuQCT
g5ub/8e7PQ/OzE81f970DMznD+hjbUp81KTO8KRNU8Sd79ul996/PWkYj9FFOnTGEX80pIdo2Xvg
SDLPx09iiNzojjshEy2R5L6Y7c+DRX6MdzpxT5ADqZwANWFJRRkqFNQGZcqLsJH1wTpK79oSuGLV
v2zHZel3s7KaQHGh/pn+TFYn3IWrUYKNPTSKEgajAT7nM8R4k2FXYfQj8kfL1yVAyNeDKwgVQuhk
dopYHfYEh6//6dCndAjW/we+yCOuA9yE0pfO4vDun2djQ24P4Z5tz7A0QLA9g/g+/4mkQ+7g+3YQ
Ayvf60HdAOSJS/HiEpKUhU1prZvniob6PDZy5onZrSckoAny6sN5J7XG/Ps3eK/4RP0KqmW4kF/f
W/rswKRikjxaqXT7wkJEC9BUdcQFwQxa4AUXQnAn0EgY7WEUyMCOxwBr6mIs68xTCVlkDwPTCZDh
86VZ+sEG9MSe2EzmdpyNVkq2is5nVGcxId+U9PobefgzN3hM36Nldvz/lqlKMz4A483xLGSgW3RD
h+kCeV+W1bOSVHiKgkBhTnuAUyLvAE9wEaTUrN5zR31g8ReOHM7vYelevMUgipSBXS5uAyqEHRwT
gxCYaXuzfjQnH0LLsTvlowFBer/kWcOId7G0Dmgd7WaKozqWQGOD1OWvEewujCmyGFpCc2FjJzTV
Zptgzho3Q+YD8/4jyZY+0gIuE5S6l6YSit52rnOEjKJ2Wu7mmSy5wqRQ8jkhsAUiD6yChYXNP4Ga
gKeqtGa/dXclx1zIp8UQZgfD4U3mOu7k41yy8XZ0yXgrKIy9oX+6r7OeIpcQ+D/8E3qj4rBSY+Yd
sXha/VLx06Rskl7o5NARPrY/OtDiexSi4wHABlIpMqpBOPYljbwD96FYx1u9tGNP9nUIe+QzgG3O
p8FMXevuKQAkAOsFhiZPjJ68/alRVMHKYk86sOvN/Hoe3tKlprEnAUK1JA7O/CDJmlT0StgsNtGp
F10gZ1Jb+CIFKCrnUmbwSxZhBVu7Z1uaT4qdT+PKPMbGrVYBWjZSdvD+jWIExLlcMEx7GMBibQBf
WkAMIvXcp0JYV1d18vq/9cmf1nWxvCg8auuyZp0TKMoyglg3ucnCkomsDDCQ9L0MoPYjV+57Bm4a
I6AfummwCt/oKI4rthF4I6Y/MokL/lnzy4piB+yau5l8jzg4pz047HBlsK/MclkfTIraxsepsFG8
v7sH/a5T8bmrr887nO28AK8nN9EemERCQb3rPCZJezSoYUEAhpjGp4RYIv1uYAThOfGSgrQqSiGJ
zjd/7ednJkGMH0LNtDof78KwKXLsq9Y6MbOSNhMyGOuOKV+6rKuZ4c/OfgZeZWgU1H3+xHAlBQPt
Q8xErGigB1NHnAmKs0GuVsdnIp4guj0FhMbg7Le9+iC9CC+Aka5s+rxiwwwkUIHS50ngxDnS+WUl
9RRJ+07UvbGWzXQ6objOs8f6mAEG0aL0/DCabMkI1qSKcYGBZqT/WSy1AewGe6eSKIuRD0notkgy
NTGHl/Zjc77p30J7nOsN8VWQVNHIoHYG65Wrty4SPsiBt9rpP6UBNhDWTJ6X6B/T1VL0EyPhBiGK
/bXzHF2es+iqJfvdMLP5dzCQ+1F+rYQsmKe9ilxsW8Alie3PlQFHPsDSOb5jXYePSIQ+5nkRxksC
kNmPRqutB/nWaStAJVFLHV85Gz4/bzRI4CMlLLb7WH0/O0Mhs7YFZ7NsoNJKHWRWlaFrQtNsASYZ
+O58cWVLas1Bn3sniIbXlPb/dnKb0NlIpJwBlLohgI+ecjUb9vQ8/YejbZ9CPqW0bxOrdtZZZFyp
v5vFS35LSD/44wAx//ie/EFK456JEl4G01z8as+IIZYNRB9x3BZMG1HDtJIbZzd5qhkhTKG+asO5
sbh/g0Qz2/yVnMROvz1eqV0puh7byUjU/6V6BXNdBcfQPNRGbmUFejaw4IO5lSq4aJzLxMzLIt9g
XzPUoUYq+bma3kAytKcF/dbyGuLYwWZuz1Wlpm+3uctZbwPU60Ytt4vTr160cK0Sbqj4u3wNQQXR
ynwGC0nCLzBZOnRYquE6RK99tiL2UDtzcwaryDZv6Wvd5UDzm64uCY5offalqPZGBpfJH+rlhJD9
mhvnlp0qr6S82nWyhLLcu3pR3oljQhFOQEfgr2i5rkO2C/vn1+mvUVouwero/MlLE7A57G93mSqE
Q8HeArhgsv0j+4IN45cAWPt4TBejqdAC7pYSqa7BnIzI2BIJGz+vu/0SoaFhonM3dgEtBpXojl4H
W2d26xxYuPALbjcycsm4NPT6S9C39ewTGfR7yQKVIs601iA6ehRJlJ6ObPjFoOj9uO1Sz1BxMNrr
afSrRit9MPRNyVameeYrmBZ112I72mGdi8iaaPjPT8hDP0ZZtl5G1ESFCOYegatJxw0bPwLRoUGt
I/VcyQ+C7egaAIhQ+xv5DGK2SVbBkVvrCd5CpqB7tTPrY3v5q1LVhJAwVeO99U5IoBvydDbma9GB
REi8koDArUIyy9CUFLl06EFcO7Kuqwqw27rn2BUYpfRDZH/QPmdd7iz5Wt81W31CT3z0g2pdpvW8
rnCb7vwRXjuPsrIQLPTTPLasTF27aOtdtNJDYej8cZqVuX7FrhWUfMNq+McHuTxAbRIBtMs6FhEE
dQMRf0h020JaO35RgEDUtBZDG4+z2N8Cqql4oYXULPrP5NRgl1bKk2HhDRJFcyI6IFT7+bc/0kPP
9JBQfGsZXnq+lqNPLcMyyzL7ftb9T5oJmybszHmYl/E8TBvldB+D4lw/sjdFTviJg9PveL/houQc
PqZhIvsK28E/ykHZb71qgFbtGDQErIwEEjOtLoGQPQci32edxH1u292Nv2PJDsai/2lH4LEO1FC+
4Aq3zC1vw/EPd0XI8P+Ic6jG5j9AdG7ZMdoO5N8J3DL464nQUg2dYrDKrH7iNkrqkLf3BxPSAsf3
wKKVrlLkqwZsub1gpzDsjd/N26a6aOee3SrPF61jm64ukPQcoN+LCAQIgITtewvHrdomY49l5WbB
HHdgb9ZixuxK1vzOlhgwTXVZupFt6KwS+S1IHZ06FdGrMuSkm7oeEu6x63PIJGCWUoVoFpzBCec5
i+qL/OzsTqnATDztC0gXHqitEc6pKwWgPsHxA4llfLUCBlnOZsnoQmKayAfizuK317+ORLICwlVj
bZahd4OA4k1GZH/GDQrpe71k6T0nERDtW4oXYcfqXYlyTwUrRfAlf8od1rrA8VND9YH/UghiS8oq
E8kJzQsOnwGVEAjZp8ey4hS0wP+wroPtoa/xSHonPUg4OOViDVFzecKfv0w8FLZWlXgObpwBy1vI
iRkPV8V06diTDUmnRsK2u4HXfYJo2XelEdwM7+OQZzMw7NzSD1aN0/gGm7XMi16F2IgE5ZW2DqVr
yT9afYndR+igMmhP5dphOKDzqZwWz6al4a57zT3FYIaeNV5IfbcV38HFsvWsuZ+c9yP1LB2FyEHO
+KlUK4qY1RfLqr3iArnObBg29DOzMoAaw29BFdhO0mnpZsKCeFoS3gqNTGt8L83yY0fM9coMTR1E
dpjW2T3Ed2bscfx+l48oOWluC2TGyC7Jc3UWprWF68DJsiHEv6mjvS66/awtUnLcnBKMOXs9aaIj
d/VYD437D+Z/4N+OtU3BYx2bA5E8WENGXyeSkNHoDLs4+5bDkhwdkwvIWvtbyYqoRErJcKJY1WS2
26+cdGkOfSgWe8ZXlQkl4uDH7PZNpY68ECTK7NIIA3INKY1UTcMx95+syZ/gS+AG89IhSeRZX3GP
ABBoto+EqMol6JPH0ez8hZyhXsHNnLEzrUcf+UsiLLrOaqaJkDrlQVfV1gTHCAiTulEmxrNuKeDG
+3BnWCDhern91kY+zX5mZW/uaEXhzh8mUkZ1+2djrmj2Jdf7htKA8mPgtS072+Tn2oOV3rdsUuuk
M7c2CLqS1CkhvW3kJEDbyvc2tnnkKEr/h2bR28AM3axZmUb2g6xhguaRItTEzdkl5YpJ5dvo8Zcz
4/mnY0r0k9WtCPT0pwY0VU5eEINaGFZj86yBeQ98GzBpDfOpSmx1MOFV8pZzY4ywSiPZ79nChXoM
InMLfErm7YlwZRlpuyiXK6dbW6o5FaXhh24jXz9B1K2Kynvc0R3Y+JBn9OCzb88lxjYE3mP6Aktg
nPiZ9lDdcd+ra7+UbBfNzpQxceYj35is+BtPWgAhB94mSrzWAXd84EFuSdV5e1DCE0yt/kLntpzT
QEZ4XE55WsRkTsWfaNrjzGPvZf7q95JF68oHmw+IAPM5MVcpDzLH+Dy0NEwG9CkvYCPtbq0Lfxm/
kVGhktVRdre/p/+Qj3zPlYt54vBtkK7o9oEy3bJB3nTuekdUJ8PpfiDDTvo/fUIETHD/CU8NXAfB
16yFSaV8NwF1cK7Y7dR0TGBh8fCLdBGh5nCW6uqMY0vL5GDX0vfQBEwgEr0r38KM2Pz9OsGQUZpr
9nG6BGKI+YNLpCYjbIvboa4W+KhvNQusLAvjnZz26xH22um6Liyhnuho2MBtALS3ouikNhdUIjmK
vxRb1UY0Ru4P/pj66cJJ1HvDiMdZehfuw7Q9DnHGYSpvcfVJa/JbcjhKLqMIgR7X99PlzpQVeOCD
AXLskUHG+ZYAxr06o2PwruYl9Y4uFA4YgZEoWqi3l7KQZLF+f70KaYmWnDnTnSUvFTLbY98zqt7v
/PCkkmzjlPK4b1wphuzam63oNrsTE41Q/H6KyDZ42B5idPjh9Sn7CK9m0ZnZHqAWah70ZdgkwSJY
4bppQ1QP+PewKl/9ZfRpcHDMVBJKjzJ8tmkK3EpL8XyWP/wLtNjiMb7ZPTYCeuNYWJidhFrejFhV
z/AHeORRNxFzdBp/CUyNo+//c8W8q6HN+xfdSEv5JcFSlLY4F7haSWbQtN4sUluGuPhbkM5tsgJ8
WMOGrnhLW4IgW3S8A9ekuhGkwkSBIvfxEArVHgw7kdI4NpgRq50gPNxa1EfxJEtid/5faEMCFbnf
m2fc2YjrNSTckYffvWt+wo2XB1anLhJ63hSMSmdQbTHrHmNEAo4HOrv5qQt4fQXdMj0ZtqQmEJNW
FfXpHvPAyj3MH/2eFtDTydAJ4MDJRL8cSgBoIioLuV5gcA66lZL7S/UR2uw5xzz4CllqVufgTI8C
vI3bnLb5MaGLwQu5RCGiehpmzJJY5xXo2q7MTfftL094ASf/yjGyd/aO8Ocu3jmnCnBCpy9mSeDD
fc44Ty+IYp0XHc8JnDH6CzVmMMEb/cmZkuSJFsCYLqAuK5Dzwy+qazlNcO5n6hhhcoS6QdIhmOe6
m9pAL29dgvahASPpE32ZEsuJOBhUJIUbHSb2ykOpOtZ4GxauodTqohIrQVQXT7acNQYyakG8RhIo
voZ7ODYBl6gyhgO0rG7Ky7uQTk96JeweprMgi4GOvyZBSkeQMitBkmAor6/KCuQhULgWGbfO7xUg
li9PpNkboWGViFP/DWJsEGzeicyhM0Mdn9u39LtVmusbjogwxgGS/hwOeyDToneSBX2H2OK1jmlg
KrM81BMeeF+2YCxfOhZIcsLI+PcG97fLA5VVeyFSPG9V+JJOXyumwypOVk9ApGX4Mj3NfRL/QKHQ
dJnRG1yqllOcj8pkHOA3s9b5lZ/FZQV8JS3/67qxRvwB1IgqY58z4ibzEwEklMrh6TxlBSP1v5tg
YXPr1EmCde5Y0WXexPD0oVX9bAqd92cWDqfHtZCKi/DSTTZ3KpjMJhqy/anB6+koKWfj/4ks3bhH
xdyPjwbOIYSRB+BGul49eNMZZwUtkKz0N3OKwm3rqOhlCXm+AHnBplMCPjgK6dkZj2ZRvZnRis8E
VvxojXRPQyb8DbWTRL/prbLzkSwEUj6H20ZJM+AwAQ5pQ0vqZzuCRMze8T0+6i2eVl6HwU2CDC6w
51WOgKHjE9guHUqhvAdj5oFUn1R7RS+OPYPPLSV5INDtkny+i6j7MoQCBB22h9993VOdBVMqaDLI
iBblVqHg4mmJg9oc2aG96F1Pj1McHblX34N4Ia3Q08nzK3p0PZ+IXaWbPbynOBA6FuuzHLmpuDyD
C6MJLSqX3MKP4WiZm2B/L8d9G6Fkuq6CM9rH6zntpfD1vtBqL4pvPItZRr2kFm0jujeQAEnjqy4C
7QGR2RYN0WAZgmrxxPCOlcBJ64I+u9/5eoFVWN5X3U19wvv8c8SZU6YWugoluUKA/ADRsDcN4t+8
xZjyAOxVR5BQJJMrkl1Jm+10Y2ZAJMnLaVyZ4asJ31jxeWD/n31TxUnM52Rtp5sN+3ETW5kZL8RY
UpqIEhrvPMGj2scSghvl2s1n7B+amt/QOJ5sLwyCF0SNMauokKFUHEBh1iO1fi88Xf64wTOeJ7tl
T5G66pcU7UbqofrpZr0Ea2PuLr6RUN+CteWH4qcsgBDEV7zABDS75r7s0aV155pG1B3IbJBzG2VA
8EwfnqjfB/cx5G+QqtNqIdmxIhA9Svi5XoYOgC4NB8KmmzG9DeuwJ6egcMOcFoUBgM6AQ3xVWvsK
TnOKYDP9jBw1WjoxfDDHWQHyfH8QKVkk8FIxzMCalOURiOAcIyZEt1P0mWJdVDHw1k4y62Cm/uTv
1qMIzCKI464jHJl4UtI1rvNSECooget77prwEeRUvm17q+N71SxC9L9wFjD+ulU6vWUwGDEwfKbx
nXoMJhqQP7iDK0C8JYx1QOn2fZ0fbGQNM1tJPc4Q7Vyv2DDd9TfSgsKQyvgaV1WxKHqv+mW4YFHW
Te4AwvK7x+rnMnkWJKx7dQS78oVcoiD+y/Fc7pG2Qk8hyVtecz1lA21wycWu7sEQXrk7BJUhKmm0
uB/SvXZPPPUQrniyBOQxIcl6hrHQLvfw/ofvzW7JNUJlpzc8EJoh6JdO0REsPIn3HVfgAzCIdQD+
Gb7J1sKKGg8VUVO3TV4Ej+il0kl8YgCzZgNNujHCD66nAEVq4igj/n93xcRzjS+FtjH4plOAfUyg
lI7bqSW6Dx+7DS3tHGg7Co0VcANYG43uQIKqh0YTMQa2XD2Jj8tcDBl8BGw67q3HHH2thLXUveMb
SFmqvUqBLTagEYmXXX0RsIwUDY3bWR9XAuQntW9s3RlFpbiQjyErq3IgMprAvVH5g8kfqU5oaPix
kZH2MaAdeRCZMMO2Rcsbs6oOYZi9aFYDEI4Z4mGAElNhNBqCl6QbBUO0qXWK1rJ/GLGQO9pXgxt2
By1/EwKY9yH5rsTz0Bh7pjGIgQ5YI1Wk4G3yR67YgieptexQ8Y+iQ/ZMsRhgfS/Iq/2tSCG+VakK
LCgDEr3AfpMD6PDWDjUzmvSgy5aj9IqnDHQBzyDy+IuatVu/31P0p076SWInPxN4ODqgfm6VGJgx
W6n+UDwE3T0CjoGOqk+2Qxn2QJE7LEbefhyq1a777cxxuTxZ+0PspBYJ00O4nAUc61drIYTK5Z/6
5ebEWjQupll3IK2PtkHBG7WqKLaMtzJUKLmyb+j5e8C87H+OV5PLNM3Q1DB7J3pCMdFqSmL7pwJW
LknPEoq4lNRGjHv89VW7sA2aHSNsl9gMRIFOpmOlNdJpZh+MndDGOUEITEID4BILoYhZQ1Q4e1JK
5yyyXuzNu9JaRpcgDa3p3teb5UvEju4m0/cpEeIMFjx3uckz48OO0QkDjTJsPfbBtdIm7ZQEWl7p
SkCESgL2m8G3aYS5Bpmsv4aiGtF98dADpLkKfgcfobe2+r90DB0TEk/EB0sWGUjthcHZjP/IllsZ
ahMyxhTNAGMxnoJdIE3YVDjb6/GktrKMtveDv3lTPNy3+sdJRSbfza3AiKWME54XRjSin6cmAylY
h2P7+RVqXW0hYP9eMrVwZLzZN6bJHK8KwE4J5l23ZzCmdM0rmzlBgIZENXCyoIrIm5qVCAL0XAN9
dspd69AqpHyyViXgj+/T/0KWI84DjKJl190zJ1Z5p+rAt26I0kKJIGLadhNKquBGop+GX8WqPTBV
qS7SPiYw0OS1+u2mGFNhtfX5woLTcLWrcCkgORT8Vizr1pxKslNeogd4V/2RqIaF9eZWJd6UBQoi
uF1Kr/iVN6WJPseCm6jU0TjthFBLYIbLIRYiSBYj3KCehztT//zOLKj+Fxj+TQtxQEiXnaNzA+RD
nUHVovbod3Jhqb8nZXGIWrpU52MsxK/a27Hy7XCFZj72Z6B4gn1HySn226T5tWl1Ka2LgryDd08i
2dUe3Nw9LRaHxTwytQB7dZo1GMFoZ0qlLk2VSpxOX1znBrgObeJta3ciSkVIvwuj1SE57JAmvhrB
W+2/j/gMFDJBq6hhj2v+u/EulUNCCkN39G2fH3fkFw0+EXNkNXxxoS3O2f00REfk9fg75VmbWgvO
/vhUCc6CjC3OyNk5CvG1AtFlSOhOZ6er0+4DJ86JS0sJe/DVBOo1Eef97CuqCcXxnjNeAs2ovC4E
IwU+Q7GNtTZ+bt5QVK3pPMu+O/uWiC8laksZ/hE6aVA1jC9NTUFO3SB6GXUC86lr16CmNQxWXcaq
exxQDQ3X715kaT2MWBOTiLNGUXvFiIQoXh58XVfjFdSpRpY02SLc9RUF8xeptUlP5+kikFoyyNhl
EiPmntm2gh94wMEg/LspSL4V9lshC/dPhFqSvbKdr/TtoG8HRL59VcAPNF3g5k2LPUGJzcibtfih
GWPSToPhaXMHECjQI2iiv/sxjeCHaz1jYmO0K6drGVIXX4rVV9l54f6lCnai8+OTVuMQl6qQcy85
gkKRT6PKILxTRvKTqajggrG2Y6ypEJ2p0hIKDz17Xh9/4VWBmuT2UOh9l0pJcCi/BEmdGjpds6Fx
spEomQeSlLv3TODfXT8Rt0HF2Gcv6ntNIa9QMM40N3zzr8gjUQMYAt/6u3hu2cGpQvZSD1Yuq/2Y
cX68yBGi9UT/bXKqcqfXDKysTfAwH0Pd5QqYevcowqfjP4tQTVpE7ZIG5iy0hmku45JLm1rFS4WS
xs0CnQUDAXn/zoNYPD6NujIJ2uqlSb8dL32PDJcB4lJxVsLchDg9peoltdPuO3U3wdLT4GEy3/lO
aR290sZ3UO5rBaSiJCDpd7DDXpq4j+4z2DPxnwjN+8nfgYxik+YsMt4eMeMVdVxCkWVS3lbKBCc4
QK1g7ZSRypiePWqtDU4Q//A5rEWKcnHdo4mmijbg/I69DZGjE3I3fzbdE8ULA3hzM6xvKCspperP
102n6V7rkWv2SG2ODjcEckW+uSn+EK7tOu3+9owctg2zHSui7bVNFqJri9qSslLhpj6H53/xSuBu
gue640v4FOoHKvybOX/e5wwadfPmfFB1qWe57VTVkkGHBBDiqtIwqlQVOVvUPGVsKZsut2C6RPDb
YHdx0EPFphe9WpSOXnZ8rBA/LV2DU143w4q1rSgamfBGtyMn8V/Fyx6bf35kQGWelyn9E1ovjhy8
ptXxmXXeK5Q/Ht9rznvfPJHJbro/xGIubfUMRZPwRCX1+PM+Y3huyFXEVbaYvTH7ABlEHmvA6XGW
u4tGhW02bO2urIsPyehXFw/atcNKUS+bFjj2ljgDuqeruwXKTj6TMgWHq06Mprlhksm7/Ig2ut52
GRtEEbkJBVoVYUrhR7sFZX0Pwha9WCQ2xBoiBfsfOjwPiyJcAhtcUs5vgBg0wUIrm+P7sMQQOYiV
4yDWGQvoqjCGEQBhEojZI21/OBsQssohLVkDLsZHFGiAOacGpFJbUP4fpYLlG3xLF6f+O3oPkqfL
+NooU3m5f/razKXN9JFUFGsvBp4js66VfdnRgFikNdOZzBXSovbfNRVKjiqiku/XU4yvBJUoWoxU
4tQZj40vw2aH6b9UR7NThkLnWe/FWVw5PC0CalixZmk2I2el3vupWq62BddTYgXaYPRvA+nxiopt
moo/sxNG5isQDdV+prf/ESop+AKCbVJrojwrLv43KTIQB2piert4ppe4yfVfJURkysY4zInY5bBM
99W/YV1bg/iijykQYK7jtvDAWE8EQTJe/F7eaPmHdBscF4pCTOCfpq0sq3SJM/V+sYUKhLiq6GA+
b69U3w4/+IuU6nR5lXZBeYDLihVNN7ukL6QXjsZ7PqsHXnRPeqc9GAO50dfMdPNdEVfDjvfGhz+8
tyAqjGdVFKExEK0v9Wt7yHe0MGAWWb8mXZgmxbO/6VXURU11sAi8eK/qZejfZsh8buXykrpnu9IR
6We3i9mPeyFpnp94/YFNMe3mwFmAEulAA5psqtEXKcVUxjjY0GUtLEvpd/g51GXtOixFe9mvEw9D
sKaft1C0BWzSTukDUqgpCF/4FDi/CCEZ7ymeRRrRP8bsdft//4uXFhDMTWUo9Ka9fA4A92wyUeTh
zQCpxX+fpo3L1AZIhPzt77nNhYIPIAFyYIEjaAywakMPC6T2kue2sQa547QotUXhghNGMVTmBTj5
sdPi0Ll1iXUEkEwAhSUayKUusTj5XOzYzuGrFXvIo9leqaFUnMBizQtJ4hmup6k7JkiEH7Vt3U3b
YJEu8wXpyxKdmNGxOLpSQaGc6Ics7tP43KeOAEBWx0NbfDyrSy9ox1vZAQzEERCYenYvaCHzgyqh
DZl8J43cxLu15ku5fvLgCFkKHCdL1LqGSfr85boU8u+iUm5AvEv0kiRk3DILHC6oL9j7wsHWYDtP
qHIAQQFhVIwbz9WUV0vl8ToWkbhiFrA9GSgBX3I9g9qGACccs0FShW9p6t+s1RfDSeZvy1lSFvlW
FMooLcQHk+h2eOOsepoSIWs2hYomJv/Y9qs6wFCyqDtQyiBK2qNGD7timsMwGXaZLtFBhpuQDYva
fTMFzpZCXna37rQXK3YR4uRreR3hnhkmA21AlM9mG0mAkEXALBQXAssKk9/K2c9jLW4GoX7hY/W7
46RAPQN+XJLVFZYeNieCLcMj3CmQ02oM/wdINnZHHgmvrFHTfLW3jgIRGY8NGRruZXp+s65PcdRD
ykyOHfjL3swpno9E2NGX5KDvFH7Uk4nVH/pOzlTaqN/Echdl/GLDjy+oCTVr1w2Kk6m3AXG7d5+k
jB/Nf9mlgCMD0rpYHcWLTvsGViUYo/Cl5CTMRc5PtohHNfboklrV80qMF3CIQ7X7MaiuCV0kgEd4
rG/y6HiZIIOzjHY7z7yml4XMr1DAmWdvZz2iL+5fkFnmAQe11aNAGPTPZ1DKxKFWF+EeduG+qiTh
gwlwJc5wJS6ztQJ5lJwa8U1WhA3PTUBxjTtsvHSF1mFhaanN/7qJHQBzC0KVm3NieOHIUj9Ec4y4
LRLAcbMw6F9IwFKPplB1hKv7JBG0iGRcfpilvLkw/bVVMoaT7KOtMLN8dsBsXvsGzTziwUNlzV7i
3TGspJn4F7u4ovVn5990MpT/YnLmBS4FJE4I0hGYqB8ouZPVyXxHexmEEaKSZINYNOjWIAXOc49f
uitKNnIkiNMj9v78F2TOdEPdwna3D9nqMh5cq4IKm3AOcrTqmIJKW9tNoStXSkywEHVtq1Sq+WOK
xgqmhhtJFv63LoRACxUaGHbvQWc+H3A5XQfcxGtjmyiIZq1j6V5SN9mn+ADJ/PIBpHaZCpwGEvcL
tl/hsLzP9jYPRuW0FlRN7l5p/lR6LgViniRhxmq5Dw+e4hWb3zljIh+nP95pKO8+g9uZA3CHajlc
eCgJHbZhG9RfjiC90Dk2FZ7nVYtjU5kic1+CVg+C7SLK+JrXEFXQWp5KIgWDgzk+syKUvbHTa2yD
Mumh0+eIFT/q3LNYL7vuripEWD3WJT5baJOIgSGNFERXXxtwXMk57+qETGSDPR9H3Ev20Ym8F1iF
/jp7gvL/xv+R/zEumd0cZVSkviUafBE6hHikfAM5NhrGHIBs85a3gvZPRhDqSq3/RzU7z0KZK+mB
TWZscZXUPGf9xRVsfvbx5YB7mc3PMBGseQe+5BBD8J7So7gD4IwjIzV/DbuZfI6CHBHfklNymudC
T+7Z31UIMYbhLsDC7JQZjivPCLqCZ53Hthfrn+XaX5OOnIj3zOSIJ9JHvguFBd9pLE3UtoDZG+VE
KZRTSViiIshC0vrsI73bqK+KMkeV/3V6vSxAcQVmdNa6+6evjRgFJCbNY8f3kSCn8I8vW2kQxXOR
kM/RMIVyCnSNggyDNM8eJlZfKlKR4q2lLRLHEWMi/MBpsnLpeHG6omWi8FCSBKf8IKnA9ihffkNG
Mqdttx6qIUDbt3JVhV7EQYg7hBVHriYYcvY/nZT+etKvuOuVOe54z2mE5jDjTHwCd3TlyojPqyYQ
7M/5SFBOAkpjALftACpRsrjBMHLrBXHW15a9kCnN3I0cRmlbF4EU02dUIQCbLZZCNeoGAB27x4Qi
Zghs3Pkt7Uqb3uO0TWhXL/z2PwYVdzzB0xZ5FxD+aSVRT3MdS890JioIDeVumtctMn/GkdzUwZZ6
rJPEV1QgDcUhH3wTbnRBu0ej83WbNAzi5FiYTtIQan7EJACvuAQ7dZGZ6qhy6DLaMGZ179y/tqiL
GRLFjxx/YRa0f9dT5pQn5qQv5s3ufap03ZUbVShHzxnndsJZpJJao3o+yXYWg5vPBb0u2nR6CZWA
lZgYjcBWvn/OY9DSTK6nr4XAXNS/8U1WcFxW16JpqyOucImSFO1CLoTi01HjZv9/W8zY1wzYArXt
+CSWBeOtq91jEwBxUq1yUCSoDWpspsoKhFaWz6wIc2Jy9pFQz0Tm3AKtn7OUPt8vHYa9B6VEakcx
ZgnOXrTRDN8N3inTx6gk8CSuEbm+RodEt69avpzBcGVtiJ5wcN8fRvgSiaDXY/wxjwmEt6jVHzL+
VpGPgEvwiZtG22hALhyv9+uC8+fjw2J9bpdfYl5Gytvkx19diKohPBtAsmOnU0dHM5Lv3d6n1It2
WOMakACVHIeEsOltEj7lynoE1xXq4YMTbEeoXr/xzC/lU1VU/mSQuqBOssTbI53aug251bqzgLkB
zPrTKgAxlQ3KH1tWdkFoCWry/k0QdhhIDtcoRuxw8QyyLAhgeBPLAbYp0nD2Yj6BrxnJo1Xnh7+B
bjdjh+b+kylydmNOe7R1Vfh7fNcyuT88oBQa8kjdF4f8KL9Gva8dItDDgcdrRmzTkHl74Ai7/dVD
7aWqzgmiVfco9HFGuuURBkJhlQHRjQ1dLyAyVw6/S1IuMVYjgCBydMD7o2knzuk1j0rMpjqKnuSE
Un1wZ5HADBn6TxPtqF79olXvgZsPXXWHSuNSLYjOyWOT8MCNVEwX8Wzqr41z+FwCQTO/qZqX4fBr
syJrPAQPToLEXRi4h6yJMuAgO4wPEj5iESPRwvXNNUhBcsLJsk+5S4kh85gKaeHNoBqdHBoENpUx
PWRJ+Q+DMZcYN05sgGHPXAzrduFqka6m1y36xKgCcIh+YyFeyN6+Q4Pgyv5JwbGXayju2oNtozvr
PuJUC0eeR69FoexhJVQcEtYU47gDFt30+1U4b97dtZzeIPEn4hHtMoFJVKPi3fRj9BRMGGjjIjgq
AdKa4f0IlI+3A1tDyLmYtyisU11EMDs28zlGauZqadvZOQynz1sMWQDhjf0r5hFNGnRnQ8gaQCOD
SBMVZT6m4cTOQTTNXDVsCD4Tf5xuhsNE396Z8NlUBnAcctB72/7QBJ31A/41ltWdaqs/ZWcp2ayD
LU5zlJ306X/IyF2jyNyqcUpMPtHrE1I/1lIK9f6YLD7Eizv+lqWMKY9yXoaMEZHQsK+w3yTd9e19
2jkf1YxWoTqFvmkoUQTSYvpUXN+EOUWzP9PgU/k0Sxn4fqs61qDiA0ulZ9fxZbrJV+7ZX63yim7A
mzvXhtOvjn14gKAlBgdOfQtqAu4YWiu4pFDzvUh20nbEDsFxuSrYQdgII00+a+bjGTbPfe0zLzA1
u6Krog+8yDv1gLPh1wMzLufX5RLKUs9tRT6/yKOOWQT/mAiDvq/7lHo4zudrRy6b+WwBmwm6gHe7
qdnvo5IVJyYU3brOfZblUYC5KHKNKopbXCq+joJgggOcGYT09lAecxFNNU3YKSsJbdnMh8atuDkB
QIu7+1ZAJobRCPPh4Hcop0GrnWMFLP3HSzAbda3E/Z7SNNfY8ipseQkcWVG/z9XWSs4wHZ2bpda2
eMOHIroV6RiwNiGrXbtnyLppoJHtlksxlOx5vdJBAKbLrcsHCtB9mQu5gufpAEUArcgNUm6zQPzw
Cu9bDBHOVU3/RH8nJOQoSdlRrnE3tngRIH7ooLIIQEMUZMUrOVdvo12KTth9it+Y6cPtwupneqv2
Ixd6iRMc/l9qQGq/3uMX9JsudFpFJbEOjgUKgBidNG+owV3Lcj3B87xKUDoZUgL4/QwjCDkJX0yo
yvh6Nsm9nOOU92L2Q8XN6Hu+rWYDh+K7LWT/aH7HNt1/IOH9qd5H38nBTkLKl7KM0Q+SDYFkbHm2
L49jyDGLoBmqHIg1cTbpoef6Kh/M7kPsIeShiMY+s4f878DLBtqWD1OA1cZP8dP+o7BUCvVw99bu
cYxCM1YXm+NR2MTZppgAK3IvGkHakDUF9KaC0jt57T2H1PYFTAbJ9zoK09UJdgckPFUCzVE0bKJ+
FsBSnX2iP/gjnuBN7jM0DFaYMIN0BDLWeCCOnyJ6pmcqE/s/hX8jZE/Esh+xIey5NqcFjGHRkPdJ
xvZKVFjBFQTgaR8hLaa0OS2qA7tpu65zun0CKHF1Pse0G0L5ZWVmMqewSi7BASCkUBYufIgJq9u6
FMfOG2grpQ9PF8j3kyB8jsnYWGX+gwGSKarbGdrsjT1sp71nZUs9Zd7FB+z+d1CODzDX+/9bVvJ+
x2weCZaC/l81NilK/qi7dvmtg9DQ9zvBw5FZTemf7n6p7El8wfdtGu39Akiu33jreJJR/AWsTuxe
l+Qv7qJLDSZVNIShc9sHH1C3gEqCGgi6yxip0gpkMXMwG1cRVaFx5Ulk2DD89y6pKD/089nhFWUr
zGUReXS+9SxND1urJxGUWc4ncfNuKhXzi01DF9Do7pi3hFSCIZ6nbb0rYg6yy2pVHoeS83f6pdwK
L0JLxatzdTd6BrjReUIs9dKQP9ZCP4l5+4JujTBxbt7NMbrU3r2OlrNXZ0P3NMdht9x5j1QTTp+X
SrjgkqlI7lpv/xzAGNVJKb+85sa2mRWQRe6BhwxAEVEzapvj4vjithVhPoGuG7iymTz2DHnsS6ii
ftKD/TIEOifiA2ANQw0/FgdcLZBp8DupGT0EoICg+RI84B/+Z3RHLCcaMU87Y8YECpb3jSMMZFQq
FTvfUHKRrEB41ziImiHi/7+lK9Kxg53QeKhmzIAWxxgzibf0tYdVOK9D0wzuqotESPSc3KO/7U8a
int/3UTrr3zFA53lkQ4X/WIqwI2qJBbs0pnELohbQn+AiFh/d0HT1lGR8CCdkHueol9StjyCkPDA
ZSdewdgyOn13E8MowMMRWRGnlmrJ0NUTI0TPfnqwz531+O9AP+J3e9IVNfeAoyb09ghA9nZd8q+B
DWi167qPht3ovpR7ttOpwzw9j7jF8yXIINrGCPWeQ4Vw5tM9wVVjeQQ2gbIZ1GdGhBomsjxJdnIS
93zF7LkR+naiV/VLo3fqhAlPozPTllkVgckL3bQce8RFgq3S8UFdbSs390B8AfE/sDMBBv0Lfthe
w+oUsMF3KtBjAR7UGtzsdi26nFdNVetv2YB+ZGE4msWEhPGDA5YJggP2sM3xLNzg1Z3SNhPTHEXa
4/hYzt3rwF7Yeiqv61cOG5fnpZqQ2gnF7DTJczD7H/40AFZtqAdLTxTs+UHaVBynQw2r6yOTAYHr
TJ6cZc3iE8mMYllglc88XTF72A2NhQeQgbKaWQoJILkv/WRwCBWg9Tn2zg6CfYfQvNM4qb4Y3PcG
+/hTHFqm4kILOdq076l7D2kXPxlETjn3+DWxl+jVqS5Qv+4C2EzHsKh2pobqt/qBpI90y0qxiOAZ
tRonH17esB9OK4gs9MKZUq4piCzf9Pxa1RT27eCJ1iFWdEakoZeTZgys/GBrmevtMgVA55rpL6BS
IM09Mqd0aIz9vQ3MWBHnFoXxAbfnVQdpSa2a9Rrg/hRhF4AAiQhai0004BREtd0kZNDOTeARiAu8
mYzeFedKoWUhsWjK1I8ys+APraD+Tu71HwwSERRjtOQGvzK69nBkGilyu6Sin2Ek/8R2NqV/7s5i
+OBZcY6ubkt3xNIeKYVTEdi517HB5T8bHsb57ZaBUuzdTBV125HAiLGvXaVRD1lHrWiAbVU1INSp
JXq2IYtI6k2y8fzShmDhkesaFy8mCJ5Tfv8yaxlddhTTjGiFtpVeoTb8DDgjbhfhXISo/XwJW7JC
MYjqdq1torAh3jOuO1oYjh5kusjAsiDYKLjS08cEQyehD7TM3jrPkjyYiYBz69XmTwDO7CnQLEkf
Ldp0L+5ewQvSdBUvelEfLKpTxPut38vSKqoUK014ALuifANAy5a/pImNhMkWOFs2IKQBa2FdOXxL
cxnqaNRzwELj5xG/6jzLh0hu2r+SJfOGKBFOLXw6GCvqdQhFLutVL6feihGhmY+U63p8rIun7eOY
sWRe52hgMbtQCP7jRINRmDQiscg7u2HB1ZtNrrFSs+eZDMrlZrvK86cDalm8Dr++m/B8R4BZeYSf
ymU9drcu+9C3GFxyGGruejsbppMPEeOyzRQ+RZaOqVHwJAevhM7/OxX9EZXDLIvrbYZjsCaliFAh
F0I8nNE63b3XWxnnVwMCbqJqoavOvDiDy5r7eq1MAUECqdpCSUyoYf8gPVn03ErJFixG/le8VYJt
HBEtZk8asFQDMSm7s8QlUiMnO9fFkFQV5YYn212KuKLJGDv7Wx0Vxty7r9rV8+dpUNHfIRmbYIy5
jhqxK5RnN2XkXkcMpWt/T25Q3Pv7sZH1/gentpMAHiQtxFu7RBlTHx65Bc7akFb9ItAVPIpUdu8W
Vq71D7qvS65oleCtnVbEJ2OcsIgZ4DoUMnHo5Td9idU3yvz065H/4ry1h3QaYeXwbpYmIdK+7DVu
SHyE4jVDqqYYU+b2XYXQJDYEDL5ZALWkD7hWMGWu1j7k3rlWmpdBiLM5ogF35k4+aMwAZJDgBFix
BzS/uLNgrtEY5b5jYQ/uEJi2dD2z/i1z1KE4l8RzTDx6G0C/HegY2gQDLPRmpzvRPhJd+fT3qdkl
YL+dd+Cw3SWtjL00tExb0flcDkfI+hk3vpS4wSw722dkS0zgK2TL4IfASeeaNzdLrYrcSCKfN9Kp
Yp+Gkw3eZI3vIZ2FsRkAdpd6L5cPRrenrtjrO9jHlSMS5RZy1CjNf58AxJ3ufkG8K5WAbq8bGLVp
MWSip3X0oYm0cx76xRokVc2ihMVKV0jfHJip0+NW+pVIwwnHD9zFN5nDZ6X1LT1C0HcxTmv6UiGI
zRd/xxcrXOx0I2qW7P4Uaey55tADzLaIM/hVrhfA/T0sYH+p8X23fQFaBcwzxAwTvtFW/Fae9BNy
6ULRYbSxIZOTY1eCul4RYcR7eVh6ZbLyqwuJIEBXTlTeC/zMXFt4VGvJGVGjFty5esME2RlGWYgo
thdXbtFblcN1cf9lj6yzUnLM+rxNdd5GPD143B0YCdJAfYrSUbX/G5+wwpl9MtRgL1YLX1Sw0AHh
RCsmsd1SvcbHSFstCj/TijixXdLYQ1mUu0eMqQoLo3Tht5XTb7yoXlE9gbKNGteN3q6umHCLGyVo
MUOS1MJE4ThHC20O9lryajrwRMtHNqvvwZccOHnQ4DLArUNrmapb/GU/sv4YTbzbmbSzkEOCO+M7
yn8aJA5WxfgPITC0S5GpvJLLZECqGah/ZUBCuRUumv2zez+icKJvDLJrMGEVp4L8mq0BtZbxXoSd
M0F1qsyAaNE3VCeWYa9a2vK+jhGPG6OR6bU1MJrVDyv1BSnxxI2chjexaDTyPzvvSxF4VYttMFkz
/fq4R2j4j5o2k6hdovhss1lL3CArDr/gZb+mErLuKiC8MipjCSwNlnEU1vEVsB+SXo5114pclcuT
sBNo6nO/qrMnVCpbisx2QUxVjlNsMDnxoZm9Tb16p7lSr+IN/njsHpY5C+id5B/bcJ4Zfqv1xu0A
1IV1S1YKxiFd2k0DmYJ6VLbwvWV5doQIJ3KgF9vYrYFwwls9TJJ+YGycJOBrsKEGtIWhnxbGx/mn
ORy+B6Z+Br33LwwTViiTsT1dWGfIzhOMCXO9RySYkDd0ohUaF6TM4soXxqKfNBHxvEAlfD3M86EN
G/lJb142IKfIJh0fcDvs4T8K80U2hlP+nZMbLiIRADzBxw69oo1Bc5W0ve/J+ajO+wi60La264zG
lGH57bWi8sFW+4vp2yF6Vj3mEJSiQB4jilB+EsqtgtMWNfqgC/M9yBAZmrTUYRVxFc3sIj0M8Yw3
KFW8MM8+KsCjnBGBCewPtrPt8HhbPbKtYztXUYxOZHTLSMFilC3PvSrFLDT0tXSgE10dJEMssAgZ
a77rsc2sa7LdmXIqvIyUVESpxgz1577s02gaYc1XLGwM4u3UCn0SdyvoumOYgG6EgFbjLUo7lcEe
6bnfHxpv0WshVFqE864q1362ESNUZx8pqscmU9VDn5u3AkvgRq7LfTrHZ51OaWOBGONK9S5SbbJ8
XeLwH21RSpw/ttuurucUyPZmKQ0pNoBrpZEBbSywIk9SEZJtt0xR4UJsGmMWcd2R/woi8xSXlNBT
PDtq1AGoODrXGplbwdSryrMEclTwsNOqZzpaiq2vB0oR7UaICTbUpxEjegjP4aBXYgBB8lo2QXLm
yqCDg94e941uhnlZqXMs8orV4TJNkbu5pxSA2Sd36bR4+E6mWjuvBamMGtNY2KvGcf2VXpiurUGZ
/3UH02iOe/U2m1Z3FHQk6b0zihS0ZcV91Csqpo2OtZHw31PEHdpCBvRy9T9j4Jg0ZdDFOKxkYZaX
R/Thpwkf2X4NEtMyFXVyIMyMJQwgt7CV9EnAiK1+4q8PEjhKT1vqsGzHn3SZLZwX9rj7gL6X6QNX
l2n1X1KjDZiVIwZj5Cvuux9auvPq6RxGroiKFftwjVDRJYxdWqfuHrtvu+Rx562FgmT0GaIskNos
o6UYwNlO6tCr5EmzTURt2J6MpqEuQJfFgO9YnqrltZWYo+sPOW1jOGnFqvqPoX3XFABRQ6AVnws8
72yf0r78hNm+X3i0vNUUy1dVjHLI0qdwekhL3hMkQrIcsKQueXDD2H2O0JR8RfUE97rwCjJ5elFG
1xVdOw85LNKlpeL3qORZzkEucKyWx51W5YncI90MsGQF/22yT3HtqGLqrjdUbrXA46K3jR5umg05
IOTj7xc4SINwaABOP8gPJp4BkrybCvusf0oqBUFJkKnDURDldAhX4+rMu0qGYrzos2K4VfK1TdF/
X7s1rj8wHirpd36YV+qHyvzQLrNnNn+da/fXzm4Pbpw7eakkIsDWHufvfirw0OrgKBtVC47ybP5U
aANFwOHJh7Q6AfRzO0wbsvCEG3K7z2oC5/D+JtRMYRIX7nkOLj9T+VxqCx6hRPKT70Ycryot8Nsn
Q06sKcR2WkiseUgrEr1xCfzPXCN1O8TyowTB426XRKzqNpenA4M22seD+K7SZn9UaoG3fQ+uv5de
I1tWmt6UzVJVYxoWvuiqohH0Uvy9fxn2w6TJwWrMiIK/N298O9NBKuhJuqnpPaRBrmdOwZad06PL
ohVdh//10Cxn1KzUTmjv48E6vRl1ebgwoLKCiQw8YONY33eJB7mgDCpeVuZljaMK7mfulid8v+2y
+vzT0quVafiMWB7R/fII7wDAT+wEa1JFiL3jUnpRok9Bo4zRYbixQRTSMi5IOAUFGSE+AGHmUlG7
cpo09IMm4WG6GslckIAsYFgsYRSVE9fkhqWQG131oPyqIIAxpPPoip2bmV7pb7VQILM5g68n7R6J
TGuhZh0HUszrlS4MHlgATNlqjxoOXXSadQBgCvguCdMg7lldogalphesdKnKK74V9WTYJhS73HT8
LyF9h0n07V/1AcQva0F5oEDDKQtpsl8Ba9aj5TQ7+ow4lSgEGpYur+hOcHw4hurfiDsyJiUN4cvT
XtwH7as17DJ3KX3x/6Wop46Lx5RwwzwbVNA8A3Kx4jisrvK8g6xDsaFSRUb2yYp3+Ql5gLKZWSFW
xyxylFkSIvS08AKhZM2WUXIM11UpvkU+UHSjyA3Q8w1smQIflzcj4CjDYvF+4bEYaMBprSvETW2i
5eSWoTX5b7caG8DxBcnaiwt5C8N4IfpsbNdkYSacOu4uZyadNbHoAfh7kluSLbFpaX2lhDfRb8u7
VQrs6/C8ADtVQ/yWaHgBjJwhe4AFeUfBohXxXOlsWYx/NMZ91mAknrXdj+McoV180R3Ypgn76FDi
2LSelMsIEGRpgcNMndvempaQdfgdeu4NviZy0u5m1ail+yBe2tWGam7uBPWQsFHACXpPZ7vdtMzq
AY1g6UMwW/HJ1RixKKVTpPGf3SsOBlZxR6VSGcdzzd4AYx/WG1jnvHuwbhei/1TQ8rUe1w2Kh237
BbS0mTQ4M21wDEWJFCqxm+BTvB5U25lcbjEIiFarbs3d6UtGO17Q1KZ7MjjixgK0WvOnvz4dIjFn
fbOs8NtfcGEJUpyrRXBOJ14HeAqTQ8wwWsTlc+YfjqCilHsfhX4vxqWvP5EhE1Hup6Q8S514Io9u
qomVgudxdMSyio/sk3aLAH6dr8fDAszMSVJ8lLR2cUVWQCXdptUrgOgmOjZE05GN/ULLkx9SzS2H
iONdbCqbJ4W5+7KxUFVX2KqGZCv06WUE4/JPfhbPVU0iyTAKBavKpaFRBNmjOwfQHbXsEwPIO35w
S1rWVtysEdpEZ14jvjrO/eJKVN9DYeYbfswG10ERiLOA63Nu5EMgV2O2khrxR2ryWVaQykMRIoeR
4+f0+yhwfPlWLFxG62bnCBBYjHMOO/sxMG9RDYQgznRqAd2dY9FnU4sGGJLmEbNHxen6Sk6Pggve
9zhOFxa8LNNcgb47ejIZDcKpZRtoL5QMK8yxyxRdogFfTqQv3Mdx+McKr4bGW5bh+/ludhLws6Bb
yr9A8KJ4hCthPEP183MQ4vGooG0kZRaUvoeaEsFNLaaDmSAphUs8rzSf292OwIeYDQlNHSS/vOMi
5vrEEW+J3YGldD0iYCnBvq7V/qYyjcbDSl2d2wprMrHZSQAPZ/BntcaLiFhrYCnYVCsimuWZDRc0
O1xoOBucYAGlMtM8rM6ShsWJ4bejQKHskTOR/Re3ODiC9GpAonTGOQ7K1aqxyW4wyIojbWQHhD1B
ZKInRzPCYZIpK4rWaAukFS08FMCaLqGWHWzSQklyGRRuC8BKEzET/n91F54D71Lh9ujBDSol06J2
mwSJwJcJOpfejAxDZUqHdfX3Y31oLZv+rIKDxfn5qk7A/xJXTaMzyoXCeRlbFW7dHWbxSf7DrK+l
K+1EwAoyuOp09HpKiswB/H9Mj22sqoxeaTzV0qrmK/oKYJ5Z83i2miTj2JL6DB1ghIjMxb3AnGGO
gyNrlsWREN/5PQ2as3FOARcEDsPAMMdD/MJOVM5fyEZWcMSC5lwk2eN/Lw28NXZYR/erG9NM8bgx
PfVwiq6Y4vreixBs6PDDcfj3zmYfic7ampmgqWu8saEbnDHPSq8bWyF7MV1u1R6ijA/7y3mCFOkn
+OagoefhJHrVBkdUq6bXyjiPxdQ5f61JeUV3jCHmsOowfnVy2rrihiN8C5Da3hOauSpZCXsSbM+1
8Rn2ZL9toWuKGtFxPrZzzJGDZrKDh5pndi9zw/rbwtksyaEWfQ3URVBIIiWAlEdsZ4Hm2sfgbQx8
FcmiG4wv8qM72KVgVC3ZB+wO2jBHIAUB5mXrXXK2r3EAF65ZL+jbDHXd/r1oV0V2w61PothVIzmd
2HHJs4U/EoMcHBbNptrI0Rks9qNZZ2F6lDjskPbpqi97c4nw1F9PUjSSm36b9tQ6c+/w4byiY6BK
zndMmm6jDmvMO5oysEKNAr8xqEQhD1Y1zHdur4EZg7zIZjnkJBU6szX3VsINROSc787qBNaWPztk
0RlSY/pHviRJvDmLOQSTx+vHZYIpu8PPMWorOC5hh80hMKWMI/6ZCAxvcnWz4aIWDl4kJxfK9XtA
KsC58eKYt88Jlcq2Q3Y38MH9UaZOAMEvRbkXy8HMtfcC0K7C7y1tvHy2dbxeT+1L+WLkzCiJJENp
UN4FrAPoxHWJ8dgdcjS/4DKFT5W5OBG51qoCUuNAg2PLB5pn9xEgUYPKYI+wb0AbHgzHwCu5dJjH
NaR6pVbEyPku0BhVPedaHBlMr3bw57TAwtqOSXp9qilJz8HOEROanlcouGkIR7wJeW8h1ZDXy4HG
6cKcNfGWvBhZNMXYACDcIX5diOknCReheetDQzOeDQGKySLVXfHyxuyr2jlcLBZU6vqXNQknhiiN
UWCbS+y7ad6b1MO2JhWY/bxE8KeahjbxBMhJoFwWs51M85wMhNcwmoWbKNagp0SyjhFrr/AGLqmJ
TJedL25oMylFRpo+xh53GAEhnUCtoxysELwSbF8IuC/cHgCR1nFu8fCdBgdMdM6razeKEhk0e5wW
4OC3iJ+yjdmEQow83fF6vUlSvN39+l5erkXh/oG5WkS0lD8i0W6HT/klR9NVYH+ebpXA/rR1GoTH
C8AqZ2FwOkUuK1NxG41QYurb7sOgfRRuatlSoSuDa5YnLWj1wqXhBj2vzjrfdXP0Mr8KmsTsmVei
16CwV242cK3lJ4u9teevfZ/wo2fsyYoChoQE14lLwr7agDF4ckkTUT2VfJzlqeu+XeWasYCrFwJX
SyTcoRpTopVwOmiwJAJX7N5iQ3MM+CDoRtX7exeNVocmC7X/FTvrEqlcJRaW3dQaCEpgHGs5ND8e
zhtQbkJAXLQqoKxyjJT0+K2b4Wj1hVUm8OCJYd6hoFth01m/QH9/6kVeHqShv4sRErMTEFXgBtwP
lcXf5ff2CXEr4SysjJdqfw6GAhp+E5lhSv06+zfL+X/wJ5KpnErsiNdWphFKNXHcoCd7cNigbg4t
/gsLKg1qddlrsIX8lOlCljEB01mPBaEvNbswxjxWfDxETvnGesqSIj+Fppt2lZLWnyk0waPgMmc2
tjtheTlSWi17Wwo16AIXdNhKn/RiaT5sorXhpXXSIV8Q8rJ06KFU+ONceVBDgmoVzFYv4dRL5WZr
cs2PvQ1g6Qgie5WJdWH1cenDIzHTEQ0xoyjmePF7K3tX1kybMV/k5OpaFBlPMjJjlukqfDb4eN8B
ZsKUIyQdfGIbugfeANirlJ9ytCRF8YUZUokkl+g0qbgaob2LTM/c5smdnT/LbhCcr/mTGsyXBa9A
6wlLWYnoha4DpmbnF8cXKTfpubQ5m2ZoYzQ5VZ90TgaFz+15TdMJbUbgHBqdOjT2mMHmSbJ9BNJB
623YxEvWhpwMg+vVNgeT88gePc/hSe14oIHenMt9q6M1LqDP/hebXUMO94dJj46NKDEfkpz+h6ZT
kSAXYgJiAdlOZvEObyld+c01FZfHHzlETap++zM6CQ6336jnfyoqU+t0tuUtIs9abjVedxs3pHdn
cucap2raOwGuKypfyD60siGYLtUrMRo0NRC0qRGqUGWkBXkjHj1Twh6tkCjQbzsW3YJE9Y5wjhD4
eH2+GXPuiiKdCEirKyUgsDFnPhyfHculHT5H0KEB+M9WiybI+Mn+y4w8FdTdGoTtgUdy1UhIfM2R
Ycts1NTdsrPrs+XtVlGPrwBX6vKQhSZ0xz5jXRT0/CsrMx7ygSAVsJ8HP/2lTL4y2TAOa6qBw8wX
MS2WDytIK9MAXZ0Xh8G5Be4P9SvBSpgwhbREO9a0WXLoys9202yrGyJeuXiSu1/tPOG0dgpwuLxw
VIWUMCPTi4qEtKfuC7+e+lnQB7ezHSjCNBEmV8CvMHI6sd9/or0T2z7yV7H1PCSPRslpKsQgseuQ
hZbn0P5SwgVGBcSztwbta1csNkim61A5ZCfCVOtkz7Xoc94KlHJy2pqLfd5ss6L0HcRxSFjw0I2G
YzhhEtaZeb4ksDymC93ph63BjZMgol4uIht/h80Due9ZO42ruUOMr9dHXTa6PCfCBhVV91mL/hJ+
0qkS4EsBkCYHB2fWQvyQFlny/lcFVAh3eBj/RSczPD20R0s/ojDUqF5Nj7jEVEjSYSh6Ojv/qCNI
iZfL+JNpYNXp7dVKm7rdbYwKAX8Kl6E/SKVgePHZ0Nb9AJzA7ZAmfz4ZYqdQM1Na2BXgqDcO1ax0
cEm+0v8rzTDhzZpun+eJ/9VqiEYdqu0z/N9Z7A3K7wq1pHwDJnZ5kxobSq/TPgUwoAqX3MQNZhxL
AilUTMAvfL7Oz1tc9Y1qPN4hgQIQZ24dqQD4wB/m1Z8WBxEuj7lrJ1Y1PWMRAA6/ANY/kuoEqsHi
d4I/i7yV934FBaaqUdvqHdLw/WWq+DtwTmCDKraK2tbsTXRqEbXWzCn2moN28Eb1AsjRXM7mRQqN
z0AmfEnN9rWgiio6yRuv74CIBAoMBDS0NQGswqf/e4ctavUmBqjPldT9GFzbG5P3Adn03iZZ8Dnf
XVF5xu8teaepa9MucPbmrI2CcKU9cTJocJqgbV6Ifo9VYufrTqel3KvQYSIxaejU4tOUU/MZFolO
/wv/YO2CIDk0Cd9HK5Hqx8OJqNl3YkoQwW+ECOYAFjZRedn2OrBTJr5UXh2Wyoj0hEmPs58gWZUL
pm/GIRRGYWReEoJisbFXk9b51JCYFSZqHH467eomP72yDRlvgO0GXtQ6MkjKNFlVjHraWaQFUH29
XvOK4Z5DK+02lCpnda5SboMUxrGJVuOCKrbvWS1rh5ipcdqv9YMCD8YEnVGwvVJBJUFAtt4XdPDQ
I0xkwIoqysal6ATqVClScm01URzDzReaoEjzmA8FkPd2Zul+gD0ZSE6kzByESLM0UqCY6scqxJRt
pY72fDChtryBwo+L2tU5vVhKXYoun1fBGLDdDDmiYzhgTJHqX3tclvCPAFqPHpEpHS2yQFUkrMpc
YNFeavbEUKp/5xxCJ/A3h1RJNwHX5QKcFDw4PxcfgfF7hDpIwu6X/TKU75EzAKnCcdE2wpWl+zHR
Q0hw3q4LOwwshZYYh3OMO9lYbFWMJgqwv9Smaqtz+DHqqWCmIazPgFi/4PrO1ari+3141qpnRF0t
xiC+bm35n5tEmUVcJ1Xj+y0Bc5Z7u+1id9Xrq5RlWufX4dO3bb97jqD4BHqVct+2Cdpt9xYycfvV
YdVuuDxi31OkFYl7HRJz6klDJAEHxtuVYa+FvDKFlr7jzGCqC97u7Or0BD+I+B2KzNwWc/TP7mLW
9YWa1z9cJoQ/vXJfHms0JQnUSTsDsHJmBmfdMg+Gove5S5BZ1xBV7N+wYjjdTB/tfMnSz/zv7qIa
MNPmW064b2T9fpBofe5t4FxOQ1kFGfgvOQ2vMUFckmmP4Xhpz+dZUYEw1C2s01XOnOr9DVHXWKkZ
weaUnJas2qa3kfZ3mqGUozAQg6nF+RsfKqzO4oe6rQrygJQfvuFfqRPvuTpHrROLHIPwesln7WnC
dWvN01JWRYVqx+sVNzZmbjFrV7Fc5U7a/lQLgxQS/dHPzZySgFdYmCXTUZLRmr3NH0f5IfpE37MD
zcBTJv4CtEkRHqmYRkRLhiZOHV32h84D5KnTMOGsqTZMNXy9kt9jF/LvsgQrlvkjxKqnnJgFAfso
rjk3rA1+Eyri2s8o+Vom4vaJq8k3ITdUn1gkkJxXKYXPYqUulUJek/+mH3yhhLMDahqRc2dJ7Alt
fpfC691huN3VsK20PIlHqlk3Ps5xULo1yYrsT5+kF1rRqwvj8FGDA2rgX9Cie+S/7rOVQodKuLhl
7KWt98/d+uLXJwQIg062gPHB6j7juUIGe15uJawjWs7YYnuHaWSlF7utR6y8GoaRKRmFJKDacn+I
t6VyGVTRmXtbroAepfoy7seslKgiAI42KVCaGafJl8cSr42KFqmUknrTXgOHy0gNFjWBNjwZkN9v
i4AMTafuDb+cS1CCQHo52PkOn/RtcU6iz767aiarE8UN5963lq1+9dBevLxaFExIrSV2QnZFhzTi
gi+YPDAiVHahEsRkl9egxWOqSYx/5Qj7td/UCofXqRVfI1cWDQEej4FEDYr4L8peCyQuoLZ2Fbro
2x+qrYNE5KJ7k7XIQCEF9cYEY+UPmGomgTNZEFBrUyYTkplHXnMs4z8EyhiN29sC65MTz/qCObkm
y8NnOdHPwZYG/Tn2Bi/MQzt5jCwYDyI4wn2WdeVWXisq7KOpWlafvLugbs7dY9rpT+VRNO+7DiGM
6QviIVyR+hb8vztD2BvrvaQNrpg9oQRsMHk2CPcAwU6+yz47GP2/B9Du4Q74kcIK/AEqlmNRj7pm
/IhSTqIhT6SThINIplW5/FMpNRoy6wxS+nwzPZAjw/Izns4QEQDeInsSVInXgfHAWrivwKheJmFQ
Uab55oRis0M7TbcZSgTAOfiyDSCM+WeAhLudX6tR+rf0/bgl9GAC/1Hq1HSDLjnOoS/yZOk2G6yN
3FoWDXvXlF3m4Zw8xzYB9gAIgl0flcUAM23IM/Va8J9kwA7dLvF6XjJNP+SdLdPO27A9PCW8XmqM
RZgqUaHoE1DACWB0g8+7TUnYrUTJEvSe8FeWf7zQgDsoZJpsljy0fSwNmVFGy1NcuDKoRzeNosN8
bpnyQcumEnyULh3q4yr34TTytmUQP6ad8YzLh4zypi6iNXNQVfUls/6Fxl/Y7EInjBQWFdGd3v6+
2eLL9BkRq410OBjQy+5WZ8B/65+XqO2qMlc85hDQAJqiEhOON0Z3ZS1WpClgOu9o3IODgFrvjpHe
i0JcddJHLMBfPea4n0YzPO2f/uKCNqPrZ7TtI4DGNDW4WSpuVd3Rt+PQCJXaydqOwY7TQBA4hn1X
n/sBy3M8iKlPKVd5ri+wcG4PGYLeAKIlnv96eTkmWv1xuVUO95ISfX60lYZpjWfhYmo5wFhyEw/a
k5er0Gf0KijskI80hqTzqq35/AWTD1LA2N3KRxDbzwvwOAGjZ2yZ2ugFkC7i6zEfAe4c5r3+yrLk
//Hd9zsS58YeR23oHoihAGgAKd8Z1S8fXgufo+5vEmRdjRy0iunInaioWCOCHZPJRQYdTYG9AUoh
fwJHf072EmC+bxclOnt6L1WJRi1ZLLA1ILs8yqhgW4vAmDogtq6yc8DSQvoioKk9ELESSsFmP0Bq
ggn1GNtZIUZAbpRJXY1TkvPazyoCSW2yAgs9b0VZK88W+OnlRYAsmdyBkjd9c9TBDNLr0NJS4v1+
7VTc2002Tk4ElHfUTtpW2CggKYf1jxZdCjU84+FVnz6Yf+YmQMdDzSozTQ/hjqxdx8J9Egft2yPP
jTCPBUxEWTXsmWISN3rycTuH/pfbHVVu6XQjANdYRWVuj0wyc557rnU05sUrFU2TvwT5Ql9U6xG0
4luPGwnKKz9ZeqT6quFbZLoZZYI5JLI0s3YGwGpFHI0jM7FljdDMz1cptsvmNX3K45J3ogliyWZe
9XC7tu0T3N4vS2BoLGK2oO7G2vDB/IxHr71348X8FQe2MOH7pFxMWeQZGQszmC39dCpj3UeYabnm
F8rEO9+ZeraEbmkSTfJgdSl7AJlKQzqXqQyEM83lgYS1JwOUnrssFIhirxZzIHDKo7hzxPZJ6fsD
C8uuxO0EILDVEjlKaQ66Dj5JBcuf33Mu6uj6gmoXS5nUb3gnoUuoyRDddj2IJudnC0Q0kAl9qYr8
MzKvl1geulWTr9defyzgyFabkApTlRlHwYuLOD4VLHdaTn3871sWAGXBNnMMLTEzG2/fbaocjITi
l769kcqeL68bOyYz0j6JdFe5uob6ZkR8eUZZGDlPkY1sjjLeSpnDfB2oGg7QjRnbuWVQXkvgjCPu
hfHfuI3I8DkL2iXt0ddtNVnrWajSVcaR+2TwJKFPlNvvdXWIbhiLyK4qTMWbDMlj2l0ud2kH3QBO
wsQcXHcTGpZTfjvlfzTZbpMlGO0/FJ8qwSrX5teXbDL9Urc43XDusblCFxinWnq6DhoLf7sspYbd
LoTr4jreURXgv7lgqHfq3+2YB4uPi2RlASs1a3guk8cVG7xyIUlJJdH2GhK4EL+UeI7UNNHWHaMP
aWhPbE4UGcbWi3gU5GePDMf1AvwbrerzYwMzMA8jKVB1RvOiw1+NRmyCQvYln7Tx52GXc7QpMfiy
IfUInGD0dX13jX+WZaDpLbaWm91kJ20TSqfrOPQn9gxEPDA3ytoT8fb3cpCX+4mJKLpjZ+4vKYDM
aRfu98kKFCtGhONntUO9pjn5MFaychhXS6WUHDum2xOyni81lnkiu2RNgzWmM2dzZVv9LQMfapvF
dHTdNSdXZl4ouNLvNwUQQG1honBeTDUrjlLuYlLdAthdEAuzwrlPiJTZGMuxh/3ZB/1fAgp4wrWK
zEZ5jxDBdWgQdiab8ItZkIaxs9I4iGQa/ZYYEb/Zc5ioJL5pxZ81sOWKN/btKxKEy97vNSNBvnk/
vM75XhBcFhgA0Y7CeL4UhUzgU72SEtNvCtnMB0+QX2r5vxinLQEOlhj5QFKfO8u/ah7MJlbEQXCM
Jjyl69607xJP7SnsPLkHueTb9oNG7kzzrzSBHRAJo/NYimq7IOqkSSO42L+nXTrGgL6wjfEMpi3u
bZ9NPsGglnUXcY0RpTJippZ8Oy/I6EghnUryuC0zyS0zdGq6QpMat8ggkYZxSN5IV8DKlnN8G27T
EQ9ngE49zi/JiZsVOfsWeGm6NqihHl+6wmz+RKWdXH/crMsPcvp3Gs5M+T4HZh85sA+bwspjSUam
nLNh7/UyWjWsybEKhxqqdruhoirTWHo7uyUF1qRD6ZDOW/TFr6Q5YONDRjITt7ULnmGMx7JhBkXJ
+u/jwEFZ+Fjk6d7qW68BsXz4NlJo1t1rXBtnA+fy2PymraWz4u5HLfwr+deYFXgzjwhrp1LjjEmm
TUiW6DWl9yWwrZwKt/CZiIeGUkvZo/ku+OduluH7Q0aY9WJF/UgFTST01sL+8z7XyzL7uGJkCYwi
gjxwSMB7D4l+13nSNLaqmazwQt2Ivvbrr8nUV+X9N0hReQbF7IMc3EwPuPuGea6bAT8Lt8oHMtiV
VsPplXonaxbH7GL8Ouf7VpiZVXoiQ65g2zGqG0UG8wYBLqP/rw6Hl3AbWWinGkSNIocnoBOoROuo
mnfrFdLZ+rdRHEgFgzc6Y/Fh4X0P5zt12FS2Nq7rpP0C4kO4uaHzcYNKwMIkjIdZSZGNSJ2KyTrd
xBjyAllBbpdi7abDe/VZ6i/4fUirKjhCtdHgJNvaGMpnz8l1BeblicZ5MzMV0wT9zzVjjIPXzIPb
rrrZkGDk56AmJitE0704/cPGPMbds2ff4VBlHMzkOTAvkO7tiKELgQQpBWBTCXeIhWMYie6Q5qTt
Mkrrqq8XSIR0Ero95VKA5cd1gSwJo9u31pvCZeUlJD05ma/VcNYkK+yua/9xdgRGBk8md0rp5VXJ
3/iDJnind96Q8R+VcnWJFcjctBUWxrKVRQq30AxYg8S+r4ufzM3X2XpP6UwldPA4KScRYvit9ysi
B1Z/BveVWO8sSm0YfWroS6PC/dcQcMFIsRTxOnk0kezkFhhNcyL+zsjUbyH18JFba9MCiN4ynLBs
C4vWezj28vZXmeVJyUfoV7IGVh0JeseMks2FWTdy84BPFxegZMw2NKMdoqe4ylw76knDLFlwzJWP
rkje75DF7l9CjTd2HdA+amubIz/K0gEMzzxhx794rF7PrIj8Ip24/nxC16+7KI+p8oRZRj5KOOSN
B7Jd1K0I5899aGpxkeR99NNHFVvrUd0eXMyD+H1xUvjdlPSI6lWr+lUm6iNRzq5y4/vF2mzKC4wS
YC9ddGJDvSKiA4oJZY6oFhDAFhl4ZVFG4Om48m4nawSZv3bm7gcMTTt7xRpCoi3CxDmR0IOvSisG
bMz2bS7UzDiAEcF5jULTWBwSUigzzukJ5z4BDstpGqS+UXlQ8ewoGNPGi/elAE3xmzG4zVOVguKx
VCL1QVZ5ResxONgRqTEuzVrExsiy2O397xJbed4exiA9kJkyB/r9j0vLqEYjR5V7M3gykPDV1UP9
St9IaRNGcqrw5SdcCq6tA2vgp3dYZIPMjTgoXPdCA4q5ZmdNn28M2sXLdlTJHX2FGhweAnpF/NIA
64lUTMbSlk55GHa6wZ/7dcbTSWTIPn31BtZpcY28covOiXwF0o7XpicqSxhJbx20JzjXi2Bu/lQb
g1T0lpnzOw5ZZv2jWp+/ui1HNlQO7awejYujtzsOf9FPv5x+zmGn6LDPPLIzwL71ftB6iTcNfun1
eY1qt4TRRAOzsnqkyCLne05IRz5L7ufYOgOn71Pc2lJgb444Lgyk8Ka3GgmK2hTIGHX159bv5mdR
l4kPAQieswNw7HaiBW0ADLTbtYotS+Tv8cK34s+6lSq0udb+XLTbKmTGUEroN7sfNxcgnsArF/aS
GdlacE2GzzXaE74fctSgYnKL0NDDE7+kPkKAIyYYc0+vQ2GXHfpQ/iyVV3IndZ0qxz1Zd81Vq5kd
In890oGLNNJM2BV7tVOczErrCQXnJ8knadaqCAJCO0F3x/XwtLkkAd4LqJJsbg1FYSoRhp2hm3Bi
5KD1wvyiFEIi+aC77GO/l2UQE6nWT3u7NTz6unPjGG7zPrJdEVd0W62c70vRbspEixgi1LOHmY52
AUh0nd57koxanpzdtbtED6DCkYDLprRTwxjNvvQa5p1zw2kYy9VIVmdpoePbUaQ9XIcltvh5b3ws
2FZF9NP+QPz7lZnRq+dZnfEe57xkFNvN3tKIQHHFt/dmXZKUCS5UlDhv2/MlQt1fJqwwQo5tYlWN
Ovwbbhx2kBOaiQARTcp4vHiVfOLhNlgv6Dw80DpYd+EpvNOhu/yEvdDbgXRSS3k3PsInUeETrCd2
LLck+On4/wiI2QQbopKLGiuQmfcl0go25ZkE4i7qxPmwiW/C1lBSq3KtQXROFdsqIkBHXBEXZVQF
4o4+30Zq+gVDImd28e1djCbu7bMzepMJk2PSLysnrggEGJaQAVbzvjzgEEBphnZNKyQA+6ZHOMRJ
nItV06ILZiMz1p4f6AaARV8uPWRFrWhqQtCANx+Qtu0J/AZa4o5JDIRfiqFbl7LjvqFRtb0llt6Y
gjE5S67etikCTUvZEF5Z1L4xQC7h2KsFZD/FBJuGrmoOFToWMht1q5R5LJdJMGcfA7+inFllwgwP
DG7f6f+YgN71Qxlk+K+nR4BOdvbRthB5o+RVI32Oa6xqJfE9D7lweuCosMF2L/JDH2THX42l35jv
Vr0cHGyu3zpurBKvvYs2eQ+CN8PT5FFultw6CnbgRxWYosqcedf56Thf0RfatyI2wjDJLGu3XHUL
3Zxi3T4UUYS5z7TfaA0kYmuoapthRMggAB/fNs4XQ7x0TxiDHQCSqQTRmidOcY8B0hXR1xg7AW4y
U4w9i7l0mngu0bn2G2UFBXmJFZNcjIQgVrGiizlaOj0Uvwaz5hk4k9HH1A8cpBa+O+wnSuvcjqrE
ghIFiZslSAMJFQ8/E9VKI39vo+NQqbFvYkeZ9Zlf70iP7nXRuKY91pkiKTD3js5ZbUH8A7F0tnBL
lXo2lTpUJm9fEb1VsZn5e/d6HpllShx+lQfx9wn4AYUriz3yurUJ+rSBAqvdjS8BJyQOkveNWGcv
T+BFaFOoGD9rAakbChUe17XLNH4hxjhOu5XXn8olGBF8V7ugJVz62tCZ+4mYMXzfnboGjW+HAs2F
8DPtRbhly11PC6SdrxzGeMy43bcEhO7ihr0XgVwQuBsGmpwjdC1budFWd6M3Kug4D5sHczxmiFEF
mti0PwzVlhBsUQMLt5665IkQc4KJW7i9qsBzoreUtlPpzgtABOGqk8bz3v+3ZJyMH9TVGD0P7L5Q
W+dmsJXHTWqFNqZP8hDyCVAP9A6cl3dvE+4uL6agJwJHi37RrdmXPJGKIH2kW5b8RB+hOv93IUDa
bgYrN51Oyy8orjT0LaY3Z80kri6zCHFFQTMT9S5X13MA1PNS23zbbTBmwzI6kLfJNKvGPLVM+uiO
DXXP0UONACIg+yped4ToaujCgYgKk+pDgHXM9HoxW6XuWlZZW8tVD34C3C0BJ2EJhvmAijrLs1Ci
rF01TRmjwWjUoMsPN6L2yIBCOFhWr8JRv/sCXJsMcfxA1j+D4Ixg0RjuTP36fNi6DdghZnUyAqss
gSWoJtq3J8iu+u3fSAh7rapoOGu3lIfS7yNs5yjdUfKHHVXv2iIjYpgMrTupmR5mIFQdMa0MrtED
2Y0utL713N27cDUZwdMWCvLg49SPb6P0OadB8ffm0qtWgP3XnPScUoWITRPaE5QXTVwFwAw52G2k
38CwvqhzNVaLO4Yo6SilbPX7FmrhVurfVHS8sfO+o/tocI+QBtSBEkV2lF4x+45eAkvefwHKZXCp
0IDRZ/r0hxOf9S1hlhNrbvWzOi/YI5T+cIsyTC6eMK3NRbyZ1JICX5+jvJ+CaWvCILxIe61HBdE2
11EhnGzrHgQJVkImBtDu6qeHQS3fqp2PC1J4p7Og3jPJlOSxk1dVNyCEXIZ5Hm4M8FXNI71x0Luk
UjvISnpt9CVAhsjvbTUABcECByfK1DQ8RavB8KD2krCdPouEYE6Uc9Z4rwJevFR1L6cv7FgcxZIN
xU0NXIR2CyCc+WzI6+IuXwHobaa1DWhc6hQ5uXQEtuEv9xvTp9GkZ0+Z+M8BDdHmWIoSaWHcHhHO
VcINodWPQvxitrVG35d5vpye70B/INbMmYhA5DGKvifPjaJGfFodBOY4oBeqMTt/iHlEntuw7zHx
oFHoYycDv7f85dNCnIxC211v9TiLAqiT4DCzmU6/E5is+P+vCzq6f+oZrwO8iZyCrQtj5gud5rG5
FAAsmXr0EV7j0zu8l/7Iz6UTufi4UY8UGUYCXW5IuqbMCDsc/ybFy4x/HaS0vzm7mPJEzqpm4su5
7H2tb37paOeqnQp4B1y6ube4z4inxWw16vSG8FBPP4OVE3Iw1gGAZgg7zFWbX6Er8ymk+QwXd2BC
JTTR9E/9z3X2SVOStLMccAOSLXROJWa2qZ4aI3eSQHKvQf0XnL8hjGegCzi6KtWzPMjjdh3Zhyxf
dr1Ega1+S9JaIbuLKcUZOx8VBnprdMIC/P5mKMa+5zL7qJhF8gYI8Ht+hsi7CeogcyTPnChniXBZ
s5Fy5+Ro2hAwjVHkvZg75SVg4BSLmzzf70XXliTovF3Zs5Lf1tzDbsndsv9de9plDdzIn+CStVB7
Gax80LvURfeqNtByzw/qMnxCbiXdrsfhhOeeVpc9wm5v8ZWdQEsfQcdyNAY+aOgVoeTCNrh6ypKe
4ibTM1N7OCfa1ceadPXrCrTzwExf1Ta2lsjCiDa4VYgNn/MX8iNlTasOBPFzn244GQxKtgfswyoM
OPEZeLDiR/xJYXSeMSb0tW8bmL/B+OuPkooo0+HpUh/pOsKpJAfECY2PmHb2uQc8wVifT7z+Cpc1
6l3yQyJENa9N7hsv19ImqYvcnDY4VUYJtqKD46bEGRY5GRdtbIdaAA8oeORDT32kdwuT+/r4td/5
L6Oisa0ooCzfr24A2tursUGRbnKUiaPLxCGrW2+2OO0Ms29HD4vk2Z2gJDTk/XG+xg2s3ZxT4SKs
eTF1RyVcQutmwAaZRNa3wSDsuRBAqdoG4VbcB9STZGERfH24YmdF7IYQBZNgtxa2IzKh2yzybWWL
xSqceVdUFnPWQIM61wEYF6PVapBRJmHsl5ndE0V8+VKD83fOYzcuJf7QtKxLglXgJLF6eB5W8+jM
YE8bZ6VW2J6GxFm5SKHse+Ng9wZpxvy/2m8bvIwARJmoH6/cU37Yngqp5h1ub5zz8oeQSV88bVpw
/FbmwneNgQJr6+nM5MdMfYxeJ/oEtQTIdSiWK+jU3GVus4eD3x5veMCo5OOfpzy7B39/s/o+IVBw
QjYwGsajvKRsspsYYhVRymFFistxqCRyf9D+Dx2mKgw01VeeNtXtoaKSKeV+BRYuzFXyP9gVoLTR
ggJY5F53u5a7dGVsqVxKju0oPozAQkHsf3cR8gooOrnPE2f+NMEskn+sb8SGYPhV+9RG1bCY0nyd
RCMLTr7HJbvAZiapbbQBHfpeKxCNJH8qWAXgD0xz8e6wJZ960I5eP4WREGBh/lZFTwKfE0pFAeKM
/xNbBdaIRjm1F/qsSfKv5OKY2M8/KwjQ+tmR896s9+e5ARMEBtqAY7D7aeIKt8tiI5mRCJPuO/Ag
AhYHHmIcdf51+nLE2k6TBbSdkXWOwRdc4wvnxQm8T9LlnYx1EAxIRmcxvhSBNCD3/SE5T+yJBT6U
swXUjIskeMyoauxOK+Q8dv+J0L8208FqhUdzsK+hV509v9pwgwDZg9P8388Jtwn5QlHR+7Ta4asG
3IudU9uIw12De7RmmRNR3WlWC7FZPai/7vM8jRpdeDGk4KzwavqTqoHAfseVYG2w8Y2LXyrGTngJ
/uRKOtAwQPPOoCLWJPCILMibjNrTitT4rgR6egM6bQWVuyIBi0S3lbo7Vs1OY6BUxn47/5SzC9f7
TYC/2hmzBuYfkfyvC8Wd5yAIuB2nTmRZqkxfj7J1oENdjGlLJHkmD5XaEtQBBPVnSnpyAP8Q7rJY
lcEkBMYtr5Il8a7CB2TthCdJHpz2Xw0m9dAtujibs61iRlJq96LabPk86Y2CBOyvekyX8hyg3lPl
2htb0ZOs3SJQDrrqSyCjsc0TvPglSWU1zHrdUbAYoMWj/zoVb3sZW12SQKe8bjAi1w+nsaDA+FNR
k7J3veHFA0qvuhvKc2fviFeyAYF30p+TtCh9zzTPsUsPvPtwRYEPUlyb7iHdCnzod5m6xBAXazlm
Fa8/KTZ/xyemKPDEv8JSHBj5rDLfXViVhyu/jiTG55zDdBReth5lJOHMm0g7M9hYHxAWjhFnvFDm
v5+aDOFJzY/t6SIBs2kRD130dSamVcXqZEkX6BABs3n0a+W3aSrCT8+bZP/2Ml7XxETJNsRYZhxk
4xJ7vQ0XHqVPQlXCNkS6XnJ3EKF7Sybh6i4K7obqpzGb/L7n1eTgT6XxJN4RLas8si/fJ+CzkyMF
gV1EE79kG+DVkI9ENEC9mVqqoHWodaGR1fOOjpi7/0ZVdT5/QadH0wZ3oR/75K1JC/wDNQa1LBUG
YPismb5D41NeaKeipBEydbyrL2GS3WzqrajemAC1/+mWTduMt3OdYF0NhaRIyaZIXM4QD9agcgEk
A/ujmtet+UxbwxRGd7tZ/WGoyeqI/PCkk2qVrXkJEIFNPIpkRZEm6hw7nNtMsjnmbzRf52kUTk0E
70+TgAnepeTCgwM1B9rVkxebQnsO1XorkqLvlfhPOQiRjD4VMwOc55CtLcN/1Kg4vEiCe/Zcnry4
ATfGuOfpiS2otzo9v3rxjYZfBb5UYN86joho6GczqBXibvnOqakCRQvKRvbeqrQJCGZsthSeo+zd
PQVGgWd1gDEJPIM90Qy6E8DJ0EUVO9tzkcnVUeHxPHXerxQkGUYUoECqn0qM0HLgR28V1h7SF6e5
Gm/W8ZDQ1r+ixoSTUzyNI0YjWVQQuehyAFo8X+EbeZ3vKX4P85sJ5FbWXDgYX+kMOydwlaMQljzk
tvWWBLG90xfcvmZbYGeeoJOj8RlMDBNnn12jW3BtGCnijBXzb1SG3fqtn6Tn9da40lUhqQ54DyZo
9GtmIn1WWxsrZpoJAvXTJQL7l6AUiDafHOL9GlrMRl0+XOT/huL9XTP45M4fof2fvanh9TGYd3Zk
nK+wsPMWeuK+Z/S8aR92Xaf+Y+mVwic4ynz1hDSulxwzNk1iENolvaU849EKdiw0G20nej5WANnY
+oj1qzDjQUpQ8Fv+g/+Xjexog8jc8139jaUJy+AwiK/xvXb6kN00GBHy27emBokuM+OUfrPbuovy
65JcFXUFzFUT6T4miqyPs4JMhPoSDDqAh/J18z3X65lqHhuUtMDVrXcpFhOvx4g8d1XgqjNOjaoe
5lEQkUufg/zGrg9XDOnbQknYw79ea0RB47Ebl5m6RSUbA4lxv+zkPgGoXO4yZRTbQWMFY4u+mVbB
rIJnJy3ch3jee7WJrEN70lXXhM+h1Tm3Yowq0B/o3YcB6e776pXFQ4We73P20Rh+GK1WfzY9A++/
Limo+3sLLOWCzNvUb9wpG5KSdAEPx/Y5CxN9yzNKTJo+2vzKMu19kJqI2Qc/W2dEdMTKt6mGe41N
EppVORtuQgDuTOPiSEdt2wgRhZGa7XT3FBKsh61qoGPpGCRDUtgnH619EmGR6f0XBNOMOyjcI3bK
DEXyoXC5QIzPZtjICInBV7LF5ymMgvu8WYM0ZWv7u94mwju3lZssf5c1tm1UtDL4AEuod+GI2hey
JjxAWNjVW2/1J+ETxeARsFG52KmUjji0lopOX54b0mgDM8lk0xhWDb+JPxM3E1rv2TapOCkP3z8C
YLZYk9jiF+aptA+3UJkO94XKzRCr1hr7RyRrY91tmzLM9WxBP0zdjj8VsOc9jbdEvUl98hnMnGCx
yEEWUtGXs6NEhAFoD+6b7HihRB46dp19bqj0Q4o+lNQa8pBcw3FMABm3mPOm5o1Dapdr2BpsR1c5
UGyOyHxeOPZinsb3285Fhwe9i8cmEVkG80gILY0YifQwYa6SzxGR6dxQKe2yomV61ImLmpoV8GEa
Acy0wn4cFIX2G2rX6vOVBIYs+c11nCN3iEvtNtxyqm7pQNeRehsX3A41EpW0WmpmNb4al0wY1AXv
TQTEyvDB/8GVdWDMEbJ4oPA+xaOATlABMNNF7mq5U8gBkUFBeuYipIu59QeSs81b1AcVPnMMF4kU
1kH7fkWz8UP5YQ83+wa3BjpaqfXg5HOA1ek0rR++Acylih1M8xexry+8znqvc1gRQbrKzejuPsQ6
rtYPSVZHu3ticmbGiC7QCWh7QE3nUm0MVf1vJ9Jq21+e1wwiGdgaDNiPnjBO1/EAPJC0NWeLQQg3
Oh3a2dmR6cDrYUlCwSSvMtF28jteTH4eNEXo8bTurZesctbydAVhOsAqOxnGoGiLmW269iWatOrj
duf0noLimNd4h8+X1j5GUBKk9dEVvqpmDjmFY+L4SaYUVAdVw9niQWuyelGp+4HSmQywMiBvZ+uJ
JzySzIA2tl7Op8Z0IpocPUI90ttbK+tepJr8jxTKLYk2HmTzXAFNQKr7thKJM2v9LNgDJ0QAhpp2
M0CJavUowte4Zf8uzolUsvIxuCuVXs8sy85hFNBL7xR+ne3FVBTpbIfmUQxLJWZhnKqDDTVcvE0l
P0urL8GYxptFWF+h/HSPh5nfcnvs3oK0o362ICBTkM6A1a2TBhh9LbHd+ZmfjDcTTFDP+EClGMaR
iVkUonWHKqRWj1sBgTnfqbf+yT62w6qVL5yuB6aEZTNhFjOFrNan3yBmnGRCH658t4OSyUb0OlgF
oUCPmSHM6fHqDu1Ypx/JjDnni09CAqmfRGkqVpNwgzDL3xkPUspj3qPVjasoqDnDWVl/sa2yoIMP
xOHttMLko2mfgxfvzxgKfOAHWD5XAO69myVzRuyt2XvawGd9InPZVMDV+KobBx2IZrQGZhOTMkDh
Rba9xdftsUyEwWsqNXnqqKZSTXYMFtdh2Lo4T7eYFyJBYnxCwlFUI2ielNOeWSJBJbQrkPcXl81G
koShxEAQ9rMIrQfdYWDDQ5Pc1BKLrHNpCC7kbzwsK4fy5vuyiI/hCU5OBgbzaSDQHRtXx0HJtxm9
W1GQ2HEJ8r8J/ymjfCvGQNpQ6nlR8jahLY9FW62JCzlaJ2wA2oFfueJo9FX0ovGOY/9AzivXfwq5
8qCKCy5+ikwr+N2i4QGzO0iC8Yl+kupFN4y62eQPJtvoZfVX0JUuQujMcUv9QnFN+JWqStBXO7rA
9cbTjZ0J82aSbBa1cQ/oHELCoSDDrQxZn9/fDaaOvCbm2S1tJfHVsvjh3mhFgRMs5O9NW7/0ON4Q
x1+H+km8GTkdr2L4CqJnoqLbRNQMLT04fuW1jaHYhozJasUqxZk2hQxfusSXj42E+f7mxtCWTDfs
8EeCeIDrKkck4hGpu7v/fO1cReYkhNWqotHL5O6wLZOrmRCJSGNt67zRPU1/JQRg1f8f4/Mu8Ma7
6UlZX9jXFUBqOuL/SmiHonUwnjFDFD5nKuVhgPVsDX3OClwiaocnPVx467BPwI3rS7j77z3nY0ha
Bs14juYxWFeZp8CAtpAc7v01XJ1xQSaqeAjc6U9n7sMwUWcPuPj6/Mw7fzZ2wRaHu+u0XGHpsKed
6/VE5VqJNOKtG/etWi9rbVRljDwq+Zxg7lQRiUooeBEsux3agtslVtZxyNfX+CNUSvlXiE5I4J0J
COhW0X2vhLGGW4RbN0yh6RKr+s7dlA0mCHDn5KUeRvGMnyjlxIBchkO3eENHglbBvO5y0so6r7HI
nPxu29QliDrJ9jBVDgsWI+cEXiV670D/dzBZJsNylr5YrW37w8a7HEUPGJW4sxC3xDWHg1iJ9iZe
/z2B1qaYjjyjszwxGT25wg3cglYneOqLuI+PeO4ZApe6Xx3f46Xk/DfgaIx2LO6fpQfFBqZGbq/n
/Lv4kRHuJ+JQKBzXeEAK+BvU4Ery3DkETQmPYEAV1lNc6mx0quzSQ+LidHP3hlK2bQxnaiie9tkM
N77PT3tZesS+5yjU0ETqzoaiEjYNgCJ3wOl0WGu5+LFWZR3ctMofAeQTGKBqK2yZFj/L8wx69wSD
PFcDascezUIWPMjHpUWVZ8cUrlwdcrht4hFgpXI1jnlihcLZczmh/oVBUn5N8t8H9Wf+TS6ApaJs
3fKJida+OIFWm23e2VJ1hl20tOWCseX15t6xUeUYYxg/rAcpPRfe5ysmY9+EzrI5Asj29VqOHm8y
a6bLK69Kd0m4FEoeIhWjITG1b09Vpu0MCfbyEEbWLGD1hQpWp02xEpMUg+KPXJGv/nnV/ncJAmRu
Uvv3cGQxzdpFawQbQSFOvzInaq9/dOYpmDtis7t5QeKZkP3jx87bU8TG6C4LmolZDWKSvVhRTwFV
+OSMIb38SJjmwb4GhczD7mj/ydlUda0Ol5PLr90KmMBEPKFghMLYrK90xJg1Pr2VQqS0zNMKYnTF
VXUff6nFvkFQWXg9fGfXTxCD/bQ0WiJPh1gSVZK+4+B0eBVu5oTFp//M7xZiW+L1ikfRr4M1L+0b
Fb6kOj+lq9/Ol5BVaJwqtdM6dSH3h4REqvgiqhOlkI7kBL8/rHd6hSTpC/tzVeqhAKaKBAjQp9CA
A0tZ3WiKIS5TDb2U+apziLs7RdheUgNLmbk8WECMgCqup0N5QnmhVdaG7dJZ5SxTjskF9fEN7wvF
spItvzaVYq0BUSGhO4SdTL5jFOLI7q67C+DIhLncDDfNhUpkpbwr1f+dHt3zkaRv2PKrb7aVaHhF
3mgU0z3i0JIA8OW8HgnBU4gIbKrfGE3pu5W3n+aQb1Ma/XUoWu1L2rxnUILvnLq/kU4VxjXqUbEd
x7bcMqWpxlhLUZjpzGa5h5fiTKVHLQfGqpf55NMT+sJa91Xdqf7SSWOrm/qDCX7BsLZvQD4CMYUJ
LH7gaJiUlG6Oy0GihG6z0t/qdDbLkDsRSpZDWXnNFHnYcdahO/qmuZDmKUs6MnQZaoxgIyiqweTO
mVuRgBO1GuWW7u6VQfbtZi6kRnlMUPrMPvPo8YXSPf25njwJyFpIWuFsj+mPUBH6JfF7+pourFlx
4T1O79UUciMwW3G574yzhqpmS35S4GcelIhw/dfRtEsJDLCRz6G3wYgqQ94UNViqEENsGjD9bnow
rmL/B8z4ROnasyzVKCONcD5RwY7skKfNyXkHVUA1QMC0RAAhBJF4JYfAJzUeFFObxRXZm6U4o7OK
1JPbg+mk3J//BJRTgpNggvIhBOYCZfde3r9/N8aoqYFxawd4dN8CUMIDdZPSS4pG/ZknuWVhrDEQ
NwPMmIgzurOGavhiEyHhXWGhIZKoDhrxehFOpp6vHMQ4pv9yMOZlwOwuIaG+4HDSVM10IXK3lwZL
AoRIj0+tccgi6GygIQfeMgX82qrFZs/OLO6I7VIP4ZV0SO9+jhFse6EnRHTP4TjQyOWzKS2afNDB
mmOBF+I4Q506Y3GLK+mSMOqZSpbLqxRanFFu4+kFW4oeuZioMdublGqZtUzHhIypn2EjbdwyW5oi
4JpIsbqhNsUhtXOklVWltTlijUGd6jgZjnveNYZjXvQyCtgmnRufHx7dffAboomywHwWhM3ZYcLu
bPCTHNG1tOuN7G18LweG2pKpGUfl/9xOvVKyX5iXQ3yeFapnjsfz5HQhFd5nzcen+YaQI4qe2QhW
P1IgGadjnxIMDJocYG+REowQMmV9CbLw3trP5dyfD4XIfjPIaaKaVgsFkAlJTAhb2fB5AZ9m0lCn
Vg2g/fm1Ca6Hhrc/uWz9trBEVz3WZZguGdEjv+xni8w684gVUg+Lxh4uuPEJq8R2rqAzr3FFQtsd
Vrf2t4CGJ/TSaEzVdc2cIgJ6wkrdTqBmbXaes+Zp7bRSrn1yPh1CyC6W6eV/ilTbDZVw6WIV8vRT
s5W28SeN9PiLgeWoYyyfNYhP/uVPCTRsvgkDqII/qzrdYhaF81LJEVBcUdZ8PvTOthTf47zFigIM
Fab7MzJ7UGCFKQg6xS1uMG0GGTnnBFqBsRTNvP2m+sK9Y5VKMlOUsGuxjzqGS+eV1JNcMREsdrpx
Lrrkh3PYIyHs7UaF87m8rk1/GSGhbBS2Lx/ATDdOmaQVm8jalLQuio9PIWGHIiD0a+fWr1II1kxS
KKYseciy12GC6y6Y7Cl/wsWl0EglTYklJrCVS8IeTz0GQOmkR3mIxfScZT0fdEc9m5zWqQqSn3n5
ChgZEpwBOxUE9usENLw3XrdIy4xAT7q5GDgX4d3qTBNGD+npT3pt0J8d17KngQO/bHnTW7Bd6qjw
PiL5AXw9yQNCc7ipzc75/PLiP6WxvvdxJbsKa9R9TLeTtgUe0/WdDrL9+mvt+4w4RXWsIDRmm+CH
M/E/AdGZXYOjLD74sVXRj59DtlhUBq+FGaKG9vDSDfj2e3LSCStYTweWZeLzwbJh/W1P9jLm9cBu
MMLk7w8Nu6CZhP2Wa+CfR1SzdtN7mKaa04e9/rHyZzwrFcQsoDUWcnmrGDfJFNjE9Gdnl4/qcM8H
SSAyEd1pA0Iaenex8hvJq1gAiBTzCeLWkSBjBjDniRl2laaxL3+Tt0bAKwAjR24rKedk3OWCLjG2
zWyi4e4bkkYQuMYiCz0RVhzs0cn699VaomWNWY3tWzpjObEgAQoAdgYx8tfG4PVMB7kgQpr1vw9B
NzuZHAy+Q5mVAQRgfQN69pCqa/9ekW2LggwAkukP2rUxmU+Hn5jycqUtLAYH/n8c+noybXD2WCJb
Hs703QFW/T+Az8jvQn+Twwikm4XfnaWrco3vQvJ025sry8AkOc9ANddDYMdcpKlBOxBE+uxwur6U
rxjhzkZNqPLNQ7ftzwKCFPHs5BRueSzAkCw8BXQ2yioR6CSxvCC3TL68wLFJAfTP+3Q/CBFYVOLF
6OUwwlocr8HLPWVQmTYOBfRzGJ5PEMZnf8Se6qDS7uAQ9ZiGxxPA1MJHBLMaxMhKn1/IqdZinzrD
y9XB3H+yTk8ZapSwmimu+SPTDd44A4St9twlegR66n74sVLPnkIeiZpWSnvEWyeNUri+Sf4ItEZ9
lvahRAZq4tmPpNZWd1k3kzt2B9WxwTXrS/xDjAmDpfXaGYTZf+HlYOep6JhQevTT6W8XHe+vDXyb
psi4bUyH+lFSPgJLaOKxV7/xZ5jhpQH2U4VLivwBqWr4ujZ+s6tiQ3I8msN6fl6gM/OKKYiIFmqk
NGaNPLdr/1dBdFbztbTMUIppRXhRlyiFKGl60hu0KvYR0vjTdCGtbI8/2WEhlaYSWFqdldv0obGz
xjvzMN9qnnIXSJcMZ7ugd9u1h0Ei9fuM/53Pe61KgHayoJCGBml7B1G7ZlrJOFbjy1e02cq/k8CF
9vxDTJ4KMMYajCh6sjb+c0yP8VymJXyJtPaFruBkxHVCE4Uq0qdazVI4xHXcZ8Ze+0hJ7OMJKfeT
MZbLIqFFPHVd+vR4+A4kWLeYjFPBS2atOu+t6WToxepZ9/cElxkL6UcX5jHwCdbuWi9HyRSIOMsA
BdaeXmkSP+JhYIdsd/Tcf0Es6fQnqT+EB0FoSY0+5xAJjFdf1nvxpTZaqZsUriTLTzLTwfNjKgs1
Pn0no3pQqxp8NWVBPPFN+264bflVx63/Xo2wfT/RH8dhAMi5Bzic/3VdhBs28y3H9D//E9oGclYW
HKUL6mXz7lXJOr1r6bRdd95wBI9e+PRUesihmJKM64MfPv2HvDULs/tdbalR0Ou4ZjPxuR6pMDAo
4Z3KKxGmLikBgE3pWJOE0LZ/bD8IJoMBf9213MyfE2vm41AlAD+BJGrC6KHYF+kNmLT8Np18aHpc
SoIDB7dUVS0jwtHgVRk+1M8CJnYhKbT2p3TFw1l6WQlUIHzMu3slmOxL16IgKG93gp4/JDFwdMo4
s/v64yRg/MwmnJHa7ze7Y4mfWJez+VryAuetjP5BNuNGDzV35Xhq4u7eL8UpK8G1g1vDO3uFcMFy
m3DCpNLmBKdKkRffIDq9haQGv4i1Ogfd5A9RPDJjd9xhABaC9pS1orExPsODzYf6TqVTq7tmjs6w
I37GmY7Mn++HZJZGIj/2unxdhshzJmRXp97815T82A8eLQmrgbrkjN4j+vMYAiKAoNYU3/8tPt62
85I2HXEepfns1G29F+wIVGz3TOFqeN/WeGSKhlAYMOPpEhozk7rrT7lyVmZiSW7vY+iMGG7TEVXN
uh1mzxKk7YkHPxaaUmSGBQ9u1WbEDls88MNnC+JaN0y2Nx7Nhsf3QuHZF3sleiuonk3YlblfHw5X
DvjAoI3o5ECYoYSWb3hRNN5CG7xRf/QuH0wgdUeaGsrkXHD3hrdA58F6gC/BNb2Y3VoC+Z0eTlbN
ozEsd4zUhP0ZVHa+NXZrYs38roqPrVTwBnkKPPbMeqSN1PUsGAcrSzaaodg04Uwwp8YiTp5zlva3
Bn5MNKj80Jmna1hMrjyMyZcwauy/UiqzXQaRpsBD0kFUw/pVNIbLbbQdQ5NbL1MOEnUUhawb+sQ3
rXWUdegBVE1JkTM5f9EotLbgTEaJSJLm7pXXozuPuv6+gOal4vZUO5RY01L8FRRpY9vXshnyLes4
Lz37Ms//nnkVP9jQ0SMeAZS2aCkY4ZlE0Pt+MiFpBaxo5RD6Lvku2aBJQ1a6Ij9HxUGnEt2Z5klf
gJXIt14UXrnAKd8W+5QDkCeGflJbCzwEbwra8X6qaGK8zFL48OyVul/7mzCMVmuAmHxXrpv2H7JP
Litl4582Jsh0tlym0mMAEM+4r21n3ojODoV0augFVqNpoOByxkAQJ/gsca1TnPmP49OA+/AxK2se
pyuNzVjR89qPRakLeonZPnypnfHyGrNNNj0OvXm44uYKzpqMg1+ZzbQXTJX94BouOexjLlm99Fax
UfxEviy4Lcry2enIyvrUzp7zvw0CPa2GwhmonEwDbtKffb25DQVh6IEjl0js69MbkmKnkRq/Wnwf
KjeZ6w7tHSbbLKqtXfe6umvFBaC3PqC6TGSy7fXAT/5l2r6n90EOlMDNoGBlb07OxAmT0KQxGV+I
gY+ufRKyEOcQDiSWjgaouLatUs3uBt+SZZMePJFREtWR/5SLVLaci9hW7qd1b9p1fjBFM3TIpnKc
Zff8vNnx03JxFPB+ZYD6z9OpDihOHT3O0tw2f0jkodlrMZoxqcJzrfnXXjL5pDhMOJukFtqRaSHg
ee+SwTJOj3hWTQwqkeT0Q+uv8SetTPumNfRjdnajzlZDklxpxxFcKoEezIehq/sHvyGru6Jvvpxt
XtqbmiBY+eg5HN1iQJ+E9Y3z6mkFLoQDWZJmcjtQVVwyiB0pJY6U0uKSi9yd2v4oyHmzWZNLd65z
GpojzZODXaGeOZj6AGh8xij6ynfB8NMUS/Qto47kGmG+rEuPXEqmweMKG208HPPZlOg1qJn6/5xK
GAwiMR0t4v9+9c8/IXmy7SzfRqP9KZbnLDmkMOT3ScR3dbLnrdBlOq+32WknMwP+OIGC1FUmvd9B
ZaPq002DGCSVH/rJ3X1KP99WnplUmpeBzQIT/flikFfq8RSIN2NPh9+sBAkrGYU+bQC0xZcdQJZq
wmr+XTABp5ihO6B06jOw2Q7pZYl3KF/RQOfnoCgZqJ+2CRHK5twb44nYv/ZFRhjswZpSaHxE7VQi
9gMj/hkj8CwTwDGkH4XzEiSC04MJJ5XhEk2Rw8xkdEAqFeXKqcVFHWXNsdpNdGNWQqCq7rzhAbqR
pa/OLjdNmleuH3oxTOR4NzTKua1Z4cEYz2sy21BOds3CAnUrz/ZnDp7ObhQbxBUwGq9SoH7dPXTr
RIarQZ1TKJAApdd4sXm+WkEEss0Le+Uv8FSBNWRxptXY8fUpKmtehUZo7loKVZvj069MhA3zwfx8
G1OGi5qiKlmVAWKhVuvSsN3XK+ul4QszffwUr31CWy7XMdp1EuM5j9DS4GOtPk57xMBKRENEKFPB
5neqV5sZjoOojsZJ9fkg9tKw/necK0KxeOl8w8SbUUOy0CFS1KaPxmAkmv/bcOmzf+n1KtBUMn1D
ZBr9pZQaTcMpZYaI+gK3OL8+1jEU7aO5W319X5fcyCZH5RqDfeiD7SueyxoYISFurD7oBdHA7h0G
s/kgS9tOTnjaH6Cc2Xe6+JtdiORr5bw497ke6E8HEZfZUIXvh3vJx0LvEEane1lBGxhTD3ostiZC
iL9elsD2rCM8MXCooF2MpFxIkY7P/FtEgws3QmupCCRAIOCh+qUgmHcQRnHhJ3k65c1Ku/4FMTQk
xoRFxKcHI765R6nIuxUZaPKAspQKBl2hW7LuUVFxeMFzmdn6Aw6BYJIz4fMc/81IE7/5YMqKmzT6
MfkOjdIsKss7m8/KtcbySWQ7JsylcE5+aEfepeVpZM3wkWtgG/PdIFkaRZZ6Js55OtPdCznhkObY
XhQMymFaCsbuIt05dHv7CUAVxvVPivdMJGdvbLsN+I8L2Hha6xjfiahvAmULKjGt+1xjmCLnIr59
ykXxwO/6+GUnvZjDPb6yTUia5pq4MuQcqca8V/cB8K7DOQbmLhsAzmYkycTNe4pqssE4fKIGiGZX
OSEE3MIexY8xGrH1PTJ66iYYYs/R6Lhl9CGs9f57zTu2U04WwTyvWqhxMGP8UARuC0zoELRXBmtz
gbpyfwZZNfQcODJlKLBlJ+1lmyRMZLwpFXQ6s2VDoBjDEk2bHkikDkMFmytY1o0wuxBt3Mja8lg+
gWph5gILnQ63Ho+qvI4csrpdahG5wEcODPec5Lcchb9QlFWoGY69TkxOCwvs9TmV4gOhrfNz0NOZ
JVBBV9XfjKOPkzy5ojLMVkAfMpBB5tcdeahODWRRNpiJZwqAm4nWV0V9KVTH9rCWvGkcPk1F0/W5
1EwgMEMe06P294rBgvBO71B+blveWPmMKAcRR5A2wHdZju/1/d4oU4LvTWeRsUamZG9pjCnrbqad
32owHhxgW1sZ9l3pZIY0CDnt3osLWnoRbWNjcozuod+FhrL5Ol4So98GwDkCAXqPbxHWWXDxauGY
+4s0shZ2pr6/CMSvh2Mb05RLvDAvq9W7csQ579AS1ue/Hzkf46yf2MFZ8A0uVZsGPK0JOKiIMbPG
diDc9dPDLHk0bP9TiFUNdrIlUl07eZ4Eu+c+EZjJk6t89RrEu31EKHtaWwDz0CEGgAOJCtv9AMvi
6Xl0uvI19NuQEnGlRPgOcfc67j8t9Z9jGNTBV9VUEU4TArVWiTIUSSwW+xmiyaSAqapdnS9J3AKu
jI58KAJvI64h8vEF14qmr+w6juprmZPKxotTcJF0y6Y3A3l3W1EvtKWh9n0aIhQO2+jskztJNP1E
VDz5nMFr3wgP+CgWac1hP62PbZZTqH9XSHrqU8Ss96NsXkmtVth1wd9Bq28KHyICf+gKOcYx8PFf
ySsNOI00ZCLV8+ndrLhrcb8pliUt0oNdsakov6hbyx64EZpwCfJnmnSxsg37k4INL7OB+sBq4pM2
u538byqKTuBFdlpDGkjffLVgelQidTraZNvH0a7uqIEtdFBwXmKknqWgjOAQPIMxwWdplgye2IoR
bAiLZur0KdNYWfnPNPxJpUfQnEyzX9TsM+pQ+kQIhtAE0t1CukIHQL6U3Dks1VmaSq/Y1yiuz6KT
bgNTHiC+g6UIMUms647vKgntDhHhxxY0Hfh3uRsVjgRaUttxcclO5426po5Z4a1JnTzkSalUaVAb
lVUT/49iIdzVANvA6tgCBwjMDYOwo6iTfVH6Spy0668bgcsW/gZB4c0CVNZxuNxa6UkcRNzqzeht
G1BrOzx41vHDd+zmTrdaF0gUJkcgyKlr5Ftg/wtVPTiUWAnQE+/YF7UAyNt6Z93n5yhP8h98pvUU
8c5tuM8/+ZtyNxkAa3nNHUjJXgDnurAuBpU4rtxN7s8sutdTdBck+BezrBkITOGc+g1KXy2unITC
Ter3F40uAF3w2IK2iiGKZqlZzQwSOSfgPyJbd3RadzvYfE1/nLq+ouU7JjqzbBCbaJRl1aXWe1jt
dzn+bZiIcC8WKwIJabygp/iY1OyGaPQdR6LxzX5ABREVGa0MMVYOt4q6xXLhwTTJb5UmOg+Wzicr
/ZvwvUhixAdkROEbTrvy0sT8WceaJIK/fSBG+2CYLUJWqPGB7l114hWl9C5o2aCDs/du51LKqet7
L5vXY+w6s4FosDkU+5QW4taFxOY6ds5rIjh5MG0McsbpCsbI+d6tS2m9RMclt9v4W/a0LaLx/bPv
oJQsv4DIyP5kJPOcaC+MH24qfu04/taGkt0Lwc5EJ2VFN5ulWJha4Y4AsfE71U311e6BTSBHaXKx
rQ4vTC4Sq8Nwd4DPmFMb6S6d/UYtjAkko4KYMSQ9Yiw5FFeBqm80EOwr0eIOHIH4Ct0xFlqd7qFA
lvjSUIsc1l7hJqNiDWBIkcReweL3J3tjfXokuEK1D2zCYPa9A14CBWAFWMW8KnbDuEks0Muc0Ktv
XUdsfG438DfgelXkuE1NW6VDnO2vV7scUWiIlfsRmhJz++NGVFv83o7v/rISMbIxnbEXN20POteH
9oKoQPlliocyBo3s3bfMBBEz73TmVjszwFEHdkmLyJkQ8QbRz1Jrw8iHBc3Q7N5zzyXhkw0ZXucf
88eJFv/bd6bxq6YxDjc2pvPL4V6Av3kVVwAD7R8WaNWQhSGzoGdqwl+F6jj7XsXq8q2AAV5+Nzz+
krYcxlW0UTbJIcN4RxjZzJAw6YCNWf8GQDOPxj4p8TteZOO+qtLN6MwXogVTsKRZU3Hp+k5NRuzM
1Sj8pfncM1rRv2KDlFxOAWR+ZLNpl10alsUsebmq1UCv49flquQfmN9AUPsrXRrMahX8KFUvcbCN
7TD94/qak28+A2XcAnVdJgJOdy6iLSgPNIqgNtiXjM0yGO9v5N0lBBrWp1/FxpKVoaxdOFi6tx/A
axVZ5hIZyCz9o9r9oye/CSA835gkp1ohulNeJrOAFgoBqs2U9YVyQh8P/NHXhlRXWffK3HEN8+B3
+R15NRh/lc4lPSXhIDH9JfzvR42M0i/jf89ILxAkMy8lIGszRSoYVBqdbdS407ON3+m8ljEqEmkP
gokQ69ZW9YxEs6QEYIPM7i2fKNL7s/lKsoOEv4CQma8l5fpx+Lx1d4Z68gPKL2bNDI5gN4cPyhYR
U5aOA0KdrtL1FDHcZqF7KLApWIAef82o5wCi/IBKXiyeKCK6JQbkGUNtQbdyEq610jelGEMFld1m
SLWT9rz7JAMCZIS77GewK4OHuOk12sHEh5UxIYZXc22zEcaP3t88kwLnMLnd1Xwjnlzu8Z3/OqA+
6dE6Mhv1ptzXpJdikMXHaAFp4rzl3ZXV8a1dimwW596iTTq6x0Z+cw7wbSLefeIWbneL8lJC906n
+uG6Y2/bTZql8z/rFJ7wlg9jhze5QuvwgkGjigXqJp/9FWsKkzf46HTOqZlHK4GHeRFHiHcBbH4d
yodQp8CNoLm3c9pak75cTud/JmKRE10H576XPV69uu7jT+YWtXnZQulgrMvkQoAVPGHgxEjNzcun
r68fE5V7fpGa4xo1I/w72uFFiVHE6UxOhMbPiP9Wuqnaz1wnZSbZZBINGO6N9i6tQJm238RjANIE
Noe+mg/A9xrkkcj75h4KbahED9AptxDgyR6Zz3razXZrklvBTTxE7QDmx0Guqb9n/fmZAiRHtSwy
jOW8OQ3URff6t2MOOsgSLrHPAYRF8fZlkXNVWUk4/t3yo1zG35HSMd7SID2HpNyprpuKTR04bYsN
eiFpNTrGUdPOKxysHJblb8JNJEJkBUKdfiMCGCeOf/sbmyOdawXt3sIVC/1WqZIaPTrkmL5zrrjY
aRwTemx/lMFZjD2iH4ugnRtfIkWBVOr1K9t/mVSYZ4wsFDGMY6kOhYw+YC2DOl0YRW3XzHUmKhaY
lHJYBR4PeWWfMdzKYyMbjGvjBTi8qhzqYG3vRpNxUuHa6B9ALAR0EH676RvVws8mQMNG6g9GEprh
Xtse23XuNcCqzsu2o83dbJZP1b/QGsCsqvSLJ/eyBQIlRJvBhBSLI166q7hR/zcxCIj6+h/b/xgf
7wNZviQMLtOAbgkT/SfAFeTClmq9/eiI0Zpr3CoJ8C4AS8ZHKIvN4bnFnKaFtKShXyJ8sfgREeeW
OXZfD1QZaH1Nf0VgIrl9C+GEM+BrVW/kpznCsueGp9xW6vM+7QzUgzum96rGO6Pn0Rl9gfJce4dP
/4PGhfYbzuq7bZZdPfg7Uvj9nEkPMTe1//Rtwi9yw+B7mvtyFu0Ce/+2CPuGQF3mjxqNPBZRYyP7
mH6fC7jRAB6g6QwSNJMGyqr1nNeCRZYHPsVRkemwA/5Z7uVrCvdsqjRANFaH7H/k10GgBpCJtY7K
jYxCkBSFFcFZQmpDIDBImaSmaByREHw0+dkh4CFA7EbXtg4PD4fxPFraOUg91Dv8Q8o9O6KcOBjb
FaQxX7H3b2mdZPqqfzDcTr1JSedA/7gaWrZYM4T75CBU62c9kgTOj1UxSdNodI+qe09hlmR9SXgM
MWOCH+dKr2FTlyN1sUcY+3LXkxYUt32VyHjvPzNs5Fqc+KjleMwqnsbCGTuv02ScZtduXBhShh1v
e8fHCMNZ+JQbnXVGQj8bwNUTQr8b/u55UQexPgNnlwnsrLQ1ZaVQD/w5uQfsyGF0QIJB87XUEPNY
xIiNUo0CtZYcO+OWWIQF35vP/7k8oWVn0amoXitGkVufku6v97Pz0j21hmM5IIMNns8um0Pwkl1y
Sw9z/Ae6q/xOI+NoHglgwkY0Y+c3vahHUs1aKAtFcACUPiGbTE9jl+m7QVgzQJRzScuDFE35UyRk
mJoFcwgxomSBisBhdbCY9agUHqGrZfeqiJeFtpn51EgP9YlxtpyFLMsjwpq3MH2TZEpFiOVKpv7a
91f4RnblPwJag4jR0iJSYdvR+1Kz4KmTdLDPYiFvSAbgMsEsbZIp9eNil1WeJtMdEgqzmrTBLjAx
+yeikGvv/6G21MN1uHJnE4NSV7paU5Kj1ueNPVJ8fA6NS5itPSDADwDI5oMQtb+9kkqmjtSVMccq
bEXTCyguN3rKa6W07zkKXTAvSFy8cwWrtw4kOLZuOk+7F+e1zr/vPgDQmz9gP8pUb8CZJDo5rkMc
Q0Q7S0N0jiWTA7K1Vyi8QkrSuQB/n5z7TPPAGwMB1uz5VKP67kt8r4/bwYJAgDM2ZVnt0dLX71tm
dwqlymBi0LKwHmjpBSvreRipfFrH4UWvYs4X+tGv4WHHqwvKiKOPL8zSfwxf7G9CA2EonF5RTmNx
b3XGuUDNeM79mrqinX5EF2AZ/bgtV4P27b3bUI17/Gn/U++U41TTNxF4RKB/3ppl7rQIlZaNFNyC
4e7GanbptHuuFlmvUbQjTm7JBy88LJhIC0y6MvV0EkkPUC8Lqf7qJnDbJs2ClUF3y1BCeax7ciiM
WU01Yfsd+vojG1A8rOqNQa5qhqYEyHpceLXAtpXevwCwV6c4tX+jHvqHGTapsO8t5lJ/3JpLApxl
BJabNM2NT+PSiQIu9EtBBZB7jIymzdDGTO1uwYsB+cqMXJfK5GlwadG6v/VIJ/tAcIQEWtSB6jVi
x2zQI5DRQXHGYvRevUnmz2eIaCWzLSHkUBBGaC5R5r+a/MPyW+ybPMV5fJ/lZ8h7xsFSzFPh/JgR
IXe5Vb1JTlW/rewMrcMalvj2noV7i2d4nBoIlaJQ1gJjD1yfd/RezR3Kl/mLANNANug+mqmGYB4u
ke/npNA6NqR0C6sBShBCEk+9rEIzkGu4Cit1CBSd5oiAn5fUXuj5LnwxLtroGqO1BFSzOOvsmmJE
IMN2U5bF76t/6a6jd/83xIbi4oLd2UnVyMVNc8E199WT35GklwQZPGW5UZZN2osXDyj7He7Eli1C
w/YOYlhmztgCkqBwId/G9Yd4/Cet3ous2uGrBDNFD8KKNTRunJoGJRpNRlP25xp4/wIU9HdgAqtT
Qbf9LachBnovXdm+9NC+8rDn/d/1hxOwiUCUfZgK1knJp2pE86Cy2oFSGoWevfeUcQ6vhNFgCccp
4VGsynhRfH+NPZex8+VsE59/1SbuV6O9RS7tEqX5aoJqsywNP7DUZXFkzEotDKD8FE+1RuCALpji
/M5fNoy7b9ujmZW6XNcGncqLRwrD5P14z/+Aw+DB0qlAwwpJtvRpB20+K8I73gm0V2A1zzvELKzp
EwpPMCKGTRxPmTMVqtWiN0UWQWUn0enmagpwwSuIPMR5pTfSAUWiYJwOiqQ4SIE+4GPfPXmRsNls
lcwvzdLR/cq7DlWqXbRKhV2Gq0clphnhySLVHUQ5eKw7pgAC9AJvJg5S1wWn66W6g88m6LFcFS8M
/wm3wTXLkw6ISTmFFEf5BY/OlZf1Xx23KgSr++j2cQ2aVBKlvP4ToKU+CsB6llE8maNshy3g1roP
Ue9Fi2DW6NCfOa8bftNPRC1AH05tuwFGs5jCO0R8vkTPGRb+teGLGE31aksX4hXuzZ8oJJs/pE7j
90T6/yIcfN7AIrW2+C4apCqHpTEAEK4FctexIF5+dEnh5Ioj2Skc8ZakeHNgWwOod3VBEq2Uy4sj
KK0p+itBYU/9I3OHaYdrDb+gkp0Jts1iMZc+7yFN3eHUxTj+B5u42wIJT8ZQku4U1usdIfgJbEwU
qLq/N1TobVMYOYgZ0Wr/cDfJyIv8C6JgCPQR54X15i60c7QJV/f7y2XzXcIlYuRwvsgo+o4iyfU5
2/gu3SocVVR8rF+7fvjX1pntvnjn/Vco/HBLGXhpChY14ybP04rNoyvAWBVetOoqxHHJ0qAnkwtA
SwY5XEI6EnN9wTzdeny71XEyySknEW3fp8zBHFRKAd77CKT0gTt9k8NEFAnzO+QpYr8XCKMXU2ll
j0BcvHEEuo4TMdlwtzxdmz4RBGiVai3qcn/RD06UUkHUkKC2e/JuG9wJ+jRKglDK/0o/5hRrTjYg
fEQxoZ4zDeXu95dUCFJvXygGlk024geayu8UVani0Vt6yVU5JP0MWdLDLuD7HGqX+QxryGD7c5Dc
K1s+8cD8UHW4e973t4G+/vVPXBl5G7RdYWbrs9u2m9MaxGrtMWpc9vS5xvdfDMcuomW2738ncVLL
DqPydkZrD10/2SOZzhNBrL4wFfpkNNh+ofzl1WS/8b6RF8TfKFKzKmG9uRApYA7e0c3iJAJ9XfWq
ZcJRCZs1ZPQ7fnhzfNGzIn3cVyIT3+n8u5+xSzRd8eVH9iaDkijdDHF4s0gStQPC1hpk3ltxqMML
AUw8TJFp6ut0453TlGoWE7jwPrsw4u5LmPmpNzlaroknpUEBZHq6D2rDPgfcLoYHmyXyf7tJxH+2
xwxCnV/xMdbrbdJYpHsFEHpOvdAn9B1BZR2is0lqo25lQ7BHWcN/9eto39ykW843irwseKy00Xkr
h3CQkTr8Q6i8tqHwcjvd6JzKaGO0y0OQtjTreMEttmKBQpmQAU7V/wqqnbw3VpdpFqlTsJsRdtwB
gx0HoA1ZR3S6FOqZ1XpjMmQKX0IPfFxzhDC8sQdZ09Wzv53bPkdTtSJ+aWwVVbxnd62wbSgP4WAj
/GRImb5qjm3EovzzddDqyrifyfHXAkvSOBz0htrzJt9Lt0I8S+Ks+q6yMK6qm5t3mjqH+sLGkNqs
vI7xkE01aHSFn5QBhcBReBHG9efDe7PiyrNlK4SdDcfcyogzlwnqrwz4qb/RmHx5jm8SN3/L5dua
ASka7tWIAp4CQO49XMxuOkEnEJm0M+BxqchJco+ZZtMNnN6qn7YQds4ghFiLJggR+tVo8ouIeXGh
2k9sIuWoXf1U+3CyAin7AXRQX35wGWSsFlS+JFWz0u2FegBo28k5Ow0/pvO2fa12pQykWFMYRvum
Igz7ih+4kceKDoyXw9JoMwzs1s5cqE6nuQI0TkC1UIlSi6i3VdRrqxykfAxMuknejCOVXXgOXmOl
4gJzuueyC5c0ZNGOFOFwnV86Zpi+Wis6ABR8SH6T+ybXwIg/xRhElExpvvOik+U7tP3Abza7t9NX
ksQmhMqSdM/XlKmdEQ5U0gcvf5g/7gO5KgRurQcszINOWy44Ur5hF7A9/jEU2c8R3ZOLJ9ovrBy3
pPXW0rcjrUmT5sl91NQ4arvdlVaWWRrix3dZdjR7uiAUXAy831sqtMmh7dQQbW4LUkZdqzPZmbIi
raRyNHClSPHoaCylV5wWYaltkFgzc0SHpnaHGHL2enKv7S51Z8yyj6bTR3KadT0ruzmfaN2Z+JmR
mwY9ZlrEJETEsXGnzVWkcdDGqDX5HA7iSRCt+La7n/2ejyf7YLgHQLWUOR/ECFbPhZ/UkfFSK+Xc
ngnkshCyHHSwlmF86Y9WYUWmLel4kuM+tGqBqeEU1Ltgzq0Zq6MdC6jopORex6a5lBtR1GvnViVE
r5qRbIglnnxwiqzTeFxuoJmql3RpqjwyZgDm4CtJ2vbs6p5YJM9AKHGJMp7Loh7GQoSV99rNMw7c
cmkcnmu1G9BxH8r1d6zHjQ2H3HQDsfTLW7k3xm3HtynzIboEtM8BzI0OZKPijYNiFRuojHsGUcZF
+GlPKMRTO997vxW9XioFyk0N6gm3v0jI6T5dV6xqlW8iJvB4LFvMStPQhiqbFf4vG5JYvEzRjBiP
meUkqBaUs51kssukZEKbybxabcQckkwGJCA0vEcud6EmFqR73pv2fxPBZ32iIPECDxxyIypmkr1P
ge9veUgQ4nAxf/1sjaOCdUugJZkit7nmuQSKnK6Ikj+ROnIpVzPoeW898On8eDMB3PEaZywkD8jK
ylaL88cl2wa8QNs7ltNZoG4UmY1lcQR1ncxAMPjxED+qve7QQcEhZnA2HDGq+vwARk4AhWTArpvK
WRGR2AO3rzYQAr7bdRqveMRi1z/Zj3tk565i5rkANfbnYXdMX5o/sywYkiHJTl375KNYtwhgV+bT
PkcI5KX15S85Qtt7mAtAd5sisxMSOKRr11Ak0IRkBQAnR1v1mEYGniKU270abVPSiBfTwlsXAtQf
V91odhs7Yvg8GmMepKLm6mXh05iJGOpqr5PxW1SHk6luJLSz//mbodmcYb+ifXHsnny69ObdqO/S
BZdfibXUvM1pvyXjUwnj9xpsxsbFf9UgvxOEMuoQFvTLHiTUaySoTEGPUteNTGkn6Q8tDzPrJdkY
M4ZPIQ83rPbBXMhKrz7Bl5wabqpM3GK8afKs8XYlrLtyXa1ISkv96WjbYennJbMO5CtuJ8zFhcv8
fNeVxLaIuyz2Nw1dSARiixPG64Ng9tPv16kGhlLCCLkx67SwfGHSb6h9afZM8DLn6/rJD0vrlx9B
/heEFF7dZQsXhBgqejWg5K50CAJA2FZKP6OaXMwl5NKOqlGCYsItxaZMY4D3bBbg1WJIs4xoyrif
y+2yAjmCmU9QIwAJZIjbVXaXGyTOqklx/8Bw8B2PhqixZG8S8e0JUDQwPe5rCUC2mPN2PJAKAWI6
sZXd0REljUqwAqzcbdnPo3SdTaUzxs/zBFmWFGNoEaZUvMFDDswuOm5+pVleTKat2W0aAGx2e2ku
CpfU2yMRIh860jgPGAe9ucqQnPG/V0qxHeZ9vCGhwZrmUAaWYMz9x1Oi0oblAEjitavrBgn7JhaX
0ASexFS0VTD3lHN3SeTLC5erC9f7VfMD07VhCgJQRWiehZ0c+RYQw5lT+aAZk+KqmkMK9GNZoC4K
iQYeC27jfk7tGmX5XNH6zj2FFjWdfXNBpwOnGfFK0cw5V8zJH2saOb5UKlqWEyf/iyQj8qXraPdN
Z99HrkqBkNio/Hkku7dAxRpeqWu8k8oTB5NjvfobZ3FhmNu1yrVWDTYIw7DatMzRfOovD6B0F+SS
Qv71BSye4fCZ2li0one0YyA1Hj/R0M08NlOlQIqQCVN+Zhtc1JAK3DJ8+KgE6FfaRhfGgtxEthw/
vsRJBPxT/yHNE3QIXwMurtGKMrYQzfg7pd9i8v3XbcaF3npfUtaFtUucjD/rmL4lrjDVdv7cXW1x
JA+AVUtaYUr4SPgpfSF+I2ecEoI1vmOrZz73byIa0wwiqZ7i2rlkKSHdJjiiDHccI+KS+/oP/nAp
1X5CwGg6TERGsjUmx8leQ0Y/A8XNVkmS3KDkfBDr5FFHLOSeLNRsj2VjXKlDYbJov79eog/TMJTO
swb4z+kEBP6Rq8HlTadJlvB47IXRiQsC7Zl4yP38DvPX+hk0wTR4ShiwHBvTvOLCHhpUKpOK3U0e
dLuQckYNaiP3pmSJiM6Q9RHXHCLfV2G9Jl+TscJN9WPqkQs8x9b04+vRKwTQZj7VBNaLQCoVigOr
bV9zRebMHC+q56AdtnX/KaM1zVrJ6rm2cTlVAqX08IWQCZD1GraeC/AQ5qhGxiRBtK4zydO7AiU5
RJVCL3vF6dfv10d4PaXGJJ0zJzN/KWAHMtptuZ0KPBMt41RqJ0OitWTP66KhLkHNN/2+BEBRnAVt
19iRQjXdqxbqdOnjpknmug5RlSEcbgxHnD2jvLhocKGo18yUHllWGM8OUiqv/INszaRU/i/dEX1A
q/7N27GI9F+G7M5+i2G8M9iGcHrO9zlyfj52LgE16Yg45B6ArflQQNoM/OXTxt5UqOSl+SY4AQZ1
uOlqc8tCf74kY2fguNueAhyYfWjzIhq7kpfL9hB2Umu4iAm5g+zXJa3ug0lu+17d9P0RXbuRdE+0
DtzyS5A8G/hACcW/coA2I29K25Czd2AN3scMlUbK2LIhXxw6tJUzc0kAGn97kMB3DcCEmDXwdOUk
OpAntI80Qxm8Mxw4flTNgblx2ok8J2GtTOeH60BWbw7B+vmMOyKUktdNKCvxSsmcK07dknkZ0lWH
JESoJv5i3ekeT1Pgpigp5vgA0kNflNkja+C86qOeFtpeN8o7tslHfaddEkPFAgx0L8u7CPWnmcq0
ff4Jm7kdUfVjkbWsRwFjj+WtAsOVn6eZDVMwL05P8mpq9ZSxJd+JwqU+jtTonRL3Xs5zplAjrwKK
/MHpovx1Biq23r8EBkTB9j7PNE533WG1tnwONsC8JLP0zzI0XZ9fYR+hQ1U6Qp6wi7hF/NCG2sId
6oM3LGQgjCtPtkVrd8v+J3d364UV2RO7a29eUAxE2HomMT+Cb1ZPmwO+K832jPjBiu8gyP86pBWU
NwnNye+k5+G1QEiYVZFOradmWbXe4iGOhc1AQEzxs6ihuqAsyqal2FbvVjWFYutysokxnm+aX8XU
1K1hUC200jMGv8SnMfAcyx8R57i5ldh0p8L0VgWDN3fkl2RKkh/nFrksVj5eqzY8ZvaDWZfenvlJ
lB7mpxa3aUkZBpK3Ut8yH8Im7HOGtqmixZPT2jkNVucThHkooLLpWQDigbt5NeZRsojzHFmqz0Vl
oRlKXQniUzf611eOu5f3PGQQGp+2zh+eCuq2RQc+QXkQgtA712bDRvdVQo+sEaT8n6iOL1NJQLW+
c4KIXxtIRn4OHAXV7y8zlVMmCUMhs0mcQoL4BhzGbHegsBgumT3U++l++ALmRoO7NovOTWl89Ia6
YsykQVtRdCLwBZcsNUXE6kiAFBn5ohcOfEqa9MIInZELKkqnIXG6xQzgULSGijWZk9dFXEtnF/OU
70nSuTrWJVCy/839HAOKYYkezYwANK2yLYCbMM3UJz5Rng+uvfPhH2PdIgaPI36GN+sek7rBAizw
9F4+W7Ep0NwRRpFny3ikRilf7v2ViDfAwYPLK5gkLbBKHzTBIIQFmcvReLol+tO95MSzSsK4Knm/
gmweAC4cC0bfrAAZrnXnfj5+X4nGpjqrSE+s8pHCv2yNZPo68xN1RF5WU+BHSDBQSmJ3o2LYopGG
AprbOMRGjJs3awUGw9UPzSVBmM6QX1OXDs5GL1OTCmRDvXlOiQO53YDfj/qdOXbu2faGP1R+4Slw
TD9LOfmi9WY8xz2ocSncomTWrisFUi7gBgtr1jvFJeeZn411OlsMedkFiBP9wyS/2Ce37oiM6GLF
hVUrbv7RXo7yOVxE4rohhrj57si8GZLJ1GpoW6yr7ySse2NpDYkxo1B8B9QppW8vGxuLI7QknQe0
8M64bft5hjtsH7FeOwFcDFgFkBZxUR5Gq89e4wVHtUAbkm2BUTYxsuv/ouvfBcSWVsY1ADJjyfAw
CnSmwG4PiUuYTvMeByfZliTGxNMFEzg+9eEX3LMdaLowItC1zxCEF5/S5eKBsRMBB4q7Ivb///OV
6O2Kc+4MKM/Sk+B2s2C0DJ5nA0kQrb2OzsifEZ1FL2GYjCqLQPUtM7S4KtGFCO800uy5WKgmFLJe
jRSjqp3Rgaszx+GfWklJNw8UMLQPzKCxI2MolppYJN8obW656hlv2jn8sRVl8Gov+s3Zkdfclgtp
rNH9M+jmFURCRotEQ0fGPcTicI4kDKmWk9SZYvXnMDQaJp77TXFB/W04mO3HIQBIpwNkGb9YRNJ3
U9Elt06cRZ2pVuDLUR7N1P7n8LfXIg0uZ6YPVaXc3xmsbIWVoocVDzW5em+ZL8BKuY/FqHBdGBkT
hIaL30ykyM4cnvUQFk+n1+qH8djnPdE+Pnu3TdRmMlS7YXus2S8gum/KwYa6R2urTsiDb3Kl9UVi
W0WXHkQAdUa6o+oJnNv1wKAHynrY3wKpAyP89lz2X02NWsAHrMErUv0yzdokbyZcYNPSm5T0b1AJ
oRMUVxcNKYYxfAdJPrpxacaAatscbE2ebCTPDpz5fD4cTtlkdKHym4JJCyXV+Bsr4uKGrYfMvrTK
U3oWm55GT0bgOBhCB1w++Mc/lV7uuoXw/IiUEDU2W0oeMrOyZ54Fb1gmZ9D7YNmvnDj/W7r6hp55
1CIDu+eQ1wtoP3C2XaRknVucStMud1oVF77MeV7j9iFq/Oui01cYOyuSJ6RQvwPIr0vm0vwcUNH8
a9qmQQq3iAAoR2RgMrDveXbOgEPFyTDNnML4ETKAgOo6TMlZiq3e2p95IbE+VYfh9ULqloOVe30z
Bm+pZI8eyhIU1cdZKH3JPvYInmVg9UotlvoFcS50oQmiTlbUstEkGus4cglW8T7UvLXlv70EtoRq
crMQ+DBe5edi9UgFFXHnLzAtdgxi3mfg+ZNwanIj31HyXxWS6exWq7bGb4d5Ls1mpqJD0P4dj7SW
4oyZd+LxOYfrvluutidFY3VNvo7zWiwSwga6cfw0AiL2LmMbTakW2Sluh0hBeyUcyNbGwnsYkki9
RJ67uDV17AJjKzRNVkgHWM7zFymEOSI5LndW3C/DNXSzrNmYatLhUNFD2C/owsqcjH8/o2R5+oRp
3bsaGVpElehzJ0AAB+Hrn0TjsIcI3pi9HtwAu5VgduOt32PaFoLjf73YdVtdExAWqdbtZ/jCH2k1
g+lgF0k0NRlatS7+VxGL5qhT/k8NJ659QRZZYvuF6wUC7s+rIixEHHjro6CBEhB/g7YaaqCHzcGj
BFHC0i/jtZYhYrUvLz6/wykHmQaa69kwlAFP7b462u0cT3wB282XgGtCHmKgL3Go/x2h+gVXANBO
31Gku8wv7OnL2OPDHqjo75Yz4jzuKbxwla9V5PbxiKsyv7W15Sj4iqDMadsyQa9nPpOwY6GRl1HN
3ogM0hNWguY6d9Zx1jU2ZT1paoxivlwId0xyc/66g55KBB7sQruR2mxdLnxwJP67mdPl+AqkGS99
3qNk8y2k/srCtURv4neON/ilQvUAOmVcZpnm5ev0Xyp+U/0rSPYSuiZaHePcWH0j+c0W+fLCR9CN
zpl7dNE+g53uPVK/KA0ZMSP0c8du39F27/eBgQBMm3mYnfQGtPPl+KY/xlqqD0O7gqb7JIcl61fd
nog/lKSE5XUBYTza07atyttXB2e1sJKpTGqi7yuZzuTQbUVAfoKzTX2BDBPyPZkXCebgPmChCSEt
ZhKIuio0Gp/UjaMVK8ATXUceza8vk0VD5S4rG+dsjWpZbimlDXGxOohZH/hxce+yBP9BvItpBVvz
wSh9KDh6+UopB5DgVMa+QxkYF+PmwcwhXzPIm9+egI8WROKyXjQpvt01TUZYe1w1sYPSLfE/SA7j
djIe9gl4O1pCIVGddrkav7ZL5z+WQQy7yHWW60Gtcphw90i1T9YPuJ1A6jhYJx4U1mcJrEicC7HP
24SCBCprPTefTmSAd/5UoLrd9ify/taYR5Ok/+wcXhBMilc3gaD6ui2vHoQ0nXMFf4i5CchCpxjT
EVswtsHwbFRybC/x5UANb4zm2G6ahOm+43nhphE9RRr4gUV/lJTsIVHou8OFd9T5NKnTc9KQE4TR
3vPC785V8LGwZtTvrnfZS2tU0+cX03jBytmF8fg5PR+RFxERNpOZ808jyyNR7XkPVHKl1BtUGi32
ze3DhyEk0ZatGPXL2KZMSECe/WNMS8scRMJGtQaLO8gRNlsu4wKromnnGhRoLOwumi+2EN1L9kj0
0fgiLb3oLbX8HNBkIRFB9+koX4yzxe4JnMw0YRTgNNjiKUrCcbm/y5ETRTI9ZRuViVg2cko2U1I9
cJSY0UH3F0JLV95lzdffOeuTx6Khf3iAxdq8HzlIqqB+R3dGIZtXOiPtEyqxVPvo9dhgBaxmGiNr
VCyekFRzXHfpxe2+K2NNOjCMDOpdTNH1LcU5hvN6uDqyL2D2wuuVXvU/Osc/2ajqWnKqJAeK7MCE
FzMUf6F/WgeUGnEJd8Om9oyqn1qnEFjL8K69KLzRCiC2ulvqM6gQ9jBomrm66r6Gz+zFVhZ2cJtj
hCylr5fakKAU0gS9YmPTKWfrBELVdjY/zlwg2dvK1BP/Y8idhIXNuaGSRYm43r8Lr2ujmAM5f//W
UuWGxFuwUa8PIXHHQFCu7lA7BITj2BA6hZTh8oZfiGSsAZ8a3yiDpsVidtu+KQjRF7Au6NCuqLTC
U5cAC9FTwOqOFCsm2Ex6mThiEPpkL+BuMeyPm2jhCjiM7QzILuHX6A2inYT+VhwOnajCbOLTntM8
F719cqi1E8vnrfzV/FLQjUH1YAbeNljJppalYoDkbLam+zdSMJhk44OQ16Mi3YOVBMovDq9ar2jL
grj7PNYF8EQ97z7kuODWIrLodxMMGdap37O/R+xWDCwl9svze5gog9kTJFW033qNYubQVjEpHFTr
e9stXDg6GzUCwHM2yompWx66ihUd5XAEF/tSZ1ybHcx+rntKkmy+kc15InBAMYFpKJNanaNjr2DA
mO5feLrOZ3hOtVu+Ey8M+OMeRZ6rD0uxo53m9Mod+2nzxl4rjidJscrbgIzUUBLbBDnYg1ZvCJSm
lNmLWgIvlXV4PPC2f5dSLqM/rgjJ7/LyNSGxsOlcjD6cHsfb4KwHxz0U67ZBwbjUKMNbZHWtCZaV
fnpSDr/oo5x3hRWlWzNmvCDQ6juJdb2dLsqDGFHgaB/cF65DvcSINMMZymQTvSOj8AijGCnZDGjd
H4M0GG/cXC1PvJ50wlSv4cMEETXthYToDco/7wrPt6Ot8rneYiMgVvFdzVJp6aAoHrjuTN/347zT
Ah5Xbciu/gW9563ZmpcZeobxc/Mwhz86zuxaDKtOyhgyPT+QiJb0gJ3pEhTzSoJBPqcnP5Gv7aTG
AjQSYwol3lB6ADp5N5p0GKrMtDY/T97F5wul75Op9CTceEUG55GGwAcLnEfFrgXqKtBCyNraZG41
h8y6ARusdhqSdH7XG12ho4i1iF6Zy0Bxk+uUFXsvFKoyNWdDtCvvSVpEywt78T0ItRa9myIkV4bv
eNLiiDvG0QLnEwboMD9QYeQ8/QPYNoc4rWwMHYDizv2E7dX1PDiDbSa4etfdGR7raKUzxxTFlrJY
b8wb8OIFC8pM5grTXQIBHmIaUPI2j37NSt2BqHK5APRFgUjv+T5TSR3HJ2YXKWVI+B6sKLEcWRO0
HbD4Au7gTD/lq6EbricPuF4mduYXWpmgxZ4DUOxmSfE5ypqdhM4eJkuVJVJpMVatHWtf6Vcwrk+t
f2hJkaZ6UxgJW5otbxmWwIYx8qIGbn828ENDYYGTMMG4Tb5rPuOsQ0UI4e4pfrgQ90bttnB39tJg
aq7gB6D6FJ+v6ZvpW48PSRCQ53yxwjXg5T6ywKtqFcscLKazHu3Dz4QwkyfUCBdcNdfjivPzHj6F
Z21B0MJ5FUSV97fCQyGK/Xk9Z2EfK2+PRRw/uBBZICAw0pdZUqWvg7oeQdgJUWVqNd/xTgHo66KD
zjrsadctb6GTX5AsgJ3zPljqUDqeiaOZmbvL7oAeYDz1nz+yv1rrz/Tv7iKdCsNDFpBIrq316lEr
4PJm5kJ4iEOLOG7WxnatQFXeohApEUC2XtPaP9qeF2HOeq0lOarbA0shKmvbLucf/j8Ey8imLxvb
lQrkLapys+/BPSrpRu1Ke8v5BsXUePzU03lz7LzxyRZN9ft3CKKl/D8/8EoVPNscv6zIad9uU3jF
z80rYghJPv6Lb75XLhvnd/+zb/kbBzWXBW2UfecGVWgvzbk328rbDPPGzWDlPu/cu2J78Z8Om8Y6
wGSXpONDwnctg/IkB3ZLMVt5iJga5egFkrByiDQx/i4+y7rzrnO4QyLjp2cVzqaZ15B26knvwR66
uw9DAJlvSYH6Tk9W7TKgzdjdvWHnA0xzbwQGmLtyfIZV22Ruq6FYeUerKUZpVfJVS60ksbkg6MTF
uCZIThRRrfK9R7Lfask+nAjlWJerZMI+wLtrP/xu68KpUSSm1hcrxljLH2NRfC5gcSm1QmtOBode
F5tZDr2w0rq/9eva0pK/3s5OG1ex+J71tR/liknMYXu7RePKFW7qJs6eRr6JgIZHesfOYQhNtkbk
db2Y9rj2IPtDaE+RMhsA6QPY7ph9njPMVv0pzm/qOc/hKZhqEs2zs6vKhJul4/4rCFKOx5NU+B2d
pgB9VzcPUwasAG47J/lnz68zA1SoemwfTsbxHb5OUqCCIuP1RNn9wbEHSBUe46f3Yi5vQcXhBEDK
roXMMxz9OgJp9uHVTJwqL8p6QkJrfbcgej+cC+qNYbEISvrcojFroxPeWtzzo7fIPZYMlxT3csZx
2zaZ67FjO7OWxtN4flra5bFnhr4XXdozSvPHw5I/XnVIGCHgHaqGpLc/7+Cx4N0POt6+8tAa318t
CezTnEQDYrD8TubrfCDfNmMqxWNlLDcCwIPsuRj1wwtlbkiHrcyhlwMuE7rpGTss01SJZxDVIhOI
lzYC4ldlT//83weJYc1N6V1Iq3ypkQVRXKe7ORAgvgvV9skYiXQRzJEX1yJRiExcPRGaEY6TW5XH
Te+j2x2M0uNrYFAWlWSqJMu7UW5H2mKXxkKqhQVwP2ROWS0Vm27/2Z2JwwgLZEWCLLgHnDtSALmv
EaTLEtQPFiP1w0FHs2mVraBTneTYeFybu/Aw2tGdHUDj7xlDez89lksUUOat1Z+Xrot7KoHAL6R4
wGRmSxGDGXbNQc00vaJg03o6q5E02v9xu93QR/tM49fapjSQmsouqjo/7V3hUUG+lMpcY++W9rAX
Qfx2fRgUGuZBRdbsaTd72mI9hV7N551oN4Ro5zER+bBIsGPohZOQZ0hEMjVNx8lCmdWcNIBMzHo/
aWCzAq0FP4iffA05IS23KFT/cAmxxz714DUcHvc+I6ZYvg/sxXvC7fRGyhczqVpQyLHVq5pf1DW1
bpLZFHxwYGmdju0ptSY8ycNeUDQEhpy3N09+G0B9WW14suCuAYQ35ZZHVIdYIR+DU/9w82nCpHEc
4vxAk3DObdf/YkHSS8/xEcR8SBy/dmMZUWOpNjnngfmJzO5svrV3vYfcoaK8en0g326G6hbo1zW4
kwt5X2UyHmaYs+b08bVEy4B2SKBuzCDsdc/E6yhfiTvXJu2lyqhrNIe0R9oWlLRpjqqBxSp2+HDB
pifL4evwcxUskEU3fsfIwMi3iIKxv6ejIBxuVIcRy1po/i54gynOtCqpIzW3/Xaz2lz0vI06UhLc
7cxBEfkl14faD+WWCmO4epByn4fXnlNqxBIKafDWwH/kmSzVBYdMhP4NiV1LdB68qh9of5fxokUp
o0fiK/7QMV+eqkI85yv5pBX2UF4UZBxFWxZm9fOdrU9yvz+ihaqqbRExync589Xv3j0F3Z1eH4nU
ZOkMDhOMv8i1U+lhqeQ1x3StmD8MFcj4dTCkBd3Uu8VvHfIFSuonrX4/rNCILjS3jil6mr24GOae
KzLmOtx66YE4hsijic7z71NpseRtfVBiZ5xJTwv3HGrB1JSgIcSD3HkKv3YXgga5WJBDt5U6DjS9
MEBYQcrfgiQmJBuscxLfIJqEZ7HSCqnceeSMxdz9GR1rr3ozaQiR+g66Xt6+RI07ezLlaeQRljQH
KEl71Cdu2TBfpaWove61u+wa6UqtnM/n2X7SpRfynX8f4NnohCwKF0yXE4pea5oHM3Zu/7ySFGjy
kS82zfakK0HPRGKO3AZa0tdQK3krxFcbPY7aGsC6ryLIXx9nbWdAA6OfgnHdISn/uhV/Ja5qnDe7
adhCDgzjyHW8td/3Q1KDxvLKYgTxzN43mpK6V3tGfDTGJU8yOWHbJxTllju/uADHrnrZ72euWXrn
VbOe92KL42hqme6lJEdAnWCJg8diIaouk/bd51vuyfd5bS3rY8yGmFGM4TH1dQ31g/IP3Qw/5wQJ
OJMbGCIKPHn5xEcgTCBlxPC18O9L0fR8YbqIyFNyx6cuii8ScgcxCUxoqmLZlUeb31V9L97GFkcT
wdFQPpsKVe497twJKvGm0ELVN+kIy11bUFufKrKCLRdvW1F/6AZOHDQ4HU0VFXRqNK8b9SlCWFQM
itK/PNzOvONex4lxX2iyxglu01c2A5ZY1MwmWUDHoAC3Fk+gl0eDlRx327rpm/1u+qEVleJGFt9p
BIuEDqve52v3B9IXSU+9JdRXayEJ3wYLUXIGfrCNoNq/E3MNnwVAr18pfnLYr2mbLJ+1evIJEeUM
9jv6SwZcSBGMymgWkuOdrkBU9tidWrMmO5ks0lXAiGdGS/q0EolfBb8JKtRGC2kLA2H5MLTL1F64
Axi9ckWufwaAQObYoEE21TlQwCC9y8SIluzdz43KSLg4Uj7Ody+BfKNub2yuqTSAcAlMAbY2yv0z
UE+XUZgxO5df3i0eW18G/f+rxVB92/M5Yen1EG7nHZnOT5AlmeelMJWnEg0h1QaXJ4iNZBN3duEG
Pge3CHWPtbujI6jcgWLG7/8YhwJshh7ETK7Ia9rLku7vEl540HUMgixqXrJfI7H3z7g7X5H85Z9O
SZ+dLSuuuI7QYbAgpKRxRHdIBy4QeaECPOjbrPAJM7iGDzGcrDojKlpLBSbXxG36m55c3m+viq1t
8+bhN9fIj8Ct1Q6baklbyOzkZ4XwzWPUjqstjgTw/lE5UzPfwZKzX2HTXFjSv3WpMaG4xBe6rYgW
Ycc3YzAOgPkC3CbWTOsxQDqt0RHp34SKZEtRuFL9pi5yY5ZG16E+3swsyJmJp2/dFYtZl3Ogiyf/
kiNRjj6k+DuQ7yd1cx3YgGy+dePHojqkU1I2Ms5hoxoellXxPjpjnCl+LEFWbwnaMNRYH1//jzV6
WgRJuIAdUIvL13Hi96ssB9TBc/eyIRkLlohQlJJtbQkX19g3k2AbKvQQETNoGW9xol/3F2o/S9qk
am1+PIcRhZI3A//qUmEKQzjgfywHdpERv5ehMYJN4ljDJ2sak92WFz3bZUe3ok+/yYaInu9ZcUbw
2JHr536m3/jD2mizZO1gLuTQ4ewgcDqvFgARhrLylH0pZydF6mA1RImjziy5HLVW6sRbbxvtuks6
Cc1ivWfjjtYkJ4kEp7D4ZlCjq2aN3p+2LNIKqhPh8wXMqpqmi+lgQgvQwC6tSh6jNt1w3zopg5AV
8yQAuuF8BqLj9NcaXY8C2MuMo+b1xy1Lf6k32V6WdpUvPwfLLDjVdCTaHY1Sdite9SJHz4FKCe27
Tdg98/yNE/55RY9OO0aaCzlbXFy5PpoqI2qSh7pXOpMPVJMqzuQ4ToV+UVX4cJwAUgxfzu6CT7M8
UdZUJrMIHMzOnoQjaovg035/pi8FAqsJoNXzAnRT5wLniPSpHU6v0Fn+2BoAK3jR3Peyb7H8lI//
dgL8ahV/IpGeOu3FHrxudDOJWfH9F5UASZLgqu7pa4+pY1l4oRf9yqXl8LGAMxDd55gieoGw58hI
YZ9FuSgcJaEif5KNR949hJi2/OnrObC/aSV/6dAwm0Nuxa1GY5NpvYyV5jnnuuzIOZOBugdnwkdK
OiACzpkNzLM8bddW1Cm/zcUnKJDooSvO1K1J2QEWinjd/1LH13wAGmopeJI0aK/7hfwhuDR3+cN5
VxyowmKxHPBq6bs5WfJSog3EBIoOmF0tkHuml4ELNNDPjTSSWgxXUylKEgN8XnZjhUZBAgQdQgXV
OO5O7KHDsy3QZBhDzIcnBuMTT/+SvMAhZptuY5lDtCHwASeXuOZgMX7pqUt9UamqWRqtn3kTC2/Y
kj57sKHOg+PhqcXW0lF66HtZ6mHuagzm3G8JWom2xFNQhizu1lc4Wfw0VtXa8knQoOmqibVrvtY1
oQbPrD538T6wclDpF80Q5OzNndPFdXLblvazwKmWQsIsBzH0ahbGKBC/68ZDyYYcB3xi3GJSrW8/
nklnge3kZ9l8tIWSkQBQgEcO6gnz+1/A3KazOQirZDyXnlBTH3bszG9Cx7wek6KqNawlYhcSk+N9
FrKhsq0plTdB/mUGW6xB3fqkOdLX31NUtqvEtw88N6uhrzxFPTvrApb/9qg4bKJ7cKQnpMHeZgXq
TIbybKKGGQvt+rt1yOS+SncOr6Q5L69Org3oYxkRcG466dJiCH0kZYMsuvgh3OncLWRgqzTf2z3/
0s5XKk7mLc29Z0WCIZrY1QgQvJEF9tyvF3q6ZhO+xR/j3eBfNNAM4AKBEaYXAtSexW/KvbOpD4Xi
ZiBVJSCu/JLZDW0iE2s/7i47Mm/xJMlAARAO3tPO+l8nbImt0R581LmoFbAiTGSHDjsd3ZEVpnm1
7fOlTpTxUaNShrNcAMCds7sML0LZ2IC1ZfXf8aIbNBaMsqiT81k3gUn8vVrlStMh1CmMdpetWw6w
RKHJLsJiFdtB+pn/CrV11oA79IFDFO60IHtWtKthAYPTM4f68kOx5w7jmK36zhy92sPVVWDS6FWM
k+NU6Ykng+Du8myNnmRbqacL4RqmZXWVnqNZ1EM2ws7tk6LSONxINYoQwL9yXDCxC4klR3+IaI5W
DOSC2MGKhT0SOHnxzKJvdq+AHOzunI3S3Qyl5WmrQ803Lxyo0jRKY4VaNGC07GZh03OecibesBpP
ouzQ3tNKYpRZmJfyn6DbY79RrjTwAN2HpfWTkULarqFGdp4Tf9JgnqWA9CoP0Qx/gI+DUHdcr7Zp
RUmb+0W3CnKzXO/3YppqqlpeU4QF3e1Jl40NmqSpFwBdTA++uXYvM1PYWHpBAZoJ3ilhRVqJCj0r
3BQxQDATd5omcPxdhjXkmRzdy36MAAZVN/SeYj0OwVTzGSC+DEP+x0ORu5Hs+PsZTmRuDsgzMy1G
pdnd84TWrwEvOtvBXtcFkB/Xk3jeLMM+xwvho9xuw8OL/uzeWXAE+kwiLO4X7VbHj2x8C7TKlk+k
YXsc9Fb7trhUjOPA05cFjNMlda+at+GUpGNoJtk5LrM690V49RfcaeOsinlzve1AubF/oDqIL35H
+c9KO57m8LrhpVM1ZHXVEOQ9eCzEinp1ydyr17O6wSoE5OxL/5/4siQ/ztdMxLfLSxE68IZwUJ9S
DeiU+krYBtx/kNZ/E/AdQQfqFcAP00AOpKSXzX8uqypy9g5j7i3TTvG6klb2rih+Lg8Bz4OdlHWN
QIaY7s2fNa4mNmpypvUb5jATeqZ3wG4fxUvIp9EqK7HUc3CjVceQ4jdW8zdtbje7EB+D/qPoX+u+
Ta/4JyckIsMqQH69KEMlTxTiGLge0olfWqAvPvnTI1+yEodzqa5ngrCO7M461iX157JrqlUURnYw
UEYmbcZ3e6Xa5qHfKPG2272JroDms4DJA7kAxBh94adJAVKlJJ7RzBrBccV/gMq8+QacEOmU7AH2
s7JjMIN+WWhpUfdp4ecb7xH72r4RoF47RU0SAuEZ0wURrijB4cnbMDaqgwJDFsGHtkg4668Nwd5V
LOhoH1RzCpcdA2JcdTuisDdZZ0jBlctaWeSbXcSyRQ95zfnrb62EUZq0PMNdaFmkXGdf4HeKniXv
5y6vVk+LzPuX9FtbNVBLdB8CeTGrsc7/jKeixc6Ay3FOW9eBV2XTuM18x6r0EN7a4XyNWJF0H/N5
9Nz3NUtJ87gHSnE62L4rbiCw3atGdZjCEd7ld4GVg0ZE/ZpYkgbg5v6hKOK45jV1Uvno4L5EMhm3
hcdrfvAsTiCRMd/cVK/V48P0sYDXV6a+Ms/W9IXrljU37IDxTgvhJmhf9nXFs2Xve7VowzM1IM5U
fZc9he88+tS2jKxzcMj3qlmZRP3kdbQC7fy/Vk+V/6tS6L66QlEhjE8SKU7rS1Y775re26l5UeZ3
zx+nsgox5KcKE+M9el5wU2pn3TKR167QXXg6FeNrMAOzlYA3JBKZLOPwgVatk5ZPxLaWvm0CfvDi
r9YwEtjOvT+QV724bU4WpdIIOEgd+Yp2mPyZLeHuXi8LbYUVapcyshiUFiSPtnF9AHIqhT8obBoC
l7rS1Pvl2hCBnvI/IT4CgcX6Qf14bVeEXWnc0Yn/nCDeWxqYzQ9+eeCx5zl1uHkdmPJgDxZ4v3F2
Wa81XnnkLmHzDUxEGtNjakjR5uXlt7Ag2q+69NGQJM45X8Vy7fvLFR49VJ4rvb8Kgm+YbVAig3dJ
bqap5VVyMm+csGk0x+sKvTTlMJ6Ya2yhBQel9cZAbSJ5Zu9fjuYI/JTEX0phV1zcTZnEVa1LxTc4
tBtUV1AG6LoimlKp23oR+bz/VeSloV+BbFpO+rCIbS7Vrt+QBkoFfFPhupmACYrjCO1eU2UgayeV
glzY78z5L9+E1mhjyNfUmY95tfFipwjlOBYo3FBx9zZIoRd4RMB9t3nBg1r4u+udscDH++g560OZ
slxIo3KTyZeJSbx1aKypWMPQdX3Buiv3dUZsqqBSv7kcVMFVzAEf4+K6nIfKS1+Av2DvizqP0C3i
Dhe9VqFXG8CxuWwGXksbeXEDQXfF7aSO/V6WueC+d6lAkQ30fjNVoeHaP3GtgiIPjEJGVSlZaaK6
YAm+5ijzIvF3NCJeyfXJKM0G+0TP9jBDwc+oVJhAeTylYCXuLIeKwAXuM+t8VZNg48/HsaVdUJWb
WlE5PWTJa07fyI+apu/xCWjZ3S2PyFMo5FZa48mBdkWrZ4dR1TW5X3eupywaIyrLkyes8PJniy6K
VW+0t9PKhGE3knMzM8AUkzVUDiHz8MjZ25PVHbIkUCJMerwCYx0Gl9TfbimBQoEjbg8bDzgKiuti
iC0gDl5ZIUD80YXg1CT59n2p7qdybjUDHSnzwJiwcGPRTgivuDydbbKuNy1aIKXeCpUj1zKU53Z+
4DSrd97NXodi4pZthC/ZTZLj1Q5QvWx1L/sNdnCS3yDvIwVM03wSRjCcxqTdemegIBFxHwHRirhV
MQMsuGFFj+o8KEhy1ZGGUvsgWfVNXgn9uo9HigyVlAYpvzPT5+nXEvnfQ3dMqAYu4iKFmcest1wh
N77OF1WzJXvUzOTJovABCmU+/NdQ6UozWggtSnkdWoZny8f5o0Rc8qGl45qlmXg0a/Q0wOK8yWeL
JPNvVkwmT7kW5tKzlNwCDd2rP6KACxsv+56U96iluEFBCP9LdDIbLDi8SkYDQbvclxt/GqXuF5aI
ftQbJphdWXSkQnErkjnP6VOnhGCRk4P17r41yNx7Mtu1fpDhAT8vI9dYL/XE56fKJHF2d4o4suwV
XTKDx5uvSAZrNW2Rj1qqtlasH1mYcDlNjH27HPIksmaWfbzSGSCS9RvPw2BIgRd/iC+Xn84/wywk
pF/dwGOxkWBk3qw92aACb547X8An3UTIV7qTLMDiBekdCJgK6d20dPLB50pnOkPJAHZGhM6ck86L
eIasUEUJv+1kqqM36XUtYMw0I1ITDN3Qexse2M97W3MPcWw87fdSctA/DptJbXuO3ZI+lHT5kdF8
kGWl86BdqHpw643bh4Q4xjwzIDngtslabbviH2cDg1iFG+T8k5xxvg/Ul70YFK9aT+SO0MXWOeCl
qC+sG/foRnS0CeiiZLjO/QutrBH3FJOBIbFRpSZRIUFDcJ/VntpjoeSLZQiurd3VUdiLuzssD9Ez
D/W1lbN9O87UyHXklbcCUtUDAamJMEMBNg6+CJkVxT9zWruwxrZNVAi1mWxUkd9AittlPrYb69wK
KgLpuLsgLtLDIZL/w76fL+3I53XftvzwcCuCxBKzu1Q/Qrpv8KXuSkEkxXaGjOTeceIc1S1hQqKK
Jn1qZ4rGJgpNzfrhfWyFmuF/6kq5LFk/0N9atmvNOYUD6hpjCvoSvX5cGQduQlnNR9UtnJQg4/Ym
Ru2WhgpaoW6EpXFeQTpBaohJ0V29iREcy22OQhoUW+wP/CSkPXkrOwAOHhD9bGnSwa40vTv7d6P9
DpK/ihNyYzckgiXenyqMIoKUGhMGEJnO8pk/i/HXJrvJKrPrh6WtBBcCe/dfsb6T31Of5sIspnpA
DmAbbEmP+aCBhu2mtZdPXrfBC3Lw09LquHzIk83dwFBJS14Ra3GjqKmhDPXt/IbjmFeSEki+12Nv
Jk+r6igdk0S5D9t4OG+NbCDvDTfcfQS8njjFGaDkHsuKlEezGIkgSz14ggKr6tMWZcwbnTQ1MFfG
9sW7MHC0EmoBYnvO6+krGAFxwfjeSeCPN+fyuau1VFjQqYLT68jf6TSmxGQe8EKYh70chlJWNB50
xXRbkRGmIaRj5fakS5xArjHGuVg5AhP4d4ZgC9bwscbis1/ghtz9gzhE1QfvdQf/0x2y+770xksa
eUZtDY7IJy/Ny+K9slatmNLSEJgVlJv9K4jsLjgNirq0Q8nZ6/sDgXjzzLHqL2WtgPYsPSxsW+nx
6bnK9xlJ4+23f9A5gXcM7Gz56s4jc/Ko1p1gY6Zm0eSWcJXOHFb+JPCxw5Jh+rohoqsxpIkgg1L4
sXyNW9Gysj8up8FJGTnPJiC/I0Ry7Xi/Ae0g1dbtaQcKVLsf9W/N2bTwELqhxk2vBBbnB3Ec8v+E
yszU4R0F2kVQwdxALRMlLKbGkSewyyZ2YtlLyugEwhB+UaHj6gfDN0L1Jisl0OlozCD5MxBXtz4f
EyghDuH+/G/Quo/5JJlQxFz/ZMgpm/5Arv8INDkKfqnicNs485/TmY4TJ3gZIya79yEd5UoKRU5s
abuZbdvsFj8w+ofLO576R2y9QDJCBecajDrCWg4BnO7q/8FpKj8gomB3uEgOm/XOlN3FnrEhoXT4
s1877g4X6GG8XYZUuaMHNB3x0o4kMFhohwaA0Crt1s7CgGHHD8H1/8lW14//HOgGqEJjmHz9K6xw
89bS/GIegh/6um5zXk2ZVOO8rqd9UgkaJdc14uQ49XuEeg6APArJIUVJF/SJAHNvI2/x97r5ZPQj
pqratxX1Q+gUlsnJEZ3nEUPEfcpSKV6J9B0v7GUQh1JcQPuQB3g8qP/H7UI5Ivw097pSCD26Mmwk
SJ0U7bPA4Vn72nkIDtfcAVA2cF1Qmn20qTVZoO9t0xL+YlGfVdaJBX8ISwEJT986BTETS2jYOd32
8Sl5yYJvzWEMUdT3RGx8NuXOzrXJVbLQTnEk0cl7rwTxbPmbI5cpVv/aP50p5xgxWBCA4NXWP+W/
UxnrgGRdvC+xlLxjjz44cgWExEhxVHyv49OCfTjxpgKR3eD7sjZSkoyksWPp2Ysnx41iUcBFVojl
obDtXqj4xKwARBMmGXeRUYjfsgAowV1MoYqI8tr8WVdzn4P68yDBZUsI4E8ZumpTaHOn+D47i+W2
NPHnDui7Emk6zktmIE/LX0/XvuHLhWdFSCiMO62ftzVXJJbuX4ZBTEbhSvd5xmRlRwCMpRd1KFVT
QaR+esPVIbS40vC5Wwn3t/9mScG668sU0FlT0dazLhb4AlwAmj0qwfS8LqBu2XnaIwd0w6TXLxVh
22cI7iDwnPBG+0htmv4ZICTPdGvk9UyN6G0rnaV+wCbjjPx+t3qjpUt+cOs/9kfTdzuIv+4biWLX
2kgybKnGgGF1Ngtgl0KT1KMcb0YtnN13wriM0H7ZrGWzXwzWWqTwl3QntAEKnPKOjKt2rOYmSOtA
J9qGJXDmrZqRxaixUIJtTlihWOZ8msEsadJhBCR3uF1XC/6duTGodgeOdvTr6+UbDxYp3NMBCIBG
p0UIUJo9ItjQwaL97jz0K0iHLn++/UiU1bd7LYKzJPFICZ8uW3yesQ/CHoLzBeHQ9tp6M+yQbQg2
sQs0Kzb3mdSOXJX97Trtx0aIeXVGmDeH3HM9rqSJr0z9CrAMsZhn4H2/IkhQ7G732EnX/k8cGbld
Is0w/zINS/SXXpB9MDfEjBjS2EHkoObUGRMlCGAKhWLGp+A1z/gGiN4lf6Ap5NjIbLNFKEJle//6
APGOrL9tmVcCTa2fxtEBnyZC47SuHfcAfwHeGQf02rLZo4X4a+qBoCihmd9dGRist9cayjo3Vpv5
2q3aNMTYcGiRV5QkOx5klWhqwfGv9I10ggW+5vdyL3eIfyue48osTGa8oMlePJuaS36d9Ah/UITj
lJZuRUoWr0/boUw/H2BddR7JQ7yNDjGNhkqUJnQ4cIk1vfeSYn4rb35q230BoCYocQdBd6dW+JGi
9L9AHFhMwNGKhR/46DlpV21N1Yx4hnX+/0bJkHBhFqHd3W51qsHebqzuPYnM/Y4kQwO06ADmFC1S
a2wFzKePiEGy/BlvWH2n7qUQv6dR0nGmAkaspBI0++NXwCcS7gCZtnM6Uatq2z7D3L6F0Ypahkzz
WW/jH9neILQDOuAVmDQLW56jmPHC7XXlWYZUEtg0okR7DhcrrBBKORvmu1HEcKlTgqTFhaEthEmV
zSJDzpIoMJ4XJyX/eQMgboqLYJNA56GCKajbqR/EEQCLsY3leOI36+CmWcT3cWdBzXGL7JqzwIog
Zg3rC4k0xoGLRxB0W4g2D0xciHOhBbxsT70b3l6MFEa0v8YuUO9Jymi564Vt8siOysd80ls5CJ5U
ptGsh6P0VaK51Y5KH/AF3VBSFVzdEybLd3aHYI/0JJqMK2nki1Uc9Oko+ickhJpnx8wDhno2IVIW
1P40t/ibBNsVRNqsbegswySu1vgrZcbZYbS7GUzVMHb7aU4J5G/h05qSa71vLYVuoT+daORPFbl/
fc+1eAhujRcDRb//Lhr9orekXWBM8iDenClF76beG+J2Qxhf68yADADkPIzownoTMTxBp/Bnovvt
YeRIHdi4K21YQ6aBkzu7E6heCtKLXJw5pK0UgqRj8M1c/S0DflAV3o/n/AIjoJpITLn7KtUi4uWR
1sEquUqwqVtN4SP9yi9Chrc00TA7wAZev6Y6SGChezDI4NtX+37ZGhBq5FVgfLeduuoXkpfAcMS3
Yiy2qXtd6ZoQ0u2AsIArketfeIcMO3jdtBAOi8s76HpvBC6sAeTC/HzALBw2fsqzQooWFel2uXJV
OYb2JIzk7on7ezLVL4AqUzAo9EduKj4WmBkkYpaD2ppWEjXU1A1V8n3Rvkx2T/+mp0K8fluQtbjD
Zew/DySKS9BZmKGQCbFvD8vZuDP0D3G+lrdPlP9fushMtOG8XUVSTKMu/3ZVRkWq4DM09hrD3S9s
YAyyBBUJVPqsrC/5RvdJUaJVJJVfvIQu5Apj+xle4eGcFwh+RDB05cYkdmwb5jro9GKplFnugD6x
xNUa9HnzckPCbMGs+I/wITon2k82zoyNrG/5iE1kCnWVXjD6XrweT9sA/8uSQXZl4Vgc+9QKygbM
Q/9lg2P/Q+tRnLBQALNYkXjnx68khYWPaHVLSF+sZY2OjnHFiQunaOk9MDx6FRVoFSvSiCpSNb5r
qW6/eCXo97932aUa4KngGAWLZkjSFX3jjcYaPG5lIsqf0dRhTr44FVEmw9NKeX4MOhvcHfecre96
Saf4jvFnShZKUEfzpguc7ihhvQVTeMI40g1Oq/94Y+61h0wa21jzkhIyBbjgYC/ek9Ymb/nAKf3n
eAvCR55RtLSJ4hdK+kuILGFDYBV1bDLYawgfqLFrOdmzXMJNDbIyhPqDc9NIezum8vlo6cSL/66k
e9osFJ5lamEtMOEe3Y7oKh2PdcPQQfjLh/BBqiOWy+FAl6WOq610PxWlE/0o/L9aI5hg0I7p9DnM
VqDKRV+bHhd16dd76vP7QVpyX54TTuBgHVigi2mCwKSkm9bbvDf+q3QCOdeKIgvKaWp5Um8muHii
C6GjCePOn74utjSQpX4V9dg47tF4xUk45YB1Kc0mrqkQhlPIKmiGV8h4N3aCiryZrqqzxZVpwvqn
yhi4ue/xWLz9o3V/NHfNGmDlFlEjrE6MR63fBLLNk4W7KzfDYnXk4drrbS5Zo5OFpb3clwrqWjEh
f0GNFCbw91nYIkmjVXGMLFnvvq7CAHAzEZw+8wIyRgjv/rXejooQ5G6RopEtFfgHIWAcmGQt2T2E
CSFE1xL5zGmxu5vlnQsczx2zdP94vahE3cMM4xJeFxiStXdc/xdO6ztA1eyDjVpPRGUquHDf7DaH
79K88rHTrBafQbnNv3G29U4lT69ZrzCAfhAkP+yICdlEo5txqmwM+w7o83SAh0OuC1CR65gu8slv
sU2DEkmBUICT1+OriZgwc7+ag73ukVNxZ2Exl1OM0q/Tdsya2ngu5xSoM0RQKAl/YC6KMDxRC4wu
gkCiQaRvS9KFXU1AxD+qs3XRHBqwR3kf4UcDGyUq3Waqpj/9qVX18xv8ZpfZUqHggu+IsSjfA/TT
/Qkr089OUNGPgMHtxebo3mqt1hfUZD8PB7C4YMvSETLaZRWnZbi7X4oJ7a4S5UylVypu9niUJozx
n+B1+mn+pYzyW7krjmZJC7x4zd4fgtju0Bb3rZGhgdGsNCp2X+31lL5QGxGsRMLEiZDc9sXbYIQr
zJmifD3Y8zEapC3dpCpw/JcvfF+s+RhBbO675wL7D6Yq2RgsNyPdGO42dXp0hThdiUMhtR9n9/yM
H1Jns562bSL3+bdz4B0j04KdmCanCiZxRqQ8hpoG6LEut4oDZamZYjmhSvYUnZv4d0/WsMZILyzN
ww42+xh42jw89iHxyoG7/CQnHWv2ZWGDJmdFDZN/ncj+BarefNBRypmyF42IvmLSdjc3d0DmlUx9
gB6QLOKIOYsezmYApOThLBsTlpAt+jr44idR3VyrqZfJtWHPnLZN6YNQF0AkzTlQoyWot+vYqulD
MVbT7ceIxJIajDddB25hkKVMiIfT2KdGIfLoB2mD48lHNz95teK9ZnHAd3Z2u+pVn36drOyIazCV
Dp1jqTOqg9yYGGI8EGuqewGDeOSe3mKyMrt1zUPAYP/dECdx6SpvYMO27Pvq437kwKk4gHq94yyS
hZQ1YUmMQ1wDykB6ZEizfoKplbw36J3PX0pUEGZ+uieUN6KNFKTA1FXi0BOg3O7sgtXoCe6xhL3H
x/oSBQQ6TIs7JoMGLscMADwUjZ6K/WlFMbvQeuMxG/WNVrwWaSxYgm/k08QPpbNob96kLfwDLs2G
h5XrtKI08fdGZRUeyNHcurQWF/QZWdrQxJU187aa982aD0kfxIYsMnragURmPEL8WOf10SxKT/ae
uneHnhB4+Q2sk5nHyZVs9nlFoJeVo9iFD87dm+TCoZY1VL/FxnrvZaqZkFrqqmD+CvT7PKUxLJW8
zJHaDX/xheC6Z86ASdSt8HamqObDTwEQgVsrJYPUZ5vjemElncyXET95HDUt7iXr6qdX2V3CMuOc
NHYoy45pX1MeO/aVCkuZq+ZvBF9h0dK/LHwY0+lbyvY2bCiRGPo7gKqZE9l1gZe51Zn4nuAJqFAQ
tVLyem9IUT+3nFqeLuhwTy6fHa88WpJHSWP7UJzmRN5AH+ez3C9hjD8OzulgShx7Q0XnQFN6tW0+
NAZ8P2b9liD0cAl7dimpHBI4Vz+8CCcW4ZVWDQoy6Jg5xCFyhbGyVHZFI/cvXkoLeDESp69nwnDq
/MpKxHeXMyms3i35wqCWgrt0BF6tDLuYRCJYaujnvOt/5PXZSVUZmqafoNye4HePnMz69+xsNewx
cRZ/QeUJ6TBTDIgKfvBx0jy1G1ZUvSTytnpnSAIhgxfSYLfyYgsVuxh8Uc5R0m2alC6BYjrUImeD
HKitiFVeLM9wPtoOzt1D8NYdrou34UpRCQ5UlC6c9cvHQfcYxqXwqg6sP7DZl1v1wl0mtIjAKCka
dxIKfrTYOzao94I62pMHItYk0Brs5r9N3wpMcK6Bv6Iy7QvTHcwm+ShIGn1Wapq5mEndTA4hPAA9
cdXh1ogWzH3zMMBKb+Vn7HT4nSChL7JOTmBYcbsf14Kok3Z1UqWnzQ4U5/RQWCsiEMhQwrnTEk5l
zcP40eDCegxJGZfN8pf5lvksb3BvSmunh+3MSY6QCVMFId/rrCUqnushInmrLxR6tW/cuMLtpC2u
aInXElAMlMryeQyHS9FzhXMUJqB2YBxs3Uvq7bpJp0jjTx13fMwFCRthtoI5xYDXfrg1o6tDGHsI
uh3Ddme+Bz/mIAipFqLBVab4jrseOMZFKznRAFWIjKS7tjz2ndPpdg46zgDsYmCxHYrwjD29d1Tl
egP1aphGJ6DY61Fj2+sH6JkGz2QfLJJWY8xIplLP80t5ROfGaOMANfR4OSN/brBjza2ukBmu9aeQ
8xkIREpP/rJizu/iRx2aD/NZfPWYd4b/rr4eW+4c4DWlR6wkkCJ3V417e8urhI3B5gcOlzdbGrfo
+/ZKIz2VHF1cntzkJ3UfpHpLS6vTEFm2xvWXrH1enFHkJaaB8yepq7NlPS7WW+IAxkp22RNtWO1K
CerVPu0qYt4Vxr2jgGizlL1oI+PUelJdS0t1Mvzeb3ZkkEcu9WrEnJgRdXEcOmK4ZBxUdwiyxR2d
LPHzFRe4JUVTfldvuFXj3WyEhPM3b73XlRW7/8s45AvQy0EYPG3hulgzQwTosyMYXMx2RPEmFgnj
/KwEhZl8TT4tXQtPdRSQLQfq+H4AKR+imq1Q5/CWGn5U/xqkEAixbDWcgQ//nnIm8ydA82xQE0/O
CuhpUlM9oWY5Ft4XNniS7CvnOwjAfSlmuTx4zpmMPb1DQ4HV8XCyUrbi/kWTljZYGzGNroAmX61b
KEJm0VBVh9qmM8KvfddnvcDWKD+F7AbUhbiV1r3FY82+PZHOJGQejKZvc+Dg1Xe/QF4H7/psQNcD
NWf1+81xsEh1iunwWVWL1+aDv8cMr4d4O+uKqEEVl7HSU4d4O4M4CMh96Jtzju1B88yfZdTDsQil
YfxlGlwMUyb8Xbzj2FzDZrJ28ku/upo/ApXJHdFnXTM52fwW3E7iNqF4SqmmXKtJQs1IxjfK5yST
MsHlFJJn6t9IE4FOP0phH8r+BC3ZkXkTKr+4r07YzhfvnXb6nNmZU12v9Wz6gHLdDJ3NylJY6d5J
HtvIMpY21D/dlhse+SZUe7Yy6TvxIjdw00qqxZYDsQxkziC9g+aSThhhxU4GamL9CVJx9pqhGuoO
o2IpaCFTDBg6rh4UHPulg9vhMCQD8X0Q+17qpcz6KLxPDdkplFX0FfFGiJG3M57R816uumTLJXwm
/nIHd2BYlYnln8T4VAZK+wFQYsuxrbEByVvjsHpIy92s/dEwOb94n2dn88eGVSsyypVdRNMHlMEJ
2hdI7luZvZ2AyR1RlJ70nGefro4QrCRSBTZ8wxjSuhRZI/8wmbft5AxemcM/sNnGtbmNs1FROAkr
XLdAeK+mdVqrzuR2iETJOk5rN11y0rhN7cINBYrmGJHoDDt2qouFH2r0IdSuCB6j87KrAJj1oO3O
EqOUWsrqa8D5b9+lYZ9MA4O6WNT522cWc+W6LQ+xHHFptrndedly23i0m/vp1/51aeBY8mCZWMRW
Qfg6TsRiCy6PbMsKxp64cMNfky+71alIC30BcOLeQ7szSD9qJbK+GpbSHq7TZUfkd1schx6eLDGh
RnKCpWPQlYnL0R4N3NeIgNf9BEk+wqcnSbyzsWn2XiIQxGqQgdDOt+mf29gQY3F7up6wrIwROrVF
O0SuxpSlh7c6dTqfSZG1lyp//9VXQoSTB60jDSIxnBnSU36zvXFbI0Fhz04tUs/8czXg/jz8uq0J
vKnNTITXzlkZNSVffx1slvkRpqWcTkfSQNaWwBDHYrc5Pq3LZ6WX47OeZyKEm6giQK1AQ/VhhdO/
+C7kfsp9ZkJcRmFazHThwS/zm+hykNkYn2YBHwMGjsu/pu/0aUgdGTNTSqdRYpU5AsZ5nV9nknus
C5R+VE0yU1Y9V/mb/PuUwf1hLTEpDevrw9fycO+5AZXtZ46JFbN7jGghYu0NBtKU5nXbb6ud07u7
+knsDLS/1DzBXjJuBn18IWPkIk8q+lthmCZRtTbRz+htY7Mi1IqwGRkOuH6JvKyMDr2DNTpQmunf
4N5Pr7ZsEsw7eV/+g4Lrh8Cl6a3CrjKzEpZihWqgF6yknjDGh9zmviRiS8cEYQELMZ6Zp1v2z1h+
gy8df02bj8E4GgqnOGtgwwVoH3gbjDAmr1voq/1vKtsPnlEApmHhHE+y+Qp2yFApoMP7uMOSpKPI
unJF6ZfGLn/dzLzQg/b55jEFBHPvOey73RnyjKVClzp+h20ma43QJDhaLuxtzL4KG7zzmEvZ71db
vRQHD+s26VFiqQ+q5upK2T8eCQF6UWZDvMUu1ndS6D0hGtujHDpLLByFra0YQHZx7I4hWf0bdhuc
7KBBe2Tmxec+bQXcKptqOC48WSpe37X1vcdOaajTBzHOpY+Vux4wxbbvcFbeqtO3OvsX8j426P35
CbAVfoo66h05f/pd0b8c0nuP6x5Rf400YU1kQ27uYCN6WHt2ixWMEYM1gDj6TyMuz2Nl+QvHuXMn
aufR7B7cVlKwNSeSUd5FfdRmwhHXsIVaY16PZguAj0F2yd9NHDp4aFo9as5umlADI6HaQghiaIKP
8KNajg7AZ7g9RVVn+RBml6dJgUe/HFTtOpm6s1KbJLBvcggoNBK2qZzrWdf0K7kLWvgyoPe3h9a3
m1eYd3IAz5sxkJLrVYSoTYCBH4sUNdhIViHgLyBeDYY278P63XpbYpDU6tvibyf+sAH08hNj4b3b
S50oBlu7y7hgedwlwwE9holwNhuWxF6oTmC0zCrpw/+HAnq7Bd1/ApXYbLTmP9u9gjQ5GLY/Qpzo
sEfjInVmHWEO7j1RvjSm6WLopMMM71r4aKweFmC30q4Mpr7Ank/GQqbtF2b0JwXZfdLPDPMjBNzh
njRdJQgLd7CM4b81cc0l5zKWmfA6X6cDMEVwAy3HmaEl9eSLULf8DC0xV+sp+Viw7FhpKL+B5hXo
4xDfee2USMSd316jRhSceKOgqGwxZk6XFcZeDWwkeoIZk41fnyhlEDYWSt0xVPsE5H82dVAcSdgE
iPEvUJxJrC9PMSqSonihwNneOnpXOm8pTKrmLPslvyEySg42uFmKHfc53h7AnNTpz9juQ757qIHL
cssy9KKGpAgfECvKhoaey4UyxbRu53Ap82YDCIhjuY44x1RAX1PN8Gg3yA92MpNt4JO0VNm4Eur4
F8tknTMH+LPkTLs2JMB0O/0L3Up1VTxtopR6MISeeFNiyxHSKUbufY/vKjTzFLxQS14p4kh+YbmE
lBlHxmamgEHULnmT5BgAg/7xm7dO1THiaKbM2R1tWT/jpHbRQIIeKmes7lq0PSF+O2F8VB9pnE3o
g3UdqKVJ0qe2M8ACmW9JkS0OX4Hz7Iqhn/l2BMI83GmzotQZPl3YCWNHwfJvfratTAGzIjE2SwPs
Fm8FZE+KLmIimNIq/CjVxw1Au+ST1XGuFVCL48kQAY22lZwyyOjz3Bfhq3LAi1/Od2E9LmQ52Qim
vXlFUeUZPwFEqWhqGc/ssGZrJXK8E58za3W4XsG9Ejnl4YXKWywjvLYUpq7OeQrelgwm9X0zbMga
dn6Nm6IKlkxATr6nMsnavsxNKwxE+lJyNJ6yjFsDJneUumA782lcizq5TvXMR+JOFOS42H2Dqmz5
7sIbYyvH0Zi72K0LXoW0hqN0WUvOXdeM7hYTv7O9glzqbs0IeplVAJznJsV59L98GDV/awJb1gLG
iY3d6p15Ja8+Df/0F9jmLhzgX3bHHoPG87cXGjD7A1vojcyl+FmC0Op3L7UF5gAHn3QIhsBot41z
RrTIxwdGDs2mvba73KZRKlTzF8TFfy6QbcQvxc3z9Znzeqc70nB7Q16e6842theXLWCnVhFwyq9c
fGbxyY/RFZGl21a9MVnHos92a4BytA9UpbKveempX43rgLTL61sITuFLIUEZnsrt3IrB0HUEFkOB
DoXtq3uPN5TP6T8CxANqHcSnsRkEp3Aq5QD+6RL0r9saE0WrjuQYaTUwb2C+ovkfZdrJd9ax/iJu
RVsRibgq3H56KR2icKvjESiTvMbeTuWZOjmeb0QvnSo8QYpUM5ECG52zFOAn2gIk8pRXnRZdpWaa
dUB/waWmrbv4ebfB4/NLAsJ0TsjPA5D/iOmIVd/LW/mH+DKCVGUXfh1ZnwANwXXpbnNWkO/FHblX
EaJllHVuVmT1jeF+TIRGjayQNziHVgQHS/LdDaZGfYu3gp3miov6jfvIWLbJKsvKjxfPeeTEpxUx
GLzpxMQhYVvFG0uZwkLC7wz+7R0mXJ6nUCQGbDhQTbNPc9SgBd0ZEZ2NH6Sbcii8u6vjS76t2u9w
6/mSiCtfGy5UYGZbfCuFgy5hQdWK+jMTWWMk03BfRBbREKEc0fRiptMzElu19riWnsRmTGZUo8Mi
gNlW71HBOemvpul69n6VBvz1bQ+OXyu7JsyKfIMTQinKUo9EvH9jW0sr8NCwxTIdfGR8azwy1MQU
HkId2wFtMaZrdsDiBPdRcOcximCsD2Jbe5UeKZ3DWxwxg0ZZybOGFS/rtU1nRXcerpjzz5w9HkCF
yhrtq5lJMqAy661PGuh+C7dgvmwDNEqNi3w9W14Z+1qrwQd+XmiWuJDq6yAifQ5+IXtzw2QYGaE3
703EsHXERFNzLALIdAo2JbEOT2k6G4whM3WwMbe2Z0VA+MLv0rDX0Cz+/RXTHFTldwrqYpe6J7XO
oZ9goVqLWWO7rhQk15KoL1M5Jf9KLx1xB3tcKcSxlrgxEFCViYaMMiu9wX6oTY7qdtJJNYW8NfD1
d8ci6qDGWzyAWEHp5AWWarhf81X3LPYGZO72MW4ow+/Et0qwNJ9kZjU6jc3vLDjW9czV8vczy2RP
rWOi7UL5OjujS3DU1ULbibdlZvT65S2lJK+o/A5hmiqGSpbcpfmeE1olSJyRM0dgF4lrO9Haj5oQ
fo07VWm++2oQEcwloRq7SZhmUmMMLe2jUBWTATSLJQJdLR0FPwmXv/CO8fhTqkPjGmAMHQ==
`protect end_protected
