`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U42dHjFaD3dgsYxtrKXCtDiLA8PYmxvrJNQ/lY8+XXSOByob0WDF3LjJED2UIkR3dXbq9wvyoGnk
QjjerbVjcg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T69pOnRUPhZMkvPwjzm1V3By8fCqYu/CBGsu7xDgNNb6gwVNzatlzudR4AI9xh6MT5k8D1F2V7Gm
lNCD3ySW+KkNwevpiuFaxnYBFxeMgsbDFklFonkR0Q8hUkLuUcyY2dsS9x08K838QgKe8nt8for7
SAy1DpnyzOmIbIraJ90=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U6u6c3MOL6GUwfoUzd0DdNPVgIKv1s1dJy4XBZl45ffgwQKwrrlHNc1A5lwO+66TD2Ds/0p49pOO
WguBc8l3vpOkC4etIcq9rJVMZROWQpsN+rD1sct7eikpG4ciXs1EDqIJv1/5q2yMQen8G8Y24NuW
WeJjlJyfRouBNvViTy0EI3+Jld5Vw14oM+tcImmRXC+x69A3qpdb1pLlbcHOnJwpRgNqKSarJOnH
d29LitfyukGDD1ma0nXVkAnsXDQq0T5OYjOIlFrutkflafcgxMg+tTjiV4OZ2kpbQV0a3lqIDwCf
Q8L9i6BZbPCEMyQHD8aKffc+Tr1SimWcGgzo2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2giBjjcy46Ty02thMXqYAQ1eVwrOypm5VY3Hc6IUa+Cxrp9DpPFPLWM1VJ07gzZ/vC7ftALFQZzQ
Dy0SyPi9aRpOxbW1xUeUR5OR94Lyic0+eA8HtOvKUg9iuihCCJx8oyj+tIzMfLgJ9g7oL+YqDQ3G
U4B6fPOS3KOkQF1rXnk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PdzNyZ6ywVmAbf9hxxaw/A4r9J6Sg4s7/z9PGORJhr33fapOisLKU8gV62XyUraqXRRZdXCf5G+G
GDy+7QsuIHbi5hlyiFO0xhyyx0NXN8PqBNX61peUb6+U9xReOSn3RHi3vk6zaOEeseucAZhdtDbX
YzhiJJPl1IFHxSYqqp/mJKKn5cuRQksMb4THrNRG1HPKG6zaUKtz/qfp231a5erkuMNxIDGFXrVk
bBVVH58Vr01EHVWdBxVrABfbxUrQ55nEfIcAePgpMzrEGCo1Bza5q0ZPCMWdHA2N7vbXXMMsPNCc
YEVgUrF4bPkjwGA8KEfP269v+7MyEL5Ctnznaw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
KO+zN5GmU8Wcz/b41HANQVYZLQ24dfRPVgcdwIKZGVyjGqDICYc3ZDmq5E1wOPy62RhHX805p4z7
sOAoZnjA/RqtLvdhMDk3w/Mb28RNvGlxieF45jGlQrCo1Cci63RmKM2yyw0vwjGHxL8BH5B4UY8V
2m0IrgGAdY9BC0nH1A6K6xYOJ7DVo/eQAq+Xp5HxD2bh2AvODM6kr5jz3d+CsV2s4MgGDL4qn+bn
5m+08y4xw+NXNUhsA8Nkd+ibtGxSPREbhXdyvrRihLxVkiJ6Uv5d+SsPajB90CxK8CHXL01qLamD
RtlAy1deA/uogFzZObpnqjkUMeO46J6EFmm+XnAb2eXdhR9y8rFAMcsnut0ETkyuI3Zfpiaz0S3s
x/qJkA9w3Bj+Sq7i2f+eDsDJviVxUo86Wmen5P9gV333NspSeU+VIK3NAIpbu4EPym7llIpFwSFQ
57TnZAbC1OsrZO2AWPOIIGf6n8htwunF8iAra5pX8cLNgMKaoRNZrNHo3uU35/NryPEMONbKHooy
EkFCZXMcTZznmheTe9OBmFtpsFMBx9NvyQ0d6dYzjHKfLmgaKhy9LychHCg51wBeTHDp6dqPbgLh
u05YC2l1tKlT19ObSr+SlXLNQkZN4Vp7equ3q8mkgEjgTwKAhDzE7FwlyT+tCCTNtVLnNnQ2G7IG
hraPtVZyqMBOFtMPMInQwCRY7IZq9rubnFmYyYVF+m/2ky2Lgm+vLr+Tmy8I+vMoLWBEGacK3zYd
YdBCdkxyj2HHW5zUJFI0YdPm5xl/XxUE1WFqCJQYYe0X1mmOHh13anmDPnKWj5UkWYWpvj3Yf67Y
/59G9g1XfVikz35m8Z9zAi42/CblvpQ7wXLjviROaq3/6OXyMkqI2PoKQioxDmPY4qC5e44DsdlX
OI3eLqc09Muppwl7miFPujakF1k6/E69EVG4kdeclNvJVmVDMVR1RUIDcs0hiB5cELX4AdlmUiom
SUFm/rzIOg1f0ni9HbNqTqtTmQ2aug/t3ydoRtavbWlNbkGd03mgVX2c12fkxyqIOu50xloNNsfp
USxn3tat0Ivg8LsmQJ5fZHjGkn0VoxrT3ZLcIATR/NYmS2gHiMPiQM1/9CBLRigkx7QVRg6UOKbq
SFVI2LrLhiuuLe4fvO95+fViUVFI/8VbapP5V4hCL+21XxJcHLcU5Mwe58QftNnCPNM13dSRC6I7
DVdrkjp9kUCdrypehnPqo/dqHhe3naUWD/Kf0D3NnrqYKoXRnCi+CPMb7pcS9CGyz2MCPApS/47l
hbcqTxbJRg5evjRHjxfodWePOUVxicts3hFvvWix5/0SDR6mt8+8LwC+s55lmkGsOFlDZ1kqlJQZ
k5NKcRAJd0AJ1Mu4POl9QC1AitzZq8CqNqpTzYEZgI1bOjwEm9pOtghxxz/dvTPfr6fNHkg7oubd
oj5sqPHgVyWs3lH2gYJJsxs3lHLtHqpKKryPAASPx9RPCc3MXIs8PNdosKoBsdvCZudJEvbm0SJr
SuqFK8Oj87YSfEYUvTVp4Xp67izfRUN/v+EUDUcEUpF7R9AAMuSwUvCA+BHXr/clDR/nItqBdjFd
pmwnC6m01tlGFYdRXPvLbDT3+6j12qKMipowHuj6InEFch7NFW58mJaeZ8cC00JuRkFVSGAA0KAI
Q5nWZgLI0qBvdpDkjQNgqWV/6OWCJ5XBJlrELcYOLwqEuIIfWqqByKNN2GlBs05ySc+G2zZs4Ea3
6I/jAH+Z+lwQA2exNcMi+sNHqZysGSdtx4vQJrnHV5aX2hjezys8mmmWdZN5gH9fK6+Ki2oV/ZVA
6A/7E19fXtSY7aDkNTQScwr1gYo+NoK17McG+X8GKWyqAdXyt6uZuGi+P0gJzZaezoeTbsbA14Ak
I6EECEmpAVV3Eb99HZ7JBXQV4Iem5hHNMmlJcNTGgMw3105Tun4EYaG5ZDaS0CYaEiKybURZ75oZ
SZTJl2XPQvVe/VFyBB6/6MES4ks/5VAXkylTNEofdk+ceQht1KgZRXFyvMgxRF93ErqnWmzF7SDg
oE7zJYTrTav3fi5A+Q52J5M1qefBvmCKZHnN8DihFcZd6d3sf091c5XVuQP8w9E7Ui2HTZQ4Q2HL
aTuig1/h4qSiXsKI39fZ6zPvkm4hnBeGbLbuLbpgs7YUCxg+EwiE+VllNrkG/ijzb6g7pNmah/BE
+jayP6Jz2WdEMplfCXtC+KLO158J/ht9ykwEYEA1YwD65dY5d4w0ho60L7QCBY94HZfuRbQ0/fbx
wD0pK4TP97oT3UO1rCmfPHROcZfPt/CKH1/FYytzrI0MiKAo5J7n4ClNrawIawFSQg81FuEUlZqt
IDfnvPS31JejifQ0B/yLsHzXbcWPkrU60yI3v+BzkFkkwVIcFH1zBrBSfW+lu8WAaAabNxIhxC1Z
sNe8TmGboEaKf2jn0Cc7JAYoyzeEmIv262NUFr0o8rQSm3sTstwDgr0+IfI4vHLYQtlwxTOx/Afm
agvJSZDeacKZ3jmprqsBayDVqpP+UEuqUjJ4ORdqJrMT1JfY+uuv0uj9fahmdwebvAW04gkhqAAn
IOivsjL2LqtNtSqhxWzqg2S1sMS8eRY7Y8lNGj25M9vg5Rloc3jxhigQaTnJn/9pGvb1WiP6p7yt
3deep/Ahjs0uRZqZmpGZG03jHP5QtSP+6mYiw7stECt8hsdE/7smSTFKkattncfjJjA7T2VTXp0K
j9dyONL4MNkq7HtvNxpLA+CqyDhPU5sB+Vq4FwvVD3B+p8CVu9NIZF12/a2h2aGGMaEoX0A4Z0OJ
ViGXZmOQ1Lh4+ZBMADSGRwHEkjK6kZvyGHDla7d2G9PdZprkn8+ToYLqjxgXfgg8TpChAYPH2RZt
Et7xe8q+lE3ZY0+UqThsI7XFpQSFWSEK7Lr+oZMJCalbC0wGoWSEDkxDTkVL3pu+7HjXcfh3FK6L
aI0eUZJ09oK7BxS9fz2Mkv8N5ThW9zptHvzqRnV1rEMxw9au3VFi9wgV6TMRdYBhEewBTixsqbg+
mpz8WPAlQViw35Ni5uBG/wLbljBKO2h7zYcgIJ56Mcbyse2heEj3X+uJw/qXOYcIcZqCEXJZ96js
PHmmOmv+1RBwU8WhcK34dv92YTjLEceXiCJa49CjbFklCaghz8zc2jIsUrDXUdJSwedzfgWpo6Ar
SDwYlpMttn5HrSpp8Z9g26uT8pMdEhptJ7KsUnUHFODmPAr+KwTIUDT7RT/NSyYFHBH3St4GbFNU
oR5bxwQWxGAD/uYtXAWLVRNnzbVTV3BRceozSjz4cfTvqn+zGvbTSH2Wqk2iRCtauk2Qp9G3QQEN
gGoaIsHHHOZyiHEFCJ9HnxCRDaN9I38dpKN1bqUvBFwkk/TIUkU+NYM98klowMpiXQ8+iNdUsWt7
NWh+6qw5Y4QjObHKkUGd0F8gwsI1++x74vXn8uaTA2eJZhTMdehquZBCrzpnibktGMT3dSss56+Q
gWglSjFVUs2zCe4YAyEpfVLuRzbZIeQ6pvxMFXM1kcnpNzBg74oidIDyV/Qb7Maqm1hHv+zcxpFJ
kFkz7y6y71xwC7xbfAwp24zlyGKZF2379s86l7PNSX0fVKBJVWbsD9xaV8MZLqHCLlSHBK/qD9zJ
J74Z22rpjp4hhCtlZSMPBSY9ZyjAD7fHObwmyHqkc3abs1tnaa5+um8nQh7GeLhLt9eJhpAt7HXC
IvqQboqih2H6Dd+VoJ0gJz1DPXkgjbVw7QzZZ7Ycea8CZMLYTx73CtHXjPZAEjiP+w6a0wNHtiSM
HTzNsHrc9lsegUpF18L0ahjzVLpdci8OWANTvCv0DCAdgCAK+Bg4SzJu50yhNnOtxQCL/unaMS5I
M8y9dYxzbgCI69fr+KO2uNeZQgOJFE3sV+bK7MNchPiRNwplB0mVYPHP4OocCWaBIomUj92C9Otl
Eat6es0CEiFDgii+y/oqc/wqs+LiHYfS3TKQ8p12lIX0CoHyu7FxYR+lRfygdr2TNyFhMwnxGHZd
bNpvK5vKOav/Sd/f4EPZAKGTrUVvbJll2yTyzgatRjKL8gBUgx7c5273PhirZpDyK1gcQVBEzXg6
YJ1vVihwd4qXR+K9ia1dlvf+UoFEdO5PABoER/JjZrY5ZgCx/15IZSAkGurSno2ASC2LePEkJMhD
4v7QogpAplDslrx6V0XMVS1+5KLKBwibWP6Vt7P5dGzOE9x0SrdPVGonnOzfZXJy+Nz+/GvSgClh
PDKwD72ha8ljdUpg7emAupT8ho1Cb9/FtL+SeNa4Wj61vONizHgAD1YWpogwXLivs7JpgyMZhlyI
tZkCQLpbcb67tV5HJLAW5f6dJa3oKhjM3N3NFG0KPsOO+4tinbCSZ6zZk/g1Q2NbsGKV96y0s3Pa
YOTDLbgqIUG482hF9wBvctR12JCysYR0iWZjWDNTJwxaZKUNZGZIdPhv8Xw41DSVXBISODVhSFLd
VxxUk402XpvXyzmSWu6GLDbtPnIkvJF5a2K/8Kyoch8dX+uefvfjM6sQYjnLKxGmWmGaZL7Ufrm1
Qg3SPyr3858yxHpwwJQ2GNSuw6vlzMKK/BNRkSdi9R2y5xjdIWoMA4qJ2Laax8Oa5Lpkohu60kYg
b70uNh/m2dgollPeeY+Q2VOS4C9yN8MkPDJE28863EEAIXtPb/thiCtNeJGyapekctaunPUEd+Kn
wANroEuaYlO2q3y+TzoVQRav8xvnqwK/9zsLCD8p0ChLCyxKl1H9/WoWKFNG2mcCjoPDHyVimKcR
Or6v0x6akRVloMfL2/x50fi9HmHXSNTp8Nv02L5pUth5SnK4CEQnJq5+4tqvyFf5MfWipbsGs+hD
3X7A3L8GksOgxgTqnlwEukKEaeLU8e3ht8kfaByVjbRqTLpkmrb5dMOS8wLhkz8MbosSbD/wjakf
z963BJCDg5Uo1UYNKXrc2/gmGSnhfaeWPbL+ohi/Swwn9QP5NjJljiNj6WlF0tvdN9m2C8PnDXfg
X6fvrEMuSvkD5WfqHj06M+Cppba2lWlXyFKa18RbJvp/xvX/ZvAQiHRm+mN2JSxd5nzZ1Ij+OWCN
6Q+jnSEXu85aQjN8Rce5vqNTEg/m/YykFfZBoN8QF2X+Xnk+NKpvlXQYr2TuuXuvn/Z+FxpNeAh9
MhtBT7ViLBNlGckl+L7c2u+iVvUyHgjy6RgWPoyih3jnDO+ou9P2mQh/SLD3vcWO1j59oGFKP7gd
jMSNgRWWhAJQP/EjFXPdg8YRXsa2BItju8K1frLryNA5SJoV4rcan7hQBlXTJ8Kjjb8B4QYgKeeA
BJzHj0xTOrJVQAmA2JiV2MErkXyghhCB/UETeyaHLhAtvlHWOzEktxdV5layXrkJpdaXzJja1Khr
rpw0JRn0h6AdpjZibI6wQvI+2dGthAEPKqJQtW9cLFuewYK3cs0653QxokSOE6iK1RC9LSfUjYpZ
Qn3ZTcx6TD7vzQvN/ONH3oVt+HI4653xu8SmZyT9ribaiSFX2x0j2MUo5zG6TThbtnvVMQ5qLjNd
m3aCvJ6XwtQ/tpDX9UvewmzyMg1Effhk+K5MYnMzMC9MwNa6TOOzhUOWEaW54v4KD0A2mNFwIiar
uxwoBpVpA/iZ0YS9ewBeIlAd7QC2Omt/Y2CdxYSL9MDFSDKtYeBZ9ocQh5cE/tEQPLt3E/3jpnen
SUwY+7I/epB5EufIlStypjz5XSHKdsYlUr2TGWk2XOO2vf0dez1ZjVCuJLOCr/fd3k3oHBHFvrxr
QsQ3Bn/6ekdV8DO/3uwMApunCoa18QNjizmpzYVTx1o+uqsCyGUD6Sdvss6CG0GUAxkXQi1JN4K7
6FrAxHGVtk5Nh1+xIH7bUj5ANg5DF+YpgCHU9FkoVZaq/8jHFKH9UUeaL19CEhCuYXXDnPuObqA0
VqQ5zqRDixxjFxAMztOgbjpQ3LgFG2na8832WyfSIxcoG/K3vgbu8sqye3OX9gAgUEq7U5J6+AKb
K+yDitOxaqJ2yXoXdAdiTGqS5sRCsHE43xfufdEbA3XH07wzz5fc7olBYRVfvSv2fou505imzMMh
3Ku1p+wDrCcWH2MCBgu2Mwl1xW/n55Mx0IS3Dpc+/OQ7RdsIQ1qmA/yfcq0I+SxPvA1cU3vi2N5U
X57Xv2dUDZMMycE3j7zSV5b5SZ8rQqKOnKSAaPzBxwh+dodYNecI3occnWi696cQ8PRbzOtR78MY
Q+ai9Qn/tEbbOmI3HJhtKdiZOPGn0kbKDFwB92zM80vXF9hPKi7rSM7MSSx+8GMsr9wsRg42YIda
x0gBkXuJ97zeJ9qWfzI0U8sZe8upriRxsIxap9DjkUR8ETN6LSawFpTWAUYZjHydljltE8nSZLZZ
EQJUKqHCQF5FAUwmEiRpWYq9LzcUcvqCpDtlo666FL0dcphnGB7Jt97ogPudEE4XSyWQbRERv6cC
zqshmcjMg8yk0W0S5b8VFMbWpCloJqLe5kvbeRiGIdMTPPyg9Ke2u7Xq8/HoGvIYV8DWteR5/duE
Lbfb68Jrth2RURL5WssIX5+83jCVuJZGHISIiGwj+bod7Nz1dkTENahxcecAWKnVAYLqcIycvHBC
bTOYeFOtirgKIulDyK9CyQ9IwF976Bcc4EQ7yTA28Nw5R3U2lU/Xlk9Or54poVkXM9+9LkSZFeTl
gdIsWUQcLp13hg0Fq87Y8fZ4RyzHCJhmuie9018PGXTJLnbLuWhajQQrhgU/RUNjfSDofHLIJ/Lw
3HBU22VtGZzy9ppauHlh0saVcznwE4w8hGIiy0OEgspJ1jlPXuGgm8icmgTFqgndOSE/uvcbDOmq
Cgk8m3RtZMLhx+VQ9vVQTeM3a7HJEB5CZjgoE3g6eXmOqfpJXDYEQuBiEr8/rtF7sUzAyzX7iyyH
AKslubeQ1hiHadrV1viJgNg9K7Boo1t5LQHu6hUc1JVVPacUYhOKuQajFfvFFWe2Yd8xXhsYDToS
6I8tdfntw03BWKcJpsbbyVnvF6SKId6WVKkER6vVkwA6bx7m2F1aAoBmXHRr8VbjY5+gF3z752fd
aGxB9ooJE6qsCRugCfmWxnTwz6+2WbhbMkZIrWCdLdDu9JICZCv0ravN9spC9uePRnra+zQeDbdy
4AkqH2qAL/+RW/ZRhzvmTIPcC0H5nj+GHYWS492TWZkOGhGUp4l5J73wc4NN/FAzm8eLUhV9pA1Z
Mu00+B8wdGPP0vajNenwF4kajUFME9PMkMHH1iKIPQ585OKCWf3wbdBWsMgzq+k3INyBsh5pFWTd
PS7UDaB2R1XNEJHMhENK1hzaC/LDvyy9IBgrldAwSmDNb0PGHV3TLBEP0KGjCIxtDqG1iGwYyhUc
7tCDl0+LED1dRA5+hY3Lc3FWRez4W2Yk1U14WAg72L0c9sPHuLlSK6Q3P6y9i+Gkb8tExhGmB7KL
98gg5a9h1siS8GsHSCbwtQ2GBx3XrGSj081sajbOK7BwZScf23DLdl7spsdreFVcPQvBeInfIn4h
h+fJPUujqrfhGU1l9TNhhen3DVFKrsjO4RQSJbM4xbyPB0QLQLw1nWB+rQ/jAczxcxFagCKavwyy
p69fdRdNBvLNI8Y8vrd0e8nAft6oJG6udAlLkQRWhDc4sa3IWId0TCum0MZQwoK7y2ruQVM3b3Kv
CMNka7qi65dXdqGbMmxEf0uXICh2zkHLkaKiOxdeJnD9hx+mR5T/5xqJQMb3U4h65bhS8keRK+Jj
i4+tGNh45j+MA4dae3BCtlh0MqOGIShM9ADBv3Pl+D9FIWWm+8cq7HrZ4dVuxDl0qcFtLBCEOC12
1THLJoyVxOs3Qw4Nx1ndjxGq3qy/UgmW7Qcvq+hBuJne49c2zGh8VGUqMX3SUyG74lmlNHuJhAAc
Z1Fsm6p760ma97J7xoSNkoEsbRkcY59H6J1iw/3jW1uiN/FDdqGBDx7juntAx3ByYnyra71JcQzt
S6G+ajIcNEIBO1dDFBLlD1F8USiA+ZFXkKI7QWonvPeW3qNGmEy102gKL8vaTF/wvBOGMaYwqM4B
61hiGSA0n870HiwnLO5lvYm/Yh8yz8+GA0se8QCxwgiuKTBZ49KdnXcXAfOWMBnPbJdB0mR2MH1w
0zvFeDMi0kjI+bvCE7Zs0xRPFtWJQTtT2XCI1exxQn1cXtVeKq73T/sBDq2odnjKSiVmCAk8uuoW
mx3lsqV3KYHDGz8NtpQpTL5gSSvKeU4b9NEyr/GKyyrw7WulkQGJOGL/TDmXBXee1ZvQ5uwEHlEt
JJLlpzzDd3dody/h/I/4zCNeQnHUnvTCS8wls86+IU1Sm22+CsxDTVa9WqC+JXJFcvFoxNLMz2R4
+x9bfWYcMryhfygelVvWtG603FRhTxAkbDI7bhzTVWfShi7QgB+4JCQURVlEQXaDI2WHqJImn0pY
+bJmR74/VSp7LD6cbHLEU5zujJRl7CkhGMdNPoKCJSltml+SVFNhZqVJEeYaAHIcRJAOObUMc6st
fY7WtuG9IQlIReNL7PL7OMxDXmOru/1OB8aAOMmxU+3ugHlntMjclumLkNwtbMcAQEawY4L6Y2CD
UcHdrLfc/g3M0mCFdKkZpSMa2m22jqTz5qOKZjV5g3AIf0qQXs2RJ81UjUubSMbWHLRXQSugwXxm
2Kln5A7mabnspVJDrJ9peOJDI3O83kF5DMlkQJXyAD4SSR1X4Ox+h0ZEjBH9l5JPTTBiOGjvCRE2
gOSaF/PRpnadw9olqnUvM1uOlX3JFy9Ex+etwRh/S4mWX57/L9gKmby+NNPoKK/jjZxTb7w1hAYb
Pl+hNYCfCDtKlT3tCVeOw3ear3MZQ7ZEGOV9cHo6zcAcqf3qAWeqz4y4JmVtnOygcPqdTs9opBe4
IaH5ChxMvNEJf5wopO0hw4w/WUz7ciYOM5Ldf9HXRoxTzypoybwwvydh47sYAgIExmlxrAIB3+21
IP/sDQCr6axw6Wn0c/ZOS5Qe9etnShkPzWrnHbzNLQaKzFFjpf2iPJC3EgylNcfJFUioFzPS8P9X
2kcGwK0P1llxns5r3g5woqYrWBPz/fbxKOdVv1FO21HfCys+NNV0Q0Utxup3NE8WCaO5PHt20e5N
zP8ie49Yji4y85Bav0ycEusPpEn2C6PyQbndNNa0rU3e78pssX1sQaImwtWsV71JTccdCESrRDgU
bx3IXJlZZLygebLvDgX8DHyxKvBIgE6uMZI3V+9cA/iGiUDWMkO0C0rkz0s2TSQbD/S2esHnJt+d
rdNujRTISaCeGsjLUb9W+HaFDP1UlNLvSWRgSNWqo7UHYoWADLVtmK1o5CViJHAsy2ac/G3CLd1t
/oFcyfdv9L83OOQV75LceBBR0l1zbs2ZUDX84egTkJgtVpmwF2s4/A+Lk51KgMrPWVjhurNJmODP
967qvwgx+KQWsUeBOtVPgbl8GAUfrRGThkoOq55pMuIDcBtKs/O/Hazk3WUNTSCJdKS6M2GYA3/e
FEiZcrWxH3zQD3mdyc9E8qSkZFKKo6tmNR6/w5+/tAcJ5McWF8anREP3dVnbjCyOeNhyjy7pyyOm
CgzpUy0tSRLE9Ijb1gxXL4TiKvF7fW9kyPK8ZbbSromrIwqEl6B85PjTh2jC45dL1EbSoykeVhFs
t4dMV3XU+8GPkz/uYCDREbHGoC6y5viJCVJrNa4uJAmI5grAZvEGzT1TCETlxZIDK93P1VzBp98L
viDUxro53WOAVvtPAKLeN3zt5tKDQywcAjbSz0HbqooLHagdE0GZFS4uP5dQsVhl1D1GSdP0a/kh
f9M84oKU0/zeKBFYkZ/os/SR8Mmw0DrQOIotr6+NoFtzADSQy1rSsu2l4xN61rrhnjPlKWXJlLXe
Vlg85uiGzrgThhq/F/6tYr7cKInguK2MWEqCJeSgR+5wudmhmHeq8FGz1t0aW//MnifpW2od1zkW
TrdBO8qq/Q2dFuwbF5otZgm/t8IGaEnPqRaiWdVmeLKcPRKA9AAcGkMqzI9dsXmEMlU+UHM/+9aN
x7qZRim6ixvLfl9/IIRhca6ZLjqKvbv1y2tjvu5KRQgCZeGhGVql8ibSoP0lc6bKVFnvCvXrI6Xg
MmK29MrNaL5wuxV6BNMZ6XfdXVwUGjth8TqUb7BpaUS2IRzBzsWHQyMnC066wybFq3KB/jPVynfD
KUqMwbW/cZ62jzmpkkY26f2sX6CD/8UauPhZKiqoyp5eSonC+v862BjWmtPuTkMXd/CxujivDbHA
yMoI5kZZqNVlJ4LKzxseCpI8B62271h0xPN50I2o9AWsUXaPBJ2NLWFbmkyEC6SEz8+BcF55NVyI
IVPfK4c9MEc6Ua90FxNojO1JVK/fqh71ic0510vCSRAJ/0Hywmkky24aqdZINk6vKrnGdBtQngOU
csYjOf2L3YIcgHY+1VWYa5qGfGfVBkhah5ceNa0Er4FigvE4Rexc0v+62XbD2rZHxXtfG7fGVDu7
1oaRVYO3yMQD0VEnGrgbJX69XkWWXJMA1BzMEMSiFImtbxp6J32mEyx7XiIUNb/UQ2vWz5Lx99aC
NzZej0Zfa5NeYIrRL2ufKXUzgjpPOqcs8HyfA3TkQOr4TuoYDKS3eruvuJBMD8SIgwKWD2Za4Az0
9BPe652G9sYfvf/6eRRTJBeaPKuhAxjXBgucMOVdqChk7EYMHtTEQpDgr8MmncYm7paNQo0gUuWr
U2OxjBaobE6dPDf+kEgZBsGl4Qa4UUlERgk09VbEeqt+30I8G1NWnXERHxps/eZrS0Sn2vRNIN84
Sk2MPdl2EwD4XScu/M0xGy70Pdta2hmNX3JzFYGrMfCe6AXW1g7UyRNqH0lYjT/jzpxKUeqzXfGi
90IO3HRvSBQgLnvkLRwVPYTC+BcuWk779m3swNeePGBtfN4LNiCD/wlKUTZdbqK8V9qLGlPrtHli
FA0u3tL580SElYEfu3txtS24G4BzvMP6lZh4kUmJWrAHBUyG/1IgD5Rlfz5O3RkZZ6v30TE32dYl
wmFBw5aGJQw6juC/P7fpOe1dQvyh3sD6dfbZu4XJwaz/m/t9RsK7x5KDmCCFYHkSUBNoU4ZMo5Cd
M1v1frZD88KSuhYXe7UbAeIr2Yo5F7Z7DK7XfheGaL8rIA31GUO+tz7Fo44ez3HpS2zIt4skGIZ2
Txxo52uaBeAFWd7AEBHRoUGoS13gWUUP6W9tT1nRL6zV409U5THvwqNj49A17e3RAYcmSrOq/gf/
mzGK915IF6LvgQ3JznAa+pnG81FIBUkew9qmXtF235HkL2t7QZ2+4tAbWljW/dY9LRP3s03yZAMI
yOvrtmaoPtqnrCo+zkwuTPvufly/emK0RcjvkXAj5KMzY5fydLXG1x1RtqQscAaiewJRVSta1VPE
4IhJznrwZVHPu5rk0m2R8h+wGgiCGgJv8Y9TnlX8MjTrjhEe3jmuMRma9q+8UJ2kHTWF8OnVhyOO
PqLfPCLc50Wbqpp/f/EPxycZxvvr4iQG31pXMT6IvJbLLvcl+qfSJ8MSJ9t8qHoXoZFkkEFtaceQ
p1iHy/JYXBAMgxq+iu6y6uiLkUoY7u2i4l8lJ7BvCddH82r7c8zrk1vY7eXw9tuYGxanidWqjTqB
hlp+6NTVjS0S+gsfeJwH/RBTFfxjOfW+SEngGIHGm0AdS7UbOOgH4ysL/caT9L2zim9IxkF+MnEd
rv/6zaulBTyt7CBTs/hgbcClOKy2gAbglVcopDiw4ly6h7VhI66f+kpJiIRPFPYI77L/O4k3gIif
gt+s3AvY6JNV61EPJvjnZPyUqIeeXB9BYl1HIte8ZRhSHoRLR9PYFI2iL9ti+s0WA4vqmgYwtFl2
r53S455LBQmCYVe/lq95/FxcKBARnGWTcHKofqZ+/Uus14CTQM89NJGndVAbvO1s3yo7/RY8IqyQ
SlVu+vSUFpFqS0RahvDEvOjlNQWlATXSCv4WNOrnE9uXS11uILbC6AvVfQQTlKyTY8wDVj56TtjS
nn8d7OnMXGCBKiEfc3xByv1hPVdeBCZFr3hTjo6o0T+Ku29HkTj+8AQ+Uju8OBp2+n3jBjMHwsSD
R00FFugki02SUpC5FCdvALk7t0hghPya2DHGUf/jShfMXzcd3A69xAmH49Sl3RwulPYogEsxNHa1
iL3XkOnyP3p5i3x4IUi+zu6bWhkYik0HdnayxOnMjyajlHDsmwc9c/ZmrXH8G/sUFSboFL0PNwoA
Kc/OYXr/3zxi0JaD9xKHjY56PQsD0C8w5beFToel+xApJrUuKMbBMQ4ThkafGaA1TijVWWs5Gfq4
CTgm3KUxh7CklRQiWYH6nJ249AVOxgBfBUTmeXfqqexkbabOFcAgA/rxRGJRm0PgG1vqALfCshti
q65phDpq+zS2+oYidrtMwXY+OxAZJNTO42EPZ9yWfnhLKcsvMr68RYjANYCqkcygmIwRTdwbxlFl
K3P4bS19owkbKjpRCfTarT439AN1F7i/27lJI+ToptbE6hDXWL0MatQgvfyojlHQIsGS3H1V7DLB
FZ73JaOj2muTOh+kl2tt6snuoBS6wgWzDoLgSGIDsNIdicw5qInht9CK6C+KvUEmHGgdHToNse7r
+MaH1aexIIfogCccoDqv2wskDUszqWjtmqcOpDH4Cbr2q7fDEibF2LvRm7R3hctVVeBXSDXDAjLg
km+/Mapte0aYftvxRtxDXoCFp/y4ZqK5Llkkq1t/J73AyzCCMi7a9H8P3Q8jJ1dAbX0PojO863Os
Qoy6MRimfJNVuVf1pN429Fw47cNHAJdWogMwJrn2jt1aFX9rIZUJQtUHABb9PYIUa9TerbCgoZNL
GVoak1GE3OOxQtHkVh5ZxTaPxcIflhKLThYdOVsIN47bGSECp0STyd5tOl4kJUN6q7msKkGq0PQc
8U0abJ91MPSsx7UW10UTz3NqgnHN5uP+wvE+DW8XFGAYriuq4OusNQS5e0bOCAN6DdpMI1o5W3Xn
cTRuWty2OUIBNmKdLOC2NV5DfDFGhpqtvC0c7G5VfraE9Gmd2IyO715ENWEZLcjdNS69C9g5Nm2K
S7/EQf6hkcRwGnzLw0rBD/XlzJxsh7QGtKxIcPqBv7aEQR4yLdN7P2wMygsuyiCyNk+Vf+ibuLZu
hhwangx0rJaTDxf1lXf+LiOJlbzhMzQYQXfw2uAQK0SklpGhaHp3nJog00ahE9D+yqWK4RnyPk7U
LQHJnpAl+xpnEGu+bRMTCZmvQYlx6QRunzpWp++zV855keUgPJN33bv2PRwwV/7IkwuE2KSrx+gB
UBwawH0ptEfvyalUUiDjLDVcL1JeZ4bYZdxjFzEkbGQTlcp39Pm/USGNoB7EPLtfvSZ/ai6ZR1oG
1CAP8X1lSUV2K8EZrquRljC6aWmRlTeqzhx9ySQBL9e23ErQ8yTLLGZDCVF34Ure09V1vH4TSA2m
YrIfowkqIoRLEIk9CkO/Q9DF0nrQdLXsOIkqRFMM2t8oFOwQRTDZ/PvlWVbu1YysYf6fCR+Snuql
uW6bF7mYkpaQn1e4b9rCSRjKrxrEF5BjIJ48+dEVIBcg0iC9um6WxvaUx6Owi3IBzfOy6Vv2POgE
m3Ggp4F5/OQkWyFbWy221lIN/WzCIn+IRW/UtojL9gFscwwwXJP2JsYNhmkezjFHW7fiK6RzJFeE
1V0io0b9DDx9PEe1E4T67A3SgxyDOPD7mbwrtRj/hyt/0oibQJwmmi0euSPDN48cQcJqZPEC0T3s
9bbZwz6hB3pNieqnFF/dj2+rcxsnGXbjYfXiia4t6/NqgCbe03Qlc0tJ/3Xlw1cVWWUoyHfqEFWk
U6itOR4fwnpn/ERH2z+uFYM9of0KWJo1K/uHXetHCMAVc9H5Da6l5xoZIRdPV2o/dopsoqzt2TQT
1GP6EXezpaw9VMbLIonx0/8VkcOUwCMD7c3irewGcPR1+6xjanO+dS9RJSH2eEEkimJuHeUZEQV9
TEhN1xjWZ9/5mAfPN38R8vV8r0WBCRKoov/Zy+j76v0/7siuxmVQwzzuLOcA0raqlzo5MqZFyhPX
vT3oMWTi0dpr1f94OdkbIeZripnyVNpHd7HfqzBliDe3OfVQo7Iukflp1uyL8GhzRMjXFa25GrxB
/Fptge5w9MNWH70PUkA0u0MWj50O3BiityroJ2EG7wDWFHaW+/n24KpVLWt01Gk5tYzfDXj29M7e
IdEs4iTf5oETQERL0BdKmDSr0+VfBtsNjJStZnD1SsA+t094f7wQ7NlRImwAdiiD/BJJZt1kv8Ne
t/+bKGjVsY/mMVvPWd0yMWitzHWPAOOUqR68wl86JwgXJmPcyBWGEm2OemEtZHLGWFvTd+hxiZPx
yrd7SL2etQPk4mnIZCr9L51kzw/PJYfx0bb2RCYLeQSBcbOFePSEDBvLn4PxEFV0B1/WQrWwtd+c
NXxOxCWyL8ITyRAds4kO5VmQHEnBpP0fK7TdGRxioz8IQjU+NP6jzKUlj16XEqCWBKWRclhVEarF
c4Dm0fUsIoTPz13ASA7iv5JEGj9+B49U6h4SHazKDqRLIf8pRVo6wCijPZ6I9sbw6LU6Z+3LGKdE
Ie4iMETjiXT5079kOatwiQSZTK3IRpQ1Z3UxiW11j4w7mKQeSIktIvZGpSKj5cScnAyWnL4jRTJV
twjNLt+IL+5gI5Hva0ed6jTgD6zanz+pkhYcUinoSbPbVBMMt3T9p3ikI6reSD2VibiVoVi+3rpP
lkxvhpwWphzKkPvZJVnf3rIJvybDACdSMbfrUiW0irpuG3au8h6f27deCKBi8qdq4b4g+KY+d84i
Lshk4bNl4uxqpwOD4TltJjUxgc9sWhDnMU3m+aO92wTh7dowFp5GcFhi6AevSwvVry5a2f7h8iP6
RrkVrTr1KWonzK4La59ogr0wBDzUXFI6xprBNTA/iO+mUp1iKxPfzp7kuK/kMcfb27MSWXtPbrcR
geuIJmkViTbsBtnK0EBMPcEis7xfgbPLWfwEliOEsOJaQ2kRo9ZRk2agi0ITBIAMaP+zkMC18I6/
cEL8M3cs0/UqiGIQhKPkQE0vHVrA71Z+BopTIpsjKfA/8M08x1bifuyuieybN7oP6C/dOe8xIit3
4g==
`protect end_protected
