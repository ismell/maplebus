`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpIeCp0eEPDTj3K4Uv1riW1H2tnuvhS05btKYb/YEbeFY3QFo6naj1wSotWcBhOEG17yHatKDut6
7muS7y6JZA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J6hu5EOU+eo5Azqym0gz1IN5zG5pxk4nC9LguQybDiiH+Z4ynYQn9eKFZYZP8K0veFCTLYHHefsk
tpngEFOui/ihqeYyxhal9dg0LpElQF/s4Y8K2ySnsnGS9VVF8XUr+ZCUtWLLsnKR3SAxUC1XTe0z
qf5mho7wWKCSRwqtfD4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BFCljXRp1rI1+Y0U2Z/ZKGyt38cgLBhNgpMeQrzoYiFF4rXG1yCthnFbJ7jRRp4vgguypYEPk+Ed
GObj4Sn6wPqSfs1SnMzL8rNbrR8msNIxK8UCbPdC5eqH8rsWiM5F+PKHQBeH9N5jA28qdyAqFJ/h
OrFpv3HWMPWXMr0gCC3SHKypr7BnrpyFG1LGkz+ZVoplJFem6O336evvaFAuW2UlM8krMZXP7KYX
shJ8+0Sh6FVClGFZsSe1aS5vap5MNAFsxCUGSuV0tSJEZSWzkn0H75w9jmLzIRcLc7RV/MGnq30/
V8tLNmYKQEWtVztgNG4haBNlXOHTrnif604dSQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KgBY+JElMQLwoy/PHQcKPX1kBJFDyy2cOmv4EzEzrfuSU3jJut1ngnxyvuUV0cdaDdHxqso9rYM5
gyO1hvEgFdXq7eB3Xt69j6Mj26It/f5wfo84y5RPoDoT9i9wkeOFFuU9c252HCvGgmVUMRXP8aTv
+Sr01GDHoJX2gTv0F9c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a+OcNnMEm68meW6uNCVGL8ZpZIpHA2bFrE5u+qmk43LRhJ2Tm96hYzvERSrOJzbP0xIgs0OesVqp
qBJA+Ye3umQ5IqW1bj3bygsOsKj+TCRG63Tf7CFEW0XSpcAhRWx3zkWXjqqkFin/hi8E6QcYWGTi
z6hxvbHbuDDlnVTaW3gXo2F0fENUkzpyM4jWQ2ZMtadGa969GXdREVae8l/nyyvC7kpP/foxA5B+
9XBUSlPyfdqN1iBkiUrP27XHuepPGTaJwXeed7HWKZw7iMfiYGrYs6pxFF2ehPB8vbUgEMmDtMJn
jweVLgCYRd2oVF8JcKUx6PbSbKaY/QUByjN6nw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57600)
`protect data_block
1QoFWtqUimU39uJCMStg7ejwnWxvxLyyGtbHgfBXwqCRtdswxU8sEWs5AhD6YW4p0xdvGcx5kUIu
7hXVap8yUDB0dgXR6nLfaenXNTSyNyz1Y98+QKGbyB79bbaw8xyxxhQQB93D3e+4j63FyVYvdkno
I0x2VnSAIIGxyJFR/zIzvsGO6VmIbIU3XE5DnJGqUu30ZsQ/Ul3IuaS6juhurZkRao98w/dXEUvm
xdkhkqBkSwoIGuCGGWC3CqxXXftLMqiuuW6jmg23GaNd8L5PlGPIyQGbm8a2OXwdaWkch+QpfSTK
uaQMPBhWwHkVGfGQfblXIccphqHXlQWJmn1vBxIQ+rOcOXDAjjQwFo0oxXNQ7CXblyvRAmhqqgKm
3cCJUJeElCmI9IgMvix1hKvaUOii6KUkalcuAOgHdJPw2BKCo47kI04H8IsR+3dpbrIO0lUpb+2A
UVAT2+5TH1rMoaIoDqdSh+xNpiq7PDoUIHhivqVngd7y9CXbApZ9766hRJkBOfFhQaKqRS45bd7/
viB8LrfReH48dKZeXljSf7ZB2CwSe1xONpnzAPJUsSH3Ep1ekdBC1mT1fry/8Hk5WMsVQUeQg++y
pwUhy4DRDvnbcYmwakYFkcpdw6S3WsNSectTvbrnGTFNLoRNccFgJpSi1P8V/1BPFM5CoIgqzMK2
ylZG/A0FkDvSOmFK08JT9+fzrFVVShTBF9NemHMXvCFl/Pn9lwQ2CLgTy2VfBxj1QnmZVoWtfZtH
lyu7Ymgbh8uoWFegHAMIHtEzjPMjUJpgqtM2XpYYNsoxv26q5cJJFjlNrGS5gdYho2/Eg+5I40oN
2l/8Ao6KBFyEYvg9G9xZV2xuVITD4k5dKiwSNJEQ+a5cpeYWdoRRC5Oira5I6+DNi2FPFws/B+5z
wSck2mXPFajtXMMw6aAzqVVY71skVApoMicHHZM2ahtuVGapXcsIzCgv3xVkKoxAaPmn38Op/UEo
JnkQJ5s1MsIG3aJVWCwI1w5z/m3QVwTvBZwTOIhEHu7/gjIPLpSk1jo9F6NO3Lx9DBaiq0qCnWKG
wYcrKrgfHBx1/TRpptMMiPV6KbwdRRO7LO0yCc59rnQdEydAzCThZLMLnQTDzwCQfu599VgUfZzn
QXAT6CqrmoTGw1LHoLOKL7T5pwzS1mh1yFShK/JTIsuT/O174hVCQshXskfU7OapZSxQ+qIm/Opz
pwEuju7apT9/FcB3E8imBAg28S0v2EPuIItKnsXxVaywm7t8GbivuLxssh8NQyDOpvAgv7acxBmI
9BZMnP8iBjLe2iWahbLPRSEdtRpRHp9k8b6lY7bSVdGcQtHt9mKJeed40Qpf814ct+zwbeeCHPHm
9NXCQH0pmABOErhHylSaE8s9x9Z7f8WaCx1OGnk5TWU9sxd9LnTG2C5VWS+Lbqr1ht0C+bz4bkCG
AxODCDNwjq87n4eVVDN0MFXiNLfp5Nu6hpB7zbyLKMrOZlPfpEcsdGTI8+FG5N9t9fdyQY3KLyhL
96vClu8Q9CHcMu9E1GtOgiGnf+WvtOcz9mVqDQkeT0oZSwM1YJVJJLZKguuX6TiwZQ4t9Q5nyvKd
oMqKT8CxC/1vFWpdocq7jCohfEjt12JUiSXi96Usb5IPQkGeKLOstFF/S/1oeoUDQXIriAFDfhbU
CDLgLSvtTT2DU/76D1HxPV3q6Ok725uUmjk5uYLW+ajRUOuW16ZAkbaaCaYb6zrUA7p3dk59FF0Y
w2piEAdcMAJIErzX5VHln2DQbNr3kenIVJmYU7J0qbMw6ARLcJDT1mF/Ka5ji9HRTs3kVDQFdS+k
c+iZ7uAUR9o+8u6YTUloIEZVBrre/5aJ7ZW8d4SelBQSOzvRcr9TakCQ0OC7jhIahv5VAQz2EQRf
wNSv9vF5liVccF1J3/D63fKAVkcqlASvVpt01yCpTztNBeplftQHXtMhIT6JSXVVMf1uX6wfbAJc
uBZEBod4a/H2bcM9AeRS1rPzqzalm9HbYk++JGf5LLzDTZYZAcllepaBOoR/fcq3FAUh132n1Ggh
IT3QEMKhdmTQCfe11TmUjGyNd8OCPMIHuA7oVdDeELt6IbNKlUYO5Dzjb3MOePEocVgc5bvumXhK
LlDHu5/0SGTKNRaCNmpS54QNt2eKkOI9wZBGzUBWNA91yCBUOMJAyROCLGSZZ37Tw15ii8RJqTpa
k1DLg6LUXRQjaWG+DKqk39RWf5nxmgYf/WQCxggJLTzUHdPR9FacdRRv9U1zJ/rGWnla3X7w7Hoy
Zso5Ky5NE39+LF0RnHoHrig4QeUJXFSlS1sJOu9grwPYXQLBO15I94X+6WcxxdwB8o2JXJjyJwhP
OGDgL+DWzxxz5Zbd2PSdUNeppyCgL2hWFsPtG6mK8ajJHbdXGzQRsuNiTeGDPQalw05w/asxaqS/
BUypGoIaqYbDit4VDar67lmwwpUjNX+Z5BGJt0aDPJdyP2jkcq2B6Y4AWjHjEnKuPkhmc0Hm0jTf
xC3fWr2tJUbLuYBu9PdE5CNPSdE5vy0DwME5DI9qlPhqFo2m5c4lli3RjjDdRIBBl2ncUnHxo9qL
ulrPwNvTFOfkPyfvNZcCEHP1mx9S8Vf6HYB+Uq3kiN7/xYty+mJ2GhSRh/ULolrOC4PVr5Ebr/8i
pvj6J+P8PPJVXHFUhpAsI03kWYMLy7vzFDPOEHikER0d/U0/hjMLuzGJOveo7DW+1p1uI1ShIqUr
2+h0vBfCyNcr0TxI0RewpqiOFwfT4e+8OHOI0Y58FtUsfYgnPizL+9B904qDWoVF6tK+sfDqcMQx
FLlgBlVilSz14zWtWROcgujiuwV6VVlRJK9DkFHxRE7yD2Xy0ojY/pbXAZk9ZX3bnH+l12Csd6wW
YwEQGX2I8/PkttLFXS8DmZYAs3Qr/8yhpfdleq7bTMjg8Fh87cbAuL4LPcIdXgPlDuNkTniIPHVG
CrSOAjsfhY8fNjWLFDUT2fzQkBozEFaISU9UV+PSDVIQ/3VwWsHrXiTliEkG7TiyT33Yv8dbRwa2
SRLnpnIuDezye1Rhozyg8h1CCb+h5lxIhNfjoJMF8ZsCbdmX1Fn/HXz8VlzX5fHVtyy47eUoTmks
7STpIPnnhf8ukUgNgcyNkDSSjYGv4FA6r/+BALTIe9k/hMZ5PBeMlvFt3rbMH05u6kEmU/T0lDAN
PVtTsiKLSKoCQcTug9cNeS3wlRGf+BlDthTsQgWUQ3M/A07VMdtNjkJ7vd+yNl7gGPM+NDdWqsA5
DrT/wCB02ZjgJbPKC4D75liEbE2kz0FANavIfrWWxHjSyI3JEqi4eT1P7IcmuEcLm+bB3H5FrXti
LISAn9dTKKhtBIKIEj95Vt9SEK+DKK4mhAzVSHPc3AiQPc4Qdn7jEWLj8wtDKUSwSIzPbp39J/cP
AqWszxQgaSkCrXf93wgbYr2j3DU3H2ek4FZ+WMWFo9C2eBEWFTcqosTX95npCTsiDMh9AUAjlpub
tE3kS7NQCd8LyhO45Ii/8bcAYQyuZRXo/s4y3orH5At5uEZMrTITtIKy30g9xi71monXRMQ5NuO3
ZrfA7zHnjnd5OZqbwRdIkEK4SHVBqLC7YKDOtX+6cJdz78nvDWg38xBzu2s1SSMen2HNIW89uNb5
5CgITK5ELah4PLBOvQn+Ogv1ITLeT5aMmYR8wmHN9pLTeaLXkm57NTN3kd39XAba9RHb4PbO0VN+
rVCNKxLHmZSITE7pQxt+pX7gLBEajfaV5il9KK2+aX5xOd/PE9A1495w+HkPk0ZOy5Sv7GLyZvDi
zj2hf6uWhndTg4i597bvxgbUC87EYtmYRR9C4yVCTi6x8sFIm5gps3h/FXjtTo1P+WBxTkdDV7a/
PzjTzJ7ObpkliSSHEURJGGesKD6yajDUBU/iVWM2EG4hiuei8lYmwUHw2IZKXpKvhNwJBBId5yAj
T25MFO0eecmvVGXJkOdkBjIBLNCkN6KHoq1jSswuipN9v3j5iS8iRwiayn4J/LO5exQgkHRqldAR
/oad4ViRRWMAXnM5es71vrx/bftdY3VX16imcQqR166i1w6/NYifzwP2mkQ1YU2Om5tUoUOdJwCS
YtnHFFszPAuLXJRCLDQTHuKczDY0gwNOJKMS7yNi5LI3c4h23PRux5L2Uw3Gx7UXU2OjIrWjiXbz
NNxQ3JTxMx+1HSYdp/yay0L599sxM2MI/43HRsWWb109J9qCquLJZiCxsDVBvY4drnT5lFlN7Waf
Z745F01ghkXTbclIYNVIW3SoauGHWr1PUaWs+ipraWTJ5hd8irXzmJLEsdZEgytL3ATyxyVIopGs
Wn0+p/pr1AH4nhBk5meLs0og/GNnObiOjh3SeXCavSBxv5j5MCYpUgNsnYIoe3JpVRlMawRczygR
d1dKPXK9B1SnIgQ1w7iSPGY2FRw7K1TB7UR7xwyLVLrMMGrmY3dVKc3dn2U4GHbQhaN7Tz7FMcHY
w8MpaNKOrsp3YOACvm5MpnLeE14Kugenaw4iQFO4E5bhrx2VU4rjGSs5hPJUU3ylJqxP0z0G09QD
BaUh1TQM0i/g7sudqlsiBjTLoWvgF2puv+XEWOkBUEJbt1spkS9SpaZTyQjNIhy53RSrx4qsD1Dz
wN7U8pd1rmKPvR0l0yyh0RqpaWvesyiSznlSYxtWC27UXKD3c7VBRBOiYHodKNSNfkiJ4qwMXu8w
A78yimh28rSGJ28JomjxrgABVRJBejINZrqaAp1gyflMhCW0cZt1O+0YLdZ0f/FmopuUrSeBjCtt
UCXgSbx66Ypbi/vbaQUCXQCLSEybSMqhNEO0AmWLx+wzjV6SHcE5n/iJSdxggA+SdB4rIqtFkgfr
Rz9m6hSJDHr6wzMXzQcNEjybTppPMDvAZ3UUHAGLA+pzy1szJ1skyGiZl4QhYCbbvzjbir/PKGfu
wUuaO2m/LC/9yL3io6UJ2YzdpihUV0V7NxqKw04tSskow2c3CaaNNZo8aNOIzWNwnOlDSooX34wz
aLWxgHjzY8bsy1DZVKetbD+Y/KXrLUM9g+eyk3ox0oG/UAThdGsN7gUFML91PdOwqNQ4AO9J3JSB
tpsuVak+a/XEaPxxEsDlcFRnNymmKMIw2YqdQ9R2nrc+wMx0sOW5E1kZ9wJuqhDE/S54A0WrY51c
1f79KAc6AelkeC7jf80U07cuMPGaiH5z7b0cBklGi64XvDbX1uzTMyUq1dlptdxD4qc2Jokps4wD
klG7GrBovEn919FFGX22PT7/Lfiah0HV47AA+G/eQO2oickMceClhU6lSyHGkA0YWbOzFeDdqE/N
YbItiFgfbk9UB1e2J4DeNPJFYRKlsdjhgceiK8v0QRfQUK2uHhdCsl96zV/9PFnBPxXslzy/VbxB
oh1DLY7JYnbMUZICOUKMerLo+BgvHs7EjwfbubUnJcMzmw3q9m+co2t/YJj3pm7djdEBb8hg3+d+
yPWx7NR+BtQsQxfSJMFbZ5G0MaWyyM2gfHwJKry+kP0SnFBw3OTjpZH8EW/dsFZ/JN+6gNY+/Wt2
+w4/W8zSltxw1Lqgw7Ye7+3svHcovzUlaOeWXBMgz4TuY8Y6BHZxExDLFe2+pj24O5PefmPMatk5
3SCIa0XCv0CwXQnyFWlt8nQjGicqLQnznyy6DJX6NLhn3aJuirndJ/NEpX8w6R/knkxiVZhlMg4B
3NYT+LkOFbX5L1dvrTKEQkWGyc4faWfDuPdzvz4tX7JuZHhJjbAnt2Vg0f0V35OAtaD+WDCv2USu
ZYMWUztlBhcikun/JKXUqchVzZnubclQiK3r12jkGdxHmLMy/f6mcXj6Ep+5HCeO5G1risIMM4TD
QuhFh+GTClvnQ7+67suk6FkgSgLzJU45L9+mTF5kdXeYzbdoDx3R4yViOYe5nQ/r/IHxQ658xrDk
+BpgXcRo3UhPaj6l+fdaSMiEJIwAcROKB3HGWxR1GCkPfM0RCaz2OAJ6puGOwdRg/KUT8PVTZZNd
c0ohO7dvclds3+OBwlgz9GVYo1CDeF5hSZL9otvGI5AtFWuN23oJOFkbK8flgjPkV/ashaqZj74h
sKAJUHgdADTlmhpJhLFs4MmFn1MtOcA73kGayqRYjpYV0XwMAdjZbKwah/LidF0VURtCSbsn8VrV
Vcjj3Dw9fIVj6bqzofvcbCTodp/7GOIWlWD1DlMnfg40RD4zz0jndy29yb341zrDrvgpdN73gGU0
FUfkjsL4gh44nxsA3YqL7pQLd7tLX6L3xpsbs4Iakhh91ZdmQtlzM+KsCldKood9FOOzjDY2UgRF
6suVIakFEVbhDfn0BOcEejAyIYAT5+qe/Ols04bEl7VWyWlL6fwuLg24qmq9NCdPDQu8CFk9bO03
611sQcmsV9/47oEbEMjLoP61pPuJNodlILcRhGUW9eOy5OVoZh5iNdS8KWGxpa9KOLbPQ+I0+3+W
kBktiv4RUTEmxL6gbtgETKT29A5zFyqk4/lB6uGWCZKHdrTev9QAjII937CtG0pG6ozA2aM6Sv2R
8MWfUTbSni8/sTBewwXhh/xPdNC6oKJKN8Q0WxUip5frCaV59VPFmG5RBnL/n7U01VAXTHBrjwai
+krzXoNtbzSUaeX0lA1vvaQ17dCvOcGB0VPakrU+BOJtzI99yq2LdPxzPEZsKL+mhZ2KeHCvfRwu
/RpafTqabRiYcSqxo9XFvtIaLtdtoEGdCF2R+czMiJeV1IsSghrTLRgtMMWGkeoy+qr4iW9hkf5B
bl84Ee22KW1qdXCGomcHkRztvwkPTYwJeBQx6K/8sjwhwtjjKsVDFK2E4ZMtQiP5DTeScf0tCF/t
wRfiUf/HyVB+lkznG9jCsxwmSygGf+1h4hMl02/QJAOZvU33ZNLrKpFdhllB0S39nRoejQN612Tf
/lDSRFkmcDLVVzwYIIQqanz7DB2xY9zkPiCeV9lrLSUTek1h+gySw9UBtX57/O/hFpTsS2j157F3
gGGc26q1ILIMjQHwk8B8Y+gc4YXdl2nvUzUuaYbwaTPCXQsBvJTUv2+MJFGaTgrBBUqonkZ0fJSX
XiPJQdYXjrFz9SRKGtL8MSHsJ4aZnxU32xJH5VKdW0mROxEultjWzGsguCY0o/9LkEL/MYG+c9js
PLQuH3koUCJ9jqItTK+ejqPTDA9VDSXdYyKCQoAd8cCmttiaem5/J39RLoRN4vvZziLoRBIx4Ksu
lnHw6ig7sjFksx795MCUhOru/je2MpmJCPOiaIH1UriDH7+7TtTHLBe8WKxaEAyU1IlDKpNMmXHD
tOtzycAZfDlSYlC3wAL2SWlBG9cbSqgBPoxyChr5q53hwBBf3v5cIgEQPOkaArU0uKtGFWBvL3cI
d/YYCT2oXS2EvFN3D8SoHfPkzNxnbFkY0n6xr1Ic1p1OxbjJ+W7y8ciJeobVaGWOOpspoQJQNavz
O19bjtiq/MDFYYrkkD2tQJKeHEpHoLVy69VzyewSw+KszoB1A0hkrrmKXCOb1BqCiIHvb1wkV8Yt
O45tJt9KzbBCbNXpTqG5rIkcHoxZe4y5LgOpoo/HJCzW3e9yBc9lMjAWINRG8LMahLBU3JYXhMBY
N4sLTK1Yy/vT4gCotwlqnjALr+Dt5S/6/B5XUYGuKF9Q2f2mEdwZFup3xaHEkPYux2RajjXY/BPG
3jdBOVA1OMMqx1igx14LViAV+wVhkKAJQckMpxD06sNLPbTOIOy6kCDRdp6tvGwyWTr8jBtPSvM4
So51z4W4qBVGkTNjIDV3n3yZ3LqkzxDuT6BXXyotZxkRvNmfUuaPSdTbSeRLiVmiT4S4LH3Smkg6
u0uJkI96+hoA9B+p1nTrsCOeCJwLDozZcYIAUlVXddHEobGgUH5o1VXB8+9+nJfwHJ56bvTlPJGc
rksyNe7phhWiGnX0z55OaMvkaoFxGTdrrQW/23lRFNrxn/b7aO6k8cfwGllN4GJIfBXhXr+IKb4o
9LOlJuaZV5BoB1LvNs9e53p2hpeZ3tUOOVGhuW274cni5dUmzG4pu6zkPaZ1OccdUQ0FmiL6fvh6
2WOkOtw6DVazDZsf62Ev8lOK7gs2RZz1acO2ckjbkZCJBOTppt16X9qSJe2gMUQIlbp+1tB73TvV
vuxYpA6pQeKBkLAIkqQILr/7QF051U6Qx3syQK4bchyc+XYYIPdQApxp0YmvI76dYMS+Z9pAvQW2
U2I1fhJ+vrjPwuN2ZbDBQTA5lSUjfIgY8Q21k+T9+IiIVNgf4smGqk8ooORd+XRlfb6kwL26kZRr
QZYQXRPbTVJoTIV93wldFbCYzMWot+1Sv4EYGtenbLH7EjmAeCf/d5BDO+n+umG/4+22ghjF39jb
BBE5CcXEvq8Tc8Qtb2L4jx0nn+zSkfjE55K8sxLzIcLRqy+//bqdCi7qaXibH2r5P/9hRYSSCt+b
LGZpi4Xk6vUnXrYhU3EYuZhzJ3MWYtr8KLdDR6qGsEV+ANTrdrjt6wJdnQkT1oeJ1UfxMKQwz8pv
797QkV86U9CuH9YLFLwgSvvQf+T24DRlVilnraY7KpGCAp6MtGTxjYfDlL3noF9LVxPb36pOwrxZ
4dltRmJLJqsW2Na30nAqVs/3k91Nx2CQV/uHmK59J+S9X+zrguKPF/YkN7RqLnnitaJCLvdKsA5+
MDZ8p3Ctc61hjIqzE5bFYqBfN8it8Px+AaFtM0d/w8iOgETbAV2+tLYem50e9lndSoTKX6z/g9pE
r/a14asgXLU7uWjB+9aBe0Wfu2XTht+EiHOGFWeEkPCg0RUIZsGqVF8OCROydhGuLoryRDa4Zo+J
XN4hklNxqdCwaidhaAYyKHb6N7nfDmrCfWGQDDn/zeHfOKxrwdow+9nyl5JM4lX6Phdm1JWQIoNe
LEtEnpUAD0RfYsaCvI6UNkpDE6OZ3mczXhLwjni2ZH7KZW2p7+UheqcVnwRmgLPQqP13tpgMmeJq
OYPqDce+e6DYcNM8J5ClJ0WGBTOiw6bPw8cv7cEXCYzgpNiQfMIE7ySDEP2XzjQ+SPyREY3xjaOC
U0OIe0UE8GVoBJhztHfuuUOtwKEaRuSaGEX+DQOMJcqTG0Jqb3duY8L6IXoGCgqDpdQx9hqGPrW+
PhuR5Y/8ykbK9pmmbOsX9LUQVDul9h079epVRCmoXd//tc0eTv/WxezVSSO4nF0wwbne38mD3EOV
BEr62R91F5ZvIzphCocczb9DN21C/K5Z0YD8k9GQBYVVIpVqEJ/DCrtFMxlxp+qsR/ncbp0HUAx8
tS9uoNuezkPJI6k2qMgcyB1JYCxeD31y8+B4mmITXtgOqIy2j9Wfek/4psTza08Dur9O41zMoSyz
3B+Em7Q1HkYbc6il2IMqn0IYkOEB9MCM0MTMzdIna4AB8yWUabcEj5dxzlMLSkRkVLITmIrIM5N6
Xle6rhOLCm5zaajKro4Ygx+lOhIsKM7sAiXyINir/NS9bmRPB6PSwo5nUsDuihbCFHxgksyldlS6
/pOKbsNZkvoVH8zNKW283VA4m/smRxqme8Zyf0ZYu32kxsJO7h9EsB+MKSb1++rZGBnrgDk3MnCq
DP/1hUR7oT66AfQkQLZqGpBrDgx7Hq/HT5bSA/7e+HRk44xd+SAfJVpf2a4NdW6wycBJtCS3xw1b
5ivJttatKvMtLNPUJa5Syr6WUStEAmumSGxUFBGdIZcg4FlUpIRIP4qIGzalTJQIYnnbmQ6jRCID
pGuODZ7hs3oij8/lWVnEdkt4E9wYbzGMy1CkiVokazuEWRiW77EoEhiLx4nYYmj/BuRYmeAGNef2
L2NBFyJl8C6d2It40Bk6UL6CuYJNmhGonc0jPcKo5GBtK0ZFpCsMEcon2H2+xlqGnlOoyRXBFOH7
z3pvHUFtuaVoYKDrxOadEfBXghsroP2XnRizUfdI8e7e+Ywh2hXhlh3SNfCVdfw6BiF3G5K5EToG
h1JMj6AJAnlVoSmpTW2gT8hNGYjoTRZ/grj7md4du6V1OE65N92OBFeBtTyCjpdY+GpqAmo5Nqdp
bvndG3gzZURMaL4utJCm9dfnGKFGw8KGwopNRdAIFhFmcOWI+o0MJVeE+gD0SBVl5oRZ+tfT4L75
KIaqIIHiqm/fpnWW9UvIJm7prQFLn+449gCJGelB+UQHrG+Szx2uo7grP4xg1HXFRQZzZQ4FvHHC
dtcAmkQyGpJkWSCVlynWh/1H1yJ4hyXK98FP7dthADS6oLO4zOnGc9XsGgoHXcrZdAzxhHugJ5gy
IbdwGxZXrrEQ7/SBBzS3bFdpMz+zJ97dH7Tpmmh44wJoO3g+KnD9LOvfzo3mj2/ZRGxNL3t/e4Y6
VHeO2aFfF7R0RMzMZRvzmhlMwUYkC16vD24kBM7ROorSAoP9RSqYlGTcDIVcUJxofp3Aibt7WxJv
0E+l1cQxLo4eLyzpPDwg9/qSk6JuKLLAZqWboNJeq/ilYrkK67x8BTqB/1vK6VupHvSDPgv9CKqx
vH2pjZL+ICUhtEJOsq5+7Vho8LuK+afdhHhijKRMOa3mVz3lb/CoYyOcvreyppReriRStku4d+f3
c8AwmBHdAbgYQbOH9U9cYFTJSaGZjQUUR3W5oK3LqFPRHgv0+wcM68bHgkyLiVVzusjtMcOq3MXf
16GjSPc3+esuAprDYG8b1e1YNaSTe9p43ypRw9grLvX25xtzL6pbmX1RUyPeCP3u+hfhTbOnPtGK
WeD1Sco5mRnLZMcmUTu273Kxz6skjjSVxJ3V8theCKvfmwkWhAcifhr91PdM0gnrntFIjuxyS9SW
GgP3SXlBfUNyj6edPHURnBoNd27Zx2BmY+ffE+YqfSqemnZgoDlUkFXSv3soVVL21mt5RxTSIhuP
GBUy9zyno2x0ZKFMW99rn18Ney0dnL9FYAmlSokHP8b3diK4q36AVYQGaDroLN2jiOCKu3qvNMIV
iyCs1uS3V6ZEFaYC4d1xsFEnxJRofC1xnRI2LXLKxLSA4nH8IDQIAt2Qh5rQl13wKGtsunGqNEen
AzJcfcq8SYwkXcShrcJNiG3nkOaKF3n5RyLbWzGYs0dWUJ9jv9eL8O5fpKa3q8BpRcIgDCUhOdUv
0q/u6IQIG6CE1l6f+P/H9RpAVYCE1YAZiH3YRldsT72YLKgE+noR0ihU9lJDAOHQzte8x44wtFAZ
E+Q7gIE4kpcm7YWVLqUdn1EznXEnxFxa+3I3ToF30yal2Qaj444PJR26E/k8qzx2mUm12tqlpmOx
xgRkVHmOp3mL6smQDq/E4jea6EQdD6/BW7yPalbJh0AnUzD6b6wqMObahnSFlXbCEz6iktQK9cW+
tsPg0WyJefQw2Iyjg76tx3s5mDaVAYyy3pRwn8M9qZtfqrrb7j4kFs3tareJfHSJfmdV9KlTpenF
ui22kS5CE/DQL+NvbfQnQq7IBrYHZDF3lFn8Atn1nKnjXVNv0rKkk5ZtN/J5p6fr/ssjTrchxQyj
hZpiA1d+JJaQvC1L7Dzl+c6amCpvQN1Kj75sj1Ub77hPLGICTag1fTuCmeHo/rw1J516wJKGpcWc
4g6eWNFskb8e0jZ0AL6JIUJjEpbsDQcsbBKgqyZvbG1HNcyhE22t4TgdiW8s/0xXAiTe9Touquqm
0u3okQ2KSfzbc1QmxOa4AYLPE1BNytbKqRH2pyarv4OglQnu6NBiIGbuz0tXGzrb28rJZpG/JIHd
cmLMa31qAPO5N+tSJEhH/oWP/qeuefGXTWjGa0yTt4+eFifbUQwQWVQ5kadqLSkjK3My2SJvzKXQ
awqIu13zJ1yslpIpk8kBm4JSGN9p+S3QX2VS2bZbwA+he9B81IQlLsrDvs59tTXLQUx4wLcvLnot
tlpTiFCyd89L1RTZp3l/nmbbNbfkxLvTwV6+sHNiiClXuL2EKcf9LewOdK8U+eoBd505TQ+aUb0v
bHwUSiuJheXz+e8rvZStA7XtOgWlCcJlgZNdWPntUYiL90INh9+iS8TKxBME7oCBCJ3q26k3yBcA
7851S7NMd0SKUg1sPQqliv4HqRyve1UbHCTRXs4bN27/ciL4Alb64ZoqkFPfGi7xi4Euhkp+/NN+
Us1sXaFSvO60+B81NiFDTxbFKLIXHfskqlqIf19f1MBspvGIfNe4t/afgnnNxkSjzEEVbigMpUSV
WSRYuRaDfHtSyzVVyLiOGS5RRh9ArM7DDPACCeAw+OFgVjPzNkTK8X5rS/R/sNOS6vlBrDi0OnPs
0JqdrKpZ2f7d4BAkvgeVeBy3tqTBIURSIeFMDPwQS+/HwUanVUf58TsqJTmm4Wrnisj3562KBZIk
IndquB0y3C87EykLZeFoUzzjdfF3gnL31LOk3Re9d0+YeXrL5EQWTVicI+RwbAPbb2q126uRVmEq
oHgUqH95bcb2Tlg/PftveiOcMPNnXSsVMaHjQeYL1WNJZGM0EvHeuAkYvh1hbofJk8TTIapsb5wK
pVCqS04+sPcsSzb1pMHkV+o8f4z/cmFrtDuB/91aYb6bJjIZ6Oc09t/9+pbF/z+tRSdfVuRbM0V9
eFTW5BDz9bhVMZnu13wP0UILzFI9G1Xp/SBrtf5uutpPU6qZbbgcLGtidh+CG/En1EWwUe9iclvS
hh8eLJ616p8x/v0PmfUw2xv/HxFZ8ewkmH3m3ycXlI3h83o9WXPDzPhd+p7QGzbav25nR35X8PIW
Vcg+bjHhAC+7bqOJ9vu1tuP97cw4Bo8s+krxq/Z2bC1kq/43YJ4x9QtnfzZua2ZnULxDqfCvBVCU
rlzvN9qVAqr+4mEkX/Ax/SuHou9rIx92umGVLiU4BTyHJtdPo7aw/NrjotPxc9sBewmdaxJ40epi
y5YXYtQG60AJLy682PlIaRdOsdz1xqN2BmLymYYTjE4xx0fruIZyWubI7sF6+yb4NIL+uBYu7SwM
TTih5mpLOBSxcHhD2rNBEy8cezR3L6Kh1lVE1WeByIvPFAtSP0yqVDkMBKY0zECK6AztyXLIcqwp
MZTa8p9TaTLRC3A2j9x+LqbgvGyRq756VfZe2EMc2RrFuNqvh4VmQTxxYxHmZ6ToQtrIUxNRIvJ9
+W89c8Jezku0A2cfEn3bPJDHXObK/Ili779oRQjTp8jhaUz6NyGFUUbtbQ9SsMzqcIU2HflAKSNi
do0c0aQqn2Suk1ivyBX5X9BotTPy5pwgEidwbprWZl/kWzaBCNZK8MB+ucEf1q7+l0MroaoKRHZg
Rd5yHkfiNg6aWRrEsD2t54FuyN2ekKPu6yMR7XQsaAZYcQXphIxltc1ORYyGiivRQANGQYWZDIMD
TzT02j/TOXUn7LeiqkZdIHZZ83Y82cDOf0gcL1CtPVKvlbmzdEBNBP2gCJlnPyutH+h+XP/KW936
z0gE1ol9RlXcRdVLgERlO/gZW1O8lKwJIvUVmoWbeQk/7c1vuJ68n8fL8LMpqSuEMUZHoXepDh18
oPj3Q81wRE6CbBTZvCeSLUUqMxO/kYzDohBB5E+566/nwn46o+92tf+kjIGoJQDNBSLxhrdNj6Pi
gAKjiwpKthjfGYHwHEJueqx6s8d32fp8tV6S/WqilxEFl24DXAKaosrRSUf/Medp5MNAH1A9uBpy
9TG9Yjs2/SpvXGPKZjAN64rKMlOC7wG9ddT2xaIokvoo2s8O4Bp3II+/8FUhTNn23UrGWphfymmy
1Oh0ytAoMqHdz4lfq3RBllyseAJshKIUI77e9igjd4hclebt9t/bg05RfvpPeDqDjoPgU/QDMeeb
3IACyGxjGQ7YNIo/I7zIEWusIq0J1A4MWrCLN71rQR2Uiri+WP89CZxLF2EEjH3NdGzT2xLnmgAL
gaJPCoXmnt7RIONsTsLwxvCrNhZ81ISd/OcyDY5jkwpeuUzz7xuxCcCYRq7Rz3TapHS4ITMGeD/Q
ExlBIEdv8in9356Py+I+XGtWjwnTlff0U6Qy6pyjefbX5/fOCMh5eMPUSULD7oKIN8/EPfEbTGEr
UMT4HjNFSqS+vIOYzLP9lxzwm+7Mc/tduENPLH41vG99jxuDdQHA9rfV+fKSBnJYbAQ5SHqHFIZ9
ZSJNAtPVHtHmuAnwWJULgc0mVrKVJ/mdTh+PLwIz0+0ZkxX//rBKm3k9BHDWvgZq1G0tVUH0fIsJ
emM7LaENlRDoLQihU72W70DghKXzMO4MMS7h+u0pp93CT3rtpMjpQ8wBDVIIOE7gr6zX+Fmiya8F
tJE9Gs7uXfAcMf8iR+qFLaPpvI5y73Zl/fRwD8U+s5YeqwYUjM8nzU1O+YLkGKoX1lFQDrBqbOuO
gK1AuqkXXEbu1lKK87MHcfBBv3m7IFKNwt7K8jAF9C1M0b/QnEJKzrm+Zzg3CfDfj23q2PSo/hiW
21qouAYv3uMxTbowAy7yllxGCmgZbbUMbhCcYbDiNOhLMoCujSiFq+87kN4veK1By1VxsOaKcdoI
9KbdfwR30zKSfYGPeEAqOiWdmRZSM4rVPKmv/o1QP8g2Fem2WDF1viLri/QhwaylD5DphYdiiHCw
vsnZEyUtk1d5nYrDfYfFpnEXqRHbdfLlVH0qUg6Chd4aytcdV62VS+oV7B2JIBQaCS8YwZXPtqqM
1dhBL52tDYs+okwgp3fObaFD0CAcLrNjvn/5qKdc5CKjRaRRp2+mjC3wg4VFQUoe0TbzviTsT8qM
ccpA/sLAX+1AVCqqfK0nUF5ZlZWEvV7T3AKJ7tlbnh7o2nynruRf2SNcbRxD46LY+qFf4W3IkWKO
7jJ6iSVTDpvxysdGhISd9EagWVtUTzZHti1oU0DhuLJqzWpyqN1t85ugBahFDvzK3oVYj7TF6jER
D5Lc+56E18E7yr+3mjOboZInMUgYjecwGFZTiZilnHJDT+BHav0Xx6r+0m2xJG+6N7NmyAy/6BL7
JTFd3ygMgmlCltnZtgMPhJxXxSuaelJH4KvfNI6T+Kn+voaG4VuCdsfjkhEv1g13Ur8yYds2jLtT
xk31BDHBlzWyb4un4rsdNjlEYhGlBng9coDE2IuVjjP51I05zWKxD410nYkeFw31SVPZNLt3Mlkf
SwI+Rwwnx8NfosHs4MdmnWl7nbfm1TMc+25FJ11xcxAexCRzYIVcxxOs7oZ0iYv5RHN4pobSMzZU
zFIWe4mhDIlW/UXaAVvEw6LZh3ylcRP1/z7uSf9pAi6DoNRq2FJjB1hV3H8xz+6qKRaLqUQ3Ah7S
C1nKpLcbzI0DR4ZPHJOfngjPH7Zra8QjOI+s9sBgakqL4W/wty+rcsGcuerdrzUsVK9a3Kvde/iv
sUs4+cQO1aF46SPpK77LR1vtO4OTClOL3y0HAdN5iqbHxoni3W+G9cpkSYLbtt4rSSX22ZmxzTbW
y/5qpf2HEPbkvqD0V2QQgzjOGkMaZTZ2v52Hpmw5YVFW/hKEfY1RiU/s9w/pTMuSHzACaJeFeQoH
AxEIQZZZwNdY7LfkSEg7vTomplFvxzQoBb7pg1IeVxsY71qcf9LCwd7zIy57FIX38pt58i1rW1i4
JrgouWf8CmB5Z9oF8iTbiLN/qwIvc9jDahd482eGWbZT0rjdPHeNYgKAIi/5Ac0mqY/sdrFOTpBb
iuLg2wt2svwKePEGGFIDVQj9vrKuFRNAYczZWIh0J3Az4is2eoQRb3az4Rk85b9vB4BleW105u2M
bsMPzyzxWMug08gMJpD2S52z+vO0zMYfs3LJIMQBOMuc10P9fo26CLw9/x/BroBhAPaAxsgJZv/8
dXv2Mi+tUaxRX14Mm9MIZA4AIRJHpadf+Io0UB888AhAFwlsjZ0Arqvpdiveomvz9QhjeGSUjWzQ
5FD7LISXE019LEm6S4391ljq52dggwtXIzFzXlNeIaX0fafphY45SAkR95qdvmp0cHoRFXCnv7Of
SuKYSzyqhOr8XnHjF4CWDVP8Cm/NJCfTLNRQIxH0YiTfqTOyCxJhgwBfTuK+UQ4Kyiz0Nf6giYe5
iIEHlbKB1QYv+HdpLP0Ry0gtK4NoasqU4/1nmHcJjNIyeA8KHBOU1IUjjbV/orj36uieQg27v1Hb
WKEfMhvZP2xNmGpnjNrkN2USyBoCEMb03Esl2rzwgq7ONVfXKyVmSaG7VocVYJhrzs6F9ouTflYA
HkXhNHBFQY8ZkM3ejGWM65f+TMkZkVgpAx5PzXAel34weH39ZsWsETucV/FapBGLqK2+KjKEfutG
aPgj0OkGh/2T+7j4mOBL9Rlmg/5IX7sfU9kMY7dnDhuR7uU9aqo2WZfGKUO5yzGpUM1AncNTn+A5
mlEPtVfUTFov2piFbdX9tjAROPmg4me3uJBVlFAKJEHDpqi91UHfGkYXa501S1chPSv+xK2lSy7F
37MPYQekV2x8ylI6aX2+bF32EG3G17I72TwrN4ZwTD8qF1Pm14Mu4MZ6GbkGKWbuCMRDgygpC3Ap
NDvYKasQdutmrqpJ5VCRjHdkjb8t3Ar1QBItYgligMrBdHEXNEUQWZ5pImJhXmza1o6G4Aq06JAJ
zahFkJSQ+1H9jJHdadst1CQ6OAwCYhoTocLaiNRVUCepHsOPDEI4yHsX2UnrZdRWVQgM60ZVDU7v
cOIOSONQgRVZexrDgM4o9NpxQ2AlQ8z7WDcHtRJJyZo8QnQjK119fpLV8ipVJ1VpwPz0+pLBEdUp
03oSZW1HoFkDBLPu+od1v/8DIS/+J6+L/KXNRBWseMwK4motQvobYE+7tdKs/kON6ZWn+2AI72Aq
xaieQWF4Z2tiPDDqVSJTABy9hgXsT/w6SNFyj9Yrpy47ISu2hF59ChfJkAkgoWNuojf8MTzhOV5H
XcVqUHSRcFnvExAXftOE+SXuhvCKWLfUEBh5agxA9d/5zf4/XsGAdvS5K5EL2cA3u2RjuuchZ8D5
XIPbyRtH/mVskrMjKd0CCCGXSGTWZvC90Pu+QbhH61Iow4n3AJDrr2NaJ3ix2AQFYDas/If3b00p
4uHuIy16u9O2iWRRV+JKD07FiM7f0/h/7HxDgnCHVYtAdYR5NRVybreD6VlC9QrzgY1DKPNh2wvt
fA7imQ5Od0OXtRAwxVw2nronUuoyK3rtH73yzqtHK3Fnb9qTnKlSnXk0OO5Siy3ubYBawExxJNic
JTtEgZ+lyrIBPsANAkhLhTOmMwJJKIMgVsz4bh3uOqegtG+nmel+FunjL4RjycmGPMBb0dsjAj9b
2CXZ3hOQHDLNPNbCfFT8lLglcbktXXP5tDl4XydznW5d25FiyYvt2+aFhVp/whKvjYbZIk05alAg
2oMomwhsnUJ26joVzzVT95Khx+rSKsw3n2T5XnpuUKRpJgYHVYaQSvY5cCVv1pId3aqbEOAtzv0U
hM/4cFQRnrJr7dmWcJiiyJkwEqdq0UIpTOJbR0pdE0xj1yYGIkix18ZX7+2JlJReufYOKR2+4AQB
ZoatSfWFq1gmtE2Brm0+Lrn2HPFXCOAsykMEKuaRT4x7eqGzSIkspcWGW4BphkZCfppxIjPPYlXq
HXwtuatUfBQUdTeqNxGb5z0ZYuKyzIlLNOkEwOfTo0z/PAqIe2vGcYMrWK5mY57kU9EnusdBngjc
EtJM1bPw5y4iHEfVcPfZT8c9cKMJ3xUo8MSYpbFaKziTMwYTasChnsX8kEa2gt42pcLPkOJLp2aJ
pJYCp58zhGqmVW4XXYzdjMjwha7/JRzazni+/rlx9rgtJXpp90dw4vmgLahWd0Jvcuak5197/eiJ
eKg1IV2yucFK51AAed/A135CQ2C9FqIPTNml8FBqO9miJzYeIPc1bW95Njb837lvOaPtxdGkdF53
/Fpqow8qeZWAHRk3A9vkM/fQ4SQiIHinYaidK03Y4sBsVrNXwSdmaYDhF1wYcnmGvK1Du9/f9E4f
m6Ubf5bT8JKNADGV353RybjquR/pgwzmqcvbCmASlBKgLe5VpUN5guW9od8q16/aRhLIPpL27qON
Py/sEEjh1jgOJ17diPbGBbZsRH/rTssplkmg5qJLfJ9JwuRQNIfCSc+G1TabOd6XRgmvJjn0Tyxj
n2RLvd3GjFb3kx1Qz9Z7uimJ/2OWIi+C+XXMb0neow3SRJKvQcck7Br4RaH+29faTr+fPqEIlz4Q
hTvsjWDpSHo8KjPAdfioTpou9vE7YmxBcGI2Gmq33o1jSx1qrcfGdykslnS0PSQUxOGThoYBlw6k
vwrkCp9b/OoKn8e6Jsox/w2eJq7MzHr8GrxvM2iyk1gQ3n35wh3kDcV9Cip97cX1BV9ZVLnKnyBS
t7Wu4jRESmoffDzaqtLo7t9zSYvLKUL0RZPv8wKU6IjSUW4jPzYettyTZqcon+N1ykPSJIrAJzkr
8p+MeeuBLBd44B8cUNLOC0qxvE07Qdnwa+jE7z6mHbnSnnZaTkMHcsE6ZIogHODQHfXZDgfud+zp
1Y7V7/xXJr3dE/l0aynwo4gGRfxzMp3JxOqciri/DXs4zUyndZfj1p5+NL5UUjDFV+UTxdnftldp
X23j0CJmTNdubK9T79B23X+q+toXrDtPI+S+OPzgDfM8Pw+zs2PogIU+DvEY/BHYxqMfttGalykS
fk1S4GCvGYsJb6G44Piy4EbVIs9+/LZ2E1MzXkEpLeCszZ0Z5Lwqi/EQddLjdoxekwXZo/zUHe1Z
xMCl6lDmTlWYvqgfLGKWlyIySp81Vq9XqYirSYyz6fGCqo+XE9EQKxke4rA7hRy/0a0q+wOZeFko
1s20xgS3VB5L6ZbkpxzBzutI6l5E87OcY2tELW9dGZPPyt0A29u1X55FjCzIx8IyToKCnAbQeQAq
TSGNT9GTcq/LOD0+2aQG+VIWnhwaD/Gh68zOScmjsHqhD7eqHlPuVRAZSVagiFaxO/YWY5XeJJpW
M+R0QCDM7Y/sl6zbx/SyLrK/Ke3Bi1emrcseKrbOvF2vaw56UKNrDc15e+G3zN34vJbuHdctiybB
Rj1qeWGCzdW//sPvCu7iWxAkzWADePuDQPFYDkDMaQgOBofcFA6ghJbYoOO1P5hzvDg7xDNZf/gl
ud8y2wzW6eFTURldTwa22u4zHphVuymbDHlnxy72UiBmWtm8aW6YH4eQlVAtg1aXgHxvdpYeUxhp
G3rtuuiVN5aHu2M9aq9iP3Lk20AOWj7qXvY/P77CKkRT/TIL7L2dPLvP++mr4uJXrc9uFf8IF3At
MNFhGCKiNtxaDYMb3OBsBSYRBHffo4jXYP4uze7UHV3i9NODIkWeU3tr+nBcqlKO3b8e2/CRq10o
iCMAZ5Hh5umTWOdRKQT/koB890NmRJPr5MCaP+7kYXxwq9fG1YJc2260T46/rVL4a5veaAVHrTRV
pxWHrOaVlYXozCvdowBFakvrWbVW0PXqLmOPT79Q5XVPaVzWd0yfKoU30gam6egOOO4+tNjI/8Ho
0NCMH5ybJHDfKZQR9bFeP++rerc7WqblS+v7kIwkoG5IrAT9iInHValYmR+LrEgz39Aj8OuSz1H4
23v47S93rLd5Im1Vr0EAPnMV8uqwmys/Ft6C5JZyRCnD8GP64JbK66SwUm/IqYbukXxovzifgghv
Ispard7T5M/tvjSAaVLf5rpthVXfiAszqpiHz9LEMGx8h0uU1CE5fwf/qPxwY7XwTEjyrbNZk2w6
jjMUPAEzt+xJ0M2Lk6jROoAkFFdrqhTiBZ6kpKlwy16+4+JB15YlJgrkycOf7HawE6Pi91aoxaCj
4xAuiGpTISlcLLKNCTqG7FUlddxn2cVSaa0xaYDuMDGggGHEo8mJBgO2k56y0t1Po3lDBPMO7XvN
/zVUj/sxM2r1P+plMlLUyYGKncvSkIZiAT3QVL1UenTscDazJOlWcye49JjlsAKbEnKIU7Ne685f
xu+OPi6Sn3qWVan6nSaaJmhmjJlG7TORELK2cuTG0DFMTY60rC5kKnTYqXt0+bjf3PecNEpXFDpC
4EvIwuc3YfiNgvF0de7UB32/zpXq8pO3Yc3estiSx7xhdv6WkfMJ+sacXvkB5/Kvj2MQ0g9oaFIs
lG9EVWGBTnUi0ofquVusNzyMKTscrCn1s6v2VRKklsLosW4OeO8+IKSd3XJD2tjcau078YpGyMK3
ybiewPyciUGCYqI5uLkPv6Nk8UWjoEqrE3GxRyA8CgXYhuiNnzVY5u/l4YsGpo3EFt7JORwSoVNG
tiw5AMONWPPPqWnpHX2NpVYEiI2/L+rohK1uOr9+Rt9IN/0qWXQbil8q7eDa8SKS9/cZllMruMu0
gH+XSA55JmFFSUBt5BzksT02HfSZn4SM04Q2MVBXBmGoMdvtHo/nD+/myqB/Oc4qVmsQ+F+iIZlI
yG8dKzpg3xcuki3/wEwzeQVWJ8wIuDIaa+76Lc7EaMYisu1vqNc6OZcQXwcEIjRqSMv9BcRSQkFE
OMf8McQ35BlkNHXpDNWhgwarNxiwx+fgpInHeUwzCeUO4upZXg7wsMvtkip/+lQ/v9J0xy6coWPi
k6Vd/jSFdlUbjAf6ScM7bKfK3T8MJ6HzckEGiaFkWn6sJA57jFw15lglb9CKz3IqhHydXOrrz9kb
fil4eX8p9fr8CNwtj3381ioIGfwbsEDSVVKOxNQNMXXaKqnm5zwopUJAld3tawQ/UXTPNyWqN4uX
PoMkdZ50rgzottscTnpQJzZ16803k5r4K6wGRDfQSKucqE+tx8XUj2X/0yAFiQdOwyPpkS5USOx5
EAyj544xCj1LKCfkSA741dHa0d1m9S64qcf6ZOoyjFcjfQ9zU2CYxm8iZ3GjAf/ShJlVIbCXddIZ
wNV8PskGdP25K0aCjZ8tZ629yM7PmQ3Cxnx5y8Iylpj5YxE0ipLLYPvYQEk4gVrRtTsOZLgp2MOW
qHk1IHeOLiQPgUl7R4lZrohljlSyhcbj9vFTn0YpWknLQ9GOQIFisibIA4cgNUOONJdpkwMnawlM
1lwDcAcuKDkZLr8rTTmUq89thWUZ0Nb2Wks9LhgmfYPaetK9Kyg0w+grIWqM37c5P5xuoUMHt+b+
NcmxAHkyx0dwgZi+dHiEG1uVKGyxHBOfGFJsJ0EfBiA1ztyl821U1HIe6r3HNEDo2Zk6k+TnFyNn
NZ5U0lyYEcMB/lFC9Xoup/8F9AG9QDk0I0Sq35xu8uWXnzZwbWz3Pmpw5+4VTCj/uY+WPWErxRKb
O3VXVUysKcUHY0+YCD6RICgLYr24pajJ3DF8Vxb/byPfNV4tsz90jYEIYmWsri8ut8kJPQ4IScT0
J8WWy3a4b6/mBDrgKd4fj1zJD4vh4sEqUcp//o1n+9WCBmlggH+3MG8z/iNyA1JDq38hKPhjt0TC
p/asvYhkUF5b/+vZ6cvruwyvQz1ynZmHx63GFAyHpUIFF2W6TMGssWS5CjkHSMj8hf1L3/Zs2zYh
Gf/rOKjb7KuZVBMWQw4fD1+QMQQrPbWca76jrMbl0+xog6eyaftoMC3mEpIzQErS+RBaeN29oWhk
ogJuxm2iuD5n9DZu+USEGVfx0mG0YxiEF/MqRg1fs+eeAj4Hatxl1frcxhqdMZHkGDjXXr1cunAB
Plm0wK3l9bwXQpEXVmaQzd6fF7dLpM0UprNWEJr+bF9u7CSVni1ZZAFc5IeH2tBzxTMRKdNqljcw
PqnaPmWOJ1Ol4x7FexCVwuELLZp8H+uZhjc0WdjZddwwXkJ5/ZHjGVtWA49Kn6enlj3+j6ubl3wH
WMxLltmlDmeC7mmWjY2i1Up9MBSXqF25VTfdUf4jtDUHYEq6J82Geo+DH12AT/KZPuXZfSUbmlCh
z4wPwEdzXScVWLWLsd6a4TVh4V1ZT3dlCW/fblskrnm7gWfn+shI2TiG2LVH7H2ovvfQrARYVVIS
1XxI4VK+i2E9tX/nW0yPJV5xJKCW+uFKHd/DObA2wrC4tnxD+xCIzYoFMLymIy8b9d4AJ+z7jApz
qUkPPhsc4tuHPvxtxNRa3Ia7vb0OrEPrVPHQ4fIm+/7F5DfUeNosiZ8DWWyGOJ0+utHYk5KjsDXk
CN9zrmGyebTQDdOpZIU72kySwVZSdULC58+BZz5EUn3OhI2DNsoNAGP1f+LYTGQFiamvTCZN9xp7
UnuSIEAypniZBwrnBhQ9trgVtQMaJCen0Df48TuFAzQ+NtKjpg1L5VewZqM3DfXsNPrJDw46kgx2
rR2p7bzruzSuzcVKJDC+uCyQ0SHd9b9Wizom3llkdsXEwqV4hJA+lYoh3VNYsGroBIt0LJTP8TYH
YtNsGaWZ6PMoszcnRfwJnTP5pGO08YQE1B5Edz3gpeiwY+B/0Mb9j863eUzTHeqx8lqGsFbLyHEY
XemVOehxs0G0mX3YQqj58JM9N3FXMuTREX9nt2Wr351Qdg2xmjUd5bXyTE4Kc9IcdfEW80+Y69lr
4afBYn9DeIjpA/4O2cfUUEeE7N6qjEkkpoYTz5RccF1UmyHAbaS6QHhBBzyOH91+bq7pVyZ3BEPo
fpQbawgFPw5pwl4l/r9OV8OxZWXPB3Y2BrWFOedmZYe/KkWJqm/lFrp5y2KCczHZWk/HiFaK1yPp
37GR1WPE16KXddoi3qAaxWyfPZPErVspLMLkj2DCCUreZolOkZRWKkv8uLDrx2S5XoouFNtarcHo
04eyCMBt8sYqbuFbAEtzTXklx4riPeysobfNTklUvFwNlD4gA178VnVUL6MMzxxu5jzs+I/Kc1Ja
qcg+pRQ8N10Fzh3aKKQUbZYXGgpDK9HVfLDvP9ujW902LOE99Bvy8D9ChBIC5bPIr9uXZjsHnBg8
wnaPvJgDpX5+D5q3b+/TMZBOKeK+drZYiAIyxwovdYeLKE7ol8W0a7rJ1DehfQUF++hB3Syk1QNk
dcgKJkzHS8ErAxeKe90+cmeTBs0Xupv42Nzb6PCgAG+ez2+CDEWXudmsMB9iNTNqj/2l9weE5FXo
vSj9J/Cw7VljTn7Tts3i+/5VZlXekedshtMEKxdoVVrR+Rrw8iszWH4SF/neeVz++9CbKK4Scpol
fhocCuiggGprWBkOSll20HKORkWzucvHPQTkMibv8rA67Q2LYybhWXJ5JCNz0PQu1Ulsxuetauld
GXpBzM+zZYh19yHLWo7CBn5V48PZ18bzW7sW2uGs+HWO/5daLPS4phmnkgnL8IdAtl3N51MNDeig
PqzitpRZoD7Cg80I9R6fBxrt+LR+yrJEwpIn6JSEhv1GW3+yJMaXHnPdnw4eKwwN7x5XK+6W/Alz
Hrs9c+jUfUysIRnf4vLkRViFditraYOIMQlAIm+94wwC7+VOEz/baUEk3kWqxD/0i9Ryen+fzAB8
pJr6CCcJqLshehZMNqkP/hEZ1vvKUVL6M+DLnZQuTV2+jgmGjjg5Y+xgESKxEbkqz21qUDH9NkLZ
LkIHLj6r9Hmr0xVb14smqsdAe27aAOHrNtpl4zOE8gKm0Y19ZRMdfq8AENNWHxN1/Y4liWPo7EJt
UVvXMs4mIJvLJz418GERgMbjzbIzG1wfiwaaQ6jXs+Fu7d8nWIaKVqdTlwQkqWQI1xfw/cspVG/y
V0Sm09muNgUs8DK7h2hDotvPbddlsRa3xK3fDlS5MKpvAFgJ9Iiu0Az0EptVRVbEe4KPy5EqVo7U
YfvLkkzKd3q8GPIhoZYV14BK6+8TQBFMXM4LF7fJ/aFgBYV0zUg8cfkAAH15TcYldQFHkQ1jpnnw
8pEbUXmEQV6YiK6XSOHGI02Zp2ewevZ5h7Rhr7xpUEjtSEIiIaUUK6XZ52w2wLwWWDF4Idehom+J
2/oyGrKT6s3cWxihVz+NEJqlBVi7btSgdEYB8zNyNpSwwm3x1MUw0mOKf3l33N5T7oTzigVPPEfo
E9zxoC4QKpMCWC1R0/MI0TeqS82nQASIuqtJi3jx9PQ1WUFeLDcV8yKH4MiJKG8eWUtxRG586Smm
zaGqlTnEFFT2MsDVNROeUIC61/AbkgTxOE9C5gUTCNZse5oTxmpx7yQcWEzOIwaGMDf0xyHig6X6
1Tmq9DZn7vJi7Gc47poROuL0gHiEvtzl3iPeaSyMu6OqWARXZb7WrThuCo1kUf/z3GPcYIhcZQO+
Y7SayOmx5z3xF4WisYbL2MUNvzXMqI7HnlGMVxjK3e5+wrEUCoZwppxspwmm4e9ASZdEvOxr5Mw0
0/cFwXEk0xb71OqIl8fFrRHh5uXRtGxSKKLnMC/Y2rHGDkwh4lodsw82z5k0s8xM6hbPnqkrEbTY
GnXkd76BFL/fYgR9nxFNiVgX+xFi4c+dcYycFGy/XcE8WUj5XuR44qVnNtr17KuhUZ+5BCf8dD7F
Fh9UcguqcStinO9FEcDEpCkL55l7O4IG68GrPqNuTl6EPT4pcKerNL4CHiJ7LpXXpV68IWxxqGpT
5OCiOKeHrLWGNIxwb115dpCEUTP/i4vfBydTZNcX+PjgugFG71VnHuYeetA3pPxnCmf96lIudt8O
h492zP6dY+lMFc+crDwSfC2Qqvgw97XaYlLM8IhKGnFaeBTsGmpVAeshNg6yrwIZJFEZzJVa809k
/Ek756QO0AYUgVwQRy4oWGh2jcG0UVI+AQYN0N711FdstPxdiB7OUlr4IdJYOW1qaTXZtoD88xyU
jbIkFejxSUkezBNLNOKd1mAQposLasl6msqG6QZEeucR75VYvSNjPWJ/AGurfF8mNbaAUM6RdRgH
0XQDLJ54bb0W2e778eyqDPMiGNox3zk7BvnzCN7iaAegzOexuKk1sMBV9rajYgHyinj5rfbiZOmi
dVIUV/KErISAsZcnYmo6vPmxgSGgGJaBopumbW27n386Ohzc3FT0ObnuSeJ4fKWrP3kRzNEgfuaB
FrZJBFVhnK7F1diym3UvPTbNRPXd7oMmta05nkmMl/FJvQWEMh7KkFgjwE7pDf0zH8tS4TmASzkx
tW+eS2j84NtCNQGAJOcix0YjD+NYkpMQ2ij9jH2KqUV3g66eu3Kgo+bwF0zIaMBniZo1/QMSJNuL
cc9L/ejQMoFCpsJp3pIQH7xAl7tK+8/4Au2QziKlL5QmJORfNvmj6cYgAjq6xS+iUpOjfzNskV18
xJg8RicYGcxRARRTUc6ZYCCInvLk1zfK/TqveKkBiDd2ilXbB6jgbL9PyPh5piKwWOH4ZmNR1e2z
qjL+VqHrs2EDBNO+9ZGnkCee5JCzcV+y06siHUX9P7IBRpn3AIws1imCU0S7GT9Gy8Oe9aOMy9dW
HMPNEdL5ahr86raSH8RPup9GyUzYm8h6MP25fyo/busIkGpNxMeXrskd1uvVEzI8ugWn9aupe5l7
2qTJN6c04HFX+bRwDNaM+Yq0af614122D9Ze7Wo/6RTXIHbEtlmWQcbBmxFazUPcPTkmnPV1eOeP
f/cUzSoj0Adse6QzSzfRb1V7VbftdTrdlK9eUurrIc5KdcGChunMzfqUwPNSAGwguU7WdfKDi274
7N9BFUQq58/f7X+2ZTOasYAADmDmNvImg6591ph+aufARGmysuETr7UXoqP7BZsfCbWH0EUexpnp
ThfkGHbSPLmqR23pJ/0i1eduxyCkgC6s9uar4NiCMSCyGY1DdyqczlO+TOBfXjnweLvj16msftzX
SaHyQ1v//dekvILukV96SnJpXMK5sqTwzfSMdLwJfzK5ftvdd/QtjPoAf4uyktz0F1dFvdZmsswl
lzBVmpLIWxea1pbSqhqdyKSQsC9bJDFTBLCZtmNNYqHvEWWokgUGA69FaVx4P38efDyNMebDwlPc
ECN7M+NLDhHZ413dDfN4ntfxMlTemz5ShcyKUKkq3eitXWraBEdptveD3gbG6JLxD0OzTj7vjmRe
kma8S0ILRsf8I623TNVu0XOWW2zrFohpDXYY9fG6zErr25xiGCn2vGslxWcoVuwYkuuQB+GJUCgt
iT7Rwfkp/D0FifTN3YArQilKr1GIuSIiGtbDb0R2aZs9oRHicD+SCS4rTm1I0V3TkohG+Nz3eNeF
KkCzYkrIkyQ2A0q4CJhJ4eRkFzUlulsYvKRnTo4Szmli770YoOCx6De1/PMqOicmk8rF1kFhJsSH
uEtb4yPVunJXJFZkkvxud2qH2+/mv5V2QG+/DX+ZYcl/C4+27a7rZ3fOgVsheAnLMI3Bf24dl5/g
qi+nfbqE7boElo466cTReZqx/mwks3vQ9N3QrVobvsWRvJPogSsWEppvnEPgqRwn1Trgk0/rtclb
CCIGcUxHaptIIYs/8GwY7WsFtJ8U1/l8L3i0yeG5bvUXYl7/+AxWgfFHVuKbD7ZWHrUcg3snqJZP
qg0OHvfPRNphb4a94D35FntW3MNfB2P0GR9dyqajH730D+7kEMFLXi7K4YbzaK/936vWxu0ySsKC
4lysRDGumKv+BEb3EbgGnSVNhZD9LfJn6f7aAumawrWY+bQFxUOVkLUyvafveVadmIqVyM+8yzPA
XQeRwkKaHT7xUQhsZ4rm4Ck0tfxSZzhz0WdHbX5BQqWCF2MtqF4UmknwZbLHs42S3OglIm6entGQ
bJpEGppMy/2+8KSHhZB0DfVr+XjWjrg91iR52gCKnHfvv6qL8sMIpxh083XUOFk0yFs3avgO8qmP
yzj4I5+oR+DNfEro3q9g/P7l1c8gKUQJ58z5kglr+MyLpQM0HAuOqkvazDaBMFETDroCbXq2f9wA
OBKMSCWMwcITLpcL2ApBA8osF/sA+xWAfnm6Dt6XlN/T0cjj7bGcSmlyoa+50cFb7iXPme0Lu8s/
9jOrkj/eRy0gFRBT7p/SSBHMSQomwLrO6f6Jd0LTJ/qUFSLvTqAq8GXgRz1xtuI+TjVcVknvmPkG
eSWTTVpiytUhdO81CTxTJETVDyOzSGD2Hh1byvoByFdvEF4fzbzenyJxj8PyfYbVOcjPZcpKLdoi
w1lPQsZ92TIEQccQ0/l7roCjMzR7mmCyeJ8a1TZYkMy5j1sGjsGAoIejlFgAdfsot+nGBoH/NWqy
WeNi59tWRjrAklN/UjhNY4LIjirrIOeXr5PoYHe4pIKyt64Ote+31DrVqM/Q8PgMZO62OcthW3e7
m8ztRc8Sf/Kd8Q3bcBWwHB/Y41nsHbfwvz8P01FwY/4B6HfnEi9BL1ai7fUl7+GWNJ2JZxsPl/2V
iFElBp+I63FAvuk29Q2oL91AB2dmfL0jlpYZxLlcNvXQjbNqmhPj99m5NIZ+fmKKZHygOWMqgPKr
o7drAR7lPeJe4HScqs0sqJiogy3WUBAlP2QJE5IbhUMKyfhyI6U32abjC13vOVbeIiJzZWitpITY
40TIhaFQEzBatYu26RdzKWv2/fK1agUvvztvksyfw3naJck6Rs032yAA7n+ycZdy3eKoPyjEVSTS
lfW7pQ1SwnwoJDk3kZVoDbt9utfw8WUCaI5EDaW7iiUVw5corPkKvy0K3HdwOKS7TcPH+vVpNwdE
2k+vjYbAYGA85H/KmBzUxQBO4p5coOg+Ujsn+nSX8/nI4Zfo8aHfl0mLMeqo2mTmH3p7tWRW1aPe
7ouh1WnaWvTOGskiHPNuW3q2fA5l5BPEyMDkmmbHrrImsiNfP7RSy5/s4b8a8+2LwGi15+zbIofW
qF5i15Pb8ycFCiuaZHPdo8wwq+Qoa1tqv6VPCHnuT1eKqhd331NGfS3muCx8Gk0WzNH9K79C16Gj
V7Mx4JOH90Ha4DLYE/5HEXnsBrnBV8S3Z8KrwTSc7aHPlHwuCe/bGvHoe5Qi4UAMViI3l4SN2E8J
yf7yYLHncR98GOZvZJCngbxinpmeX74UnUwenoglYc4hbin7kcq/sJOEIpphlJK2OdBrukiE2WzG
fv9tk17QM8nSFBXLIB35Wiz6LuUH9eJ1LRDYOlA3HTlZF+6tfnIRp8UbeFxpqENJ08Ge28+E8xHm
cTxE6qtTl3AHON88edgoBmjlRWN0JhpXhpHfeDag2NqlMJPbDg6nW0X7dRwenT3kY3GS225QBB4B
5f9kvw9AyjHOwlB7WbDdnmkh7tvRFgNHIyhDbzGnympiCA0Pkrrs7LCv4tAuDlGQEwYmjxS9USUV
nNfbOIQEXG34X5tyUyD7HuWxI4cMbGqBwgViYpokAdJZGhpLIQsrMmg43TAysDthK97+VkXN1nD/
xlvuG9hdC2IKaI0lBInkMc5hLgeAx+1xsR0V7xtOJgS+WYTgs+9LYHkgHjBZ1RpRywRDrpst25v9
Eh9f2JoMt6yXo3AW57cyjIeBaOwZhbtrgTxsfzBYgeW4ipI2+HDLxCxcRniDhcoYffwDxb9rzWxG
peFONUvkKmt0DSniuffgZ0Kyc9Fl6RyiXCsthdECN8PvyNxJ3r9WALc/Nt2YppSiz2szUf38TnIL
gxzOrH2BL8jTs2JoEc+9Ij2ZstfcJlTKQLkQFloOxsmz4b8vmFIDsFud7kbgCl7z8evAxFiJ0i6o
PXzpYymX53OBbUYN0WHhmb6I+fGxBDGMDC7i/xq3MXPWWQgl0TDmksteyq06d7HDgj4jZs6NYqcT
ahTvKR2xlP6/p8KyEMbWQVBEShsn1TZRP5YjH/5kFCzC0pPTcXPzGaCFFQ7xW6pbjdeP/QvxBgip
1RNPTkkErEMgKvfVPTaJgmzHG0fZZFWZZ360Qk/JmTGDeLQ3ZwsfOM0+O+SOOmwMgCzbuZ+rqHmh
U1tIdwBIhuqK3yZmfe55uXDOyZhjwmf9I1FeIORZIHGfl40EcYe3cUZnn6ZtYGE5tsD1RE5lWxzI
jRzP/OvU2g6Qspd+CPBajXXuGR8TsPtE5Mbdczvnu2R5Q2qc7IOzEC0eVy0Y1NEHE2zZ0+DYR7zx
/UofZaExnX5e2A/xWJ4RU9d8oF091YNYeCKRcZtVMGUgOidmcj36JTxhNm102TIeSlZiMZS0Z88E
KTv81UNDMozyNxH16wHreSOz9KlcJd6NEIv8ALzXWCZHhQn/D2xo1rAyenpH6YyKo+ExpctwZXET
xJRLz5vTjPadKNmbkvyXQqRaQG3K7N89Q7PAiQJS/F6BkErjuaIc4Wq+gPRnkzf1BiQCLmNqPh8I
vQIIE+VYLPSycGBvCAQB8JtbjEK9rgfLiLshYd8rGcCn8AgLZfwHVfrHeOJXR+ybtq50WhYAm2bS
3NUkG+AtxMoSMnaxu+sEAzOPldMP65AM891Y+S+zL28dGHk4Y4uNnckIA8ZupLO7apLohxKaH30r
9w7epEMNF+/GZzFWdV9SUWt0IUapDJC3es8PUxkylX7nr3l5M01q2UcL0hYj58F1S0mkUC079CpI
+czIy8kRzm6vzWea67mAf0bGgFvHCXLnYxfSwLxOvV0nPiJhqsFWkU0yqo5MJqUKkTSWa0GCeA7m
0mbIVRY+g4tQpkAUQlx+UvSQTmndNfkb+Fwg8EpDLqpMfhy6zdBG7XCiJZMwy87f6LKEkRl4s1Qr
5k97Q8ByK0z4kel7TAmowJlIeIx29l1UfXTulxJVTXJEC7ujZJ4e0fIEZPsJMShEfckjyroerxP2
nDetSinOoBGwYR/mljBEuUGEAw4U4KyCkf6QN4cVHmDyHotLL0MWbLA35kaurKLd58Vy7SlMDl7S
yby/G5/tjLfKqFlnt4mMbgrND/vwWmkIF8MTFWxk2nx/Old6ARVmSqfD1r/ZMUTG66x00Db1q0l/
XcJPitrEdJCrB/k8G/gV7a5d9T7Eix6awOxWYaBljNZUgKnpgZ2xVdpyfnJ1bqprhqX7lmtlnG+g
15Mpwu3zHj8tQ+nagaLaiC84RRHgNbB6FAcoVjHHkzNiSE1z/+zaYfXMvh++bO7ldSOZrT9P+789
kPa7QbtQ72hPQIMU3ydXwqo2hFrFdC6iirYdo3rDnChm2un7bw7Q/HAClAqc8wi+KWlX86WqiTjF
FlgH4Nn/5QiNEbS2vmf6aM0IYO+vajFdUFx7H00pJ/1H6GnroGgm2FSt7qKtjaa6Ae/Qd7z598/4
0I2u8j5OW2RcDH2IYJDffhZeG0HanJYEwZTSvXE3kmE1/05eGpcsRH5eHsDicQ6ItpoO/ZTpdt1g
Rmnl+oC/dxqeI/CCqzTK6ZwOhFDXLzVmzUpepLeDm3fbFNsy6ODwIVZireLWeIb5Oncz/IEvjplu
IZL97km9NU6JlVUdvL01iXUYKsQ01ItS3Qm2yBzTGKJgOQzzz5C2t0RVp+G7ErBr8A49z0FM7/ia
7Q1mno+Nloafdv3lNADkA+GrLvElgo1ZUO7m4Osg/J6Ha5/tHVVSWDrWUBP9HS1DM6m22S3a5uni
DwA2sulsXYq6fdu9TEPefSJFZD5r4Tuy5oiNfFkJVlKB/piogFEa3Y0G9b/z/My/bY38F8iJLDFb
NqNSVTUmvo2h1gL2+CwI8EtUdnwlwUe6i6RxVQzkOeiCjGrCO6C1QYopyAJTy6vdeTiiRcnvr/N6
Uods9ZRFe0cabez+g8sirDll6zXEl770om+hDAmnwj6MPqwP9hYR0g0tkW91D887sGW5AkovdS4B
XxJqYh0ATy7DgLcnArZ+a3QoyS9FQROqH/E54GL9B0IYp6o4ux+AjeUqg/hSRBNzzrncaoHA9kIx
LXpp3jVw3JNrGBkMojg2wZAviVLWxIBNu27ClgZQ8ZKkJtieTUq7clLD/gAvL9CninXg+MctVXCw
ukuH6uzG4Tom4BQh5ZPPUbRoXiVICv5gKPZIMiiNhFPQfUHoTcafH3VYZlY1o3NFaMYbvSNbUcp1
EIDTaomFJ7HOeFciMg/RkBjaZSMGz0uximce23FBp5he5MJHzJ5w9B8dWd25pTn+RBR3lIxGbRDG
QRLVGC4VA2Pt6fMeAa9t/L+F0Wwp3mdWEcTBiuPh1AwvdCSWBAwwSNsklgPFk34psyBgV6zZI8F3
90wcogXc3Nt7pFdEhrcV0x+NyIuZyDHRodCDXwWpxgNlu+SRaQU31RdoMyuHRWsnDln9CosqEcMN
pNm2WHowx3MLEyJ3vpiR1OnJjxr5Cf/L1g51V0oGD8dKJAYQzFBP4f1NoGC5ONx8jObz0Z1e/Zbv
SFILHmejoGamzuRrkKisFmiev+cNUlbhMCUrI1lB0WIXlVAkOijZUbLjPHN7LevoWZ/WWFW7guOw
pgx/LS6VdhU/mCj5WYX9G9tJKKEIs8AJK97iwuh+LMAEfyclKcdZnO83f6BNwpdm6BGYDkvuaWr/
7UMLbhu15gKRtb0fpqrY5s9ow8tLP017SeZSK19zG/mdeHhkevU8rB6EuYPHDc7sNj9m5rkl+R3R
hKPvJ8TtG9oTRdKUpa67HITVMHXPtbZV4tlD+XEyjLBzCK3BJk8+Pi97zuFCeWuyJO5BzrbN7HPd
R2FrzNZfKPH7cgpCWNODVijpTUhf6a/FM7a9tPFkv3vLRkGEvKBH18lUeNGHec09IrfvaKA/DxGU
IFEanfqw9cU9y5P/AqHmFdfKJUk4GKAq9/uda51xSFd75O615iTftFoJLRPs03Pj3cQ7T9kTILMA
5wYdozZbbRB0A57GFu9XuWiFXOPsUztgavSxkPgE0dD0Oq8ydKgevfPAyPvOBBcFxIbTV1g3ea6I
ORxDZTy0hEXwsV9dfaG8yp6LHthd6RcScVccCqdZXCfDbg3gCg6XMAd84HkMhFD0s8r6xhTwH0Ck
hIHCvlZDOzekfI3kZYqQTncbikshf0UpVNvywA189+DhRJil0/OFoq3V958ZxhUVxwd8i351exKL
VkN+J6yATSz+UnhH4zIDS7OnW/6N9NWJw4J9fcWXpVSHAULuUGClkKj+o7khcuM3IUPS7yqvPKqa
apw8zk9V7OUHOaWR1JRdFhzywczFslvxUOzGqvwWTW/pgMjarQoNM8iFY7CCMJf1fzhVj/YIXDSr
GK2OIwbswLkdb8dj814zA1bdy4ESrnVgAha0VDoyF2Z0RYoRS4wLAgB4DkoyMNbaz3rgf3OzKrFH
Iv22EnD+4hobmM1wH0xEg9bNXmiv8lRgyYlzx66tRLdUdE80Wowmx49kZFeervYwjJTyb3iaOyMs
fgp+k8rdVg549DyQpgcy4r02/sg36xFCdOGMHIyRWUf/Z4lVtQGHqfnAERpyFwRhBolQ6dCDuNmt
SgI0WREYnkiclSaG8qdVw8j7/vJG5sawhHq698EZuJvB0G/oB7mBx4KwlQdK2HiePjkWoQdh+sr2
cijJhA4EXo0iIP8beata6FROcCNeV6eLXGMS/YhOHrue8f5O/xHFMpmRwMTuT7BnbgjAqHXGKsmb
8xBdJZ1tYnqcCpZHN/ae33Po0C1KMD02LDBvOz3GPmd44Y6eNJLnZ4gC3f2h2PW+E1jfeJMve7Xd
/4jvL7GneK1knXmb6M0HeK6+3SKsbEVVWjxpM0D/9tkCQcUynchjdP3VHiDIhN6Q9ts1439WQml+
CZbFZ6ciiwzwIWiDgnVEZdT/FCdT65mXHio47UQCmyAljhfcidzw+gU2E3KelvvlOOW5KM+9qpJQ
G6n3uu3K4g0zIh72u0dhnOSbeju1WpJsBBcSPUBPjcWjqWBJxEzbSWE2tSdK15RgJoJw6L/gv7OE
fpD14aA1TcuTKoIT5oly181xcMrfEDgsTeptdq227+qa7lGYdnrzsT6EybHZj+ks0CYM3WSaD2r5
TZ8MbU6ieXxuFwWYj8l4ifs5CWaYd3155GkT9CZam9GP35COmfdD0e4+rcoPvRJmet3lcMGTUCVv
ZBlg5PBt0riZGjNlH6oNyTLx50bWkOOeUw6I65x4vQU5H1XAKnjDw3EMqjOgT7PchxTrImT/pH4K
d4q0zNKuLq/dV596S3sG3SPUA5fYh54y9kEYBjqi6BMey2LnL1ov3XPrtB1rZ5AK1WGzxcO+Q8Sj
9pcq5W+nTvFd5bUyzhgzG84g0xrxHwcGDhZlOyJfBIgb2UXhOtdNydqz64nB4PEiA/ABCuyBoAcC
mv1rfGnTA1aJMg7czo5E4nIISt81PECkTMI4VWZD0Ib0nPA+LP8yma26hN3lbjcmzu3Urcr/V/JX
eDDrDcibX0kQAiK99G9RCoyqtX6NkWRKUM9VEKFr+l3zcvLbgkNGhbPsK4/P0C5NLjFi9kvJK3f8
zOFhe/9xg6AknMNoXWMVTRw3d5w95vZJYyzvfln86h9Y/d0EJflMvn0MTrYR3OBlZEVvSgFwLO4q
cbznI33VYTJ+i5XUH66S16CIPtsx79vrx3UILeQBcdlvsfUACaV6qtKlIHE0woBTZdw5TSiqI3Tr
PQv4VBBgArNcQYe2cXE4PFyM8G8I016wVIUSeLKWjAfGZDVRT4aF1nnxIBXXjOFbp+7OTMotV0yn
9U4uSQOWYZiG8IXhh+7hAw5PcTHpHTlgjssTCrvtADeYijBC/TUd9Nr8D0G7nFV2VFAZdsMqwPZA
1AN+VbifA8OYErkPyf5pYmcjkT/T0NhZSg1uGt8VfJRPaS1kSoJqlr3frFzJnXQsisx+ygIE8CJQ
6MtzqbZbmYOSvxyid3vFJRydVuLc/PD18o33FT76OeMQZccP1pBUiezBzYySirxNuR7wcyiJ9aKI
GWiWGxyisV6czzuLVm0hoWRxAGUPCDn0mXUidpjYFOF1j36iRbTAUGdsEkfUrARRT6ecT108pdnA
f3XsG8jTlv5xKId6UPKSzMqI26VfYXBMlJxXLECHgBBf2pYaqJtfty7ijYHm9j/vzdBBVmYtR5zV
e0qQPvE+wGxOMwtje5K/AkO/GBBjIr25xYcsAv+rr91i7QRSWemwRI3OKgh/D5b8AGKDxXWXFNhu
fVlAmulmSsvrpXbJkatL0BN758dme6Nlal6+PqL4ySPxqaYsVzREBElrwBcRxwYp0FLqqdE8AFNt
C0zlDQHeYMsSspXukoYvvQxlZr8I0Oga2ir8BeM/5czBgsoH+PG/676rbD3QDgOfwiOyMJU9nch1
YZSlTosriJNruaOQjPyQVO2kh9AwWz48tJavh/lyU69l0wH02wYIY4uvC4X2OqNuUZ07WW0cqUsT
K5OEIqeSuehT19mcBiFqk/P+zSGaPVQeBNyC48/3xYqVJZHw9JQAfLT+ZYB+FWCqUcsea6SEdYtI
t6DQfTr7//pvU2tGDIkS8h2LOlaxSP6Xz0Rh0T0oKuSbwC2f4bnPZ9ovBDnzhuUPxJsZSiBvV8vg
qS2rSDp7dbgGr0bQ5VGhuKOZm5YlJALrTeA9QYcu2A5CQf8CDL6BtQ8MCapLsPnPvOdgmK4qr/MD
GFWmQ5psHHiSJ7inDplsswjCpXoLydZ878Et7XIVyowwyg1yYhdLWp6FAXqxFF5H08PwLsbknEA7
22sTw/yA3LG6j3/mjjEwEXDX+HV4xf0ccmGiaVYkTnIODvbQmCM8Dg4/+DukX3BnPacQ4P7histM
6CMYju7CEouCUrffdiVE8netPIsxU0YXsUXbsW97cp+hyJaztwNWDQJALHPzGJTFwbds0lU9O4f5
ByvooMH89ddbZTwWrZK88Ic5AP3fyvBTz71bO9p0qQ8MmZvsP4A+aSalF9YPDoomj5n7FAsjrAsu
rLC8lsGEaOkmr1S2NKHMqvM6aEVsA3cxcW4Ar5o1K3k1PFfuU8Or2V4m/T5IMaCAE6hgXbmJPUnS
4HDP8IwHzoEV4vf8rmQQUzTnu+knpOFBJP28dd9xpQhmGeGZqLHGlZYT6kVx/Gr0tgxJsDzmNipd
Jei3C8mxYeJJkOyJG0I0bw9EV99/9jbafVIE010d8UpnDkAxcm/UeOelCf9g+x051f+tomcl99N7
HE8VVUAFlK3Hynnq5TOK4lKtsVcJVCeO7h4M37SW+nSIF+QCRRyoc6ClAz6jqFT5TfTE5OObu6Ah
9NSZvAgBuDVctNPBKxcna0ubnv2J6rwTk7WK/XxzzecoWp1PBPSuA4xoiIw7F5CIbhCx1vhsj2U4
PEgilk8L1ZhcvrBwfPdm4uIEAHhWLCw6bJdVb+0Us2le5a4I4ENWAuYJW2dyFrUXLT0EX9bDCHso
oCvA9NNgz0S8992OhVD/5+2nYWF6iWFxeKycbxqPQzvF7PnuH4/2fJPs4JDdgzv+6tqOTRjYYDOX
9wB0e17PwBjaBiQ5HfzuYaz0uiOzNI2HxcZ2sy/7rH9eW05nUOlXZrRhDyedZyfBfayfDK0C8QmZ
zSPI92+KV3gtnZcytokfVJqabp3nV1nnvKCH96csmBIGOONtahW0jQYKop9k+p4BHnns6c8LGfzV
XpGF61eR8abQWauyOf0+ajBb9PZNi45DI+EBAiK73G9FCULFIYfXlEjAAMl9s72ekmoBZLeNOwUA
RfWoPq1cydg91pPQ8k5OpHvSpU9NUHGT4gRivqaD5JNCbFU17iM71x1QUGqA8reoQi2on89wbQjx
FOLmsli0kYtCBjq7AVDczu2YUX7lsjvtOa+ZF32XIKClgSIMH/S0dMnZzXVCJzXPgZsGZAoMZ54r
z0QFj5d4YBHHAxNPC3H9sP8XmMMJRTHyEb+QDjF60oPX1cnz4MQCfivMQRGbhJaZ2qXIvyorJaCM
ujuVRgeWh5iVDpjvZJAhVNtqlgBU44gr+UJJB520K38Sd/hHcvrjktr85xtqDxdEySufXNPMhOI3
bY9PUpz7JVg4efrc1iS1tQLxn0CLjHfQWw5RQ4pcM1l4UCsMMxE1xks9/pdv5JwIwopuqvz7wrqM
1eZOccRETd2MynV7to4opi/Qv0xp/XfvTbXXsYG3YMLEdqPYmEDlx/IG/TPBUpnHgxPo9+dLbZeU
wD7lJ7GgSIXm9Hz4/3042Orhap9zXggcHGnvT/2MLOQEuDQtCnCWL9TSXiKDnoSVdjTPUoplxRSY
GJCzq0/zj0bZqPx2R6UnISKTw6JgyJv9EpiNUkGQcx30SXzRtie4JLZa4ag+XXntEtVvsf0jiPnv
d0GZvIGWaOk1/hO/UGR9Y/0tC6Gv7toQhtZRCZlUFijD4CyNuBrHjCXlYxOJ2r3UgIBmkOKUJJO8
FrJOI+vSDjTYZuKKho9GAkLIDGuAozad0rjKrEX8E86j+2X3JWFpRpXDBKhoA7X2xWWcJZL5M0s5
9m1H91rU/mixsT5goL3mankehJb2ThDtuq2bX7S/o+U7y659RkPkRtGDZazaqWAoJ2ZWoHQVy1aD
gYAKNuS8Aa7dAOAtCZTQbOkbMOFU6+NpBnpy4WLTnhBZWwkwX6Mci9PaRg5GhU7ggM0aQiit2hbL
v7rDrS8TWJNAiDfKcS7Ps/s0bNo8v93XghF7KJMahCsY2Wn7MxLMa8sWrXhFN3qFOjgjaZQ/RsFk
+1slYfRyn4nNqUyksRPoYvE2s0CIU0QRCb6EDt0aninBhWexV75BAplgQtfUxQ3P6XfN7QW4kFOQ
zD7lePnUlgBob5lbvn6znRCbgeh2ApDHyMZw5hxMojGutkFBMpUNE15xvdc8lttmkrO1uvQt0+2N
pk+Bkbjk5RJEErydPPnvKPbUWYyCUTljUDhnyStTnH8DJycV09h5Q4uWD9ITVXzMAxk/kgwMVg5S
tpLwTIdXpeUZAaxJ7gM2SK+pEn3HB/zcbkPl09ZckqbrYORit3cEheA3dPHxjrKGMTpfWYY5GGo8
TdC/nNxqHCiMHtdjSIsG6/l2b5ZvtFdf4Ce6dwWCuUoTi3ylWa+MWXs/ZKwDs6a9jlhxz/WSmMdn
b6yksEeT7iefamVYaQC5iw0KuAAVH2L8OOWDi4YKm7xQti2JfRWTtXWXl7Dc+m+qGydY68gmzTzh
5m8qknqG6gRDD0RtDAhmckbDw8n2adyMWabxQn1CNTiAu4ftsJNGWniJrl2DHaXYuCRIxXJvP9QN
o0iOwjIB7LBQeoQndwR6xMXIHIAr6WLDvyTCzvw30hhz/3l2YnmMMv5zRDwQeufYDrzxZuId6Vb8
/ModIhh7KOStxmv+hnnj972tMnv/9pjPNL5cBEipmWFirckUye1bppsWjX7XkXijMN0TGOdWAIeq
YJ6PCsI07xbx9iXdh1h0ne9l2+oAANgQo1RplMaTBs/zo9z5yUEgOKYzrcZw1pSLaOqnIKVoPn0O
9B+7OyHZtm1D3ZZ6X/I5HWyg1QwhSlNK6X3twtnnlcD5e1yh13k0kIwEUKZNnx7p0996twJZP1yZ
Gs5guEc4cw/kmCZP7x2QuiI6Ez+KlhReUS4id7WqOP/WT0dan9tgGS/rTfPu4JXCBJfreKR+ck8x
S3EFHoVpAJ3NaByJN12ULYDByulILoB06KCNJw9GLwt9g8cOyx9DyPZhvayMQGXtEMT0yB/fVl+0
gZn6UUDx+ZjQoXvZZYnvh3TnEES7Df9FZXmGcziowSdBpxC0wL0vlomyVOX0wXp1KPLkoZs2A6Sv
UGMSZ2hy5iUYai4+raEbLO34eOZc5rxXQvJMtD7//6sDzQNrrcJ91fCfWqRKHlxq7Dj8W8vBZWI6
xLhBO/hOiYZl4Ri5SQMW+jgG93hiZXYVhfH5vwwcMr+JP2maXG5dc+onVPg427CP7W6ZuccdDcOy
CEQprlK/OzmcK5hcuTY33ox1mscn9/G65/v+gQiF33qK1a8Oa5ZaPcul+3iMbQjz/5h21OjQQNLd
w1xE7p4HLaXiSOKsLFa1R6QJL1GjDMWd7giFqOzpNUcujy+FwU26rk+Rg3tQin24HQL2B0fHtgLx
JhBCBlJvJWQqccfkn1XbCimbGYNeEj+rmQovWrbuM/v994fZoIImfmvDjGqWLuUYq20Mgl19MKd4
8yC7BsL4t0R3Drqv7DciIabL4ONldNMUBzb5XCBJA7fvh+IK9c4/l0iXT50KC6uyJWctsGqxBJwX
MXVrX458euYKN91RmnWG8AMavXPas7sHGvItRDj0O39mJxNtYwwMp5dCTCyGsfnHxnPTR2wHhuOc
3oQm6HWLfpx+/VLVXsOt+zH16rpB1r4/+Ep38An+CL3NxxB8jfJ1K/RT/R58YkpHu7M5TwzAGGYn
4m2SkWwLq5ERDgx0M25cKVK9ciG65dB4xBjehLGuumjLSCXkZUGQ5NykXqrT2hvZrH7PdT0Ea8um
hYXyhabCZFHIyc2zgHt2vuUuNCovydBOv1PY2BHKqM15lr64uYkD0/x28L1FPWergFnyOIlNJf3h
GMa/NhRHtljRlsyZgY6GhMaefWDgTylRBM3aDhrGVOsjqWBceyfgCgjQZKQdOCiGtVH1jLh9j9pI
Tf0gfNvxSpSy7G23b4pKLVcc9TrZWuXdeycFfO8sDlaEOcl80woDgG4wQ6wUF72foXqLytatSzXb
LdqHCNALFxsT23/GAQXIncsBEsn9o3RObOhn5To3h9opL38/Y6I4pdy5s1OPce+RTdzJwoJGZlmF
BqOMeJlGmX71YrNg/wypd3xz7X1aQPUSocK3Q6fPo2JkJJ4cRkMxg3A6Hn4lbfFS6tlTKCst3NN0
j9p4MUS0RNVuhIs+7v8ni7wkN5+sf8tUr7jzxLC3vKz6Z0xiFzo6KieTfIbqLAbwqCH+7O13qKzF
ydmtrlMV0vmw0EwznnyZEqGGcS3zheBuGc7udklzDx5pe3R1Q2RszQCocfS0KSgBZfPsrDdICMkW
kLvnfbQTvf92GL5BhiLFDvbmSEFYHy6jSZWaIqTu6YTTDTdOK+r7fxxv27VIucqRSqSLCSNDZQci
xav6QD1y4j67MSnx456d/BtIF0k2KBcZQGqVwn7B4Rm840rvgia7oEDw+g0vtF7jv5nhMy9t4LtW
VW1YqtjSFIdc7cVzZXdlx2hdPe8DROhJG/ZA9Ot8t1R2+6ujqsbdoyEl3Qr9oeqXgviBoVCt8dOf
vuCRtBL46PvVbTAGYX+b8gaGPXHDuIPWstCi6nsxRAS9c5XMtU5F2nSIURpQ8MFShdn/DY/8D/t4
Plyekk8tzdIsnUDKq7fNRhtxMNBQc08bkd7/HxByQQpZHOeR/+FUinALs66KNS0AR5GldE65V0sR
Kew0FVod755WOocgL+HUA3pStdaW9aPw3GsDwGn9mhkzVqdAs6JbZZNxKF+rn5TlzGPBSoNmAG1j
6qjVUfX9OrDgkTjeqNM+p/Wzm+d8zwXTewxb5d9l7dfY/6/RJY8wSgrn6iiljwbZnbNnIn5jEzAP
2hKlYJCQ24xPPFF8xBpH6xWyksyW3tv5ULngt33ShSIwDRy5oR1Tv55x1+HEGzMm67tH7Xj9U8L4
sKhb6MBAhVe21avIjlCNW/anHs2+ftjUt6CNmviCkhg6lBDl8ECcbLeUZMTqg6NS7Dmrh/styMm1
QKHpmDfEGmC9DzbV6PIz8ZxW2CtL6EhU/gQq6u6inPpLURJcfaAadjbysP6cw0cHBRZa9T/sUThi
iDow7jqbzp+yYpuTuRM3dcFBWaBpetkJd5a4uxTkw3fZKwYfCzrb8pHdD8wgbfcueKRXGYrlb/IO
C7FyF3kMJHJVNP4mJ8jWotYKrf7QvR3yRieHjpPNPB8u9o6wGwhvA07KYpvKwHCC1kelqbsh96MP
rFDV4PG931ZT+HqTSU7cT40VcgM21AGKhox8DircH2/1wBPCYshNo6l+UXHxm6rpif1PUBvnbSvj
HaXoAxX6CNdghfuMbCrmYIQ/ntPpaBzrC4TfGFrXSXXNHekioe5Sze1ZDJoAwIKDz+/XJYHTzmmK
Z1bTojWRMhCD88efI3CV5niImYBwAasVuYyR2V+Zw6HCaeZtrVcIX/qP+BapJR64jULIkRDcwlP/
KtspdKspVQh6Bj3JYiQE80UAIk/4szVfeU9u4m7GqypuMVM4Pdcddohr9QkzU44sbKT9HZRlYsel
T607K8RNhxCH4CIH3XxVnKC99NnwxJKuwzNb/ANwr0pXZ1XSuzjph0vBqhm53IqdBB9zc+z/cc09
zWq16ZDxIOgWFVwfKmbxiIa+9yUVSxq/NILleByrzoagPL9Iq8Ke04Mm1T3REWWJA2bT/4/sONPa
Uj/uA9trFQD1w6y8jMm1IVR/UYGUsVMgDqZGaxD9Y9h98/vg9tJOO0If/lKv0knmVtBvREbuPNAX
X1menDD9LQgfW1nHNssk4vqG5EHMWrCyyIrnwxxuNcwCWp9a0hi1egCmIDb0lSQdtkUq5Zz+vJiA
GpNrgTsPgwqlcvCPwAnS3dbNxWR7hUWslx2OtSOWe1LjBU6pm1zMDs6pHmnMMgA371zgD3//mJ10
sw31KqhtjYRnnDpYaWcYg4gMEzZRnEYYewrgd7acgGkDIHiQrsWOMgRHpAK2zD2AJ5HP9yeD4aGK
I2EU9cTP5HMrAXiKNl1nfWBTCv4Kf7nSXX6gxiE4YPdmbyuePdDZEyMKftUZGdE8fC+VwmZIlTPK
Veq7NTzqB57fVuCKuintc+DjXG+/KGMKE3sGocqYgNoH122v3Vscwu5Tr23k94+9g0jjd89Nb8Ix
+HLvbR5muh3J5T3876jRfoRU32zR9nY84v0hdHeYPL5BsQYQ+ZwVWK+ToPOxDqlvvQfY3uqHHNzn
LtNU9kuVhnK0CHfpyXtFxSz1dG4xkSFbU39mNRAszyfNr90IffJFwBQea9ijcku+4qZy+9OtMtTK
uPkDbehi/iyj7X4klyhSISkOvaMGvNxkfK/0ZpYi8kVFVt0jbbzhH9KHMrW1/iEbic+1eOhMJw7/
BxbhkedPEr8bffo7TyIWMPy90bYzUU4/AvytWe9DbpQ/7pYYs4hIdm06uac4He/OZQjXz1wtOHe/
cn8kWG22eS9OrCuZN+2s4kVPJGNR0liK5MreDIs9JJGYvLLWiKVCqDiDYoyGcFNkPEWvNBMA2heg
7XUsopi1CLsy7XAJqH48do0omfk0yLSQvSrw36EbEJ8mQk2tbGWm+8uOEoGM070AcoD+VLrSKfF3
NGzApA6AYQquHEMnxSxBxGIgMgZBEFOWhzG1c1+tkvm+vBTrV3kzDfK03EmNAFJ16RC5IPB5bEGd
/XhXeY2HT6lUD0D4GD+dmIHaATcy5djjkajJHP5yuo5dF5OXOiLFEZ0F+slnvPGqyAG0pOkATwbB
r9b1brNGD159q6D9f6xFBofh0PpnZGDe3fYV9y/OeQXvw/YjtIl6gYg+NhBOFyFsGXjK6PBnnp5B
l5aOYFWbUHHKBnXEQY8QORIPLCX6TgNGAwY9vbUuURkABIVAa6acnNRJlQTUpQ2qHV8OYgOlqYle
i4jb9/aGFm9xvVuFJAlbdmNJ0fsZZedBdJ0Mybmnhy+F4NB2EKRy0EI+lT/iCvT7WsmalNUPhPRQ
mEzRCtaRe3RHTTnxMdUuB+GPqis3ksg1TjlDvgWlXYCsel+Iib3jYWxVlaF1EOLYDZwmcwDMxPhY
gMN5z1QRvaYiT5hPZXwwWmZCq0ZN8r8cUT3jQwMwvDGaVjtevMg1ciqD4Kts6ZModdpe5SdahzPb
sDa//fVlOJDS4iQKI4XGZEiV8m/vdfpHnoVYUL0iJ5RYW1ticTqHq1En1dVwEBI12faSd4mBY4P/
q2Qf2epFBa/B/YWKGO3x/CIXFhqmYRDs7N6N+NxGziR5F/BNSM6X2Hm+f360+BXHu02mvSJRe2o9
2ACWC+eIEvyWZXXfo7bU+nPfw3+CSbfen4AkRHqiiIxEB/vgPw1kE859AYp/xLrMYPhgk5gIKoKk
7LkgY//9SWjppUIMxnFZbGRp80ZVEqBQISCdPDGBUBmeE4pAPe0KKg0+V1H3vGtD6VosuK/HTvv5
uOw7Kg7z2srbKycVguyiaXqQC5NZ80CBPvBHq0LuOgh9ySN8rflMdqu/TWZxrvYmRgrf+oONluCR
2f25371X+jxQJRnpvLf4QF3ljVRErDAqs6MOjktWz3xGSFHqu8AW9hNPL4h2RbccZnTg8Qrdjm15
7RE6rtHm+JKYg64wSq6CdElYdCuTjZwC7sEfVjt+LrHudHQEsCwhplKPd0qQcMgMI3C/XOLR4OOv
5ac+OOSJuHtqcHmZLOX3zll78lfd0u1+/zLybFgF/cUM3tvIRK2Ab3TQVh4IDjgqF6b5ryL6IuSd
6/1y2BhzX+v8a+eBWOiLQZXdfV2M+82btQ2IvDy/RWH9xeUKw9S7cE6y6wyzWxw9rPtQ+Dr/AlKN
ZKbBu8IFMQABwQtzFxShntvkW4MHEAaxhjyc4070BPWvBGWyNXlRxIMBPUHwHO/pOnI1nNiuqAig
ls8uCy3u05j+si2yt2BTUfopxxE7ZWxDdWzWQ5+5ZnUfR2eBQlmziTYZEyCvFSRw+lt+16lwF9Vy
v41Kbj+p4U5o83X94qsgvj6r/AvjDvrlwCMKhnEyrs6R6xTynR90J9yULQOWGnoVDKYfmD0Lc7Vr
xxNXEqBpE9GcFCFK2DN2+3F49x6pik6hJFhg/jk0UEq1WnyKlSEsA48WobE+aGzvK3wz08wKt6Ax
L03M3/vAlOm055YZwaaLdODWQv/ikdVhhjw+dkkKPc1ELXP4hTCyGsD+ZZn8XArez/PSjeilx2zW
Ty5rS0B9HW+h4l+5L/9T/k4BFlcARDCicmtru3DicPaQPbcvQ5GoXawpwTRp/+N7cIsn28z7qpz9
D73IvoH/mYH5hUZpVe9CbU2kHiMnOIvQtDhwFJahfSqYF/W5CbWuJI3ASJEgk4iX+YarQjOq8egb
yxn8b9cew8mMURK/6C0rRBaNIBAh5LgvGjiIujgurTYShRVGre3qRtw/7qSlF19Qm7NAjnsqLQeM
MtbrJL75cPXMsyGKpugpjuAh/rWmJLZMTJ8Le50eFL2zBP+vC6wvt27qn34M3513TTl8QlKGuFkT
jKYatMZBzMbUZJoMM/MJaEA4k1L7c84HkV+K2btGCkj5LZzqBNLSBSBBPbu9y2v3LysPUPdyBLil
0ZySngpGJ7uQHluT44HdpAsM7T7ZhtFrAwzdB+r+A2dL5rZggk40H+Jl+RnmYPPBmUxOgkVIzNb+
BI0dj6prxm6yNqyOfwxKP89UdrbdHw28pfDt2jC+cph9pCfPqR4MN5m1PnCfw2YbSo3q0Hu1e9Dq
9engLnK/6rvfyuuHTVQU0IFuH3R33pwfpHtstJYLao4lzuvOxBznFw5G1/0wXgcXhmIrKUwqqbHq
pdqfQQ2lMEla6reM3Q9aTG+olbj9hRfcZEvLQJWXgMdhPt6zfv4HhgkZEMygyEjsZGr0M2k33VHh
FWBHhFDNhhdOGDniJyUkoJlxGadYmDnPenlhdrZeHnYDeDFGxCHDs/WuPHXjGdyBa+61KlrAGlBx
Lstx4mZsn6w80Ebqe31KIuZHIpG/Fd13aCKyAAvrpVbVPqZcTkXjE0+xONlKgm1EISkc/6sjU3OZ
5ZEwlapnNk937UII36aFxZcX3D4tzlz9GT6Sbsc3Yle2w/6QSE/Nlgvln2cDgmH/aT3NSXxD0e8z
w3uhSFmL4xbUk+JLN08sbzTQe+Aa3xuVMpg20xjkNp1zY8zl3Ge8Y/HzDzWdgwoyPEafaqEGbuS8
zs6R6zTD3F7jiEZAx6qOqY5K2zzz05VbQI0QaJVrgYD7oA7G5ujdV07pSfS3CDlKJgZS8CWy97gb
of26JPszW7bfQ9nF6bzDMz2uIA4L/bCMG+FvMM+AqDZAdFb9RxhCik67aWsYzfkp0FJpXW6/EXJT
r/V7DdVeGDetDAHB/tWN8k1Pn360+V0KtCZkJqwyiVst/uhzAx88SH967G4UEFsAojSa6f2AcWcv
lZpagZOatTZWWOINYZLSiNgds9UjguEpfIWmjvUndb2sgObIct0NgqI1r7oZ1jwngexIZRFBZduf
VOe2sDOSaq537UMdPqGBgKI8icHIo9hsKypnpEUzizJRAFzXjX7gYqBIxtRtip2POG5aV9qJAlfR
SgnDSeAaJxcOT9/ZeEaPevt6Y+QaUsO9LnVHVeC+eVBxVvoWreJBKltYTk2swRCZtDBm5POlmXP2
+Ujfw+WpSNMMQXxCB9ZiOn6U9eeFFPEYvz8Fj656Amwx085oyJJtzyIyCNOYuacjiCQ4VOlOXh+s
DKpKtNkRd1M2yBeGyhjc0RmaGuypcQmNYwWAOHMYpQNEFRgPcfAs1XoBvoaJISwvZcaAzF+k9yM6
u+LEFPtYGGl2Il3N2Rk+EdIzRMKWr7CFfxAg6/RIhO/Bn832cWe28unrudVDKsFQ75LRxVBVVMq8
WY0YswgPEfiB8P87nnXmDxbCz7SW+CxXd/R1/Ia30GiE0T+HrYU6dBvpHyl+ESUdY5dww0dsMmlP
nBnHtzJDQfVMqg4GsWSIKUDqKiXWx+NFk+hjuoWC8rtv+jyyISFWX7b9JykQimi4d0gy7PghVC1G
XDwTrAF5/YGhDb3pdG8UKl929sRlUPRQZfNhBpcuSCqIUr2Rg/M3J8fBc3twEVYNYU7ibr0KnIh/
hHHlmOVMqis3uwf+bbg7u1j7ry0gWRN8+ZN0nB27gyx24alBFcuUN+qPh5/94IRStvfRicfA+9f0
l8AgPwH/8UNsrh8fspvLRdI8iCWUZc0rJLcndi/k6lXyBAwZMHafwqV1XsAVxTP175ZNWw6LA2do
zy4QGXilfDjqIhSZg136Nht+1CfDUuefXIaSEyO6vEg0lfHcDPUYsefnmLITcsnyiQNHGnXjNLC5
kThqVFx7XjascdXJFS/5lDiarvgnkpN+s3Wkf5Pd7N5GeaYGqckvp3xFH7YnSZQijK3zKdwfd7qo
ELHrd4sSe9BlpnoW705O04r3n9LLQohLjIBmcSBHgjsfuLtr7EZLX+Gpk6gt/qHeBkukTt9J/f3p
+CnwJVkHl4GnZfvY3M6NbgFoiFbc7JTmVK+EkcoUhvNyFEQD9mpBIKoAxIyu6vXhPGcb6GojSwdE
liNAUiZkKWj/JWLwpeMYTCX/4kIo8IE7AgBWsmn6LxBPNJ+GNqTSuc0zHS0VjA/tbTlZh/CSLViO
UmCk0AiGwnaBFMVFG6mXDvfNcpywvknVqvsvZY+YGP1gLDrryzy3SoO1Z1QOLSKvmKQGO09/m73P
WxN1qojcyIwuacOqvwCegmypdvTZHzvwJBr4XbmIukO0ENUSOVjkJrVv151qR+sGRcMyPrazCTb5
UVrl/lAYxUop7bAJd7HDpXaPXwTfaVQkaCjNySH2OOGHsCCY1AHZI94rvE8q57jtCMrdcCSwZPKr
DBBNno9o+4QUefWOSiWdQh3PIAM5C7VaztkEwpMZzw1U4p4BFUh34fBrmpJj32wV3wtWmc6gqT4z
54mVPDHQIPiHKWydloa+Tr/71YtwUJnyr6uCDAekZL/ge8+ZkBxu9wBEI3Obv7VlssvfJ5TRE+9g
6WjntDgG+42Lv+Cnp/OWvKYcaOBqR6fiMFNv/OZs/vJtHkxIP3/UHIE0/nHue9WW7FpLuOYvqUwC
La6XIaUulwE8saq/AFsiQqOshBmJZK2RbYWGDsfRlbLub+qFYpoIu75P1xolKgPHyNmjAKfd08IW
WyJxMGkZYPW9eYpnLlyJ03QJNnEJp9wrTAMRaVeTKDMLRcCqW9gob5UNx8MjBzkL63no4FngVX8g
a5AODYKGdTNn40Jr3a+mDHHDnMkne61i6fKnY3Uz0fASAv4n0P7nnGHyzif+gnQfYAFFt9ginihK
udUTw87GNjP+9BD4AAytSSB+NdSy7A5+ZB7boEszRzoezmua5VDVfjH6Kquq9FDiIC+l5IModA90
d6gYPQ4nrEmzu1KftZ9WuhTtY4qOE7F716ac/sfgtLDnV56FRkdiOSuwvfLVUkqtzBWhIZILIc91
M8ZLd/GyDI8C3hCLk5iTtVGoLlCEGlbrOOpD/xMpjOQczmLlJm65F8lbw/VPK2IrnbxZiutWLStQ
FlaaH6/3EEv+FwihUBvZPkkL0FEa3Ae3yd1NrqnqNWqbICteVrgXvntks5u3bU2/VSZbme3OR9hF
ton12pjUX4YJwaUn+tt4oFO0oAf6pcULl6FiwKt3bkrxvO1CGaB61KKqDB+hrzAQEeGbw0RA8wji
w6hOzJUin0xbBTSCIzrhS7IL6V+v3XU+2b+4WGRgkwe1ovdIMtw2VBdxfPAg3klMx2OlQTAsbbWO
XWzXHkxgpckhpe2urAuF4ey7jnxWCM8JT8ivVPI83I5dV7x6WILjCo4SeWda1V51raYNsOnugRsv
hSoyKAya/8xtqoBd6QAMqomnQY0M2JcFVoRYCW9y/X5M8XyiMiCEcA5OwxJx/Xjy8ivjUYXnWjjb
bnNVI7FCY8AeAIhg5CVdoLeX2PdLcAofUEZuN4VkED05P6NrN9X5jSnZtd4UwH0q6UPnQCStOsUK
ANHrYYzoHZmbhoCPkL5IAdT8vaZV0WgzS9+jNIjbF6TcV8Kt72srnQlu+OIN262Rc1+Qs6yNZJbh
63GkJ/Hj7mrpTGym6usOGfS8ksijKkCu+q0/vEEBoUpqm4ubK9mZnbcFsrseMSQFUoBX1ic8vwmt
YlGXCSxGOPOvaY7/L09nTWtQG1dAoRlj8HN090OImTksKkOVUKRLwKUnmTY05XbgVK4oWej4jw+j
MMtEZ0lTjksk1WzffmIEkCafk7i1aexey7CR7NVGiidAU8oESK/BGLTepTpER0xUg4Nr9gmBPvHE
mEfZc/J78Cy6YuocNpu9VJGrtkuRUuleg0a7y2HQ6fpD836V22Qo9pYgPo3HdETeQeyKIkTVu17Q
AgNtlp7eHe6OsYDd96YO3QUeRRdBsLDVkaDgZuVgFIo6xVAz7h5SYWQJmQ7az3EeBH/DXLMpMXGp
EW5KEBqy5bMJTjq9rHcwMReKpCzjI8hWYfAYoKF+LMgFC1Ruol6USopPxAiz9R8+YsXH8fNntldC
ZGot0mkN5ElTbpMxs2o4MfqrI2BfvscQOYimzk1s1gLl1d6t7j6nlyFHC9ZIj3Zpt06TgYeilB50
msISyh2wtRzvQJ/VDPH18RJXL+mIM1a1w+AzzxBSDAV0Fv5jQ0MEFrntQvj3crcTdb9OFxFn2cel
QSlfZwsdlbX9yXy4ReN3AbyCrnV7mXakNeXfAPGOutzuzHMETo/IuoSoPpD5/Z8BiqxtwVOh9Q2p
SCqia04V/Z+6muxQLgnd/ZM6cFJAuqMxbqMG2z7RPvSg/DvvoJLU0z4UoisRyP4NlqFUyToBr5/0
sZHkhRWlWNHRC5yCh//Cplwi3Ovnn6LuOMWCg+eppq98ir0f7Ctk7dDP/hF1s+/JRK9hIqMYelrU
Y/L6gffElM+GbYzuxr7Ko70OVlkkoLNubaEme4dSn/8MEqVjG13F6BRUqW47eKFyx0siAQ/+x+NV
/dpBMxtD6c0hMs6qtitnvNcbp2DP4Rwwv588LuLMpXAJXKZlaTX73xx2qOPPalXQyGEUIv8UGNdw
e28GX3SJEW1vnFB+9u0mVg7ysYxNFQ33nqVR23jf5c8i0z/MTOQl0sOVzryFgXBQqleyiUOyIb8Z
0xBqQ9vaVx18CM8Roy14mJ1/PAhzDMyi0AGNTAomC/9OTHgAigY7mXGr3U46ymWB8hJyjXKj1Ou7
2s3M88FCx8Cud5uQXLEzYAUDrtsTuQMjJiKx1yM6qQeqEAIcEbBZylN2Z07efDAqqINXpRSjLqfO
LQyd72HsWPsdya7q61dqYjpia8Bp2Div4LDBjLjjI5rHQ+NzRDJ0pbXl9G+anHSsTMoZJ+8LLGPn
nMmujh/UpDtljZ3vFY2swR+KdJu909u185axPACv371JSpnwtrONdLe6f0jySpMe0cdyESuCLMka
CebZsVQnH6t2D4gDKoMpc4tSmbpzg9tPGqfaOyHTM/eKosDzqdF0JuVgLeyLHmZgPs7lO0II9v0Z
YUjMsTpP/V0LfvIxB4HSBnl9AQSyYh5ZuQnAKezblKAPU9CgKdnLd5QUBUHnvy9m9sBhoQspC5Ft
6oY4mSDjtgddoyV1wm0LSenmpXRtGetPoVNo+ZTMVka2ye6RbRk0A4uEcoOQIzVcFUDCwY4DmnMR
jyC1XHxj6GMsEoGg5kO04zP/iFoJLEkIjFPdDhsI5Keprv+064gjyXzOLjf+tu2v/ZmamcvKkSP9
0Hb8ImCm9DRrIgZ38O5egmzFwv91H831UCXsJcBx1WHRMfl34pURxA8HjLvuPxivOLCkG/APynUT
WTxcUIOhBfyVdnY46l6gO6Q4vhPRVbhrYw1TH/z4zGkGI8hDOmhM3nIajHmwPfL+wo4DMilPxV+d
Es08V6mOj7zvOst+kNQsz6B+NDIw5EkHukxyUW3VzPKkJEbPGSNTqq0oy2oxCV1DVtWV0Pfgbi49
o1RG8HVIctiRaEroh7jFkEoW+4H1sid0hPFmHt89gX4WKvsbefA/VsSI/y3TFKy8IaLbuqmp4TOi
Nw5QbyFNIJ/YZ32Qk0cEsO6C5Pg/sx+AGOncZ1Yl7wNnQcjbS52agpDMi6LkJGMj9l8AKmwRMkE2
iJS3Ymb5CtBtdo1y7T5lmxtv0sZHrMJMQTUbRmDIa81FW84u5kxPSpjRi9TJUY5Wg6hHFTrxt8RL
6LbIo0XL0H+zy1YrU1Rt0PcF3W6fz8i55vgifyh66Vw9P592q6zdxgmL00bSNcvIz9Vv05AxI5hC
6e33xvkGZdqnLg5OE32T2ZOAbxBfsLmtEmj2HFbRsAjcAE9yD3jY9vGqs7rU7a6y5Tq1JzXvPdbC
aY6SEXXE2bImACFj8vqo9aLstO9QrtibFu2vgMluPzwBrKS/Vs5240+93M3OC1MGvAtQm1kpbfR3
OFoyxv/997ixu0EssvjjypwaMclU07tv9xzh+R0hX12YzmCKlviEqJ8ImMvoAvc3UklPf2Y5OZzZ
ekWDAdqOXbcf+xADS0U63lw563l2YlIXq6+YDugRWAkupiGUta1qXpMfxWSxXSmrgqi2v0g6RhCz
JdpTpQZs7ac3XztkrhknY3pzEQdIqAaCFjPhSj1FJEciJ/uW/xZkPaUHzdhwBtHw+b/DKLxZMaGY
vP+vUaz9LF8SnpPVtiZr0MPXKSFi8q7iIes/uv7jzvJrbE9nZ2jRdf6bOKkvY+aWAWROzpKtIG52
3n5gJBQV8UidV1VM8cj1L6ksqOX5manXmypUFLd6pB+bFzdyN7b/tuFyIMQGmRMSOvPN8SBqxb1G
5c2V/JdRRUhkch3nMxOHOjYWQYXT51dZV5n2O62+W5LeDU1tuKh7ESOofgMn07SHWQvzoXlPfPFv
k9Mi7Gem/gORIppS/TdePDShztKlcH6oHJYpgz7x7TuEz1Ghu8/uiVyVqTXbYkv4C0UdiV2nRMgj
PUWlgStOpnbV74+JRg0jIEWw2Dh1ZGemOgtFWHWKS/hFIkCJfwkN+vxQNjRA+m2rx+K0VViDVeGu
NyJptQk619UYNLp8YAf1ggNND8eQow4B2AvjX9AsP/8r30Z0xDfQ/6TxkdD6Jm1fpD31LloLjoik
7Z/bORY5K3Gdt1RdENQUSHOEgAHvw/qCOc4i/Rq30Wm3zDk78dLLI8bPM5hx6j0UemdvMJTfx/xj
3v9AjXTlA6GBA4Vsf11Ygl6wxWDlru4eKaXXhq7RJnmlcssRwAVLvwSLR22GbY2UxASC663MX16X
5TELu+sotgqh1GDX3YaxhOkJ4tunH1qYq34VDoPWWEuc19vt9Q2C3I2kgPFOz07+7t1Bywul08Ns
6a8Q1O3Zcq1aCG0uSS4TgvxYWickktmq7YxaI03IYkGVhzU0HgPCh6n6LmScgkqrcKT5w5g/rAtR
i77xGJyEN1Nmm1ca8hA27o2u1O+phvFFor0XI7NT3XoHHbOM7zM053WNCjYMbvbyRx3TYq5rSoB3
UtYD/qiQCPww6CINgFaVjk/60vjVarrMybEAWfsb5v71uL1Ahoo7lmLGxzdgNMzYXMLVWNefXzsl
YzTBeEKbx08Kyl4h+2IBnNyr+8X+Ak9+Vb0q0uX7aT3hqzvHorqWSoBG4/TfLKLdjXWabGua9mT5
xUeQPb0v/vXxEVofro4zpTVpFtVoPhbIIJo8wc5dVcGRRddSVuaIJ2CRWZRfkifvsJH7m+g2Ve3w
17GXoRB4nYNkpd8a3W0SSfaCoJ+uXNgSmC5iThVyGQcaD/ATKafHF0XK1L3C94qn53AQICzyyQc/
B94AOu2jhLgK8iKJBPlon3ugofj1uLkdQEdhvKTE0IISMfDoabyep49ZY9Z2BOqOypEiQdYB/nYp
y2ZjYTArJLJKfcb41qB1CZrw4dqI8Kn4ERE9EOtvBJ7GNYL0I4zVmgatZFEGLGsle/VTRa1WrOEG
6VeCNptE4EPve25o9qqeeGjyvQ8GMPgn492mtRKm/KC83MYnaJW0pUbcRFutuYilA5iySqn8QVjd
RFSMS1m3AZBrAWaVVe4yYqXdmkn8hlwi3yuIw9+1gRd2hAbxkzx522iwBJnOGjnY74rjlF1FH3BB
8b0yT6a2DntBgCx43kFeGqRtbnlutvlJSCvUQkSBI2eHTTKU2GbkqzNarAcCOr2pdG8dl1QSb89d
FxgTCZz6xXQ8C6YzMg8kYEi33e16KVNZ7imh3bkVw/H8MiW+aM6aMdldAuvB8uHksVcmR9oO02hs
C6z2sKolkY6tuVpqvvAD9tJSr8GkZe0K5AYCvVH9q7cZgUw91SN1RU2ThZtXqEDpwZS+WGqfy0w3
7Da39ArdexJ2KsRr/ysvfIe/BGSEHhu6Lxd+fq4XSrUq++99hvyU3nGYYN3QpxAEs6F17xIRbNQb
VKtctMGgRh6gEGWJdY9rGt+Gt2YBrxAl42quQess4cVQg82KuBNXlUU2YcHz5a+G3GCFEoOR8TZT
Y6c7eLm/0hGl3apPHpunPQx8h0vkg8SpCyckFCr9GpgZtM6ZN3Sm8jnwe8IU3jPOqNAzH18k+Let
/jtTHTFFhvykNlk7R/enPYKv5roLwFBCoHTJm7olM7MaenVK+LyYXqulMECWB7jhYkVDm3mt7Qnm
WbcHyjaPhYP/jwgK5j6g/53CLKX5uwUWzHMTZ1yfIp54B0/T4kfBC+sh7P5CblaPhuWL2A0VkYQO
m4Ox57TRiLGhASPPDSkqwvyPxWyiZo10Kf80R5rhDR0l5uttPFPIAHMg8rBKJ6B4Q0hAYZvx4g3/
Gh7QZNHosCHtcU+RHZeGDJKwaNUsMEDdvecf3ywdTdMWN65xolnt85woDz1XjttwKUZBju7sJUH3
WoIn60Zb8DEouY+QaCu+2q6RWAHseFjrYcmZPHlg7VaoFYuiqLl9DewK3ZivX1fCeVKPKkxsdVL7
bgH7eM04URtX1j0VFcaVb/7b/YShpw+wMfZqO0Nn1EOlt0W4r/j0VGgfJcJh9YyLfTx2Dv+5BxJh
esCVh/UBNaRucarihQERgZ6IB6s2T/4eNG1Lv/7CSL9TMwLsLXc1LqZz4jbbWRVrzSqgtqsyQ2kS
X7UW6xaXLPIV3LivTDaOvv4QM93p2J8TTBOj+41j/EBksmrIuETq+JxW5fUkAjtWOiz0x+llkVgF
d31izQa8CEe3B2hELB0kSoyZ0SbKZqBW2KYFv8qnVV71L6b6zYavvrY7swGQCqZbZiFGwNy1Dfpe
AUUzgA/DCjxSMIWDVhfXkir5oOvbz8ehVixYSSBWdQAMzuwp5LEwz+RawIVIbrrm2dvYo38nel6V
MPJJcInrkxB5RpL1aXszHAz4+VffVkongNwAKR7wAwZH+ODmGk7JuawSQGfWNK2rWJAX9W3f1SEW
q8WA13pYgSMvO5GLrZrQBwiFQKFbvt+/fHECBPi1NtGE1u45kIg1q+IHzxsQyLkg1T2wXzJY0A9X
0VFQD0Bjuly4tbSjRXFJodlgplfACN8QduQzeObGhwvHiNnzoov6XFmKOOUIhrja+SuzaYugDJE5
lr0lxeW5qCqieDaAdoID/EMQuPCFulj06Kawa19GcEuab3LQuqL5zirqpG5MnlPrxFriU23lfAWO
0Kzj1n0zU/18z758lX+AwZtte/ZGFzsW9J9jHVAfqyGbj58tNItH7BFzjlNkAFcSv/RMxf+6x0CE
xucYJc6QhsFToJt+hyS7+T6MCsPdUVg6rZBpa17z4hf2X7Nl3wzT76dGEoFssjSh689UEEuGVa3r
LnoA7Nbr/SCeOtq3Sy/qRhsxgZyHjTsgCIQU2h/Evli5ulCS7A8GYTLSHJ//CK3pOHA0o99iIo8z
LMQ6cSTSzjWuo07MLXB+C0BOUhMDIyt/iqFvetXEr/VK+5qgh0PfKn76kdGRq+1+sYaz8ShvHqCm
opP61grv+YXOZ/mc6qnhF0rFAL4kPLMP91hobNWB8CrZCEZtGTNRBIBFDOn0gqZqOTuKjExwmA5M
yILFW6EOXBsuqOYLDrAW93Hxjnvxx/Q++wMuUtjbY02idqXNc6VJMTkmBOGYA/reVdneEOjtKpjd
XDSTz+foPeT4Ncg9ukJ/U45w/XQZ6DQWwOJqKwioA04vifZK2yMYsIqHc8XoLyhc6iTbNzR9oh0t
w7n1Rf3wwV+PiIobO9ZR4SkF3z+qi3fss93z1fwps2IGU1fK2Xvl2zan7I5cIdfKnTmMXp4vW0QT
S5ts2mRuBsJw/mkI5teRhN5ooK8psWyk5UiObbzj76eaYpRJzq6C9A9YQRV9B/1CYzbQaxL6K30J
5I0pcnCuHCLg/RwuNt9Lz40JICqSFLGsjW6nXeHtYlatuRu2zGLgIj15sSj/nKQAIld3eevwdEx7
tUpSdIDJViMD3MNbkrK8MGtqQ0vuLlTu71mu4RrZ93Wgk4No7d8lv5Tn76LyFSUpJypLrQrIGghJ
OlmEXTvtTcWja293BsqT+/TkVxS/Ssm8ZhXqgGyBeBQtA2TmLC9rq8Fg8xrnrYjCDXRIiK3fX8cD
NIt83RX6q9IMjvjtGPOqVVAqsZklxJ3k0to81ZxA2grBWOQ5Lf7Y5Q65UisDO3uKk6G/7CC/y9AZ
KjS3ehCe2z1pyo4yP1O1CQV6O9z7PVnE6cnxKEuflI1eJ1qZ0A0VltCYBzsrXNNpn1McV2kVnv8q
qmRZxJjCaP1wbjNlQQT/V/fsYBzoxTZBZzs7EqQKYXRHAtHeDqvxoSzwdp6Vhp6GlF4mo6K042lV
zQlXvfghrT8m9JbNcM4cSG7EYh8pam36H2zVO7BLwxLJDY/S/gdtFZX0TQRW4IoQOTY5GWNFQO95
K4jU42TUDoySMR78kHajnWAf6VFAlv2i81VNiTrtv5TnDLm4nQsu4RoPlXjNiR5FJbUNjLp02ohj
EKJTpCHAh9Crf6WxmB/pxCtd4w83fgfR0NxYBkMTapxWyRa/kZM7FgenJcMDW274ndBrVPR30pdh
iJSdxF2W6FTiGAUJhzaILzD4HMOTsCRQnsdLx9HCpfnXsAOV5BedZv1yemk/LJBS8lPmRNCxutXn
/wBNQQ7rv4wHgK0TqmB6gMeudoYBCavwwsbKnIAiz28/49ro+DJ7uqGGBwYVsQu92gxeT6E2Kquk
E8sY7ZkTFSwooE1g6p0660VTdAIyrB3Od+aoko9ayUgKE6uf/CeJGsN+86Qnnwra3tdj1Vj9Pluh
WUhNbcAtBR8UKyr7Zwhz6CK7XZ9bakYgdZq+A8NZCtxY1pH3C4/a0EWocNTOlu5YP+uihfMANeSN
tAyeIemSG0Qkj7NKssYuuPcsECkdsyZa0L4HnQJbC7WkZImhbAQdIc9X7WHUFrYI9A7uZY/aWUWu
jnxx8F4c/wOK2y7FOwbx67TmzxpIau2c/YtISF132jHsiBFirL8vNcQln0ohxYhVmEFe+qd7j1tm
AjOQ6LSKzLlwxHmMbTt8OKS0YCfX3xnvO6tXI4RPMgTZ36KzBGBQ3R9HRsPkm7Hpsc+nDY3OTIwN
gCrF3pmUJMQnZdQX+5lbz0pOSLMtDjw7zyOFMtl0+wHr1UXuUGJmUQV5OSjlLqpi2jwPpNkmrncE
KUqArsBQA7jAZglNU3nvoHdyId1DG+D6sfh6KA27gIsAIDCwF0I1moTbUsGBi/F2cm66RW7Tmiph
gJP2ai1BL3GywMUkuVe7kV/JPQlk2OjyiEvHzkjVbWMBFVUahVUqKKxRpg2t4MRHFHGRnuvKvCj5
kECsDZFY3IPazUSeUrbXbkr8ME8RPdmvy1eSMtLZizLZRMlVlLx3zRG2Wr8yw6J3aB0MQLs1uGG9
X4N7UORo1jYSw5I9swDuUV/ghkGqwJ+spv1TlZJX3vswWdw02HoIeW1VQgs079RtIK1eTO9qNqwA
3jJdiN/fcCPzsB0eqT2MAqNnUuy+IN1I1KSYIHlNA2H8Fq0RBr8hd0CgpD0zqK/zDDuWB94Z4GWy
UotRD2tZq9zB6CghSUizMJCGzsxxzzfqC7hyB4RJdWL8jl2Q2riyV8bGJVHJptYEJ0yQZxiwrkN1
ELkNdN8L6vJDuXR+2UwKmXhLPeI8oL8Ur5ml8HPWv1A9Ow3TqlfbLPnA5+dLgq3JFcrKRYpnWZgU
5QyB3cZmqZHsyikZcXLuADbOfRS5bFE1QROLVdcurzni9p3mtzLWm1gPnm9L2sldUchOyyqlf08+
FP67xodCRx6+uDxEx/pzeZgAo9XQsJHvUQdes8QgPanfHm2LQFjpyqBZI1rGATwlaP/H1UlFEafV
aXR8OSOw5m3UbG/8GUQ+GTEIKk4QD+TTALtIg1LTYsgG/2wftyKk92WJMoMPGQQCigyqiSWrIom+
FdwqAHXrn1zMwj8mL15b1utQd2amBEX7AlPTJvFIpR/o3O73R2gfc7wSm8yMEObDtGNiBhfTWzaI
QTIKXK7QF3qBRTv2LOqx1M70eBrVwN39iJuxr/xviaH7VP8frEEYESxKn93vSrKv+m7U+q5JIAtk
fyM5sWmY+yYId9a2k6mUuy4WFayJ2Wn4wHabU0rJEBPThDwxoVHD8HElI3bRAZBwjfYN5gjROV+M
VHSWVIuGXovdODOi7FaiwWGOXoopNOjT62Q6Y8TeVgosQ8DwFzAxchE4kMsXn+z21HrTZcPlC6vb
aDqvskIuv61h/9jCetNjzJO+yUFvxeTHlEnNdteydDdLp5wpXYQbw4ilzzSZaB8Ky0LBM2EgNhin
S9aIHR7T157x4a15RN8uqHESYqL9uuRiTi7yS3D5ajYxgWEKY05/A7vM1BZxEzX8JA+IhlTXUW9m
45UllAK37xx0oE7tFw1K77RdrCrbh3B+VD9pgF6H2JMfZVDCPaM2Jv09CFo1YwXs8tAJRc6u55JE
QM6BErdLUVahjkmTqr/miVKZnjRVtCR0kzny/TQw/FkgPeudXyC0X9RDYSJAza/OiY1VUIteEDSE
XlzVj/MM8JvCgZ2kTmSUXC5S+JHWLqFNy2p4fB3/gGNiJCqQ2Zyh+l199NlE8S2D76i/JYVhbXq4
M7YXEUDkugF2QXx2WnuOtSvSqZvl5Nq3/aTAFLd1HVf3ZLUKdeenFfNkaeVH7ieWiROVrU0MJJ2Q
ilKOMjaFjthDARNSOAxwJXt5q0ZADP37MbeL/YQTjffVSFfC1+M3HdnK4OtVuPxN0baJPWmCLyHu
0RHynbaExEA4k92QUq0hrbHF+bIYcmj9Q35xkQkRP5QjzNzK1Y/PAv/xGqZxaLy4w0YXTVEu+SKI
JPNTNb42G7MIi/B6XU3u/nxAB26qn+6m124U9puPhBz8H+X6oWC+8a3Dm27ZB0V8700TpiiVb+eA
BgryGR8ZnmTILy8458gETiBadgOsTBmdAwfQYKMrrx5WClf1ixxALBkoUDzDvNsi7a2Lt7jwKFrO
KTGVtb93aooNI+olAZSrJaiGzTRQJgbWkrCThnWgfL+pdhanpAKAVLKgGglk8I7qEV8k+8wCFVD6
OmpaREf/fAqPi+HcIgLR7R+c6hdZQWkjGP7j2qHSujPu9ZsqMxoEgEt+VsIJXaQ/JLT9/QZBm/MX
cyi2CR3H/vo+3g0kxKx7hcYkryKg65o/+8k10brpbX12zQlt2ojdunTI44U5bTgfBpBmKktlradS
QYdJbm3gP0Uvh/FPTK+QgLh4AArdCYS6DSDIMyYQ/f6IMXvS08IWUBFhnrca7dJ5sK2ZzlGQfrD6
YdVLNVBe0kdwpEkQBUW9YwPbfZuGxM3LuUF371fkszUZlVta4WNzt4BB23Qpv5KUDcWj0nL4ZdK2
ijaUBONLsYX2daVfpeW5Y4ZOvgD53UJO7Ndvx7L6UusvsMrOvIaO+32R0oBSl4DmzJCdkXU88avN
y1PN1DY06tKyHpI3kDNzk8ZG+Z3SVQDDqErdz3j3IKg9scDKPmDVHYNqS668xqdut1JfRljBwVTj
96VxZZ7DxdUtfMeYATIAJxXNtyGlZSPzjIXsxjemJZHO/eRa1j05jhi2F96jn0PP/swnf/khhVuK
MwzlmKS9VtzBbRt/lVm13OJODFAGXvxkv3LfHtiyBffa8tTveSYAWWz45wKGHtZL93JPXoxFbfOG
BB4GSFuI2Ll5bvfQ9wqOq31fRgEMxZ8QPkNeS6Vm+7/7UAXkxtSVB6U7rIImMkpe6T1eCxLPemNF
qclfg5WPZIF+ZvqUKXG6Fg54DgpyvquaRnIhEl1wk1QKYZx+kuXqKL2Ow0lYj52NuxVja8nKBMQQ
cldn2gZmkoFl5PkcLvrPmkLo7QmTiID+EBpDBPOCIYMQR3aY7iXc1ib78/5h6xymVLpCtTq5sC1j
o+ZahZfyLhn+Kj91lwJEqlMazI2ckBDF6mCc6j3/RWO6jAXES00MqjbtLFiFPJi+NM6I9R/rTL/C
IulFIw8lDYDPXVuoMCuI5jNuE/uQn8wN7azr8cv06LkXX0I4iMCrPnhU2+ekDRMnAWSPWB479LHd
Jqu5TOegS04n8+9nnYAkBFgCWRf6DHGSMBkejPrI1UBHpmnUP1DHrkTI+ZbguxBc43ZXawtA5buM
9GdGhX5MECnXd1r6ChjNQEMzNEg1mTZQsMskbnMwY/1rLJUHF+oTMXr5Jkh0qGEv8mDwoZLU5A3F
zOzadY61ilZI4Cw3kDzZXAkhDIrXQO2SDwj0VPEK1VC8I225yNjneVffREX4PhNvfXetg5M5vDgF
gjjvBvNgrlxCSWhyjwPfU+XX0tgqOtxtVC9WUGyCxak7D3bkwxAyLrBRurw5XW5hA3+Bd6iFUNHN
3zQoq7abgqm3dk2DzqFTr9kcVGwLgW9u50OZss+pfGeyj+KxNxN59cMhgZbLHbM3UVCVEzLcYXWg
203ug/N90dcQ0RZqNJRPINhZfCkX3YifSFxhu6RCRzJ95+v0IZMDMvOu8FBeN+eCEaCNLPRMZqs9
7vdJJsavWFdrzULza7kGHZtiwFecN7Qb8Rtvhm9lFLQ64qMqzGN48iiuNmjGL9uNCPGRKiaRPBU5
oQKb7C6paEkiE6bA8SD8l8+rhP/0Ihdsjs2bUwJpmSfdOJu4y+d+7T37iCHudxboIeKAUQqBUoLT
fdL+kxvRZ1Yv650b9AhvMCB9E4HKLucnUVhKL3Ftb7K731BNtrHNnwhvSUKcgiKN8sRHpZCGhRbx
piC0fjHUbNpc41iXj7o1KwMPwEomK8d//J6JfhETy1GjBxFMbiYmXMlCfVk2S/D9HqAgZdYGNZR5
MOJnMl7MdCik3U8kX0iRuWvaUAVRxEr1ITiREZQkopOoBptro/gXhr+Yam1NuaVnvDjH8m9H5SLQ
oIZlJDEOkX2lomaYx8XDfdKqtrXQayDR0rSlYbY+pMqSTJCGu/ce+A+Jn/Qvev4ozsNoXHPNDjK9
vrUU5zvUupv7OyHD8i70mGvqFd/tlQWmGeZCnSpsemGnH4YA91gVASsfVhJGgyV7Kj5uilR1g0x3
RzLpEqFtBPcpZpqHZqUPsl4O0sbeDs5tWOiHOsnuheKLW7vYbVso+aHuCRedKLvxOZqb4ZX9ZdG6
b61oMm/HgnkP6R1J6Y66KGysigEFc4b94lY+IEbTE/ypMZ2a7JdQOFdIL2MmDzdpmCh9hy6NQgka
PsAyXVfQY76f84vxMz2dOdKYQotFDdonvRG7dkQ7qMwl9+cf29vMAGQsfpbNFgA4U3CQBTJh2VE2
IFA25YSaGxFJVO5+VbcRftOqdj0QWldCjOttzJifwzB01+NU9PgJSRY6JOn8++b2PmvSNRuYJ3s6
cbSn4e8RSaFcVT1SeWT3dDd74ptvrMFDvMYx9EAA/0FiZ04ou2jG9hAKecsRC5uC6urdJa2WVXeT
LgnpSL9owa1N11y1MV9VAa0lBRQR26WLOM+WNcxPjGt3X8BIQZaLYVrTAOzOto9r5xSTE/tj3JZZ
ig1FGA/h5XYP7/4VOIV5TRLjXTO5Ku8tY6Ak7CiIrPvnVmoh4Sx0PnUphOJovq1Gu5CrNsH1/Smu
FrOJFtFntiH/1uFZ2wk8MCTqY6/Y425MKk2Kafgs+WnMJ7sTHLJrle0qx9IYzRRuGl/1lyQO/nLA
g1yTAqJP8ZHyuV1Ir4eJedsYfhxZZoTh28Ue7bM26kvDIRH8IciZqEdsniERwLl0ET91PqDznCjN
Oh6LW/fhmKshwjniTqSWofvqCti6LmlFaBZCnG1amIHcWmXq2TGG5mfBK1akAc64Qe4Rk2SPbjHm
MHFOQ/GncIiTFeN0tZsP2EW3bUxS2kAW+/hniAf46W/s/jWXDGcsoOeko3dEVW2Lz9BVZOQ8fGO0
v64C3HPj394/ocGYwLdsAr/XVEWtoBPJQ6JbHwqtpPgam0mAxQ7tRGWoiDcILt8qrFEP2FnA2LSY
KcwO4PJJT/bY3ubLq/U8/wy/cpCd0jSLidjikMO3jRaJo97YjYY3Uy6L92eNu/wXZkuDrXGSjHh3
ccLaqwG7hqN6sxTh/1BE43BOtK4crtT0SZnVRP8Zrefk4zQywbeykDj/OwmlZa+aQEMZxT9ykZtj
hyNsxU/Yk8wyfBItFTKaSuEMBggUTMxxNqMC92m5Yt/GoCreQGGpoy/5OW5V36LPQ+ZuDDe4AYKP
AdRIl1g54JX4peVxd+Ox2u+eI7IHJl/BUrUr6KEmvHyMZByWx0biKTSPTPqi8Mn9v5QU+s8Lzf+z
SaptGJuv82qQb2BIICSpGYTBfJSPgROmPyk6fLVZfBCYdtnp9UqA8KOsehEFsl8RGQlGYL0l2nb2
nCukk4iWl9EjAd0rzBTszFQyli0ScFg/9y2ns+ikIpoIdCA4KIN2QuTSw6GF5xhg1IARotNraZTD
MHVGnd7Stz8eLh7+MQjhNvOVK3lVZHvG56GMPDG6cfwap4//gObIBiUD6qoio4FaaBOpVj7S107I
5AZee/qeBYZL4O2UMNiJZdHSYtNq9Mpnt4m+jNcAJetWWD0yGhW3FCygffoYyrshApJhABZGlhBn
9ha8N804ZHMipe/ZqKbmZhR8FuUc96W0NufD4aSRPFJ6lxJZeDuheimKOIGycEWmYnJfhWQflH5O
kS3oyqRyzXf15S/pQ4Uwh7TzH2b8tO7urSc9/6ypPfioFVHX1zAQSMnBQD9XlkJDX9Cfip2WJI2F
MNu4yhThUw7gxHnKVHedoevUZKaKbsQuKk3lNp69adCCuwqEUR5Xqp9K2BjLyJFAttZJ4q2W2r8x
/HySIL48PZtbEwRbMKRbC6NSHjTveKoRIgWLsF54uvuyEWRrXpdUUtKsCvtAiY/JeaO7C3btbd50
CXTN0adN5eAbsPMGJqJeEQqyPV/6sby42NAFLXPnezH+GU0AyKdF6hJd3XGxp1ifPjwFDBsT1fVt
slGYpuFU+419lVKwv2fbBlla1oUfbKEZruixd9OdZtkWk9Fu8vpZT4LL3ILSq2tUiJ3PnjQRcDVv
LasiVgAUBFDPYAk3KCrEDkkej7Cc1q/wApqbnJzL17cD7yawCQTudNn+a3PZQ/1QS5so7Opyz6XX
18hCBUPyj9fKNoiZv/tsZwxfMjSDq8uPNnPOrwaKyxqGvlUJinIR+Qd8rGoiy9uM5dNb2N/Kg5uI
KdW9dC67V4akP4rJHJNRFpHap5SLOr7MUuDWrqb0Ov/5dx9aT43RXVgYVBUvY9hfBoUibnL+CucX
TdqvLaOpnie9wsrKV4bpMCyN58zFDeToNKRM2dR9dqcurzRYq7yDjlLPwQe90HOcdgArEp5aDfc9
uTodXfPq6VnIpnsnGkKuGLpGQGbVIi84AGVwODda+rGDIfkD3Ph/UuqryoPfeSHdYg11JaK4r4Yo
vJx3OnUJPWz2AgjMfGCBAanQytzPd9Wy/aW1AM0dsiwMxzBEw/fH/Ea04oEb8Iw/Ys71aMEacdt3
O3BL5VEydgp7O2WpYBEdSPbTX61GXKWNvFiUSYFZimyQdu2rtDQdmU309coVnLnYBo07FeUo/SLU
HbvXu9DBw37xMcnMkYUWCY6sBy4MYT2eD3z06IKUb+cysb9SXWPFLebUXy24Y77p4nF6B1wpSDIu
A+C7spzRjDHcRyct1USNNzeLzGKAdzWjo9r+ckwg7xCJS9UDVuaczIi1VxRGGxDAAOnTSRVYT/gc
5gPAtldW4g4G0mdCgHBwKoHN8LBn35IBnB9CXEwTUADD8huQTIRs5CjYSfLcFW7BgwhdM/Pgp0CU
Kx4h9b3jB7mAeV9fiZtMN1L39I/32LqrZ1OKctGHUzChIBFtAhRjaEcdPHUSYLcS/rPYhtzYNfP6
wuZXqCFuZdavuo8EqhsL1MfXtMzAWMPv0IiArk85m44ofhpN9L7HP5W3C/D8naohktwk1fKDproB
cVsHuESk8b8x5wrdGHhKfjiHJGv+U6sRRRxx5N/vp0LQ6QD6h78f/plxPpSRMb0qk0PNcToo+IcM
OIq1dlDcL3FoFd4gJfei/gLBt7OMcI5HodUiYf6hH9AsLRw8+GiBH3dMj8v91hAUkKvVt/egR+oc
HaiiI8Ty6o0wnTb2hNHXxAHMtj+cMZ/arxQHve6mfDjHsisoNkvCs+nQMS3sTKYxrE5Qlp5SIA0o
U7d3UFXMG2W4MduEsb9ymOash6CRpHKbCO5VoLkQUJU1pAszABZTPy55a0nwp510HrFX1IXWcPNY
Y6BzsdESb1Bz1RRVcq5QEy4dmiHssTr3qAdWOVlhRwEOyxfwqCW82Hpq1WzXWhqSP62hNTVVIRn6
tzqo4mXvrWjwKEmR4qgave7FInGKmRoraL0Ff9rw4hVBW5REeRQzOofRcFOKYRD9ozuWmmQvMPM1
zanD6S7PpLKSQGhc0F45ir+M8Ahns7qpI1hk0GM/tFo11SsVEUJEvi1Tbnczrq/pFxCI6pAmUmlf
+J7C33Pa0FkOjbkn2YAiQNX1cR2bQPsHQFvLUCuMnuPmuKgwImlQYM5Crwx4TOgYakh7PGMxppSB
gUImzD12jxySzsZFUNUlm6XPi4us4qJNdYm3DQJ1ifCzWYY613/1EavA18k9/bgFqT8psOYJ5sSC
OjQi5TVBvZeTwwX2zhMlWAczVQcDsvVpeegYWWF6hzha9qlgkuFyUIfJAqbSGwyjUodM6UKZGPtB
/TzK8b9ch058ZhXvlsxP8GsSNcVVfPGFDT+pJWFjUHi7jzVZaoD0wfLqfLksDuyjpmpqeFDLs/46
B0vQZzYuJT6fkhP0odTc/Z0ml7ExreB/epCzAXBp1MTs6IcpeMlVE3DLTs6KDsxQEAGQml/Js0x1
pcjYRJX2YAYrbv610px2wskyW5fY33ZzhSBBZ739VYHMwglKJ0a2jhh9zl1wWwqsVEKD0eXYNlQS
Puv7FrZnzY5Pt6tHzC5bouHa856IGcMjQSGuAeP6b4/3QzSDErZWozr6Pf+t3EDVVPa/6Lhq/Uxm
tMSzeRkaHgDihXdfyLNCqaXSM1++rMVQp7K9oBq1RARhf+90fdUg+x8n50k3JsPvnlOwCmxXzGto
l2+IHVzF5KorJCq71G3OCd44YFJx3d4lWW44wIstI7dYfKUO0tWZNsUCm7WFccItSHWO4k8Hb1qx
8/A18uVYncP/cJ5z2qjSNcli1B87/8wvzkBFF7lvLnrRo8wA1tppwmohbAvFLsJCepH0sRGdT0dn
7vFP7k4blakH0dcZfcse4THJJ7sVqm1DFRwIL/b5PC0WprmYAApqE7RRAVN84eKxpi68PIfWLx2H
Uui38orpnFGkk5dVrSN2nm69jl9NkjtvYNX4v/3hr3OAHLh804PUqGX0CgSXSFybUDcgrTF7ndFz
jdPXJ2uKzbCHJhSIVUWPF9e23em4y2B6zzqR6xZdH1p7LgDyDNQkJIrjSA4r6cSfvqIJAJ1fm9Ff
d2EatXRREnUA3H/5PR6lcVLTq8otiq3ALbsgM5cGtpWnAcwDLoQTU6M9MnvzAQJCmJjT3k6ZVKVS
K2mnZeXH3K2qt5d22Y88Jz1bcAz+JxSWhmn7uAGuwHCCaAg4iOnzuEmRg8CiTHOSQIcAfbdJ2bqn
MNsjYa2DqlS1+FQWETM5vezJeJqwTuOQAX9nZahSwC5U485dlqHpviJns+0cOrCXhCrelNRtixvD
ZNxiuD+jZez4bnCIu29jZ7sZ4aUua/Ycd1/18txNIyJiBe3ONLtQ427Ind0NUdeH63DxNZ2xx1DJ
yxH15DAKoTwwMXANEdbvQhmuwaYuW2avrdnt8wXfZauu2fNiPipu+oZ9w9TGGFARVDzg3JAfdq9P
Jqw9jNyRgURfA7xXZKKQKo18cdwnrHHjRhRb1f1Bu1ZKCI/JqlTqN4ZYXF85rjjNue6ql1PJQ7Cr
we2w4yLOS+t7/xzx72K6+gS3vJXO0cC7GRITy/rYX6X+kVkK+kYnArEIaa9m6EOovsfqSF6Z0Ipc
YeP1qciW35DebOq+77IJMGpptLVEgLUcBrae6yM6QSjEzoveISYZwTpy2CXkKR2aP55rwx7Hb1z5
jqPf8s9CNC+0rLdbVqj/UmQgENYw8XZ7/HfOYtOKKXuIiqE187RH+Btcwv8uf66cBXVvl90ELAjI
zypjl5lEUqzfaVvMRzq8aQCQ7GD2riDuFPViQ+QHwCk4KALVU3kz1cagdrRaOVNrDKTVYpJl9j0Y
asu5WLITNjitLOhEc/VM549l8clk82VetGU9l4ujSWlkgOO3sOp/VnByQGVVXgB2UQjJG9QMXccr
xDSAwXAKLVu85kGGKHgAufKaXuwo4MCJsTEVR5QhK3RjwLpcjeGZcluPyJnyPAQZbEwKxrO10UVy
UVUr3D9zBViTtdzCzT4ZMozSfF4N30PHn+A3FkfLLXz6UxWghaj0ASWDTPEq8j+mART0irfShOO/
BMspKRYTz1wPV9jKSgYOMhb8b9kRg2JmrZL18q85+frYn5DflVKulOqj/B1uLjigzjLRncHBqm9o
K6/OXqfxv1TD6qaWBBM0vvK+8j3GhaKNo8RDQb90G8wfC6UXX8WHFELZZs5lq5Dd53pH+UAZA+mM
4HNq12ncHTtmNX2oLI/QK12naArXnwXhDzheVb0osXZf5FItl0EE5of7acELv0WDTXYwKiWNFlDV
MuGWjP66OrswaM5BXUDFYrAW/L+7yVRXi6dz/S4FK+VTxFY5RtyqxE3OEapOXvr1eOWTFhzdIezT
egM3dpq32HH/3+ryySDz030FyMe5pGtQooD2GQeH3l5Yz24ZRiOfCh07qEm4ugW93CVWmzalTb9q
lhCp48FS3Nhua9cGOKlP6aCV6DMwdZjIWtQxfOMKzC/HLojAy4wqrfd/0T8pyzp8IDruU0AEkMsu
QiYWhUu9ErVrFKRBrTRjI5Pmq6JYIycTZ25jptGzlgi0cFGbCpZuQ2PXTkZTmEAX6YSaI3WpS/RJ
nREGuEqkN7tmqbVh8FTd9xk7LgzIW1ASxtWVcyRwVpdpYEXplVADygA2TCTesOw968FxArkc19pq
InZTihBFpNQeaR8RFUA3nux10o9O/scBToOQDMI/jBP4CT0oXVjf7rXMrsI2JwMUvUZAL5Lqp46u
bpB6RrmQ2SCOY8DV7jzYyRzAqf0f/8lSbipNavmyOq5qVRVlqqcd3qyKzbjP7Mvgod0nsa+gC+vH
zs1omH6FSZTV4LKQ4rWml+SYJl9odDjCs0aSGJJ+ny0kYuuvcQsda00f619imc7LctFdZK/JuqkP
RnTo3gjYSX53UGYRpGb2EaP5hXlhUZvbPlaVn/BPwjdKMC5SgFFMf4HWF/kCwovesUYW4Jcljylx
oE39/RaYv3D0EN9QPoLCiQk4VNHT9Wd0mbfcdfQTlWBbL7i4pUBJ2nDnNOLdgAtAUH+FsbP/P8kP
1DhLEFYHaH7utWxmg/47SpYqwQW2uSCWaKwoA1dpPk4uaIqeosHmuSoqe2/Ia+U3nOTV9snbG70/
o1ujwXExRCsCOq142sKuVr5xwxgkpuprvxGKKCpVjhSWQSWEal1jZbzYuV83s29db0+bZ4Qf6/8q
1orYXyi2NoAlSvkad4kzcomOJrBfkoXbCgt/upyptd8n6wGKk9GA7rgGrbS9NFx0Fdai0+5S/sud
u2Si7p73a4ws8C4nw8dcbZHI3v24wc8j1CpDhgj4rmLgekvOmEwhBHp2UTwN/SmmuI5e9YyCDZGq
2tTRCUHwQQgrToImjQ9voXa21DIKlU+3iOj+S/RThw9UVKD+ijD374w3QUEJICQjOnAi802jR3Ib
gCgYVqLg93fzp51eAZWUEn/Rj4iunVl9/f6TqfwygPrzOmJdFqkbj56R3xmAD3oNISgTP8u3ncoL
IsgYfTvrc4IoPJlF5ki/qz4dnHlM6OSMuhMEPvLm0R8eXew+1M+1QNjgEqux1ZjkOuy9qxguNHuP
A+tuQdQKKAff3W8AJTgYUaCLL+kJzqxcqoqGmO2tFHShpVWwk7spC6IHZsV8ii5CXIaPCHr3bez0
8iFduNuzX/ptVtFrkyBRjv4SpKV3D9SbfMVxnEJaW7u3eXSxqOnRwssG7sthsvCKGG8lh9F6bTwN
+ociJEjzabdnHUf8TJZbm+DG/hTb0/zP/OOmqlgvYx7l6eyZcmvksfigEVLuIzXO1puGrReWBdH0
YrzPLvq1REZJYB6hhBxVkEcdvERmTjXY2zRlKb4sQzKjOAskxGrGnWdQEbC1cJ5UmTy4kSTlPqHl
bAqquRQdVN8/VbGz+JOTObh0sFs3Jb21qiTio9YBU6T6/3IUEIKJvISWRRJyvJtNgDBD7ZkuS04V
676trRb/yiC9AW8GWRKowg4uMCHx3BCpoybjjP4XPyjhSdU1UoAPInY2HxihOfaBmZABcl7HWyd2
kx0vbwUp3B0M53/40ArmdorwbFR5TWplORUzwlx/BnSyoecOP5UBEbf8PC/VpYK9l7wD1NmIaG5x
MThBWM2S+tJtEHAU3Bi9XqDYcHi8YqmInDnDFb3QnK4M/0OX2o98Jl2FeLOdaBOe8dhlxUJy8iCq
bum7J3cCxTpaiU1i2bC8fw4RdRQPpVNeIWzhYjhmkAl093wfQZ6UVYkpFvygVgo80ZyOlwLYfo1U
G8304bcBoEfFalUJc04gyTK7aSC/NzVykG2B2wWwwS5sbDEOxt9IuBJX7prHiDIu1pN7aYQlhNrF
QnSG6JT0saqDMwbd5iaibIVMGYzHcU2seSleVoE/mWq9ASHfCbaV0Ur6WkoXP40cWhKjqnGN0B1a
KPIcHY3Z9L9trCRd/iQdm5lOHnMNIGW1tUGyzLKoh2PuSn8YTiu0kGqQHYAYstdc5WGD+fEIXhOM
u7ZH3grh6OXNtP7hdMkYlBZrPhT7Y12Toglx07TAMr/hrzjhXxLVO8wHB8RJZiGKS8qu2NJMO4Wd
P+duE6Swhm6HRCSnUr6ndtXbgY00csSihtpXfrsiDsqLG2ciAlISakNZeDSn3ac7S8zYX9hz1mS0
QWu8Za8W17c8suJ5KaYh/E855Yanxl/v2JSqXn/HrBD0xa5kUN8quFdCbkslJaJGAUebrBM81ktW
ukDCNgbQGDggGIp932FxuU30Ig7GXvHfv4NRZmaDTVGQZfqAMXEX2811yT6wUf5BRuqrwRLuMJXo
2iREuDm7MDgSm7l/qrNNlMluPUxLDOnKKwtsUg5/OQa5A8nXmJGvBlsyTBfzzgl74b8YRpTiVFVf
yOpI7q+dahV6wfNy6csbJdI7Kku/Z55NK2S2hFlmqMf8mvtj1J6tArL3dvGZ547jZenSmr6olYh0
3zznJiLSkPCNp3Gsi/to764VNUUO11jfbnVvBEbGrYdMk/YK+3IFcioEGwBIftbq1Xmx0/gNSIZ5
FDfG081gVZrJCO0bNlfGR081peyyE16Hk93//ooHsjU4qNdA+DK9cqp8B+GlGae1Me8kwBjgvqZy
LI3CIMt06sQtK56FzZrt63A+jdnSuY1uGS53QKtJwEOZFAU1WEW2l4dduvh7x3rUkSZ1vajVY4Jd
hog2qZUZzcGUAqQ3jrHT6oaWvxLcqbYY4Gw7sVc48I78ppUiUi6JFpXz1suumGJxue/K0+vCQEub
xz7Z7EDvyq5d31ZHMg8+pnnWQ+DhOD2j8bgYkxSOK6ucnDc8sgD3Rpte7naAoSpm9VX/GIgG1Pb3
XnXRpwB1dff3qm9xWRuapazF0XHnap1YGcDqicyCWpA6PUpwMUYsMI+3osFwK92cocQW5+5VYcxb
N+fy0EPXK7A5hzoa2GI3o7crcotg7+U+mysRVv45jvJgvFHTU/3Hr2xBu18ER4PAMT1xX2O3RomV
da3OLO2Y0WtiarsULzPGMpPM4T7Rg2E/0Unyf4Rtk2pHpPTdMYH1xBdIz0+eFaWajxYL4X9iQZvq
J6QzwMhr/6Ig0AMVTHSf99iKY40QSuLOLKgnmTFB7/QNtHKmBK/aRYJpRpNBxgpLAY3dLtVqzVfm
lvenMNkW9eaeqlcZAgWYSBboyPPYInui1AqmtNTR6GDkpnaAGxGByfxPWDGeWpVV5gCLRUXrus7g
DOg5/sO1cbXur1VujptukXmwWX+kPihWIGUo7Y/u+fKGyFo1qVij8YpGZEUBuXtJyqpRivHMNaWV
FMSMqh7Le1KIHUc9snMmmCkEwTofD/fVQa9MDOYJIoSv23lNk/cYEIa4UMD8RSw+gMszlPz/Eojc
f7VnSyJBuJV2eUK76B6iNgaXGCiY4nPexEEpaE+bwARa9aq2eEPV4RL2H6MOsm/2NwSN2TBVy/V9
mWX14d9wNevxN0Wm7i1ULrV0YLOBbIVWWmgz50oQxh1lBpv3clcWA2XMecSaoOt9/j0BS8z+ZGEY
P0HriC7pPDj56edrQ8wd5tCoBZOCmPLSSwfJsXjee6WVf8fXqIVuDmg90lFAAi3q0OVk0lBLa5CU
uq7gw9Delz5vWmXGUBAUkPim5M4y9zTa8D+NlC0OxFMUnaE3cqJ43Opxdk0eZoai1o037f2AOx9E
mKFpvRezLKhvvtcM+NyvIwwhkvu63j0dNjHjcBQpHKvwzEmjJp2ABOdpFq0EH2i5VriGC4AQ9ywq
3Mm6xMuxeqqmXyslkFz+dSq0LfRxXz0N6RQNE54gjpxbCJUgPtb7PMnXGO5NQFWMIMuZ5+h6koxb
e1QvbPDld+GDmEwSXAxEf+ofG+5P7ZQ+RiwIKChpycLxmgq1x+PydDjDl+k7yqWpkjbXk5zJg4WS
Sxb3Jxwz4v1YU+eYWhM5VyDObxOseHLk2ifZ8fBuDauKDUEyvuVLRBJR7EpzDXR/4P1UbC3xhdNU
JDWGYnQcAtsMJBR5kiWgMhpb2r4S+kbisWz5d3ShRNk/ljCSwgQwyVfvwoS1qicpxJ2kirfexr/E
2XrUu0ytSFi+OBZ9kK/yhRYAF8d4gF7FzzKrNfvXesok4xVKOZld9haZLF+AV+ikGlVBZ4v2uXGC
HFhZJYx2wf99WaHeQzdkJ97pDXgzOOxmvsa4qGHDwP3Wkwi2iiQnn8LLJBbChaICaI8U0eifkg+Y
RaODmOgGMpfD4KEr6yREb3z38p2Eqi1FhnyKZ12ElngZeHcBNce75/9H/inDBII9leR18ZGkaG6j
CM3WApZbTI2CX+RN1RJsmRGKeVHPEe7X1G7P/VmcTj4xbuE14HEi76sRsua3Z4j2bTQDWrS3I7ki
Ti464qsRELySeHmyjxsjT2jr6PwTfEDBvLUIu8QvdiggbYrqiXVp4PlvbeWMrVXMC4h9zAfoGcoD
BSlX5euKHVmuN0Hou4DOmE3dYtKCGoHH2fmIq7ztV4QyGmFAkYTYKqzsblVZyK5e6Qlt6s8YatpP
2NVEit04SrERdgtBCvKl4Vph6HV5rDzkjvb4fsKqvClxcAeS8jrEUPM3D8UxrJTUYX/tzel4JGat
c11I7UUV4Y/hr+th2u4bHtl0a6QmXMabK+T7eTky+uLkzfDHTNu52mlY7UU/y9CXoWNkHYloHnlU
/3I9XViACXZxs2f8NSlrFZlyKJXM13JEvw5dWB77mIcqyuUzMCXUSRMsspw40rvwlK+sIeoNICoP
sYK2+Eyw+PqyfnD9vLFgtxFS2XLkMidC6Ii3s+pk5/FrPeUI72/PTfZBejmTyyYQy0orjUp/lb6h
bOGnxFwepNN2+6z6SfPHVU+lo1l+fpSIRTVxcwtHMaBTZ5iumiqWeZFAuTo/ah559UMYXn6eBch3
1d5dU6485S9I7g2pEc4KFVEwlNeDOMYRtwtMHZuKCXijZM4Da/oK1+2zfuCIdg3ofpJRwbbUEUCD
UfU24pTHDSPI6MIFLZtY1ddJ+/Z2tnEiFV25fb+Lsub6WsRCJ7pm80otOgMq6+3wZyuj3Ylgvk0G
Myz/GACyyC63agw00fPWuakn6C1Xydnsv/hY0j4/E7No2Oe9ldJCCzn0VFlF4VM6muM16vmJXd6Y
QwNscfxq+W5TXNkMoPWs7ghrz0H1wytlq3U99Xbi7dgvkJJkfgKfI2NLdus3Wg6L//Phe9ZGahC+
G7b8rv8qfAPrlVw6jkTk1K6k3Wv2TFITh3Q1IGOpeAWbJ9csHbtRELyVZ8VHvV+p40ekqS+kb6ww
2eFvjMY5VU37KvOFef3dCdmZ1YtT0wm/f3NXZjUYeBksrOD2AaevEuQYtUH02tF8SY+6bk5oA4pt
IY0DaXO7uNtz5+JzgNQU/bi9GI5jE87T+6tOeY5JHuaZpTu7XGW1/ryuCV26EkFJPvrZAjqxox+p
DDkU+78eHzVJVyW0fPrFFz4SbEuaMyAb4loGRVHuYzGxrtAK5RxTppNdGdAD7vC133R+As9b/m+7
crLCVhy+cyrwoGh/cVhYQ24wf2D94E7R3o6IgiepMLzEus14KGhsQAEtR2x3kQRJ9/a5EscuIM11
D2ZVJ7ey3uXzsHVLI1e5urMvaZTb0OTaD5cLKhkLHSdiE4u5rs5FN1D6nmWKYilmYtknoHfZJE3d
331NYqDAPkWqmkED7QRMzNnfw9SDiBKUe/GqEah1K5r7s0P4xy5guACL/G/xyztp1hviO3GE+2Zx
OZdFU2KUY69LLC/qxfKn96ob/lWj3i9jy6ti5EUTXhTE3zRpjCXlAaUSQUPaAGcZJpFJdbe4q3Tt
KKmw5aQfIRdcP4VQInB50GhmUkfmhgrL99dXtPWpR427KT5xSiStgX1tpYm/6TPBcB/m58icqWb5
u/gXoEGXIg4ki1M7SE3xmlj89ap4U6Nx7RZsAE+71FSHiNEGS4TKXYLlSZ7Z2MqslpeSbc9HKHUi
hO8SIpf9TZGBcS0R2xwV4247xNHJ6AJ7dws05L7y023LvEshrwfkF2i26vFVDTMVFy/oTllBy3VO
ztIIE06JLC7VpYYwUDWTKRrMIJZBbNF8S2yZQ8dUPnqYWiuzTz5AjHXwHNEAex+uQbNTMZGdxExa
T0kjRsAv9+e/+EiEafeBMMdwfAorC2DnC2yXqvuUI977a4jRKmMBPIHAieIyoAFMINXeAHGqPzv6
/IzuiBNr41rakHiPKpcGQzshSLsHME65b+a6CtqdqA8B/hlwpLGimwvd/CgQHBW/Y1s/Fvq+99ng
H9O30HGAaEfzHmWhxA+IpYKYPCTFVzh3M2SKw4ZGlA4N/5cxodTrn+8Sem0aD0Dyoa9oMD5PzTU8
g/Yv6cxjldYGk9xlYX4qPwZKvJ3gKiRiSJme9riN5HJcI00SJA2qTI1xWwQDTD2mJv+TAeBdP4nN
/PSD1g8CBjfq0LBW0ScKM2me0XO+jw2+o/Uk02uEHdh1dQwclxjGmzmSI6LuLrHBviu7uN02MfZp
H8rFEWoAlxWXaZrY3XcnnJNoVWpayf+w9vQVVwzf8iRgUOHds/AxL77p93vojGkdEnXpyVO+1d/m
xGac4pkZkpf4+Hmg+PbkyURyQKzVq97C1VjXtJ7ojQNnOcdFZiv4F2RtYkLspSRnX2OrsdC25KKI
Obu0tRU2QiLhjvAsvRfazfPIdIoKaqwNKFCJ/OEl9G7xhK9lgVsi9u31CoxuRSdfVL7GAKHaiInT
aljhpTNHe+EdR58tUR00EgfQnCD5IHdqq8L6cttEOu8w1J4vpZNdzknFx3VuT+wEHp9BcI8jHku4
uOiHV7pEzlqTkGiBdBm4HxWLXbuLgh2Ilsxo3nwh7qGbVMfmddnbhkdcZ1wwfD0iBCBhb09uikoF
PesumlyQG8ft1WhMp10n9cDlmKkHHe6ZmoXLaQxU4P0+9U6vM6PmWwkm21in7/nH3rbC91sQBqSx
3V2GAb5CUCjfj7i7dxxwFktUU6ANjJndOo1IEHPMzGU+X3+JHdb7AVx0/0AFV5ZknAKEDemuNBpP
0i+Hzl3UYcNVfT4FMcZktDZRfguwDqGQKt1s4+Ow8pIzI8SexR03UqoVQSF0zJubct1+ilP4YbQg
TAZy+yxQl/poYyzCxIc0hyWz6628VMLBuzsnNjg2LwGdaZTNKj5WehlaJv6YImzgUuwN9Qizr6/T
U9Fdp7BFxBhX/6g9qWJJiYwmpVSDOACMkVIrjWPXFHEYJZKB7JDxTNZil4NKRDDngcESAPnnztiu
Sk/hOBGgD7rHdHfL/Z7GCOcz4qaY0ulRYPSxfRzubhfOhHnxVKc4uRJzh6kanqNnDIN0rDEgwPaf
N2CXqMVJNeHVsb1fySnZ4W14FONRKEdQ2RUb4W8+b9qHb5NKM2YCdNwbJ4o79XV18HT7iU1ihmJh
Esz2mHfxjTdiA5PULPhNnkrh9ephll/os94WuFPi9hIzRrqGaGeQ3usJZdJ9wj8qO5N+ufC4SRc/
/SehxBzCUIOMF+Yf4AePn2V/8V5vHjitI35Ib+kBtkcE175NhMea8IJjo6dnxXBbXtqC+uIbfWRf
vKwXjNcjAHbMd5PJVC/g+nSS2cZkp3te2cyR10aUHlLGWmJfGQHdkDK7JQQfJlgddfgjM8/ZwzBl
DBffp9uirPeere+05lPtf90+P1JALWi6gso4nlSAswSRrl+EJlJQeEnCOJ6uVWWOh/Iv2Sg80+rG
Ju6VEc4eQsYQbxdqpHGD86nf4eZ7XASrhHh9rvr3vqtar2RxzH3j+rkuPFcQ46Rv58mKAGAy1cAf
TZCKPoeIL3DDKl/7C3OZ0mHrjozeZemjEKcnM/xlPwFieq5qafGJj/LOKzP3qLGIaan2JwO3HgA0
Cf6ebFL6D1r5qiKn/6YQSo4xNsXSEPoYTzN9RcHEeYpbK7p3BGwMMHVuJLi4Jrf14BNM0F8hhuO1
+ciRLwByLbjNFDRExsRl0huF2CX0H3tIrvVLinUpsdd20Icm/JldhqXPJTspq2Q59yENelE94pIn
BIqzSPMBw1BlltQPEWOYqB8MrS1+/Ep//SbaGeeiFGomghAg4ehPmanwaSEPDsTgJDvvRpSTHszc
ZzMJM9oNzCPxKhqKow3jsUbv+1KS0+kHaLuikjULOnbqmcAK70v2sAAiuTM25cgj8DKoPt2b0y0j
PKjz4K3v1dmP0HH8WsTzcNdQxWxLepoalkRjo6nEYptdAxqBwefCiSD92Cg3glCgy1wZkDiS9x9h
QGSs/aAEo5q4KL2b/5AfphyFuLzMpPaIYLdMv2cTU/Lz02Q5HOFL+Uga35Cl/kD8VCRo0jjK2YKm
vQ3uoNEveEGeMFKV4OrHutKmgefvYvCo1Ky7OlF2dSx6XprVi34C8GJvjH5tEcNIHomgHL9gHSh/
wwhVV/BcIWSpZ0TErMO+PtWAB3od9zI0aa9D5sSf2wsq1ckPeekDiU0PgOm25KZ78rUBVorSAlex
3jU8d293rFcaNhnHjM58zR/EpcL5l2FGwKrCRpkz+MW1+m4Y/z9Jw7vZp/kuMvaWL5qaVgnSMamX
xHQIC7d9oTNVu/2LmCKzXcZnz8a1y2Q1S4UexkC759L2xwysj9AXFjOwCsC1iwYFvWrpC41g2JxE
GucNbqhyXtlbpunSPDvyXTWg4COR25DhPxnhYVyxv2+iewxILk0zXbvWwKFa5k8okVzlu9v3tcTA
rhTbJwiJkT5GJj9bfJoLboeSy0td1Oj7hDNOepqGGLVvsQ4r8gCQPbVMBGRN0YBeZG6Gc+fLT/Gp
havPCBB9Rj4bHo/1XOSoGriKsmlZpIyq3sViRk71195n5pz/De2++JFQ9C3yYCxCdjRmFXlwyTqu
orse+3C/tDJOwxOcfDAiyREcU8tPGjXqGF6Td3YT4NVfIyfVB+KUJevSM06j3II46InjV/Rbv6Qk
11wSollCWMnskCABPP9x1D4QmEFThqgXo2b7EOPD03Veh3FcwDd71DXxdN8xV14DVfPMdKGWwW1Y
ONzHgg3OO3xEmqLcVjgYvbS2FuzwgLnnYygzNp4wQpwcfNs/NgQdDwrHiE7jBBDIkc9eoOJO3xrI
2PgaNe3sa4LDkhqGRmjryZfTPm0ySg07PY2NIe7MF5gMAS0absETeC7Dym7HC5tTAYlijlrWG7B+
chWEtCi0dyjJbCtiMCkwKeJ/NYHosVKVzMXhuHFTQy9YHCIYyioes39BSU+EySukcZcoDY98uZ2j
QF/xOQkVvw3rgVtSBZq6hd+V+AK2J9hC/b3ogADC51rmZzwy3SnwUSv969AKgDgTbgClipKUcL5N
rl50hX3i31Q6blzrGotXswRNpmsVGws1HQk2FijzvHvmC/uFZBXVaGudN6ZyCQrhuxOS+Wbi8s7W
EhHNTv4mbg+ZAI7QpFydjYRwIqkH1jgRcpONT0EChVg0iHyQXx1eDbwd4dmjGATldlOI5bqAgH6N
8udMz7IijfXF7UlO37h+QWDsoMSDxgVlotJD0hip3GabeWSEAUcbqPBLvhztHFgq5acV2B9esAle
lkg791HzfC160yJbQoQFg6hn5z2lkk+V2rvZ8x9dlKBlo1RURkHusLw+auk7Q7msk8kc+ZFUKTDw
IabfLzvqi2b12HRM0QC4OqWGtc1jWhWMJO/y3zxpQSXfBSCi8ImOmFKKCebddZDmSH4JPFbtBBEG
++2An+SOyQOJrA9yHNuNDyH7vhraES9FnSMW0mv3acshFFA1DPAcw6NmEpyyDTWH84jlmXpC/5lX
K6xv2bb2aY9IFajX8qmTR6OzFCXWg2b95CQmMBfFIqDwYQ/p+a0zL9K/L4ArmVnjW7UYX+W7yjtY
WmncgswCxRgMv1psZhcukC7oNoigaChbxJSkzcLHzPG3khOA+vfA4FrVfVI0Bra+6O97IEQfNTdq
441c0zMm1styfdui3h8b3fn8CpFdcT+uRWDrY/rWDKM+Olns0YFbQuLAhJ3wwvEwmKYXJoYTu2jg
h1p+CadDTh2xYhpPW1h6nm2wo3Fz4MGN1lvTTX2hXTSyy0GbTTzkFk7tgb4HwDtqd+ZifmFlygF3
Gia2IrZSZYbtMTJmkWy/HhZUldh6EEtVfI1EwofVUwGbX27VkzUP7nlNWYEpU9xdqwEYlpWvxIcS
+yci1ba6zLldxQk+dKklBl8KOevoncL1HkYxhZEVivGr1Cd1KtLp9laQTeSjJauRxdd/QucUxWAr
/N9DUAn4tXnnBIrdoSWE3UUEgREGkQrCUoTs/neec71qEnN7wcEodBxysew7m7yudUgMRzNt7rlH
uPZHa5Wc1ty0uRLxPDxNCk8/qx/UOTSDhdP6vt96qijGkTC5Mn+Rqz69LXQLY7DlUgdWY6HR5SVn
wUFU3CbmRkcz1gyMDEZox1OAYdP58LSbyyTV/0f8U9s91oPluq4/6BVrhOde2Hjz6Q5+MWJgOggJ
JXoq4kXTR6eV0gthBE9i5YPfxAZjNQ3E5pzfhxJgkm+eeTv40RnGhw/n/cjklWHU2RhEpER4SFqQ
4klCn0bMMO7JDJtzPIe2jsAbWT4pGlK72yrZuDZsXBM8oPBDgDUjvjH6sJepKVJLS2BMdObH2zCL
aWMyVSEfbq2ck64Q7imLrDHetD8Dni9+asp+Eu882PJPjQLyjUwvR4uYS3d7CVo4DWO+2Mq66I1y
SDixsZMWHa8bqjUCgIGchFgvt+uqkboOJB94X/JGsUBJMJi2MUVvbBv5as7hElxlYriAI5BloCXY
Wns76d0GHy2qEsKvHNUwICp+0EMARockXV8pDfTWtKCPf2bidd14E3La81NBVv/3WsKW1lnhIHz+
ZQg+P7ua/hLCfsRsDyerBQDsBmlZapIn0Haib3LY9vfHfu64xihPuE9XqU/Sk88Wdu6SWxYwDCnS
r3HBu1b9HNzo8J4COWL+UIAH9JnvFXZKLPeu/oKJZ9Azp4Wut7NVCiokEt8szWUSRV8nBuFxuX+e
bJDzNjdNpeYi1cqeg2wA9pSDWGkI2I4N6wFgsY95SkLkAV2fXqB/O8MgfMAodBCv4KAgxR5l8dtA
mrQ0Zl1CRzUTqtk7YgVbmApiP3+ng0JyaNwPNOO+LZtp2eVTNBmtAqIudjTxEI6KFqLdGEitLRyn
6HzdyccfXnzQrZGkmFT7SR932/dnBh9kZq9GpQTLGMOEqVrIL0yhbplaInQuAwGduU8P2TbfYG1t
jXEQpD6Vgwr1Jjgk85u2zlvc/lQDcD7u59Z8R4Fb+Tb1gfAHBDhi+qDZW7Svr3+LsV6QpRCkRCbD
WOWjlrdsJ2qegXcu43oHwkRf9cNAGp69wp+/xIS5qqj071YMpylOZ1iwfD7pohmSzICKbb7s9nvj
OcPo1TRvMeAgzu7fsazPZrx1Bq+7JNp5n2PeHj8Q6s5eq0gDLbJpGvUUj3tr5O+yinKVZ6YC84/U
0fEzn8dIZUEyrYC1GLoVz3X/zxIZzCvpiQ3VqouRLYOJniT1A49x6+RH5TyVOdfaYal/O7tBXhXF
0VRk+d5B9f6P5btnFbP3h7lamSMH3DFBPgNgFAqJtZn805tyJkgCOu7ON92UdZOoRYmxTtNp5K7o
9VRfPPbvBGYDH0Qccx0+oZDaete4GLSxgD0zL2Rl6Us9Y8fbaErc2RDlOeKzKawTauVK5Qx3e0yT
I3ZqcJrFb0fD2cBtrr0QnHh3ofdxrHQ3kfaoPwBU6+1t9UDEmJ6USVvNtoprE7c1gXuy/nUNgKUV
8dqKgx4sKuDnzEmoDcpl4M/S7UF2V0ZcuShfBM1ueFbhZ+JFVEJeJPfipFVUnb/KEG7XjaR7v6Sx
OEH98NoHo8ITpgA/YwXw6dzx+Vx06d+yjpyfmUT5CD0qEf/ORzJIUSJw68d5czq7Z9MMV4ze5nRw
EocxW7W54qpln6JWuN1plfqPoSYs81LLh4XpxLpIDyuOJqWfEwqDha+JZgsG5e2a9SElTN4DJEws
QqtpTVNzPg5mrYX9/TlSNAbhAldDBXXxH0pdTh1gQb+EXJkEyGkfmnEaU+sY3sisXHN5lC/BkMfF
SqecD6sgh7iAaTRa4QNe65l02LvsX6XeldnWQ0ytW6DkS6iUkbe7WPhfJX0/MGwN6l42+jTXV5mY
IfzeQWDLHk0yKhKz0kJjQvIhgPohLdOx6lXjUUgC7AWSKPtRspE8htQBdxaApwemoIaQm0JW3HDY
Fs2a0E5bd9U8Dxp/PaSiVWkglYsDqfFbi9skvvmELqtlW6NeO3bWcN2XPL0/gs9usCi92tgDTCIa
YNxWZqLYb31wOdWxjXaKerILVCkcCPBLFc9xpN/Yap0Nk6Yns2P87WU0BZvws3FIzMs3z8K7kJzL
3TZ5hlBeIMZ54qZtYGf4wartVEULpBYf1QjlasXMn0XY1QZMqVkGTFF3+9ZGwIIqXdLpwp38doap
p8IxnQ6qcVAihaKliPIkY8IpdQu6FmF5zINNdL7NKuwTfUmvMJXDbpVhRGlrrswajcpSksii8IW0
VsDjSCw7d1RX1pbemia8bTx4+zYHdTOo8qoZCxt/LRj/9TrkZg47KPHXajCLV2WSBWlwFNAiKEwF
yoFE8K9XBA/TBPSMKUdiDGgZu6qI7QilEaqLLZUU/pihnnSarIo706YyRtfiILXAWfXF6Jdfhldo
VkhF29LJsmmdZPh+9OXcuxr+dw/7V06qhgcGx84z91zdfi+zkkRd2aX5QrS1jCvw2n/shbDMkn2Y
fxirr2YxEh9emxrhAOoJV7IfJFAiFrrMtT32NzEd+EzOPoyZRTMUvaWQv4X58zSGws5dS6amdnG0
LcS3Bv4yIGr/hc2I6yuscfIrIm74q1ZfjMTdJQGlwkYzk30lz18z3WQ2iUKQar4pMTHyTFUNZ6m6
k6owxG//byKahckpw/ipL3gL7UwZOGVtFpgIBRSd5jJKL7UBPHcZE/MFlbXLETQyrHanupsec6RT
pwuy5c0lst1VUVZ2v+QRhcCJLaItgZFI7eWKwX3x2pVgBY58FjjkSZFljw/wPQxn/39HTQ5tOG+U
7pcBckAfvnRVWtsYueYRr5Tbvwori6jHwjptQyHLtde10r4BiOOewRRdzAqY9smE7TZc1DWAP6EM
PWGqNYZnC0s9BQc4vc8GHSvjmllSc74kdcwvZir3xmjCh3Wji/Isb/mWyT4QboLj1QdcqxqrHGXp
FfUCvQ9vnef1xdKzVxge9sMnodzeDeZLAiwYoarutH1PecuyKYEBUiFmfK1VDnZ/NuMZOT31L/jQ
L/f8NW+YSOWG3ocztuIilPRrZOX32cffhOnLTNJqSEJj5Oo0YsmjBA4VcM3v3FQv5vWhEwMZdgb7
vRPMqly2ZYOZ9NmQpxYm7uy0bUyrydn1Xri+UC13
`protect end_protected
