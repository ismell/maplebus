`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ctWqyJUUBfKRcUDtWGgYbZiwcQay5L7BHTx/RoJinudRYb+HoZhmDhFBTPkMO2SvIxqsAo3nUfRa
d5Fa5mmDuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mi/WG4nRQA+Kfc6PLPb3SPpgqy55aEw94m2SCxv24LEBLQ4Tth20qa0WRZ3qwCuPwtJnsP4dJhHs
15UU5sW4qAuttJqhfQppkwtbdc8AJFETxEQrb6/PLYKGkR5NIR+n0tQjYfgwz63LAXC9v0j6zMiv
vaK+7VXNf/pU/180598=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LIfr+GJh9bDB2zPFcM3eoWcAlWtj3sNRi5wcAAkCX9i4+wOysat+DiftfdSZXlqVVfFfSN7hduJV
X+r5A7b5RhEcvQQSGAUJ9hEBGbr9PxqjFfkSYFJmJCbZQ1wUQIMisscOD7SPWh+L01eiedMCMdxA
IWXQg9ZX2rvztg6Z9fnXvYIvqOX79kva1lgZLkE9TITCxiIP6E3lduvk6ZA9bTggBigGdZC/LWT3
cTEvYX+Ql0gvvN1EqWBqhXszhSLLy7/SsJoqw8+ssYrHjsYN0a90ZAp/jpYynsG9s52fhGj4IYMB
/Cr+/Hmr2UAQnrvRm2PTXPC+wBRisbrIry2bGA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HpvPZUvbd1qhjPREbVGtlwwVmpuvrGhaP3aD9uiXoKMinTlxg4Nt7Otom0iPix42/LYmC+Afu1x3
WJRLvpCcHNOR3R2iImun8BdoQAoaEtNmkiuEwTy/uSyonEHSqc2E4j6Lb2x1t8AdYzEd+uo587vn
YTGmwp6L8yaLaMr1zVw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rXPAw+1BjPdKhomZ5Y4Mt9ZoSw7cZunG+Ov7A4x94mH0sD/DSOeF2K2aX5bXMyFCGWVBxT/cbV1U
2vDbjESYaI2OM0+il3UWd80fLxeh5FR5tP1MprXDoTcd95pUJwPbxHR2exb7VGIrFlmR++oH5StL
SotkC1s2IAKROwVyO4jazlPFdgLxzvwwEvig9uEyntRCuHMBEwOrLLa8SL5h7azVZ/2qz+R9U1b5
ufMnmy2tk1Y4UhBZfvT0sjTI8ZVcnjtiEfRhq/tKaEeng+AlTf/gIftWXRSX0xdGhPqnfbHWP+85
6kOJVlvsHP2iy3+he7+KcAb+mwFSNAFWGLW10A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8544)
`protect data_block
KhAvQfVwTE3lLAcgRGu8IkbZgFvI081C0UqQcU4udvpoqrm/oj2Gd6TUU93nHs1ggNSpkiT7vbHd
FiSxIyQBJgpagsHZO52VvWYNQ57TeMQOYlnR6gm2ly1TVoJcqWkbrO33PHvY6SSgiiIn6208Q7YY
jij4RNiG//PpoyvJV+iAWbcis5j2Q2G4lusIKj+ofQjlnxmf/VmUH43O85PM93VpN8LAOObmKrMi
90ha1EljfpJHUG3R0dd+gWUB3cSHb4RPu4yQA/O64FZNLV+Pt1xJoR10qqh8nhyTj35BOGr0AUnG
dmGigvOOMc5w2Maw2ALEwv27FvNI18+J6fEQ00CkV/05JiIAmDcRUQLWpQ557ThCZEKA4bDFy4Hp
2oUjS/gOO2wQCyaKDPqwA29OZHInxGLpxSgMrqsG/7vCRsjSw74syFM21q22YmQ8TBuO7CpSf14o
57fHyrPYc9r/xuzxJ9azCmysqYv82hf0tJVWM3lfi2/waiJPuxjra9cz9aQwhKUypszp7jrHtCSL
0SAjJbmVQLo2THQ9SXvQ7kv4FuDac6fFBfKMPuMw3N6JMFR2/w9tHQc0vvdDbIo2g+JNnTRIW7oQ
2zECZ4+NVqEAQs/YNrgnmmtQQunLu9/9CMc2sPagO1VAXsteSzFptGo42lMXwfJt0E++diWjKOPv
kvJzaYlc//4RENqtIzq/bniJHbNsR0CoYvhyXHn3aTjqsFqUoFWEq0eS10kTFIiccNNHrOxG736a
sl82MpYPGaIJl4fJo35W+9WB77k3TRBXaM3zou/YaqtmgS1rBz55IpBvFn093F7OtHyiLuAHjarB
NZSpojse+TX0mx7yHK9VmaqwbP9NmtfXeh2p7ouBtU+oX4+D+i7J1JvccmIvhBejDR29izWwG25f
dI93rvk5ymqNlrwo4jBDqRwFOdl+qFucUe/MHSeQxyS6gDkfJawslwQY9lhKshPBezHpbEEtYhqC
IYLwZciDzCuF/h8YXyghN/saFFTmNfffDXstcwFHw2YQ4kK2gfI63kCPBtvie9FsGQLNRO0N7ga+
FK0+yjRlwfBnLAhqsUehrCXGesb6DzrqWeDXTPvBWFfZHBQPO6q/HGnKRHcaGCWjWgp5N2AcL3rc
tDgmjaovVLhiyzryiOjN3H72W/pl2fRV3oAcLJ3IyxQv4xqk8eYya5IHox30EZc/2/mN52EcYIMu
3DZP3aRN7mfzaSGPhbLKRrOAZzp6m2Q0mbu23vlrdVlgq35xY1AEt+u0MGCS2VTkDYHd0fs0CYrU
/1wqaiiZB6RwQLvFRqNWyeGLyl2XZCoWk842xjvUMAYL0EF1xUfouHb1WC5TmxpCcSAXryORu5Rl
QqQhscoIUbj3gxTY4iBiHEhBjUQqKRmcgH2iMT78ybN/ZrtlWf2LJVZ9TO6SZxUD+M8mdDt/tLxW
QSLSdMAoA7OO15d5OxTn2GDZg1wbUAHAeLme49wkEIy7zcWLVfE7wt8yGXOFNbD41gS1nDSbLb0U
Oceo2STEd7rHE03bGHYOhhayir9c06Xy2btzuZ1Ft3t7aGJeGx8G0WQrqTksgnGkKz41Ds7t6yV0
691PXMLreXyI5w1lp6g7DEZkEoYWPwCDtUODPrP6MOS8qFNLE6ECcgxijl5DX4z00knhTSOAHnCi
KhmrdFyRWtDxyMJkmSmQ7eWOQlRhfay9ejADTPWLVZWrESbcbb3adWu8URYapM2AJP7y75Gk2h4B
Io+0rYP3yGIUFJPYUiVjo1xwi9mj5XMHlKUPcH7QSAtlZZ2fcB4DCTGsO09MhtxU+Dixra85OC/4
JSUDLqyabcIm1dbEKt0YPvflFHGvqGZqc9wzTclav50TXbH1eGTDfBGZaQjMPwGdvq6iyRicNIHm
w/PaRE2Pg+an4sYpgHn229WqKNBLETbs1Zh7gXEjxc3Mg5dQmG8d+fL9IMQ0eReMcynlj/dNLb4r
vZHBDzAhwRdN6BmNWOBjHnVjLRVNok6Eaf9yww7e1lUftije2jNa2yayky6mslQHj8GPfgQ+vPyu
BvxnKRRawH0IUK/xneEEpS2NxitI2oTk6HaDI4/HCYzLVEygk91PfoemWck0T1Xxo3eyeJSXP+eq
4VROSITsFuN98l1vi/gVh4a5CLB77Tewd2CFt/mA3pbzfZv4lGsMU4gqcb5I/hObzObmKLUKjFjE
ejrNhUKQkwJPrvI/oyzPcFXivCoLVqfD4dZjrHF2fkVgDIkHKSZLP+VuccX0mN70y4duWJ72ePTk
8FfmMMstwSX6I47wlHmu+bUb2+EDBP+aPb//3aU7k1HeAle6Q+7/JwjRqV/ag4/3K1kWEQuiLR3I
Ay73bJzX3GGgo2hy03pQJFcEwBFl9E+GqdNJvbJrE7g/4Qyqc9D5r7YQVjEzTIGo2Cx/wdjTcESY
/+iulDCoSGo7d/735W6opEB0/Vc7I1wXQ1GXUXxpJ6ebLLSZlD/dKGmuE4iSYTpNLe2CCtp14t7k
OTfibgcloC3v30Kq/wsm4hTZwYqAhw3/GnJonIeyttf7c99vZK+xu7imExeCnJl13EZnBYafSAvW
sAUUR29JSNu+G809h9vaEU6Fj79MfrQqhbDc0D7gz4iSnwm+LaTvVr0OGoP0YtPwb8viQg3zcg8l
yn5W/MHWRNhXjBKj6RHDkNdoAIBB8b0q2EGeQi9tMs08i1nJ63B/GsTSZBB3goM+vuPlTDn0kCK0
AC9Fmx8WFavgetA1+p/vJL8ZFH5ckOtrenk6Soa65Iclb9xXh1vcXC9A4S7AiagTrwBtwlA0JmzC
vXgrLfhTOfwqVJZ4FQGZwnnhHZJlFHiHFIjvvo/2GE832PdH4OTtJNAEUVRNvEqo2reC0Gi7oYu2
4FoRLw4oHYv9FdRpxZ1gr84wYgEovRvUKxe76atA2dCQV1Mn1wx6pHUWgr1/AdPqzzLCcg0aAgaM
8rYOGEI/k3ibUz0IckAsDF/2Sa6l9+LIS9QEsZYDL/rFIprXxpW9gO6nqTqCqE3CEM7EXLzTS8yp
DoO7B/+6ev+N5rLsTtc8ycnXmXiIdB+2+SSbX/7u/Ov7P3YZqECjwcVoacIPe5zEa2k6gNqHZkGC
LfBxSsGGeJ8OiMaUnUkn+reGIsFyHOUcsUSiktclw3RuKjufMVe9icWTKOpRK+ADtyoGhQWlbMSs
ERwxrkNQ1MAyTFH0MvTMEUY6s/noLPHlgbPqMpHhf3BfXkJGNHzjc8hc1ISkjHw0MhZgPORH2ere
a+/caYOOgDMUa0WItLqceWO2pIPf3JT4IfROf63x4g8syfcMl0y7BgBrMY9CMRDsqhjufHqlfXyu
+5jBgUqJu1t0qmPYOfPrDTM6LuACW7TLfu225pOlJfPfBYtTFLkfDAV0yW59X5uPSdYyIvU3WqoB
l+co6RvBH0ClR8J5S0WDbEmttIemgr//WNz2dpEeItlHSK5qpBZdTuQQBzTvIz7CGHQOBUY8aUZi
Aj0pLxepIE7ddPlF3s9fhBy9tvNmI059A87ZniZ7qOwQndrRyJFNzzbBJoDQW1Z0svCnyrAgqD1u
vqN23kDrIdJU9ObEK89Kd2Kt8TMhhl+ueNa42armbOZBcpHMWUU4WnqpN3L7Zr3148dtf09g4KHq
cMa60hkPtx4cg8MIxmVJzdUo/nn5W4C680+FhpGmlz0g+tfZKiyBAb/+Wm0bX6aKG8/axpypU79y
TTofvulYw0Dl01690fyCfXWHD9SJFm08fB5S8ltfoBNk4xBpp6fP3P044p9ru579uIyjcekyOYaq
IPYy6LJVELMR8d4XxGsCRJvRmUkufkFEVQfrUELERkLlLL2R+Vuwg3O7l1YfFWiFYKS6uO7nROws
3YOuR7QOEtuiZoDbW421FgYviHjV3VloDUEfLaBTLvi3qRoQdtc8ysy+k1rlzWewo54ocQzVNNOr
/PwU8tAHVVKyX658NsuQOuaeJBc0HXTWJirykrKIvQAGcQrOCw5m7CqpnNH8JJmIGaY/7fycKm8o
cLFvA3ggaXCmBaKVapRaSnTf+djxecVS8aADH7STa0ikxr/oLq3al6P42VN0zpQ9jpRKZ0+PcdKY
ad1ltk8x1C6Rfrd8nM5DPnoSfDOAb424EF4No1JdlYKUW0xQc1m+1OQAhoAwrl9M/O4TWzuUT2dU
KI+DxM2aoG2XsV20xDxkMyTw5F5pn8qnmvcgFIYJt4pNxuHAfE8z/bIQHkpXKR4dF94+k4hW2/OO
l8HCesxFBZzza9hVTXzIZ/YGGIpe+bsNzprQzMz8sDFnTRqA3cnOrfEO/ZSkDlZa0gVDTm+03ww7
i8H2dBAsit8TzBIDEh9Qu1Fsm7wPx5BqdrNYSnlyDk8IxphB61/kPvs7ZFSy88jIUclbN4T+JPBj
5oXw/Bhr6lJJhgsWSVNTj155GTcpQU6+xLyXnRIei5LhFEzANshiKAi2hLSbna+KGBoZcKky5hcr
r7ON/zUj3T7NFGYIbpB08FF8urBtc/+/kh6Dv2OO1UOIJSxD/gf4XqO6U4mRRYalN2KoTI3Sq5P5
8NBSK2AuxaE/dYMPiR1eJ24vpgmRg2HuLJtoVJccWJAH5lgkdO1dPULPc/RroEHLXWhuCv/zFzqL
Rw13y0HJMMKNAbOokFJFtJ+sxSFcKF7g2WNWOa3NYDa7eteZABbSTQWEaWfqWxr5S47NoXXBrwmd
LMPISWhitaey9XpO+CM62lLia2kq7njXwk9Ky6BrIksUAkMUT26q0EbbidwuRgtJE3Gw6RFi+Dsv
8mNW8vQQpNt4RMuaba9UriLeGu3oTP1TUvn5bpBG2e1hF6e47S3VEFF/tTfehdJQ79MJ2vlXVloh
kpsKoI1X78lnEiX6NXJgoIqez6uVQ2ddBmLi5RR0zY9NuKq6OmU4ul/Q77C8Ips35YmfdHykTkeo
1KxYYYGp4I6gdOujgSVfvNoxx2BAN7ouZN9q3a2LQ9njMvEb2fe9oBKhKfDxuCCRYhHVVLy+hXFb
7XERfI1qCXktRMW4hoBopwbNajVxyghURCfljPOJw0LhcX8734rE8gvWyM+qyux0JCUWgwHQ7azS
uBCQ0NoRALI47+eYhnIFPS2oahct2s0+l+bNbKTckWxbhgQBqBE2iXBeu6btdgiIRYY1Dm4ILzW2
pdkl2IYQIBSA8SAsR0qnUlG9jKLd840rHUr2O5xoIQpjtlyN6TNqfgya/fBu0j4+4WbTrkQMK2da
NSkBKdzAXWK5hJAjI8ny6EaDdd8o5Ozw1QcIOR0gD2p8kiIQ2Kl6AMrOLncSrLXLl51ma43WTmOy
fQavuk4q4UG9+ZspZeAoDmL2mdIKB3i11sncG76wg9+2JmiMGSTdwKa4kNVDFLC3IOYp+Lf98F82
ntvyOWx22k9JiebYlYJt1syZWrI3gkxAhTj4fdHUrAzn8N15ixxzyPV4Ynu7in6E0immDPdDsQ8y
qq07iLRpzOdeN5t1CP18nSTfZUVhIskiVNGl/a3NeowNgjqIRkF1wtR9mfOkSkE7TaYhmrKivErI
BpMJx+0njc2ykCkbhwreoolqgmgg/1ydiqy8amPDtH0D9ECXArnpAC6j8zPX09GT8kE2UeaKPGof
DMMUbZ/8Xs5rHFoduQBE/A6lYakWplvCtum9F9jJ4brWjw3FuvGHyH0rD68ub3sQt4eWBpd3pD07
eP2TbhkqWZ2qBqsbIOE6KDMcz7sVQilH6NfrUh6m076aUr4DEOo/tqeuI8H0g63+gvGEl5MbtVL+
4qQWSraQ3taFbqyMLKgsOarRgYXc+drPezd49v4Wj+fXvNA8xS1Qn8bzHCAnbSbQKOKDNgisI08j
8ei9jIAdAV/F+LltG3bDqCjvZOKa/INtbQP/2Z4k1Bif9rMoLtKVogXqhEbgA6PYgjaHUmAMSe3X
I9y5qcXmXjro0bU7JfQ9aajDnuOGnwGbhDgUdIfDRXuIjbK657tXcE7kUqJGUaX7UCjuo3l24aka
6fMVzttHCo0GZusq8ZYUoUh7FpRI7s4a8ersnIIgCBljClREkZCLnsmMOQFgUpsvYa+8i8vGXTvk
sQ1COk+C3aGk8ZmDhNVcQcXEYjz6Am1QJwYIv0oIvV7SpSDQeDlQlLbFtYSbc3zfrZF09roe6rZJ
KX//SFKst4N/GPmIOVqSfccyGBsRiaL+yIeneOGw7roddJqH1gCPv7AWV6vs9zuMJus++lBoaLQH
5O39KGP7xKQ47+1ZFhc1P4LtTd4t98FCQTC4Ts/DgvtjO5GxNLW5ww3OOWx+GBoo+0vUSZpCcH7i
5IXLDMuKXY0KJD+FZegA768RpNaaZa0+RkbUiNZ2AMnmm+y7Z4AJZy9UMYhTLw1Rxm840n+VNY1R
12VE1Ob4FAjNlz6ykhiDImrOZ8+ZB5VMxvZvfiP73orK3gFHpSSbt8fdKiCXYFZEu9DypDMmeK9i
nft6Robb5dNrknG+PsAv70lMKp6PmsFoR8fXa4ePUh4zsUwacuGuWEglW+QXSCMy0eDncN6N3dlv
i/Auq33rC+bhPCXa05u3o0aLT8X9wf1J5n4WU20WFMXGuU9YDRuJPs+GOwAaWXZYAaGoh/d278q3
HEEsO9b5mo1srt3aYYDVSpaVnyA7ozhuuTYUW73dx7Y+TxeDLYJAR4tsqYXtMxCwMcdMTcmQmKI7
hXpo+YWuUQB47AQQit6f93uSC7j4zLxjS52laTxXx0LHxXn+xxjSNsYGzdzXIGwsqQhmAsu8Jr84
AIn8nUfAEeCUWW4nsBST+7KPLANqHZ3hOUE5vQvSwlrhKuyk3I0Lm0A7VJOQ25Xqz8UvBXI9UoYh
nVaWQujEmAnJRB17n/HqEBgll8wAtMYjP0xQAiCW0SQ3nxRGvtoiIydAeey8TaaUyQ0UFkzfTryE
Ds2749LThjmYqO0xGcHBMOvb4pG32X2u7k/hP1pE1bBVzjXD9Ax72tQjBGdsm6aNc3fVXS+GSSDX
JZUVf7mDqSeMlmut/oRgFdopzY4zdSZDJIUu4zOTnY3daJY+G5YlifAFUJnQsta5rhj3i0y/RzCH
J5BTE8GNfDxFwzsAC2i7HQkJdqFVXOza0G0QKgB1wdaucw3Aw5Cq1XwRmghFk0Ah+01Fcr38ww5e
ZFWTZv0uGRk9upTwvcIqkFGq7KZEhC+gFCuJNN0mXTqyCiigv7GdwsHGzVvxRhgNdYoM+nEpxuci
SA2IzVDESQjJdN/pooLJGCMp/P+s875uyffALNKG5gzLCap18UBjJpoZY9lk+zdcGFtFaVhYwxbw
kw/o+LG4wPRg1FHMbZdeMKw6smEhWKcZxuCodS/nsBuXoYGQVQj4RdYQzRxpVw9ujxhCCPZsMn0s
GRzTWLbYsNnG87cVPY657hJoX7Gx7VtXnYndomFxJK8Bc0AdzR2OEGsNUXjMdrZYMDLBToyRAZgJ
RB/7ndze+kWmcCDM6aRclDdPwhn5EwxqfFbzVxF2pqEsDkUdMWv8td5yUGWSZCCy8Dq2pxuk1Ksh
OL0gjuesCTZ/fYqM9wYvInZ3rLImt3MuqPZxbJbL1m+xekWFF1cncry/q1dUtujK76mtoU2PoWPR
Bg0W/ROpERID4TRUh1FSkXc+ri/maPljUlcXIZMQGrkBIPKf6G1LaeF117H0cCrhbHoqU/XsuE+4
60grlKTTdFY15/LhYAylRkwOiUuFLZXZrfEuk5IYBBpIo6HILgcOw/fy8U2CBX0/rIynB31Fl19t
u9m/2EvmojSgME7mXLmOfQxalZEheI9Ugg44nkDc3ldaL0yQrBGsXH4E1YyCPJUGhzBsq0GULg6O
uNzT/aXE8WTO0kRrYLNe9PICdbTuL/Y9itV35vw8HPvrGl8v5HEM3B8Ce6YLEoS8dygmyXr4pF/j
OGNM26Bn4paev3tignxI9SUbuwhIuQK9XHsW+olMyrU6KirVvU0iS03zoMtEuz0jYzg0a3GjISkg
IbacT2zE8QdcgQjqZMrc4jj1FsPQdroJ7nmZDlOhOtL/DxB0Gcjx4n+ihEkYTxRsF5cOCCTGkdPw
8Hv+BCvIznFoy1Vw2QwDiuVk0khbelQQTO6NNYlHkwoVGb9j2Tiuu1GExlPUBgcKR2noYGrRnjjm
0fAB8uo0Q0cROP/AOlyYzWims3czVNK38eey6zYp0Y7Vmi3usbBCzOC8umXMABWE8vQbJIjc1ZBQ
i3/s5BMTdGnfXQ0dHAtYrNXi2ivSAJBdwJZmZkedz1nJFeYyTXog4zNydCfbGV65wsK8SDlyhZUn
9MzXrZWce67/awP0KGiISpLzu2hR3lXR79WCyv6LFuPmXkhiC859ltjaduaXg9HiMrizzZB/23oP
a3qHyFHEGra5Iccne0TDKMxV4VwCbrUfmu4cB1rHFb+o3l6I9/2WLy3ZgFJxF7F6Vcccxg3rPcyG
U4JgnR//XThvGgfITCx8PRgMK+P9oZHd5wrseQgP3pGeFZeaBcn+TI450Tf9MMMQ4Z2QT36K0Zvs
2TBJCelOnqtmpY+40IYMxRQaPNBzdLbHhKC+nOXpkzPlotxV/cOCnkWFUFhY6qiuRYGPSIFJI0fF
qz/kILFBZskLbNoce9mHuRuClRrVJ8OJpMds02fWLUes7oy+7zrlCmjWKjH7QC026QjSM3UlDyzP
JzjIctAYV171N9PYVcFqYUCuLFKjoKEnFkUySMeRekgo93Hga18stZyeXbsM1shlpOsV8VCBUrFa
7Se189hfdnXoSgtKEuCLDBBWvLJpfVF22GxQkpvuznitxYHSuTUuipXtefr8tQmHvpLWGHlB9I41
5UCqlCSM60pOzPBGrh+wZRGSb4H3tC62tbplxToQ7eRD7W6TJ48/YzFKn/zaO9jtraef+ddwp5+B
4W8fb8HrOjUbGjhcqcNZv2Q5WOLj1n+H9MBFDz8/YyH3SAod5Ey9/xuQYY5rtXFA3pmWpqeChGhl
yiyrYToqsXRaCGpIjeEun5dbZ9a4rjz+wdjnm/+ieuQWzaRVUeb2/Qg3/gLeiwDwHfmB5kmFxix3
YDKf0THHrTHukNI/2MtjGct3aTkAh2VJGPHg6oumyIpl+QcJJdo+TGOgWd0prcZ2b14tAgsutopK
BGZEf+hc0z3PlKOJ0qeE0l8dmSxXBIaha7wDnoaxTRWOWn3YGBDaxSIkDo5WuQ+vdysPJeByTZUw
+fGknCcZo+rkZYweEcolFDUDz9hWYd+E4pNLDda1aN4ItPMFvpEZlPoS3wxFhoqjJBkBW4CwSfup
lc5/pCiQobhKN77Y5pMdqaoeIGnzSvZ7iN+pFtTblfsgG7i+0O/OdWyDCSZeAhqwvhzmdS9vk3zO
W/Bk5UHacPCYQtL6DXyn3NRFjBYu9ZTeEdsZ+kbK5gfUcHvZoPdZrelLKa8uA35eGyXNjRdg5usz
7vK8M+XBOf/Q0lbZlgrf7hzW2ZvMk6dT/AIPDUL+Nr08DCE8y5/XYuwOwDf8nxTi4a+44EQ0/AsV
4ceS49D4LcEGx9AJmqvWde/jSYwNQi7Wzsq6oSSS57Q4lELOvvdvWgxi16VGqZ77XyXykF77APac
kEBrnuy09wEWX1gwFzPQzXkkdDtJR9rmXaG0x0nWNBlSpAX2zZxSIlpA3oW84XOSfDJ+xVuNqACA
N2Y+pejaPYXWGkjfWMxSWwb7/w6hVx3HRAW2sYoHdU98++0ViRj66OzylkARoYdQpsxeX6Ocyxja
HBM+Ku7ujaMDVJpb4IP9Z1yJIkMQ4jfllEuz7tjdrbvzcoNMarUb7qZWrHis0fjuCtpEIvqDZV3n
/xMZ7ol9sRWveDusdByNc4zmFpHFNMqu66kpWZwFKNikEmYiX4AqGf24G/5DRTkpD+m9vOCzazzk
yuWDuKAsHCR+OpdclpPrUUhMpgCgFDko+h/gYjKAo9nOr851VVXooWQriM5v2ResEz5sQiPNf2nl
vPkiXEwBZ1qwpMtXW+xTBw5uD5vO905ZVp6nmca4z4WZK4MFPpVGNuw8wOpX8zGMrpl1/nJBiEM/
Dz+0mU/qrBW8MAcIg9b2OEqzJZaNuMIWdUnSwVb9JR5z5XUqlnCLEmKPNGVMoC+xZJbk7Bd4lXo9
EPUyFKz86ZtXD400AFour5WYfa4QmHOCbZ9IZAP9JFguuczivigxqcWaP/fISihtMV56xku73esp
eZrWUcgkFc8H9p4H2lhiohc0AxW+azT2tTAkteiaDKjTsc68MP7TlmbzWvaqKDkB4VCTD9FK8cji
ReTUOi3zHiCcTkAU1FTKyOq7xEK8XU0bfNjSqxdUiLbOkTplOIng8yxpQEhWoPNHXJ7io+2uaFMT
tcT+RObT38PeyvxORAXRJgYW4VXZrnvtpNg/c+Aen8SL8LkwDBTkl72/wwwEtE02qOLk/A5xQeJ8
xlsBF4F4JwmECxSbnzr3inwAloBD3bFV9nTqvhCEyLC+d4s4cEXBBoNTRc4B8gYg7Bx6EZ/5etGG
iXgnbM4Rug8hJ3sFsSfgEAWFBXqWQUK9QzLBGbEets2V7/VLBaSXabpUDxRpJ6T+twfpGLg68ZnE
UTAX+dk2hJ95w4z4ThsLaUpdt0FZztjhcmcVTttUjnCOIm7LdQFnf034G2VdNqzXzJBTisVao/go
2JibpkLiAHhksZZw+bUnauyDjyJpulWxM9byfe4/f0vsRkbvXCrSQh1KQRqYiRvuzbuvYO4HNvAg
wwfS2Zj+qDDgwsWQVpt6JsgLwlRtdsKSk2+DRXUrwAFf8xRuON+dTbjeJVL8bounl8YFxjS0WLh8
nmwcSfqxN18jBvlhy7yssiSKsLwBAhGByBvB/m6GUtueXGjvJPRiUcfB34YP8WaEoUpoFLACa0mw
vNkmfDK+qK59N7QuoQhXpCAbSBiNRzCghGPyrYrwe5dvX2EOuAn7Rd67Idp0i6N5HUClT39cM336
KaLSp1n3VwDIuTvZPSJUPlXVUM9l27xeP3DuzJk0Qkabar84y/Hl21jeSSfvtmBkSbqR1h8s+8SZ
nXXveTOcKg7AnmzOBJdayt8k/07KjoFIZUT8JJuYkxdKNG1fTfON5Dus7CeUk4y6RLzmO7GU0R1Y
8r2ms66vg6mMRvaFvlyfVLC5gm414SD9xmIU6H1ZLWLGCLCMxc4t5zl5UazXF2ooY4dcWzekOKQ4
o4dXCVv3AnhGAcybDTuPmCcCDCb6cyJx2TgelSQx24Z3hD8NrZeZmxHc6Zit5ZGWY2I4+EBJOe7w
dby8Dr+emKb7LTLo5uIyHbqxet67m7OfeBC19qnsig3tpSve1IXtTnwWFzGVsoxss/uZNm6gw4Q8
LScYmb51rTIbfiUXUo5RCz4Pe3cXZsbEq7E5CClgeFEGtWOZdqy58jBq0IJNSEy7V49m
`protect end_protected
