`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Iexpss0RUTco+vyA3yLROwgO+5v2pur8nFSqf26kW6VeFH8kesWRABsxXJG5I5gHmzQftxOaBWZ2
miSdf7B87g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HsnSgo1Q+MPHRPOaf++RGMN68BSS9uOnshBY7CUnJqC92dBiAHJZX0m4yHJ+wp64ANU/dTku8DZp
0CUDHte3E/nzfzlOpAb4bScwr+4Re5vqM0f2wMRuxZqmHo01CRkWym+73Qp6ypM31hKK8D+omlDX
5KeoViww+8WNeEPvc/E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nauM+SrtCBUMbgauEPy6g8d+W+IciYPJvXUjn7MInGqG28UJ8n74bcGFeR4DyG21vWOegsM5ud2F
P1rKnkFwbZ6AbX4DXpdOCcfkBStGt7wpSWYCmiJC+tUMLji+aMnye3LcRjab4U0tyLZnLru5RhW3
L82Phu8ZZWSbA6JaTjpu9t6wdZbyZyRQnUflaIo87Ly6GKz7/4vGl6NwRw1fbbEePwpP5/XR8Dq4
Ou+LxBDj6LclKitvuqBhSacZZTsLTCyNIEsLjWvx0cxeeTVsfhrn+eVDh1Lt5KwZUdMhfPb/qgSS
4axJbfToBwFei/c1lPPAC1yMpmsVQto24L2kQA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wFyfrlxs8YewConRHCB10oL3SdlLIEEcfWkEF4ZGevncyMVW8dwA6oYPwlqz4A5zzU6PojTb3xVs
wr1eV1uriVpV9XT7errwMbIGqSWKfsroL9045b+ONh9RXvwWtvC3G5GBXQiNt/U+q9mQdt/m/4CN
1XrMbWrk77wKf3zuei4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tuQoLNj1IYFLAV6jKdU3j0zitXW5Rv218sCrB85sn/S9y3qgrKAEh+cCZSSr9fEfClQFY/tRvMAg
lMS4Ww/pau9q0kk4rtMaPaCLGHQQ1kYcB8liaKKkHSt5wITsTEsk3pcZEuKpj0Ozll5O9Qz3csqI
bxmUBjMOG/demQYN3N+OYd6aAVTDOA7HDG8g5l4mf0YSCBaQktGIR5J0MU+qL4KZ0hmu9NoAfeY9
zcjDtOXNUBGxhknRotWQShaEMbDZFXC5JYWj91rm8NyrcpX/eo+rLAzAenqwLyGoDThPW8+F1NKb
thPxfnA9Yde0TJo29YbZBRozuQOT+AkXhVLLKw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39344)
`protect data_block
r0wVjodx0/lASIwrSefnB3S8As/0z/LZYuD//jVMx03uXYM3BD6zptT1k3q4gs97m57+Y3JpgoiU
vXNM3VLd2t+l4tZw52J2b8rYtt7E3vWBafDv+YyEPD78Mjk/YaSq1YDaZZfodkBo+oh7C5quffnq
FuVIxQoqguQAgyrrNC3lbLMs0xsJa459Fg/6XtLW5OjWJJowXGz8TBZd2GHoplokg/drf42JJIvq
a3GGgYh7Ii24NNrsIyJ7qbsCU8PvX+RZ4KIckT8YTePWFh5BqWRG+fgkX1NS1c0rH8gacALPX/kx
EboIzDa57bkgIAv+2lXWesHDaoO7x8h/4nIfdUsjwBKB2laT7/bcBzxmV900DUIcy5hN1Kamq+wZ
bfz9dtFrKMW1lNqCKiSPApwax4AGe+MKCfKecmIVBeGm9uY+7kTxc/mqEXOjm/zzbz9dFiB7GIrF
lDnEPHynx+c1OEeUp5fvHgTkcTIF8a4hn9HzUVKWZWQJ/tmNNWc4mB00Zda+h3wdXYbwFI9dDs1t
wQOVI5LdN5G29gQ/SKFil3OftvtNq9qR8RoHD0Sv3w7DvkA/tYeg4rHkJSzynaE/FRwKgADq2xM9
sgr/Dv5Mez1g8MtAFad8K+VQEx98NavXtn4SdVQ+rZe5BpWzFnoTRTWDe8DrBz/RQOuJhiEeCatI
VKUjJYMrhe2lRshVCJoY3duywg8oKUvrOT1Q8KoezFwlWBUJWQxuy9AKygtTy+x2oxtvfdbxpsO3
byMMTkA77i1afx2HwrEBGK/d5045fPwpGxWQVshGu4RfkqOk//Q0ETnka5o1YMga78hirpveGGE/
WhFHUkj417Z0MFk2yYNJRrlr1dBZlB1OcAkX/ox0EZiARzvG2R4w/W+P+vPJOgo+kFr2fYHRfeNw
F/e2xhgi6TRMQqpmi2V58on3DfkEZ0pvAKFsyDIcQs1UnhRYp/BF3s8g4z4GPctF1zt6GcjMFp00
iVmP4FupwedARmm0LHRwB3wjgmcRx3KyUwfd04RhtAZyhxV/+mP+kiB04hP6OqFyltpQnQ/9v+sU
TVOjQBE5qxbCe3ewaLHWadGeKpOopJ3xVFj+BncNiExRsRVPJEUXQA7cedXNspaeTehslPXdkCwg
rlXpUxCp6gziwV7frA2BOPzSkX7DSHG7sn4C1EHhqs8rxOYIjVxUMz7Z+83M1BovLrCqLZegx2a5
kbbUa7dWTs4Nmalsf5MFf9n3k2dc+TM8sSI+8k0112gNDUuLM18bS2mEAG+2lsuypu/dswHwgiK3
EC3AUbMlbBQ6r/VPRUpgrxGb+a4AeY5sGTjkIK9AJ9+x8LsYiapU860WXUzo+KnzIEzY0Jr7vHXk
T+YTboasWdNdbHESknGQWdpNCmLWNhAhWJAlI735AdftkOE6LndqLtDSACYuUscr8AxR1iZLC+/1
/Dp0ZJ+h+HZDVXs1/YlLGcMWq5RWrGoUExTtSjltZgA/kRWTs5HiWQ6lVW0ANvflyjXWW3eXCivX
InLRRPjZC0FYwtyX+dsbcs1bVvL5h8+srCAVOR7qw80TGGnRgjVBJwtUdue8QZc+rNiqkr1WMjYQ
Dot4FYLjBX8KXKU0FwCfir1AglwpHBbq1ibfXQauU8SoPjfLoJojX454ixr5z+gKoBoGCo1BSLxV
Qnh1GM71La4P0O0/C7Dh3fUuBOzSM8l2PG1OLFcsvz4iySD05Y+suaDbZ+l5hdSIgZwT5WhlAaq/
QCVLe5wFERSU9D0890D8URF2zC/ZMtrm16aJGR8K8tTIGaALxmgUE7BYAejA5MfDBJZUkRbEpxpI
eUcXmDPhJqlmk/QzZdIZ1aaCDq++IhqCrFADTrXLfqbRmukY9t/pDc6zCvWovXqW9ZF5dRheFcgj
0UichBkjEnoLYMJ2aCDA51ypODPYO1X049kTcY2G6bXbr88J38ROGZdABaG5U1s2G0UYmLtYQmcD
81m7zwgTtVXQfyPXH7UBBnOGIKkT21TuAjaNqTrzaxa2KO9JXS1k8vuYSxJQ/u6N1kigLbDq9aFO
+q7+e/Nc5Y3ng3Tlv++GGtNhI2Dt72tDpknaMpbtZiDFeqFbCfTj75affwgranQjciK1RrCyoZYk
vfZKnQESgZo8huTyGpccGQeYsVsVvB6OKdTvy51a250RfEje5lBnBNfe0+kynqIiVmnIaSqdG5o9
gtArd08km20tI/sQceXTwr31Eh0UTdHpJQK0aFijNk2UKfNXEkoulc1kif37M4XW48ev2TYeg1+3
PBRA0W643b1XdyiKWY1GTwjrdmGApbZVUP+Tv3obsTAAPwCdObY32WBK5xwwh/qkBggAvMJwOQjv
d66Wv0R2nwZuggnVMFwHPY79ak3XFJprPDkPQuwiJoMjFpCBBD+PbbIzUg3EVvCzaQkSWJ+VdGgX
Kd6VKMclA/BYYVni+VW+BTta6p9a/1enaxOqYM1meC4IVehXnSmCiYp1ZpYojtwC9smHc8Y1sIMv
8LpyVDbpHJdlTOgHgxzw1rYzh/gDp2KsjfOWeZUsO+DgWzEV26x4JAuu3sDAxgyx5svTNXmaI5ta
EkxPwNzA5jR3xaUgh0OM95AdKRzQTOI56Ib/VqXNJUPBKaGe78pTVMVcMgHv0p89F843zmbKIYoT
HGNrtMx20DtXRCbgaZBge30c2mzNPXwehN7iz2tEfUKw1EGY5OPn3A4Jk3IioefZOomxrS7TlsGZ
kVxmAU4Se/4PfB7+aJMWuwHOyG0XYFWyDlTgSVhyVve7CDYXemW2CiPsfmq+EFVVHdaUgZl0oW/o
ltxcYy1Eh01Dp/1uo3ZSPbqY0+oboPJgsmF31aNoxchxPpYEj6YDD5tx2ImK6QH6YEhR9E5bEl2a
cptoW2G/Civ1Zz3GL0+fp7x1KwsGJElOJ/fJCtBo3OXsGkq6aVIb340ZmovZ3nI8rZ99DC+hGMRP
AtkgLkcOsJEEeBtD9bdW48i4PNaf8T3pVpgFZH5bg10PFA+BLFDIcFWXJbsWPepD2+J+R71D2Q9t
dXAud7r1tQNRrfa/exfm00cNjCCHNfc43pojL08FGvaH4cGbot9mHpmXRVZdJx/e3w7As1GYkYrz
uGzKsanjS1rmYWZJqbvphtY/e1/knQj/Q6z4GqDWXBc9NrcplATRcVLp5/q/zS0B5JPLGOSnKmJA
RwHAw2DF+NN8Wk1U53GRm4kAXQB06Ceo9o3wt5MY38eMycOzRaPYMlddMyevOqE7uoQQntN+6wUp
OGR5nrCCEs9TqPj5dAYJIbDbPMMmTEnrIlnsquhiVWwthmAq6dQH9V6b1S0+qLOjEoTaxnPAY8zm
/gTyS4l4vAqK+eTByHBb5fjNjLaoWOIIRlumOZqDgQK/Ob7aUfHoMwDnpuTKt7tlywWLQTVJFZPz
tH1cQSNLAPUDV9/if1yNAhfRnPR0m9duZyAgbPmlXb9JArzffo9MVHxOyhRueXEf274yJ54/KLbZ
QLHWZQRbZ6fRrQNdE9NMm3xq4f7on9YJIZP2Iw6zrBwqaMdSeHCYYbnW8fVEuKX0XLSmQIx/UEc0
tQzJoYusjsHbDcOjldLHfcdiy4MY4wWdvb3NgBvn+1nYmQTmGv/XF7o8GYu4oRpGEKgDs44oN/pZ
o7CTq8GiyU+ltcIn/isuaFiJ6wi7wXyif+graTMwrAi20ZkhH+W1N41eOLtIAVVOslkDeMC75lcy
l5sTfpoop1X06YjgWxhY0WWEzrEE5qkuHOwOgkYEo/n85dda/nJL0xcT0vgHh/JpzhgfZj3JkPQe
yBg7lsqRQr8FUzmuKOJNx96FcInhK/izFY7dSaV6tPniPCab/kQgKaDg2LlC78Q8IUNP0Oc7rk/l
ve44k20pIje6CXfBjmrfzPGZ1f095OYPYsKNVgT/ocvsr+AGIpOtcWWPzlxZji51aacoXaJOqv9C
o/3MVbUWjaes9Uj1b86/C7HddY+XjtC6NtZpKaUs6nf6r9jlmq7FHs7nGP3G6z2vi2R2xymtZvlk
lb/DmuCbXsEApu8GOShVmPonXVcECvq1CrRM0lgKUmTKl0IUstzx1qoN654luP1K3l0MkHdMnDWM
pzvs3CAP477wQkPHcQNSASiW+pmB+pnuC9if0jEUA281gHQe6YbP9JtKVU5pdS1pBjHYmEYFTuTn
GMZLFJGDLEEPfRbx2Qtb6miTohrGuVlYQ9iwXbyP6kscJTzxUCs944rSdca0dB4wEtHJWdsYfyuo
zr1CcYyU9QwGWiH4HfBPdI241nzQZqLi2sC/goEhIQSMjzlihY8HvjCBB2w08Y624g1X5lGzBU6s
D1PMTIH/WLUAhFa+lFyhN0BzvR0eWnq1YMx7Jipd8ir8qv85xHTa3VxmUpDj3DvRGG+5tObxHfOJ
rXrQABLaeXfPj7YFiju2beGDs4XQ/Af8fOXZJSXnDB/OfCECcaW5qVmoOko1Qrx9Rxxs9BdGKjEp
c9/zpl+XvTTRy1pTxgxuuI0dTWoWocDp80IJzKxVeyKrzIktDWvnrdmqa20zY/LTACATE0l8d6Hq
s37Nsy4MBTbGiGB0ZoV6Chl0Ol0uLAYQCw7SaSeBLKy/EqJqqYY88QBB9KIFnIBB0tlhfvuk+jlp
mJbWuhn15HHDKr5Sxsse0EVVZeHetEF0E4rSrfujTcfgTvwQQgQjW2VlTW9QM9KalW3U86zas0L4
A1cWWy8nFuxADCn+b5O97bWTyiZi34QGPF/l+dX9y4xLr46fUdmWAs3GgvK1fWBbmUFja2VvXDVP
v9mq1OyufNiuzJURVi1vWMPmll04bT1437AGVG2mooOXmWydys4hTvgaO5jB3Pp/6kg7fZmLmxya
NvY1M8nQscNg1w6i19mUmINJYXfo4PCNB5AdTqyx600SQhLi1YR8CM4nCCqw3KQdM8eGOS5Busbq
FJHBjByYbDUuBHaU7oS6kLP1Rh9xR5aYVtURKOOEtcVfshTxZwxJrEbSNJiQejpK217UvYwzC4qZ
ChJoeLSq8miUYNA7uRlBhsaIw3kdqH5mXS8olC6rJIjg1jOYEWpkM2Hv0Ec0HomYeFVZSzR6rCrr
0LlrbVdhS/rCxOueIenLDfXLx6dZJDcUqkDK1vod0J/iWBsRNE8Xm0RgRXFRhKm1uBVTq3WtW0Ho
EzGC3JvB2nwRH3NDuqFLtWjsA0iScGHCulwBAE1LkS6ITF0hI8H92IuuCjfN8b5QRMr5KNPcmkT1
izy0ZCTrjytuhlL9wOJj7TeChmblw7sVBXulpYPmCinMjcu8XJ8GC3gC8owrZ7pk4434BU4tCRJu
oUqIbhWJ5buRFTF/Cj/k3BJK3QQBGabUd2yD8D9Y81qEMIZbLwRPueYfGRUYm0IT7+fiEcqW2brM
7eqpQITIlZ0inB7oMyibNgnJ886Ky4j1XLt5QIz6WWa/rHZs8x1ihkCycP5v4J22mxQH7hjMW1/b
torZTxHBfCQ5Nsp0mprpbbs97fxo2iEsTlcjul1JvpHjsv0ozlXgZwmHfz0ZiNML+QG7tHbpK0o1
A7SAtOKSh6+bwmiBs1dWSr2/nT18Fk/L1X+983OnMoQ5DCf+Z/4Qe/RQtTexSeH7mKdsZbSWDz7k
/FsT2uLHuJ+1MRHB0yxFmhv6vRAOU8xSRQv+/h8NmLf5gz60djMV2MtIV35T04FoAKilDinMRawt
zKXzFN1cSmQBd0Powmen02NLfcikD4oGU3GLmkH9OkvptOgisxPrPjoJoQd5er4Mk5em+6GPOUhG
pytxgYjQbH/08/CWvjBtTIzn2gRveGmvlcweaOXUfOV1wE8gUzLUXfrZe+DG+cbnucSDW31l0Zyn
20lVOUbBHbFsV/1+LdRlqBkztw2Tp8a4mHvkJsUrb0C2sLHN9b1h1QaWlkO/L3OkZD6IUIE7t7ok
J5aGnK1XY5962XbtF9IGNape29MzajTmsuzh9YxG9oo1bvpIuIhj8yi8YuIR4we+qXX1Y86HdIXV
hPftjAGIyJtka+eMahpUQnLJhj53cr9WlTU3PNBAcl6LQYSd1eK+W5BZ+YkgV9g5u2UxMTYZhHmC
wYPm7HslCRu6BP1Br8wDnnDWmTRAfph5jxudU+O+WUBKa5Yr4WJzc553Z+HemmZ1SQ8mU9Ntw3AM
l9+krEoks26EOKMW9vWF/3FACfCJepQeoimz6e/0SZB2x+fo4EG2SFnUypep3o6bZ/lyUMJTDr20
VOsoPoqWO2bUPTgcBuZAhbAF36yke00Ga9qEOqBb01pToM3QrB7h4zR57IKWgUWprnLlWJxU3tzq
g56y9atUyhWtOXQASsoGPlIb7LTcEVTAnF4uJywnIxpEasQIjTp3ru9djVZj0omvVTKxzM36XE5R
Q463n1EdNXWplaOYR5FQiihUvnmHz/cFoME4sqH8s7hLZXFkG2T9DB/dsbwBJKEb8kW10R5zZT3D
0+8vSFctIPgwav40simQzgPtpyALi/aT/s6bZTtudA6U+JbW5E/adkEkDRZ9mfqC3E2qcdAJ1z7L
S4supryaBw6nkNEjMRXprZXjCe9fIWTvfUgJbXU6hl3Cm/fDlT3TddBHR5Zxe3cZtg3Uqer/yRB4
qDqOCUJbUi2vz3zdIt3QjBdNNBUuTgUoH8hzkWgGJcyGiL/TTmRQQOZpww6rvxix9BJ8Z3Y1r2nH
y9LHtVyaxz7GsyG5CmLxSezf6WvnWUtVugWfqdUfwpARC2wzwRnodSTahaIc9//HUFmZnSO6pj8m
5L0WR6EP9LLE3KxG/awoAiM9OJ/kUrovTkp4MUvkGPuOITbvSDMuz6zUuQJesQ0xWv/5+5kP2js+
0cMUXcOolxHSX3m1oOV2xSKeBcdiATaF1sH6m0YVq/5eT+yCKoJMvDOQNhewcLDSsi5H4M/39zpm
JQKF/LRYeb4J08WpXnvvscygnMrUxS2h+y3fG8XGW1OofYhCjcu+M886gq8vCwXrp0Ayo0nTbNhG
HB/UYSd4i7sVy0c1UoYMLMH8yxaJUWhMz8pwZTpJriXEL7IoGICRwzD/M9m8O2t/zUOCXNjt9pdt
+ZiQdqJ8Ry3fBZbp1c7jfyxInUy0RMiVDTZjl3mJA9dx/7dvqvoyWGnGWF5hvqxnm1aDyT+pHwuj
XV3YiwpfrNvhwqN9PfgpOHR+x2Wi5Nv1WzAbQADLCNkVmFl31G4HqrzDVXDHHfBfom/oyECLS2zM
yB/moMmMErERrWsAKtDsUVWn1UQsUBCL7UnjgWZ2+hpcHcVS1aFeOrwrq8Aq3sfs5cEXrw7YxkQO
AtQoCd0CMD3QJ6+OV4hPNIfRirXxsRLP3rfqbyiJbh+XbSCnL3KHT6GHXPtA6x8tffb1LWz3DChM
B8cSn0WMNHDXyAwOWaGFQzoYY0zQFjQHM+NWM0FAbuCcxGw4tHFPiKI7JCaq37N2VzZBuc3cwZaN
LF6pW8bc2pdlpN5zbtKG3PKG9WNRKIByUddkadhUtIS1LIAUj1XyQfsvQdPoSP6cteGy8Ph+BJ/n
uZpz/ZGkBjFypWBwHOgf/X7sydR9NX5j5Uftyc/wCyz8T4wH1l4hQvnOAwiZbohslG3xGQUio/m7
ov/Lvofk/z7VOQhQrRglRapgnRH+ZhR8aSFn6IqtUQxyf3gEibIG0iVhutidA0sMkCdPdnGNMSGK
3eLuhUrBEfWN71nu+jWCQqsvl3akwkPyqxD8u1oPnX8l0cO3nGgyeGW/J/WPDQcFsJh3gDxNN3Nv
eOlL73AuUjMcgzV0Tjr0lfxVCGxT/ohwDAzULx9P5miPwg9ZdttiT1crnZBG33B+0hIQplrVwFOa
6u5XpLvfO8TY5rdFktqhvVKevg5J4t9mTAbXTLW3r18cp/aAU3b/UEmePe+PWr959w14ehjSzafM
jN8LYEpSEp2yVHK1Og3YKak8/yfYDmVMZx3OtGTGTlIjmEFTZjaXQs9FZ09S1F2ZAS0kz5RDCel6
b+h9nueMiyX8rBHiJAjoxZnNp6JaFGGFwfNcXZWgsj+ABynP8Ft+1hTaFGpoi4NJ1khyo5kdZ1dd
kiJGOnK/JkKWnoMBT2yv/4r9uJUmjbL/L6Bc9vxAgWaU3FGdCO/sYd8zTePANCy7RdDwtgun6BMU
T5v+fW8V0pPtQTisuRZp/aCQr0LCp5jiG27c0+U0tnW3DvMPBgjP62KFWX8yWbvlJCk1SE3VsLtv
IT9gqlMCVf5fAVBWctCRFN/5xv7Gr7hiLjlGxno8igjsoY3GWY2JbKisi+WCE844ghuHqRIQ5cgW
qntOz3HHox1zZpDFiYNUk/Tl5JD/cPTuPdhMht8ya2hlxBYNf+SotxDQ9kHMVdFmMprUVhiznm0L
xGIHEVwmIzxfQM+SNyAZvjCyWjxZcnA/ApwoU8VPAH1OOOB7EzZeRHmE66M7MlDVBrCKn1Nam6VD
N6SEbQP++jEEtIVnE5drVCr5VEOBfZwOYPaRzyACDCUeQEJzDgBBGZBhcKZ1HLcbVBibuKu+I72i
19inO2wKFzVGE2H7Wph9+A5wkQuTS7rdpTOkKi2kKEtd6cDfqxEg340s7XWfD0ZDldDb+S1hUt8i
Z/LBgyF3zqdQdUcfTazebWIoWP2YQGFdrgKfhhasPWkqEaiidvTG5PgoCe5prsyQD8Ys7eQFvc10
2XUqFCHKlF1kHqLfxhpf93/vfMu0dnMzO/cY9xPSt66BSCOkNY1mqfDMN6rpONkyeNh9TQka7KMR
pnnDsylAINKRQ8m5Z7oe5ebE5SrcSWcXt/+DVkxv73rgPC5wuVKierUF/BA2koaIxuV5r/3sK9Po
PIYfZglAb0b+jHnb3Rv/xvG3dUNjjl78mtEPoP64p8Du5GUvT/pF7Rw9ZuxnX7WOH4j/eGbIDNIv
+SDECRwj+vzTPBflvZ3Q8ErBkirL9N1CMC6b4pvy+tVYQD3qVsXVfwc4gokDLLyxP+4JLHwlLrcd
Flu2YcorC9WyZnxmmnI2GRYZcPlh/8zyub+xqwhPXqACbrQg9VhAfD3c3wsje4nIuNUuEWbGtglV
vi4Z3reIUMsSuWI2YNc0mmQTD/S5n5IAJJ5BdnWgMCwPE+lMN9GBEtIywUCIZ0ukgvDwC9fNC9aD
gcf/WzvNQPncmTXVfIVQ1ki8J2hSAz/dbcEeteI4meLlzA7QUzNssHx89LMH9bVHD6nuSwf550mO
M9bpr0xK/9GqoGsShoY3FG4WW7FmMrkJ5Kj7nPzy5bo4FOqqAKA1EOhgZ8RcJf8Z7yJTx+mG8k03
9vgP84F3HopwCRH6lzpUy81cOskej+Jy1+f7ZyIAuyAoIDtYOG7bG7js9lgANpJFfXsXza1lKisY
vX3fhWW/ym+PB5Tnz96EmIZ5EqW2XtnUPbArTdqybbADoga8ScPkXBQSPWkj0glXrND51bA/SuXb
wE2zkT6YDrNhIgF6Xl0/US1LmfYoLJ0n0mADWHLk7nNSTTmoAW5jGvtr/eg8waUb33dgFUzM7BGV
XdB6tFtYGfzFZv8f1a4M910O8Xbsno82qlLt8QGfIyBdlUd6lxC/LApUhQyKf6PpOo2HjzkG/2Oy
GtDwiRylauA4nVXnYBafiDuAfcIZLnlVH76PU2xGuI83L7R8ZnruQL47gNmUZvZa4/+E/C1tKR/h
UKeI4MQkRs91UFjVoJUldWLE+E4FthUkFp3bVbBjHKSzD2/3cy/FhCbmZQaWfY4pWUbQXRjXmPeW
5aaFIDkxET6I6eONPbbJCnNNpHE5tTanxhQo9LEGeX/BlNYeI/X/BAPKgyRDr59YYB+SK+OlVxyy
QYSl2kMhtMV6colE2zrRoM8DtgkPT4SELafQidsNfwW+lwQ/2v4vsa+EqpY10PL9ka3QWmYMtTJu
RsrMvGEG8WbwGG892h2VVvRGNK3XKOA8L4+o3qD4zF0dyjSMR2vtRBvt4IacpCRECFqGUNTPpVXS
G/jnOxJ5cQYt5usYA/zDwuds3CF8USCcuvfuuxW1ExNPW5nfzUwqmd9UQkSyQMoGBl4U4BgbFBOJ
tG50sNAUec1pFc2tjmtcaqiKTc9T2K0r5PRCZDqeoi1sxKezfzfbvJCOXxg570/V1PmqGMk3Ojj4
hnZuBmzhMPQ18Ev0Ns5z6Gtqhjao2dMEgZLsGmbfYh93ImVRB9bLeiYa48XrmOgz4S7TUh9eldWh
ZB1q2i3T7tqNJYKAYuniF2q11NlwVCOULfTbLwaJ8syphGId0SzPf850VW/YMB9OG1omxY+oRGS/
EJi4k/YZfg6euyUBbxIuphJmYsr3FL1YviYM7PLBgRiDD08ePHyjgM6kIcbkC2sVi8MLVjBiMIdq
enCV77WB4RinrdAXzCj4RoSnI6z5zZ/Mmdn01fJj9TYtm35zDDMHBsMtXOwpFTZpoL+ZC/Qzpjn1
knxUZLKKxy3OXr/2pEomkQ838N6uQRec0Z8urUqK5vDn5epM+VUPqF8+b+ME68l9nAD8bXYrayFr
+vVhqYl545DmNjkNwkIS27BVo1utup5cplUmWXCX+qAsWbZS34pND/CXS/q1IAmkaED0QmJ10VJB
v9emzx9g41fQPA2JPkqoGoaPETuu0ip/NGEBKjxZ+PNpYDQhlgQFtUtv4KfALaXvezj62LJyPMuK
FwUwv3RAGyOWlgZ5EZiJACZXtritKHkSy/i3VSWphbTQ/TCwFutD9cfyryf6tmHC6c5Ld2jVhKh8
oKC26bQr4nUafkh469VcogYX3vH1hCCmc4OX/gQRhAOZqsQkbq6ziV78mWj6SGgaxSV77YVQcQXN
AwY+QK4j4DZ78Yl7OBCDiHNh97RmvwIkf0IcA1qS/vGCbI4M6MVOBA6KL9KVOZXJJ3U/8/ThaZpR
aAP2QXFC8tpLhP2VU3Ueg1jwf5ObUDrNwT+8NHpM4z8RXiHcnhmfGYUW484nMYVLpyUwX7UtgFhz
U17SD3U7gxS+3MZWN9+xjGCpKjOkxEp61W53JqMW9qoqFP5oZ80VS4uQK8MobOJl30CXJigfLewA
hHhDSLYxuWHGqHCUyTHREsgPTtP4rrdiwukXaj90UgyDj3OKv68vEsv4y89nu7w40/ULmIwffhPL
qO4G+lAyfLh/+uXop9bdeXwqVw02Uvv0RxKpxsWs9oP01UHdPFGWnO2xouSinhq4bBLa4Cx8dN/W
Mo5zCAxOQQAHUtYv7JAT3RXefSMeC2GKlSReZWxaeQ8jAsaT8JI7nse9nbm1cpBJBPmx18e7HM/y
uou9+nkbokXvQMPmWoZdgX2+S2+rOZjtfrq5Cv7EYXSed0yUL1Vc1WoQ/+piDgX+qtaoSiwYrhJ1
tVT3ANcSU9LxcAgmAiKPwjYiktT32QyyiRJ5653U6FYeq1YkHurQRBFkYs4lKW/26F0qP43Z2Dx9
TYNagrROOJe2ZjYKhpus/VuJNAK6l+Y8xGf7MBdIQLvxiQx7flwCDzDqdX8HlPabR9L/3jHan4ZL
LyZmxIbdGCk3CdoScnOD2B6W+GD73+oNR0fB9T1ghYjqcnB0wSmiLy0w901QxCtNc72ik4A4WC1/
nb9OONzR1qbT0a2WDn1fSyq2IQaG43Rl9P6y0D0tyhgSSfo9hVirgfYemAYt19xjNMjUruoen2ut
1n/wUbyroddfqkQtuqvBCqfXxpCmpn83x91fbI+s35Pi5RSEGIN8mTuAjucjRmqDqMyACNe+RF0T
Mt5ktuC1eTygK4Fe+1ymtBWS2yp3fF3EdFEEmuyCZA2KHsf33034YU2+FDhdONptN3ReXkqcC4/l
qV5N3IgtKKDgVoZPOCEtucPMV8tH+ZI1YHwTVkQqSObUfK8ZBUx5FRU/jU9CkUMj9fouXdmr0nUK
Dte+0/0/4Nm9dwiCtaj1++hCC/zrmqh/ph8ILuo4QPPX+fp/l5v2zHjSc7egTdFowlWqzX6y7Dnq
IwG4wm9wcP3fbSqQNdABit+eqJDSg7ySbUx0ixFrCs0v0/geyi/YCaOcJsmatKE+wzr5MqYqTNKA
P6+v4SoNmggfzpnQKYHTWPqygdLLcM+nVXiBDMaOa8iEDe7c/oMycfvLPrKcFqT2Hm8MXUZ+Suxf
FRF4kLPaVuIwNhHWoRyL+Uv1+VAtIFPZeoAL538ywJ8ds0Dv9dUMX/sJpzKijqtw274B+fL++2vh
XtMWIvYoBJ5K52XtM+Fuq8GU9ZM0grw7IGMRSeB+wf+Zs5AKjsGPwpoCYFC8KBEL6F85Dq8ZW7Oi
MQ1axiOV3gXDYcvClZLKQIuqdFluop/6WKOyTZHCQohzx+a6VXD1WiAM91CP5BIp/pXJADwvENPT
VP2JWbND7iKVQKeWLdTreMex7oUolN5pE5KTZI1TcG99U984bJnviEEBHmfEpkZsJ4EJi7rcOxpz
x9RbzZJxh+RB6J3yeFe1wQYjdZUE99E1HUhVX0YypDmDtg2k49UN4UQZ97IVJdhPKQdaZaznXOr/
ZEG2HJHZq3mEiLsWbcA8na1zqgP936UBUNAZQc1K7bjhfGaKOBp/NDaySWr1MgyVD88RNb+utiGB
acG+Kfdbm55DsOpsq381qeUvXCrkGc7LI2lL44AjvAFZfni88BUSnhfCdlZy+ToVYER0WYUMIczQ
/4swefadaFNseIqyQcrXWT6/SI1Tcg2sGqfB9GxFl4SuNoEi1ENL8TYCaIhnXeUx1VS3sIOgn8bk
qRTJxL/OeU3LP24QlTonq08LWHPUSGWPQzj0hp0H2o4IULum5CrBKOARU6jQBIoZdYWu9dmjte2t
hgitYj+K/OTmn+lCArzDE0MDIo3DOLzinhYfDeTLBeJGm9Z1AR3Izn+2IQqrOalNkpmQfaadcFhg
Dzo8u5sRLqQCj4Jlgnx1Il64ragCaIUYjrcbrCqJE7YhL7QCHNCh56n6lj7KuZoMmrj0o/RPpx+A
AHLin86QHJvY+5tTE+5IXA8lw1V2TgR9rVVbA7xFYAt96LPeG/fo6ctyykBNeT7oq+J9E76ogXBt
ugm0ImvxXv4+ep4QYvKFNpnvtOR7EL6pUCzD5T6MHEvj8NGr2YsPpzy0r7ZnLW+xaOrzL73gMq0I
Ky2nT22iJtJf/Sel6sgqZdWkQeGBIeWQ1orNbOxX7IgamJlEqk3sLiBaG3hTpoZb/v8FDtqmxOVF
g17gj4+ChJLSqoWbt8HGt2VI+PkAkmlQpWe6jThb7lAzU1TVyVJ5725pd3qOLAOtLLdgWqc0YLzy
/hdOIwTbmgrGJc9jQ44AjsOJuPlzyjgJ+gqfAS8Vm4iYXlLKe8fEp+RjmbkHCJD0f3uo+8jUS+dt
ds9h8qR0i4WwIv0QSoOIKtJr9JLflOWTwleSfEIFp4YSqxD+qWuePCPnGuqPtaCZwX1ZGyJihTC6
j32iQPhBdtha6g00dahIwBN7sBoOGynWhZKTwQSN0IibbegaXL9SudeC29SfUVPX8bCCLvW4Vh/o
jnFPWT4JdvnTO4a7OKj+2veoP15iuUmAN6suu0PnZ7E/REsc5tOqqarGvbPWpvNVFYc+ftAACmLi
JL97PhlULBfK3sIofEITSMD9FEtpuQqR4RHh4FUB/qo9+fUt9Spyt4Zpo5680Jf2I5vJB+KBkvof
caoQwqjOOgM1W6ljCwE7RBpe8+ouJla0n+Wc2IRdHWrllY9M0W2Gms0Kim6c/mRX1VoBlZyIkwn3
OI/YWSgQiJON/8NasEvvR5qZ538vVm6XIOjqIycVpXyER/sxejywW1t8+JXhK6cEljkoUoqP0oKK
lKdCtWYrngokhc0ON5IPwdS9C6Pui6dHWGbg65pfyxG5BI/+xPYjTW95X4t8s3ruwmAm9Zd6vhn1
3/oWWSoa/qc2jqhm/SlWBfZKG/v4qdqSWhxHb6hEXn1V69vB8Qtf/QoVuuVgyo+2Ghco4z2IGkMj
gSW3lgvShAqX9YdWs50vLEWerR7G2LYzKkGYrMmVEv2ESGShymFuVIhRdUzMBeuI3BFgIMKwbgtZ
kokzKrc1s4Y3DNaih1FpzsD+j8mCsWAADt5kjZJiAUuy/zogqRtoCym/REZVIHA1s/6oF32yszp3
myLwgwZsfiDh5glv0q3HZv046QXCaWCvCBq0vN6BnpGDLgZ0q/afElTVaiPnPHKI3bSP67a75SV4
qg9xaRYvp4e3kKD5yHo/zft3/xMnJB8PtspDOOb1uRvXduwEwQKYhlMe00Tk8q/HJM3IpYWlpuc5
+SuHOGIkYKoQeb1f0YwQ2Ca5w7oj3sDPFv83QpTo4bbpSo41a2VlCjRGnBn+x3Yxbz0lGzJvo6Ge
JuiyEsok9xuh4IqdDjbicmhLvQwIrCIC5YDKK5k1gBgW4sz56ap5NfPFDcVEX33nLJOf3mBq36ZV
b+b62k476GyjTAneP++0Z/OOIPL0x6RrZt1n9bDilLNgQwT0yZ3Ft+cZsky7Wjfz5iSicH9D1lmA
Lnp13kx5twW/MV8jJYoaE/2Z9vy2hOt7AsQvBcvb0H11MPZJigC5RzIZzxIyjxgZ3QXCmjrwmhzM
iGEPyksAM/tseP6kYlVZoP6k3aL+baptc+e197v90iNLRoGhrEzrqs2lgnBKAyi4iVvefLaVvtqk
DyoVpOJ8v5YpsC3Un3lJG++po1hQprbNnVcG+81RsTVzkRHVpVBi7skxPZpQubjTBg83UzH8u5N+
LwT5hHT5kxxSaIz5EA8N++wr9kJkNOra9VPHzb+24WP2738LhRY4rJFD7VN9FBiKP0nPNDLw4Ehc
Ktka1QWt/afYDvYDSf+z3v4pQm6Aiyv7kb7cdUyATXtJurVRJ1cu3Vw3BIP+c2+HupqM7fkYod7/
128tK7A4JVMYsJ+qukZn6ZTLKUOKuyFXtQEtOqQNrFRrXj4xZ9DantIiUejqpHC1R2Zzqj/k3+/9
CSYtwrdyOjgid3kR6mQSI+H5cUKdj0BpqD+T9FuounWK52YncXdcrhXrIxMrjw8IAmLRJxn74WE0
NCNPzyvk2s6UoW79OSMv2FK5+q+7MEoycYESCtiYt9glIW6jh63D3+9CXrlRboWBeubWtidM4/Xf
A8G2SaSsmmVbWq7eFeVuKmPVX4dOGTjSv6KLKHCqsirhv2LJMEOqEsX9JNqlaTxmmcgaEmZ/FfH2
zzRVSyhKsMA2kzBnbE4H9ZiEUZU6T4G9QxTEKkyefoQ5LTXsAlvJznGdKoUXEO5o2STKIRKT0oC6
Y1UFv7I0UblJiqKi+qQvl7Qh2KW1TSvpmei7wkDb0OAFzhkZw9hIexfej9nFjWpASAt1Lp3o9JJK
/9O3IEWSqtfbQd5eMJZdXeuz9gOiaIJhFF0HBqHve66kTcaMAONYjH9Hi/Jzh3+rDvNTBB3t/4vR
tCpBU2UdoMH0iKeZYaQNbtkfBkMLFcOS27Au11TrL27SSfBGS+lHKuVCvDm4L5QYzpdWpa6e62L6
ny9gALxft88Y/WmDma44+LHYS5lVPocFdjD/xGELTpLv0ApaDchytVKBfYaLO3YANQ9RiW4q1mJ4
qcuTig69lf10jkco5jtWPj0tMmC8jYoRi6sabEkbYLfmNKuvnALCZMjv7NHhv/iQmdyP6i+AoD6o
H5sajaLEbBvv85XCKLTZl0sk9aiTVD+TUURiH9a6fZ/Bzuv7hGeBGdx50mgriD8GfGZSNfBOcxao
sMTTYPi2OmPlnttOyMIUSJ2JQA3CHG02lwx+uRDhtPrsocJS4SM3SMj69rvWham8he906pCHUHsM
iVd4zq5mqeQy19nqPZ6LuRAHwd/QTxo6f4DPapb/Q8VERVmNMJVoSNxiOkpcgW6GjUf1lRcnkqvI
nmfbADsZa919sVSHY1/Xsv6Ppdzb+JRbVsrFVoMmMBrvdeCzhql+uSm1eGbg1ACMcktsXo3qc6mI
m2Hw6EIEUBjTlwkWOojYFLjEvYk1CzCjOmVrfmSGKumDxKHx76Xi6Vgkels6WmF6WIKvqAz1i/rg
UxjI6StIccegVlNktpxzkx61Ud8IrXK/ZTjxj20aPiMG0SlZogGl6O+og276NZxV0mYMa3OXe/wA
NrEXIZF2c+pfwS/pEWP9KwD36obaYxpYcfd1h5SW/k/22c4P5FRvVx98zCDBoswl4O5JjKTXcckx
X9mz8TRbPlD/y0FBzuhuCvRrIRMOKD0THl9a5y0G9V79niXN5XNZTLtx1+EgUKgbgUSCa01/vrOk
ZzExiGsYIILOMiEWPKxPiC62+5sylyRBDkQSAOnhb06ck5jmbMO0DbLpCHQBQaDmjDdiz/VJ9Nuw
FULCyeMG5s9g92+bAsV22DPa+2QrQPwZD+nLOAXbFbAN0i3FfAqfV8rKKAnI4k3q4t79tqOFyXai
TTHly+BnT8s7/G3+jVWMSLk9btn/+hgmeVQrUJ6kRwm9zDdKZUXgbtPGAUKdjIErHxhmIgnCcfzR
1un17qBKA1BpGkoL838xOR1IOxobxeHTOUCkQbsh3vpn8tluD0vjH1AwYTUNt0B99+2VUK/k7qwj
QkL1wy6DKU80REMzgoE/AsCI/1ZH5HkEwfLl0RqMQP4Vj8IptmXB1zbeTtawoBCOoaeMBO6kK1Jr
hDhYChRHd0K/klfleBE2rO7rfbZAMpEtG7h1h/blg86akjE9nwuMD5SOtGIH6D4zcDRkT/0iWHQE
YuBPSGUnXhOCQKZTqr+tE0/e0/0yF0AsDItpZJC7TXsLLhS7qZ7Ii46Ch7O88Rpnxt6B8J+GZhFF
e7cNhO2r7yEkbgKiMI+6d3j7aIYP9lj4vzc6p/OhFVjNUvN1h4/5sJDCEMMrw9MqCUWj+iW8Wugp
NfpYqVTzuZlrVk8L4mHf6Uze5PJ2AjtW5TV6qyDUYTMboqY6wYCZvQYQN6+I9lp0zKJCWhpUhxAK
rWzvqLHSOs380+0oA3VVVQ7U7W+NDbIX3K6v/YkrbNXztNNb+IrtWA8RNGH/0uHiw/gYEnVAXcRR
E/sLFG/R1ggHUFbEJepSwk6sBFL77mjwNQ9pZT7L0J6Yl44PNRUZ372w1vstOTJSt3WaGPxuGvZf
TJAP1DnrbZ4C3CCDCzCSNS9vLIkaumU2OulhVvMIVwchhtQvGAeuxVVhjaCeYpiY36tLOv3GEzYf
cONDt4lIiZX/aGEkZVQj3uRsK3Vv7UgJJTB7RPNf1vfZaHo1zRkzHhuChv45TitK8PpN6FfylTbC
l4cI+HU97DXObgf6ASQH4v9su8ETC9t3qeEKAy0TPdTB+gJ8uHq+DRcxGfM2PoePn4c9Q6FSMvPh
Wy9dS5GXLsHsvy0MejBGMv+mzdrGr1uzG8O+ofn45KHFWesQarIkSruKm4tVf8e/rwaV3unV9s6M
s9fK7FZvLSbybRm53Uq1vJtZC79MdI04MRsZrQN4RFA6rk8UC9D0J9HZOKG65aBcr0rJkpA0qYH2
+2Hx0qmX+mNwjEqhB5whLZ82QG0bw8IZ9Uuu099rzXebDuExNIss3XLmv/sDgu5tR9Vhm07iCPJp
/5OQEfum5CFW13UpODnDL1pwpUu6CHfZFVRsNKY7E9k5M043bLaqe6SQRKzX4SKDiSDX60dIpXGf
TXHXIID+NXBHrL2uT08aXrKraAipcNMfdOX1KyDoX6SfB/2NFnE3hzA27KeW1MpBJ31oOtU0c/Jv
TWCM0Zoo132bvgzrpGDyk8GiWS/x8T2euxp1vE1Ik5yS394jLrLfTjyDw4hXAQsCezfzAxeQa5be
4Zz4ZqgMswmqiGVucFB2ibvQvcmHOvMZE4HfcH7zvq8JJI9wQhQzJ1ulzbimQYZmZ8FTWW5CgdmY
o79hfF3WnxsYxklSRwzg217PPpUKSNxCI6SeLWUnOSjY4okD208fkk4IAOB2/HUlNys4q3r7lZD3
QI/Mv91sBnZBfXwoN6C8Y3R5YMfFWTW+lPM6pL+6OWvWc7y6H73oEOxSvcW0ALpF/wJs88vYgS7I
/FNqBGZ8iTtVu7vy5wHMSRFbZlIbZtYbtgpV5PkDRS9DZXaKNskZpgUTs8YvepBXqoQYegGYvny0
cNjiRFMPK2HcJwM04dS0v0PFl+gVgirF/B5apWwslsEVbCK3lXTaWr8TfZYP8jFicBcZR1XI8mX7
sImxx26DGFjZwmjIeP/AGIGbX5oOr9OK4iwm6w9KvttmPVDz1WoXJz78Fzo4ZrifF6NuZ6rc2aZ6
fIktf4sKE9gIIUPJPKUm+SBqvZ20gPzQzEvMLh990Hz037h2IR8Q8gTs9olsIPBMZMIQfNRuzw3B
NFoXOGQ3he+O6I7O3E8p6rkW+A55BcCtd3Lh2bP05xNETL26hHD6E+0yhLWA1xmJvI54xpX+NIAl
5YQETrtUMcCmMevwY+LXMtil5exkPbk52Jtz+s13JpHc/zL5CchLoKFPmqCGYhL1u60ttTSX8lKF
++SJnUZt/pSfILoFJm/siHMIEn90RUTuYjMDPmiHnlh3yy0fM2kju6FHn7F0yNJ7Vu7F8Jlb5OBI
+pZQyd1nRE2vFt2Dbpyior663TWJa2O2y/B8MNcG2X8y2mQpw2TH465DczasaVzLK1K6y16H3lC+
jvrj+dvys6YZa5H+hBNfya02WE37v2hcYkveMI9T37CISnO2P9NH+wZFrT6YvDUAwSUI4oyiJwuS
NJ2bZdgdkVGaPJSb8X2eYl1f6AHdwsMHxNitdzIWHjRWpMI2MeI+71l+Ud1hCxL3Gqe405s934PQ
v95nlTqjkCniznQYVPk9eq3oGL2AlcNOTNOmnJ0d0wC/EOrQN0la2cnThgV7MumA7wZL7KBTpibt
4H/tSJ+2VSZx0e68Q0IPsFadn0MdF9j+Su1N6lCiB41dVVXfDJ0jLyFTX70+o9uvRvoscLl0X3kA
gAu8kNSOFC62wkASVblbA2knfmimQl54BJrmQyphY4UKZp8wP5D6N9vJpj8YjjIa7aPapxgmZPY5
czO7v5sXac1MTfD2WE2hFxyhX0sKK9AjGUgbKo/SAA75gvwnZy4IKKn1UkdWnqJ6dz03P3Ks+tEe
8YyALUEPTlWokilvmsEpvnzvvqVmQ3/rQ+9dEGd0fNEMRBTxk+QROS6E+KdkUH4i2+iz92A4PJSB
JwTgzqS4swCgMZbJe9tStncjfZt7yL9kSfU4KZcNJY8dzFWNOFWWTcBOv+GyjOREXVHPhdXt301f
aD9qKrjnsUBaOlbr6hW6I9025q7S8U3iFfudGnxqvlPX5MeF6AbrzeK5/vkR5/WRmhy1I8E+fT6A
6XUAwCihltpi5aWIIQkMaGo7pFj3agjQANybDBeChV62cm+vWUoPIQQzGrnJnbNfBBtqumH+NiBN
6hX2zzm60M7useyMJQPfXvcxusTfCa3/lg+GfNdm70/PqPlwZuE5a19MzW/AR3KnylAJKoIAguHm
uQ9ehIOLSx37CFmc6W3blIqWUOJeICWL2scKSZ3HxeyFUy0+LBGFUIFS2Tbe40ewHuTxmCTdSwLw
ErP9p1zq5YLjntfT8WOFIWgtLUpGffS1flCU+DTle1+JZAqiglNsjwzzQLdwNLjeZ1RQg540euEL
5uVuxuSpfZQFMXFEIjDBPOZN+gfOfg54sgJTSGWYGRIT7rkEvsERnXCA8cTFCq3/nCY8uekFpEm0
ENIGVRfnemkWi3SL9Yx8f4EwFv6VLes16UJcdpsIYm4ePW9Uw7nbTF3/26008BbuPsmLHjMjPNLn
qunl0cPnir81RV2aKp6BPm+8/QUG7UEDTGK+1tt7P0N1C79ErA8ZCz/scyndGWmKA+KVGg+Tq/Om
LPio/yjdud+WPDHVzeADd12uZHzkKY7GpKUN9sVc+6zb+fKDm3HcTA5HnFumMu1wnwAm85Rbm4nh
8UussnWn/xptiLhHX2ZMhbtZshZMoGrWwy47X4b1Z0tjQFmFl/Z5J6xE0RWWXpVgMPsvrJNpDE33
fd+/bcXbbdRnQeoYtEKMrlJIrVQT56yjlrHKADiAH0IQkjFpIUf8SPv2Y5pWFXzUHIUgaByzWggJ
2LEbF41PbXcx9vxLeRRL8UhNR/bXDM0YcxCJK9Aqpqz2kYLE2gvo0b/Hp5cG1dyCo4abyNgNQkgS
+srSknHeaaVfaVukFImHU6fktpBQ5n9jInHuyXpr6vAIdUiYE9IUyBbd37cpn8NnwGtnfR3A1pSw
UtDnGonfwov7EJuc8ejkl5Gx5oP9qLHIQBGD5egtwHYSdmfzx+EiaYGmSU4AZRNhTw+/oN1AeP+T
Py0xq/eWAIO03JJUO3KGAVyia7NHzOjlMBy/fPIbKsBpRrssheshmv4IIbUPVyHSYTnysMkn+qVG
TkOFLiUhrjQ4osBnj1s/Bkv/haZQFw+ZcgVRGo++UirOuDfYkhXdN707snNB2JBDpMSMUp8Il691
59gxMXr8S0bfDfHPNeBLwjFK5lpVoBC9nOca/Iiw3OeSXHmtRwnD9w0vCA7Hkt1uJRYPNBX/SH4B
4zOCr5M/ZRBLlvfMKFBAkkV7+N2q1ezPPCxIkSKclXaBqrpHLRKmx5aZoDWlvJEZQD3WDAUULO0D
IPABcwigdjSS3YtM20Z8k8k7+/yDjkCWCF8PnF7N84NWcx3oQSsVvBmvb56Kqy5TYXrMw+ZaMoBl
4Z+dZytm7vBapQl5Rh++MPghUTPZ0EKPl4ex+jsBWId0JOMZ9Mpr52L0wp/YKAjxfbfSZvWJYqty
ekfYojESkaLfZbidb5l9ViwEujO2UpaJ+FxV4IJ+1QgPHZqyjpHmnzHpqJIZRLZjBMggU1Wcz81t
QTISanARITsQ+KhJAkodZEEx14V+hKHa9dWs8kCGEkuJwk1gGaKLowiM45JG5f2c/ywEXg0CHW8H
s6NWerjJ6GQLJnQxRrtnQFQdrn5dcu//QesdzzLnhn8V3P70eo3G3XzTo8sZwm9CkYRMTSBy/MeQ
SLaMsCgOnbTkBdBT3X9MoLWWGu7FYDmB1hHlFtk3XiDlR81KE0rE93225iVX7PwH1uza4+Y2dBVj
FTsySymi7ZhbgqfgV8mFa6f5zchYh9lQa6rbc02zLFkc4OBXwDSO0MdLSLgJQrWnfidmo7NibFtt
bcOVGPX5PIPwk5dl65UNl+VD9gtqpwNz4wAIE9Gj7VyKysxi7DgFfx3ivCuqC3pbAsazRTpk2/fY
LUTjFuTzRHslAV1byBKhqLkG4Ggyr/0eczGSyg0Ka6fqx5SMa+VZZFWHB9WqHwobYsyCbBLl3v4n
8gSSkP0bs/I5C1SsLfy/mcnBG1/6JOwP9N/UBJxgP7LX20pIXyxrsYz4s9RtcetnaPk4N3Xj9L52
zVkGsqKTc1QTrUaDFJKaL5/bQLH5eSiqqjwFqisnlWAK6awoOphy2uNHft0Uk3decUNqQKB53SOY
Wx4AF18Gyk8LVl6NzGSK7mFhP2EKIObjeN8UOvvCVn/3ouS7L0lavASu3jKbxRJYfiNdeHSevcSh
VuQRyRyaubTHf45gNSeW72wYJIQKG/V0HhU3ZhuYMs3g01+g1DeUAWIvS/UWTYyr14bTUnN/bDgb
lws8hJLHlHNLEVNQOhvo6zMJJLDSfiKGypnfsborZnWdz8+peFhA73MGpS/AhlUJ6I8tnD5J6KLj
cyeXjluMc4CH4uHMgGkLYHszZgqAqhLefEsob2jdphKES5ohPu/mbFFjIJi6OqA7igyjyap2FTry
H5TVxalPxuVwdSg3iIbjPw1BaZs4En2dVX8B6Z04FBi+z+uMzFLZAl1NhDZ/lgDIuofC+j1SnRBG
YqxSCfs8dfpBrq+Rm0w6Gq3unDPRnHivfB/riVf+SfM7cEfLePJx9oKf+HpKaJhZh2JDc8OklhZt
kDX4WWU1GcA2WTSUhx4ppRxuPRg/MHOfzSo3/VSUgtH9Yj16uDWpt4ql0AgtJ79mTFtx7DrdBwOh
nSkDEVaIEe+CN1WoZcZR3k75NFd70l6lR4Z/+rhupw2ZDz4aB2H/A5UcUe0cf3ndZU4CsznduuAd
cjKsZ4d7OYX/saKNwQh4xJN6D6wUcsdNvT/Snt/CMQ22OTMYILYTBS2rFGHOLh0ctutipMKPl4zN
ynE15L8BrIU9Cn/sXnEjQQpKZnfaTV1GehlR5mJ+GGsdilKYeUiPv4FaWf+AcFJLX1YFlfE585mz
o0PAKyK6WKBhjECnrf9X2n7rtdG/VPDo1o8aj3gvGJOGTtCcY2okhB2dfFkE7pkZqJcQm40BgJ57
47akWIKZPoZiHmQhHPNbNFL9EDUjCa6HK5d0H87/YOzDqFAHUyZWe2hGAzYeqigXrBqi+MYXtDgV
vhJvKeOkpKzj/+vD8zmqQuQzLoMx6vx5CzfgXLEFf4rm4MCV13D+we3NuORbqQhMCPp1mT7sUuVq
JpFWRGLjjSk/a7ML5193RJ4aV73mBEMzmSVO+Sc008HP8F2xlDC5sfVhq5htVat2EJ08s0SLFAEC
lLsBeL4QSOnV+hB8l0Fi4TS8hpizht0OzUolK2ci9i9vjxfX/mBWcubWS/EulvEByRiU4f+A+oHz
NBcbQsEoocn44dYUTsr3KNDD/bxYHzfQ/03V4MkXHW1VeN7pn2mFs1duw9tN6nuNxBydgU2VD5mt
BOGeRSHsnypXY9SS2ghxMxG6CNSFBnx+lGgvMHQ3UxwlPhcbGkItf0hrJCS0Cr1RpGkfiCHVKiog
Y/YYTdoxIm2nDjZ/PSu4XuSDv/DndO0Bg7C9IooUaUl4+pD8zYH3sgVJtWdquWp67jD3/tXoZwj8
+kVa3dtzTswgvDDXy7kopHDvp+fotrokm6gRmyZ8CtPgtrpRQ5FekdA7mQygISiYuNMw8kcO8JsF
Aa7iZAMZ28x2PT/yrYrteHLsr3vqpWCylGUi2w6agofNqOSa6xjNEA4ga5qxIyd3L+lpKK7K84v/
RlLbyy4GCHz+F77lxzNqEXQhbo+JCj6+gaAcAmYckdIyl9nB9TIDc6CjuuJDxN6yyWJ9QKCPnh4Y
iinZReRERfTWGRHtXvYy6mwjVQJhXauwiDmbH8UelrJ21PlP9e8wUStBB+wscWWoVP6qJZmuentE
iQk/TdiHNJAp8Y6sw0WCjTcnAsP6uWtYpZ1lCM1J8sVioZKgf3lBhcTr1rz3EI5sYstB5UJrQEkl
xt0V8HLZGEouZElufhbAoARl9mPCeVHGskpMXLZ8O/zQE4P/rt5g1zLHP7NbFIjGwCX8DZE2KQz1
/SkDTow5HFai9JyzQfXjse79Qb602KD+XVb8YzXoB/h64hR9A5WGPmifJHGN4RJE/akweKf4h1q7
nQdlOij9JUPphXMJRZwBWBDxv8sFbZTHiRnTcoXAEhuFleNPWzzfC9WMtAcPexLkIJynb1nyFWwa
skaTBqWKgAdZok/0ujtUkNNn7mK5Nlwuzgt+HycucaRrRgLvsJwkNtgV2PIw+1wlj53kR6zvPRhO
ZojPiUU+imzQs8uKTieLbd7EScTMqLUxGj0XHnL98NcKRClNbruMqrmT8HQFQKOEJnURoIgpEv0a
hIB5ezxnthZkeViRYle9/8puQao0CyK2m6m5vta9XuoVjlWFEw89SWLoswIirgIZsEzvWHaHz8ZG
qT9RyvhtkrgrcGoa+bhJ62yzkLnNYB3b6R59dLlrW98U7ualhoUI8/Q11vCkXPF14qfBbsAp/vFv
daLIdgu9vmWTsl4WRZTVG0wUnlrnkrY00e8gmSbTZNGGS3V+aVWPcQbVvPEjargWII7zQx3KCvRE
TXVdY9NW8qsIFdWajtFDphinUZClAj1liotc+fCpCTHuTQEkTbjk5w4dczJdt5NfkTU+GkcM1h5E
fx7UxLQVCYF0VPmhrQl0UYMQOVo4ft51Z6H1mgBfjmiEtIYCVENnyhWzyRA5ARwMKvexIh6nbzLA
KJTiqViKwYcp1s1vkPH+NoXR7WMvIkMDC2XSXh2PwfyLp/FsDul9ei7ehOMfXrzqjeAXcR92f4M1
X1kFeO4krQ0UpKHY8IxO6Zw+rll5Gi749fW0VrsrB2uBIxscu6+I7B8VBQr6UX+dG+5ZXXCPov0g
Ib92hnADelWQpWkizlrZecPnIYh7CoeUS5U6699dz0IC53+6dY21O0uNgKO5l3VUtoiTD/mcGdin
5LUjY3xSYLirX/0KpWKz+dQ1px0TAfKhMbnE9ESTobkElQ/A5AtCPkdDIaiF+4/88uwXoevmV5Jg
cnbOq2C7Oxhzo7xDHNJ6TjANRzbn3az74hM1M7GCk7CxkZv6kJRJMhjYgCT/ipjrQY88GEsg1d/A
yMEIi0v4TK6JU/FCg/d8Yg+kiWIDUQVfuWl72xON+TcNlYZXrnnQRNXzfPWSxi1V3aDSZ0aCtt5P
f4RS3kRimFBr2AAeq3oH0Ez0OfoQhwSfo1KM09K6KQwWR6fENqlopNWmjP/eyY3/DxS3XL8L+E/v
l/8iOZ3KXlj8E9elqfnGELJFLHsxOMO4TTnR2L7c6LdSJ2jRtvJjCDaPRH4YNG1ROS1EC5zwF3Z5
vklqBTDgq6xqpa72IPAoZmpX2x8LPsODMQN3R+G1q+ZMPIBI+qvOXdmD3kEg1Tn9/nqdNw40bEl1
E1afW3/oZQfcHZytcRVzeNOwuMLLjWqkmc7HN4vZkIql6A1JR/MLT8XlL6+oAfjXY5tBEc91kpbl
Zjr3SMM8zcbvZAOlusOhyP6TMDVlVw00cEMlPQnNlPodcgV3qvMec3jxhJ2O7KoKi7NKlFk3/iPx
UkGllGjLtmydfm3dVDgRHMNpx8AHPr2W/TZTVL67icggSJutQwd2y+hsSzudOswKVaH2IK1hrJqe
8VokU872RWH9sFs9qk04+YiEQ1EBTI3jQUVAVi44bEobubESRbNVn3O43kZsI5C/y3UQ7t1Dquvx
hT+FCVynx9QhOSMMZxRNp6vm/XEih6BFEfZ0/fsqIenvD0XqM4TJmErkfSesde4h4kjLQpLMFEUc
y2R0C6cckXGEXWONtj4rXmTKYknRas0w5mODnEGq4SCiVstJFBN18oUlEm6Q+SDz38C4byaqvrQy
w+6dtxcj3WOZ4aXfSc4UE2Jbf/pPzK3C63qgMI908brtVS22RyaHbY1ANftGiIlCBhhtnF8phIbv
ozmC6IWSlLtkUUnPcxJvQwJk+hzCQgRjMqugf+e3eU8lMtJjaZKMuNC3/DafAvFEmCNbHx0bkDiq
f69R9et89bMBzOJpvpiE7gwUu8zk4aMmBugv+c7rBPWpQ0fixk7VTIoeQ39jHcVsU/O40g2ljs2i
7A0h3YwqwJuDanBefJBqwAkG+88A5Y5ImriHnXAO4MgXxP/FVHCk0spu+X8V6rb8KCAHNo3+6BjO
7AyOUqq67dhglYW6YHYat5r60/O75armZiHtbGxIN1tfC0ql5EX4BqanljzPzibuGfBe0IUPJW7N
qnpWYv4dZHo3Ygai15UNg6LNd6v1/RD5yPhVuHmKgf4VhjH7Ji1+X+Vd5ORCD5X4BYHPQ2h+5Z/5
tYvLECrNyxjzGZAElC8kAThcMJ2PyMVa5k8FdBtLXsfjuwE/SemFv1+wFd+B6GmwaVO5G6muYqYv
KKitTfWTEQKo/ygTjeerUiqQmsof1ne/K+qp1dm4Bji8Xy5UXwinEbBxAAfmyLut0x3LfMyDlYqA
IyeT8sap5HIY0KHCGHVFYZNdjg4DpQ0zp6ba+gKilSeJa7lpyBypTTn4K/qGNG2NEzaZahzE7q5u
CReSaZlcfAr1W9jAwAYae8Ujz6Y7XdnhlUYISfUqDT9VQXuN3sdFctixQFSU/DGVLvcuvn69mCY9
YVAoDOAd2SW5THTS2+pSOElRyva+UdoYc+eGKYy8JWWADK0Z5BqYsxpK+nXIZIMAwE7jCZFkTBJp
3oDLe/+7VHJy1NmbkRfgkhXTSLjgqETrsS1kJ0kPh9siDrM01Uexq8Gi2gIXrRsMH8+P3LOj3znO
6Lydg8FW9HCOKvoaUMdMjQQ+Xt6ht2SJ1FXu1IUMYZvrzPXl81Me4t5uDSYKpmAWPHSh3RohLBJ3
t41tOycfOzFONanHOE6LOtnYeRirB8DVY1YMIuATX2yqeHhdJTi5bx4WlFuRxwHeKS6h/W6XOmjR
e+Yw21SIbPuq7WiM4u0UAgquuL9HBiK5CmDIbJXdJaKEnxVU9HG7QTK/0RYCtqjkCpo6eyN4TN1q
qI34+udm398xYJZ2Miyss70KPRNz7msexC1FSdhCzw4yQZh49xVvK3UaJCS4scyk9BRDu8cg2Fxj
VE3Uk7Wz+tpMuMjMxVWxfX0iSkqH/bA9u9m89XPe8mtfIrx/kWESYjR9Lf9siN6KhxqcPsQ/m5N2
C2C0kRjwXZ1nM84zwVVj9ihewuL3vUU9dwxcdponxykQR2K6FIbUImjn4DGDi3Kfb+rTeMqcSicA
A0yIhEpBWGTlQwUR0d/Ce4z3G5NWt4hl7YplCmRFxyVnZnizZA6ePkB2vbAKAKb7FpyvLFsCzBQD
w3vOkDVaLLbMC6OOUpjxkEIpvFNSw2XCkkvn9Dr+v1jt3NozGO7wLvHCK0muDtC2pJR3hBgVAJ4M
8GTjKNYXewi/ju3i/eSCWDZjNNoWhSKlqnzcy6I7flcrTti7Cze5hVL98cUN6eMoBhTy9NmjLdfo
7nUAuhF6/4kM5hplIRirhw10LEv4f8t2FeCYaxYPxpDS1Gb7EU8Jpo6jmih+vzbvTkQWJjAtUZ+j
IJN2p/hSq1xYcc/NoYT28x7t8LDcQNTgwIepQmIl/x+vzJK7YynVeG2OzsQMhT35c+L1Jw1MuoP4
zS2vv74pl53nsNzZF7xurb9bLsn82lUaOVlzKAdncV7OIp0BEmARtUhoFhyIkb76qD2dy0DH5vq4
z0CRwDLtylJO55v/sTcpgmBMTKzh48wLDQvi0wc52EhkTuL0aFJlCkra7ZjvP5fgRjucq8agetPC
80JuCKEuEQEVc1LrFBOqkgQvYqRHTmvIRUu9j885MGk/ctc0QzMbTLEzBHVoalR6UIOP0qjXU78N
S43+te3u26HpOVGYzgEqD1axqp2/zOWIU3fMZIdPk/UAcEB9x7dAzBPAXMq6TUjwNoGz03h/DVc4
cmCshGSyM82X0UwVw2Cf6SWEIEHMdN+CzpkDwzkgK85oeCvbuLHALGMcmUcPyAbFIVCvomBitdC2
EaWn/3+I/1x7Qhkd8+KnSe2O4KKDIikPb+A/a/lqiyj0nWfZyZy8ouUwKkO29dkOt7lAx/AbZ7pu
ZIvrzrr9be60x7C3ftjDYtxlhACGaurMg4z9z+aspdQgAw4IVMPfMjyhk7Yh5r9FKVV9MOzxDDZx
YjY95KLXjaXEtpIBVNs2+XHPUte2RJYqEcNstSTYNGpWK1097OUFxv+L+OwK3sspMbBqZVqtSZ+b
4jP68KMCOfqtpCfTEf6tViHQ0LBxKclT/v12FXbt/Ju3Xh8RKo/1iQbaO2HHiTtZSkgcH7LHf9ux
p/AQNl112HqkWZFoIp/MRVB+u9EKHNX26YIewPdZWVypse8wRO2bxr1Drng5VENSX3Gq2Nzvnkts
lWdY6135bqoB9SX8W7mnpangKHEaF8tQDm5IB131RHDIgIm3/RJG3SDPswcMSuLIccgi+ogqvxwy
N9SYKEpbguxLDOngHoG0nn0/ZsflEdfE8/Jh2pHjzgs58+gan3Rdco4IyiAG0B9Ib5ys/MtT1KIs
cjYibNvocGRX5hgJKvFn6xd2dNCjzxl9NOg4ztvjez5tCZUwq0n4k0EMY6I6AawkAFkmEUAqBBTS
V5HlBQ6NUqRsxiERbln4Z0+kW4V0/in+0yEErr61dYSSKWrinwKbQmCtkPupz6uHqUf/4oBqZ5UX
Z8zyXD9f7mjW5tBAnl7PZG9kw6EsyPBUuZFSMU0yfQ9Urigfh/lGoxtYNNwOQ00gmB5OvzsFWf7G
sOKy7jDPQ8T12tgxsamSfjZWS1MfBxWVAbOc3+/DCoxbAxH7TwIYeoYjZ/U4L6FzSpFzoSlTrPjk
4p6gFIrNKNYnhyYEWCCPdCZXZFTVht8Yx0Wl4YpmqPCs5s48/qFQhK9EKz2x1eogylxnl0tUGquy
u4K6fs2k/lIvjd+pesoBioYs6cUZkBbhAUo3plHv9M+Lr+IYYSeJgYv/blUwGgpgMEYanOCDHl63
ZqNrQRN57d/IhJSMsGRU90d9j6q0IbYy/ZRw4zyRsdI/wRoWWNKpm6HbboKEwdNtSsfMazxJUmtK
QAKTAniKKG2iDNPguzm7FoqAJWenDp+ISPgnSPdaVGCu9k4oyMMNmOb7wo/kYY9APH9R101Ao6BD
GbSqiqZY4YOh8TTc6/d3VpB4iqv0ZGCWaPW5KR7Fzf4UOCTQzXcnrBfLrGunQc847PDoXiQ4+q/h
qZEUSsyvQk8MQFSDcyEUNZhz2ReKojE2zaeBgu7dmPOSk2JLth5aYptELoEPIAd71AwEpleK3Acz
C5GKXo+pqTrFbwTmhNoq1KlO9Y0OxMrNt7byWiBeg2ElwOpuE8U0D/sTOERhSHiy3lwk5qFB5++w
3SOzYLzHhhhxOAXa45f5hReQZ2AHxbqph3Xb2PhLEnrtxvY6CeSlB7lnxKpywppBut2yUYK/etKG
/A9/iWniLbK6FwYzTsQoErZl9VDY2pidQ2KHhQekEsr5OV1hlz26ODBOBRz0lMEb1/a4e1yy6vYO
q6KfBF7XLiL8ygGbvuBxXdrsJ7vfMp+l1D8AeorhF1p9gFzuOyNnwxA5BB2/pZXNk2FENg9bxmzy
/LlsBJ464mxvtgzKGwNRWCq/HrlJjwk3MnUmZpTzn6epERjmBv31ALNNZ3P5EkPo6CL8Aw9Ew6aU
kKaDtZpt7QTYsPCLN0zYjbilfuLIRQRR3mWn6/2CzFVOk2fnHqAy2tcLmMEU1g/MF3kvHtTzZ1Cw
TEy0QlzMcea3i1j7HALbxZsGjhnG8iqdqgN1yISjeRllnxmtyOOg5zlyRzqFkc8kuakjeQv6ps1O
Lnpq0Ju/aMEIMPOU60YdxjId4fZ+RaJ6wbHUzKVMz2/K6ixoUaxLbIvp2MZH5uRi0UsamMBPdZ+5
xeSbbgIJjjh0Xikt3Dtk3aAN81NYX4GJY0/VO/Aw3N4YCrNcVvj2mLRH2PW9X7zOkPYXoDOvltmW
Xu3C7vRxoBgb4aLUQa2y9kHuFjU++UE0KmhtTQz/dZq36VGhwSgp5HCL3Le+hobYCyYXc8xm6ZeH
AwQQOGbtuoKykhWY3G+APrG3FebpLnrhPgkCX7ZEHv826tZYDzM40m88JClnG5xrh6AxA6MYG2It
akJtmY3z3MKgaGVhqcM0DrH/II8eAhGL0K+DzyNWo5XO/n5I/bgRDYEKOGI7u8IW35TkCvB/RcGV
qXMyAJoBQVAdPKSwTr6wq26TRx9vWCv2htTFre6LSC2t1yRrhM2TcWMuMbnsODyu7y5zENbg5IaL
rbUcjyQaDolLDgX6WI6CeuSxGPzpwwC6ZgjAG0R6UlKkoPP/MrpNPsmnwLX1pOC+HsYsxFuTwPP9
JthiAAPqFBYU5NDOarjfuDw1gKOW/gqYgx6rspjhclop2Xpg+pbcUygHQ6E90CoECgIlCKCVpcnz
9ut9/OTD9YwHLMOtUU8N3NgTwp5u4qsIb9joJ9kQ1vvMAaElOTrR8rQ65ItjT40R6lBnmQRPwGT5
bj+kv8eJtNWCF97DB3aXPzbct72fXx/jaiQK8wtJY3xj5tkD+4lmjJGjSqAlXuF+FFcbycMWbfz/
5z6CyNU7wiig5a/Z91eivcZi3pzFwlq81xo5xMqdoFFWinF9Yrix1fVK/2Ge6yPdkWLFXj04+9mI
cGuHF2yUFiNnct+B1DfZ1jHiJrWWA2BBwXKpRW2Wz2Y8fGG3lgXQa6YBsQP1/PyddYXRgfhhltXB
fhYRO1BwBN1U1sOimfRmILq/syDDaRvOR+ovEK2fg9xSEmStQmRJ37obCW6GSmpaKnfXfFVOvVmg
SR0gcD8p8Hw2jB/YRwq84O1yVz6/L1BvTVlXKIGv/BjkZCBGot9DWyRZkGZeOM87X16c3jtf6ZDR
gWkvrAsiZ/m/jedm5kzYMO7VSU6M/4i9vF3sW19fvGzadZXAUXXQ4jEXlKH//WNu7uhU+tPeabdb
rQoCh8nvL0VW0t2jCDkAmeXYGGWcneWXCaXeM64vfFCxZvUC1pNZ0VDaGnyv8EZPkqcxRZXPexIq
oRU6r2ikKhgJZC/yJPvmXIiPScHczg7uvHDsnMmpBLh8n+G3BXD3nqE64ygqiQDhJ1o7Vw+kkScH
3q9iWqCYfx/J3OU2rTemGpE27lH62VhvcEDOeXMBisyDEZGbUezf88ASG2ElvjTHlf7besoy5zVn
QlrAx4Kdg3XO80GTQ/rkLe3ylZDF66AMj+lMfS0EF4sHEL+qHEN0eNrxhXm+nMEcRvJXzzs00RVU
OwICiNDDObkC9NW0bNxOp8dNGlI6Y9Zwcohr2a1zSwy6uOFYmw7bMl/lyk8yQMyKLfcYO7pbVx+n
jJgAGqe2UIf0J/SzKufXHvDeyZKMDyF7kZnDKhp4vzxuGGh/uY8FJUaAoaTJpkjVxkCIXiA/3Qd6
ZQ6U7ScQ/opW8p7UgbdOWzhGwulfH8pe66Y/JyZgnEmdc8iYC93wVEKl4VjoE0qnpEyNOPYhHQTS
uqhFPScwRTtozc/F2/VZHd5PLvVTs6Mps10N/u0V1lGPsQzj70RyzL9AFT6m9/rY7GMuUwr0xKzr
TMsZbM+ZfBfnI1QmLGZHigRvJYSnqBUfb3ETyO3db5wjh46mMfbpu5FM3E/TcEQFfIh6Wq+pCfNp
gWrPFI/NZWkJ/SrmOsRctOJzpZ4yB6WRMYxz1zzv/hgU/wP4U20ucAGUJVLSKef2zoqHbD4eEymx
F23C1/NUwdXq7jBjeOzS77mXpTogY2A3aDUbyKaLnRk2EbJ/3ejclU2ClTL2133EqfNAa1zbUhKb
dC/iukNui9em8QG2U7ZnS1nB/jUb23vkxfu4JmA9VDkupbXFU0c+kHjOrk06slpQ8ckfoPzAdOjE
jQRdOqJSB7oO/TTk5tIOT/MWqmpaxgybJ7KUPfJdtnrAOWlXRElwgyvj7tYCHBNg3XzxoRzIgsiw
v9fmuYxX89fnCQ7ZCvAERpyVeOmnnzIW25fR0paYe+DfDo9aI+w8i+fxaiAEGs7rH1BoT/AKIUBG
NtAHlwFTSo1ObqiNoW932ycluCcE453sA3V9KZ9Qz3a561K+Yf3vd3rGnaZB7KF5xHtacxpiqrwd
mL6oGydS58TBqOqfL3BlejmYppK52kS4ujVRs4EI3WBaWok7XhFpAlazXpO0kyimC6QkNN0+501G
D6S/zHFO87cctrIWmR4UsJecpHWtNy/w4m1wT+tp4IRgC4RcbuZk4dKO3Q100/ZtMTQ+bvG9U5z9
sedG4OF+VkOw6dgK0ZWw/jHFF/iB+YBnF1D/IljebQy/TgYUNJGzdfJFXtaoKSgZqojDuAhuKLSW
JLPpJ3HIpwS+GfEuOevUD2rI7KsJ3H1HlaWiXlCu7oXTtI4ybqHYiDJ1uZFA9KqLIIJGzI3jr1NC
4oZ3s4OBsAcdBqrdta+gRx4bwAeV3isecoBjRcuOX5uOA0wRnM10pM4R1gmzaQWb2BUB3cj87tZU
h4iv3L2LTzVgLdtXcUR9tpm8yZmNi2BNq16BxD/PDSQx4s3ujQAZPlyUpjFoM2f6wCqE0ieR6epg
43UgDZFD46MRCC7EB6QB6QvHPLt7IIZ6AeE50z+U3ZJasACQ+9Bo4tr/mXev+8wyZ3O6u2p1zqim
A6jMYjlKiO8l0J6z5fFYi+Qy6U1mxWK15Bd0LtL3u+KRHLwgobBOMWV1APgL8ckfi77vMguMw2w+
YK0Ph5nWL0ECJJV7W0gGkXpVpdhBviw4E6BpGPVLMyXxHx4sipoQS7gM7bn4k5VHs56z46IdTnJa
9kISd8l0JDewQaCu58sVb1lIfbmS9zRfF9lFjtBQnNEfK0jwzOgN/bv4DjcaQ8nH8lMVzBobm//L
Imgrhv9FNkrt3TELeVT+5oWzrF3NHVJvkbfBzcWFIXOhwpWaiBpmLYHc7XdpJZx0REZko8S1rnWv
XgntEl6RS2e3V+6PbeSAhD+ZY4JVdetZFwMOr6N+EcMClC1epKQy0AcKGa4xi9d9fextUjlp5Xhq
ATI7Br5Ejg6ffduYDdPTi+aHkDnBvYfJmVCbHZYQEWAxiNQetb48XM43bfV2utYYBAgkbICb+f+x
CUUiBBUrgZZSiJI2PQ75Ax0uJqkgt8iE914hIPiTQIixpTus1JuUGkrZI6gARD6hhYWA6mlBMnxn
JLPei6+2DsenP1vtjkdqUKdXLMYufhfa87JagbV4rGbGMjWl/K2IrpzRHqVPIu+/CDEpzoveTTad
rclm6jptlnODOrFpkGHJqnWILanSIA+N5H/8UYeFN67t/FuBcH4YsstpSQaNBpdZDkeXsw37nY/Q
C4Md2+QgEUxUmS9RR3PHBCfT0E7NmGtz4qXIpCD+DBE0Vbe4+ASOH1yoL0KTbZSZcOF4K6PjU8dJ
FzNHsuz9IXyNFKXbxojBTd9t3dFDLo35p3gCXWfv/L81ytg61SS0DxrLnzZnB6bTSCrb/veasdww
h7P2thlLtyncnmQT3/+2SUdK2N1A7QGLR5ACmy2qomnKyvBanm738FULXQbLDeEHJvGIKhUqjkku
7Atxi5WF5DsFgf5bDtXSIn/XUBah5HNKUk+Bh43SWHrYO/f8ysCoX9jNzILQDCKsjhmmIo+4ShnC
OJSeXzgmJeUA/tNFzaOPo4P9zD57qdlhyYBCHOCIQCy2iyFMPr3wVRxGF5fgVvaMdTeSeQGTAAt1
zoz/hMrxALUjD9sjSeslscF28Y/+p0V7sweAOTPoU1eHExqWOIxhDsqF1PqcBcdkIJcpc2vFHmiT
Vwl86mXrhIJM778Yd+/CDrzlJsVZ4XPaMWtHxGUL5c5kJTGbvQXar3CSHiIShe1ma0g3qcJmZKoX
1uDUBGg2KumckgmShrTsDBDFYSQ67MLXWmvN2dZq1ua7T+vQhujriSxZtg5fdNap32bYaSX8zLwc
VzVtwXuLjm57g57JhxeY3qZEeem8okDLZQXBRPPAE/CbIqCks+zb+/5Yxp7wbRV+yAC0NpPA91sf
ZLpsD6pgtxYgIiWsWfxa1RYq1Xq15PGyuhKzjEqKgzyV0pOUVxAJReoUI1axkpPTHk155/KUKfIJ
Z5Jwu4HgYxeN6zI6nFfi3Xe4i5S/Fc5t9jbN4DVakH5+Dm/imgg/93bUpWRA2/vgTInKJBLNeM3c
4L0oKiXWV5pCIIwE718gcQDGbZSoLBHDoda1oxvnnEW/lenw/cXOKA1kn4SRCIccYMzUJB4E7BWH
/IbC50wOg4mb+PBlz1PQCzAQ/6lfQGNliputizu4Ci3pKiA0ELvNZ4F0ySX87AogSu1VbXtd33mZ
MNgOhz4oq+FSkW/DcYRAGmbuSdbgdZkTfx0HsdqSAGsShpNMzqz4RoT1sPDeCyZKK0gJQcyr4A+a
muwRYwD+E+iSJxcfRK2ZwqbgE2WmuVG700/547bv3zuSkHqe/2ZTC/0yT9+jzU5XZnFSxpxg/4no
CrGoKf+9S7KHg7oZLQHxiU5XV1n76AeoPArfcxSMh5GNJ5b0PxgNhTsAmiXXdA+tSwJduWcmPdPu
2AQlU1QYifRrNvLAatUt7JeK50y0PCqSeAH7QjiiPUqeGD+XSCj3xoD5oZ844MC3oKkYprKmnosy
QfmFXx72csBPsLAAv440XXSVSyjG0iMiM+ee7QESTCDy2S5qW1ON8bT1UHP7tKei/Xz+FY091vPU
2TAkmK45+pCitSY/DEvlt748zqidyacXhAI3m92Kw+rIYut7jzfq160DJ6cSMJw5Oecuc0DHIKqy
LpCll3dWmG5ACq58sv0nh0w9+6dqLaXSMHCLSk/vCJ9EnYyhQa3ghYDVZZoznW9pfPqEZZEB5L6W
h7pwHFVFiCpUfGjAsZTdGCD2lguqjJy8KvqacHEQFVpEADI0V/3hyRtSK+7NuxbGRLlXpi2Os9ul
697T6ehg89/yGDPBpcH0JZ/q2Qfpj10rLgQNuJ2XrI+Fjcduv+iGjB4xITF3PPMgk9QwElM2TBZY
7gI1FQceNxbwIXSVvIHvsEIALGnvSy25deSBN7YQ82UfjTDYMSfPVUk3U3nqlCXUj1uIH1a164AU
Ha/U2r68pjTSaiEzFMrThub3VlAX2kc2jn8jvHcAxqi1yoZ1EQ3vL2B4tGjroGjK0jG+kiu0TYVb
lNKP/3tEJQWyOM0tbxq/WiBF8PqE84DP2sDhvXvHXXDIV0riWkeqFFzu8w7cpdzDEdWb2Cd8omfP
f60iF4HwR23GHNoBOTFHDjQpLBXooe8p1zfPGc1QVnfJRdzzEZzU6+coBT3SEVtF5Ney91pNWEYr
b41jCN/2jdVWVkF5MmOrBlM+2Nltzpli5KazSMC6hLpnBQYXlDWnOO77LX55vxDAq5+3nQOoPapT
mmfaGS72qeshQOJszg7dLLJ8QaVhpf19jXrqfph7FmLetKcOFziMI0qt5nSLjBJJXjRTSeUfD5zp
hmyk3pndQHOKqSwgDvY4xBjHrYUHBIMW3eVhL7aRI25WBcymB8wkD2s5tNypca3z0rOdhGq25PB3
ubXxiKIt+K5nWl9a+95lHhp9TTWyEejRFoN/4+l4d4IchxneGCwsq8tBgo6Bi9jDJv/a5oJkO8Me
kT0kCUf90ELwIX9IEZMPk4CYENu8g8PiKtlen09OYLOYBsUT0NPH1W8llOC/xwcElpcabPM/d2AG
fnPVmVh42OxVBAJBvH6LeTf8qGfhem9bIO6KaBvGMTAGeP7/+A/FjenpHbziqqswdrFkf9ozjFX6
AOMJNlR0reHBVJifPcXaPJbXHuUuqx9jh54ucELCHoHCoHFhRjTBA/ysJ8KyRbZYvTayLEEZWAzL
aCOmDQ8GGm7bCkn7YmcGSXmg56MI+Fdfdmj0XCtGWWZXHFX4BpzOFR/kB+Whg4sEaHEY22lo9bXW
x7HKxHDWpCeuwe/zsP/hg4nfHwcFVi5uihEn7MHdtTgHj3C9FBClPF254s6tnGlOoJOZp4GOlJ28
3KfFqObc+BMFoTBCAkGeMARz7EqaDnvYnKc5TtN7WM4DRcsnOA2rNZe5qYDZTLd2gjwZ0w5buIH/
rvZMM0KMYTOP0xqgu1dGZyA0SJhbpZehyeKJqxXkXGBEIRfqFSgTYWCbl4XPTzMEQgNEYJN1qV6E
SUDynJWcpsv5WDz1wafNv+PFLojmOMMa8KS1y/9VyzilIIMQ1cgiKPfinxM3xUFsAa/OPjR2MW9j
GgK8uP/vgvxJXEWFu5p+FPghhbQ2+o5DzriU8ata9/nN8xH2cmoDDLwUEWhcjL+hTSYIb/DCJy0q
iXfSNvO4/DdwYo3Wqh+FTeyFpyNPc0j48xUrNMbKzQuYtzjaK2utWI4eFOrz5Bg6+u3oPdB4LDlR
pQarwg6FgNobHYBlcghkxXyuBcvSuNECew8hg2eaq9xbbzfedbhstXSFbluX64Z9zG0QUZH4nY9Z
/cd76mqNQj8QRRFZSETjNL2XThqhwuf9jzh/d6fl23UkWA270PtgvXl22rtsJCYoUJ65l+IiFOK7
NUBsQrrmisr2/qbPGiqrWyfL9Ae8uTLlfdM8fG8k3D/BtYP63RuZs0GSVHE9tm7xfaxzdwFucxDP
MHvWY4EOjrrEadpvnfhCzNv3xh6HQaf47tgU+1R9P5LdqpJQEyH8nfhNjuGpR+R3gQI1eqQeN+kn
FTTF7ZQlqLLk+pjb7e9a+3PRLcWr+wDWW/ck0iaEZIkWI2C5DJWFcPPeU+41mxCBwibU2dqgPZY+
6pqOxg8Hrd2iS4tFkg7Fvt4+Q1q99x1W6a+YXDCVvR7g7aTZa1k177zQ1JqfWxi2uz/6gAmj5zg0
s5UKJzcUhHN34Q4k9b63CEBuPI8L4L3UtKu9gCMPUWl+3FIMeyQlwf/OqBcvEOLh+Viu8w20auD+
QzdoB/ctz4PKq0hSI9cstDE3OTvI/eboZukxGpNwswP1d4V6C/D6b8j76r1I53U8IU2Zkv+CbPwl
2Zp2cTBHGCvGepCRbzccoGC/Ef/FgTYyeF5fAc7HI4b/1gbKhGxwo85zpPluAwuHKZgqgmPnHdX2
iF0yIpU9YmxvH2WC+iGika3v1XoOpXmwqsN+XXpayOTPrWYRFX7HLyPQyHod4Iyd5vnqoQ0VFfkX
u1btxVsFFZkblY+khcueldLUNTYxVhqbTogj3E24OZ3xCxqmOddsCbrQGL0boZ0cbCa1px/hWVM0
08+Gos8elNHy1iBwdRypKW/jFEFMOBcdoKrznZcaX5lML5GvEHR/ARkBdB+WEGswyd3xxYmTRgG7
qk41a/DF8cKD+zs94pqP1nYu3pRmz16CUbax4/uIZ07420rXW1lYodGdlUfd0xXIzjZLAe2v361i
6yIdX45TuH369q0bzV4gQ7H/QshGaFiw0nOTmYSKgKlhuCK6l3OJMM4e7XzTG8Bpmrrn/BRcAboD
q2QqNQZoFVZy3IALNWor3CfQul5uYP+HCwDWZ6oUFZiveJr35/p+1QQLotDSToqSuwg7Ycjhx0OP
GphfnDt+vX4nuZkshROWaNDC5dV7jbVEvudhBSIdd4RIs1dHMWMIQKdEnZZ6tDF/kbMqd/OIu4Lq
Ae8oUeBMOIxM27X2Sw8tT9Jn+Nm4PHjoja2Ssr6yqPWdxOktAWFc/zftVUtWqF42vfpIa/nAEzXb
KV7Y0cWUoiqnj18oiJMdT9gE6KdHCnRxRVE9+8zYhvr5c6IDvoPBzaoWg+aTziPFGQ1os0YHdV/x
aKwRUw2xlvtpCjCafnUF67LQfBY6iUnaPLFygYYqnV5u9UFSD52PsinVHgevoWqiu+6qSZX5DmDS
53Q1t/Da2nAcHKrLlamVjFbRRICrZsOXBJ6E1JUxbv3nQxOatelHMr3yHMEZ8IZC0V8Z4CHbPBwe
5K2t77xGZSGnUS1Ham3mWu9QMwQ0inX3QW61EeOk92ePO/yfl4HgqKxnghVDYz3taIZg5eea08+T
FLjTp9dEi+opOrmX0vWnLfVeas0eU4wN7ZzTgM95tj2zTTRSe2YymFjOT1Dwed5gY1WgUtvECT7T
9O8ooVqiRjZNWQMCvgAfU3psfPptk9LNGV2xIZeATcxz3PtFVe6W+UrgKc3wThhV/6L3guftAnIT
iRCu7yaL2ImB2YfqAOFkvLlL2zlLkNMUjObOuijzbyRZmRago6ue4R+ZMF74dcS8+1XywKFLmjlE
jp9P5Koe7QDnn70EBHH7pjMAkIJYwoNEpFja3jzZdmGL6oPCI0viqDeJhKa5WKTv8sBMVX3aVKzX
HqnQX+1hUjHO44ddH2T8dTMX0D+NFRb6/O64RCXTmlI8m3XFK4FAicXL+GQynik2RySHTIqFODcQ
TNf+kJRS2djv7d28yY5Ut6dir+47bi4oMrnreVtxDUDf43+IOkeS/Gp0INt8sT+gT7Cktm2Xnc9Z
pAwePdc03uMG0jCqcDNNl8wwdCPXN3SwpiZBztJnJCNXNkBmTKdVPgZkSXOTV7nP0/9P+8TwJobh
u8iZ6Ep/PhdBXbWJyLlFXtOB1SmgWpgpiZ1I2mFHKxSW66xov40eVfiZ/+PCmHJbBNscWxLaW+gs
aG15NmwK5+bYiOBkMAdR6TV69sFX2eN45sxxmbUQrUtp5LsQGpyfaKpWr765aYqdtgHRCtZFOHAJ
T33c3+5vCEN13Rn3PPphDM6GGi+ovzuD++wivsATzJtTXOI4j3GQ0iWqe5Jwx10nvBuxo1hmbIWk
PHKW2pqlQrkaSlYAN0cjM4lnEKmk9MxFTVxEUSJ5WxbiKrveA3t6KgCrZo1Wr6TZJezdkQ+A+NRV
41lmg+dq2evXnamzuCRc3rhy37jHksJb3oQc6wdHvt3m8xFMDejib/nbEfp9FccDkILQw06uObkk
nnB8ygQlf73w+aIOHGm4cdDEs4n1bpH92p9kR9AgIuJFRMVN24isgG8rvO4lY0luy/y0E4kPfSF6
kkZ1oLEQDYid9NX4c2UEMUCtDBys0JudiIWnrY2kHof3s8kYlRATMK40q9cU4sGgR1DhDVegCD84
7AmHnATg/4QL2/0JF4Oug9xGY749D9Fqye+VQspA1cUoFzAL4HZyZBzqK6w4C1fUoPcOxzSdECHN
XOH25f3zLb/ygylvAaoYj49890l+P0UwtJKYzc9gPHFSuzu86IdsmjfnX9/BTYVaBkoY93zvIe38
Czj2mz6SoiyppJCIpnLEDNsESd0xZm0ctG8jmp4bNxGaw2fTqGfElo/hiBeec40+1bepcGPqyKbJ
IQm1UrSnz/6t6Er8jys9RnhL7rHNhx4LeaYoZZL5OR51g4ZwUjx2h5w/TPEnGomDvIxst2pYneXY
aEdoE+T7s/BgqCxXubfB48t7dbPnQ7zmPVDLMmaX06HTlzg9EjBPz6VHUr8W+jCqNQqHwcJsp1jz
74Vea2eOSqW6/34N2W9+mywDsDia6tg37oul+/dg5RFOOhPVwvSRvWO0V40Sksrt0n0L1KjSjGhZ
hJt3bGQEWYwAzVcqC3TiGQIWId83+zoS4Qhnlon4Trab6VsPolgcltgY/v+J1AS9JPI9XODfHbff
vVwlffwlgntCXkXlYqpVTwahLuQNVGWd8gzgV+Kti++Xu8NCEIKzwmpeH24ICt6R6GR3YyPmy6wj
oKUFOIV81/QvDL1gXWS7Fe0NO+IGK0szSE7aMhojOLm06EXa6KaBkuUC8ArvRNbVJ32+DLOPlBPx
rneCrm/hiu9QBO+j9PV4DktVHRcmEm0ESq7GMVGGa+tcaeErrlBtneUDJYQ1dJCsTf9JdDl5UO9Q
41RUrNM1E8leqyR4ncg+RVrjo7kUgEay/LFtRs8CjKi+Tz6dZZ0Q1HjNXfprDgcnwdhWzjgYrBTF
fxGPhMIm9vCXoI+Nfsz1m/dVSKpVcUeI82VFJORsc6s3tKsnZdLS4TgGkCpNFgjz6tsjx5pVhVt9
Jc/9jB3Dea0SyQ8JamOJCL1cbO6Hvpd10/rLdnaKT43+8Fy6rbRnhevjKuNiAqcfpZQEGFIuPhLz
aQOA1Jvr4Ungu78CjjXOysWeXxiPr6QIEwGoKV0XyAf9C35q62c+5LfNfGrP7icueOZGENsX100q
6CFvkQ5JskCFgzmwkDCRpw5ZQM7HiH/d1If9BNZidMsE0IPsW3YEInp4uZbBSzGtqfIWVkyeWlCj
kVG2gaG9cB2meM2dfBcKzFPYjt7FEc/+izdiBu2MsNXWA0dn2fvxGMntFLkWYQJxZzghzBGzzLCQ
tV+MqZUXP08/K2SnUROj6H5tpK2YUmHM8Ha12uNHkXpYlcAkzJjlr1LCasNQv2w1Oafo+ovkgRF2
GvdAr9AaPQl2UfLX3TvGrU0y41YUP/71EMY/V7DSNK3T4Q++UAI58EjKe66FGd+l+eFRbxckEhMj
DfPDhFyq9nmZrCrycpvpZWHbrzSvfBGbMMfv2oow8Dmg6WRlItGNU3SsOIbj9kqLGQwVsZY0YJGy
ixBDwZGQ04FH07bER6q2RyUcfRzTsBYUxq55pBY0zDHvEd/FMFoRthKNK+EoegyQ6zHLU63neZMY
gTU7l5rLK8sks8Sx6M8Qr6R1Xdw0NXN+cPr1EDuEnw92k41foN/GEXuwWojen/daK7xJc/5Y99yb
/ghq37tVzfXw2OrrvxMZyP6CrGEYv56DrxtcAX9ShKbUIJtkPdz4y81qgYzk2mE23kHw7Rism8VT
PrrlgMs/ksVfmSvKELJERjTnbyGGx3YW7ZLhgp8xdUfq6CIJdUh0wu5t2Kwuo8Z1RL3al0e9ka7U
VQfu7rV2ljcyAu9FiberTEop20fBEnIEEdg4Z5jgn/YFEucKwgHFSO9K6CPhevP7I3dK1FGwaB+w
b3s2GmIMLEY3dw3dhQehUm4Ij52DL/wq4LvxPJPILqAu4RT+q+HhOx32fAGqq+ao8H9tDGKfZE+y
Rh0C398Y8Rq/vhraHQQl1yfzgFMgUAjipI4TxqpL45Eix3aeQNEIXuMC3EXeY0xogC0BMqDxdXNa
Rh21a1LEmN0txUbMVeFGpqxpKBRWFz2tWOjE3uDjchelgGiz4KeJckT+e8UbfLvFN2n3U11aRZmf
Qxb3GgJX07F3c2gKCdXOepJly/YG88Acg+SyABJDyzjN0wcNTYM1kfBgCYZxGgMXtzMYW6i/y/UF
nK3JvGhCH39pEZtgPpR4xaSWglgoI3p4W0fRBG6hvNbHJQvAgQSx2GVw1v2jUfmS15kf11dbCWWf
ALNNvhsNV0CORlAtoN7NuhYKNMK7U8eeLF72Uk1ql2lj/R0o0zW2hJRNVCCHMvIH5lO+Fq1XUHkS
qeuq/z9P1Ym//aIEtpdrRo485t25R4x8kEeukdrVzAGIYgJArTqhnyt/oSGqsWvX4TsK6psAqjhF
hN4S7CihMQpcdivMPHGkZIr7z9qfoSOFIegF7wXjyDoBRYH4/6R/0EJJS+eprl3qbF5ymXpCFGsU
BRAdn8Dfqjo2bWvEivq5IcIMdsV67RCZqJ+pYbD+69/tVJGVoEBRMLj6svW8xxOapwYJPSTYuo6s
OJ16Ycjcx4kY9LmUR6u8lfjbv83mAQL5Fn7ck4vr0ZwmrvoETGruaLaUsdrWw1d/QCRH4Grdl3Vd
prZf05PPcGnWvuxehjMds40PnDp1ASL1NJQIFI/+VYpNuk6SoJ9oDdHIcZeErH9M4KcgNJKgB9eW
Bs8kEijKB9U6OU7CzWxKKswlo+nkTLtwJteq+lTb8B7WBCHzwPvWb7YWklU2RCd6d30X9A4OUZl2
FSugfVrvIss6aTY0jvt5dJ91gxLk3q/LLXnmRuMpenVeKDqnameqzDcqtm1/BI+08LQLLTRRRMUp
GezMehlJzrDgOO47dAwNwQkh5Ot09AFJkH6033NeAypNFjqojEUY6sHHtCpul9RLTkRJ+F+Ri4Ks
UKlMMGHiShmdvzV0n1VVpEZgT5umF1VJ7/3Fet4jHq7PJ+ztCc7ivGgHhaqb5cDwmqLrCeOU0m0f
An9VzBAqBcUVDX/RXE2jzERXrOmLxHVn+mi8JxASwgSnbEjhLc2prnFo8dOve3xZOQziHS7ixvtB
Xi0R9COcz0oysZIsoyt2gH1ooHTb01JsjPiMNxPmX3jTMvatj2hQIRJcgdiU4vAk3nA1mJlYIt6/
wpauUH4FwDXv+UPcpgi9c0duDm0NWH9NWRZBrqYzUpn6YKlUdbCJP2z1HMCLhiKll8U10X4Fj7SK
jcyT6dRJ4ZPXDHkI21lCmhWr9NNvUZsq/Hf6S+l9OnuIYToUtOOifYNglcZzI1426lU/V6Pn+yoC
Nh8lwEvTOLaU2JtA7grTNb+Qtlj61ZLktavHNImuJ067PezKXlu9EwIYeBBVNgKufXc4CSi80D84
c8IIT8YgHVsiDcCea7i4VXAA9rlyrY6YR/nh0nUTZTg+asIZ292980mUYe60BPaOw7JyzMRXiLY1
VGv24A3yehNzMyTKc9R6IwImvEBMPX9CvC4rlUVO4iPEN0OEgX6/pYXEyxxnlQYNx+9y9dI/uKP8
gC8lKUA3V850ZhcXMMcEEiCBW2ovS+9tAlFx1O2o3MsrF0hJMDjPL+kWpCtEfs4WgRFHgqnRNPC1
VCKYlR1NGl6UyJGX14/ttyTJ4riiUbwF4B6Ok9jXpDymOCOFfjZkez9TPB86IM4u2iRtB18JfGD5
Dbytf2jc+0iyTZlBEQ7x6GjzrTvELzRwUaLNEIor1hQ9RyUIXI6OTKUsiXVyiW/D3ixbDkZI3MXK
kkedpI40MOS8ucZMLe04hOlWYFx48SV4XihhFz+YGS1qwhk6kyZ8k0G0U+fHuA5mQkn85QvwI65B
te+GTR5sfjOXamE5D8AgrXHSoZULQAz22LNJxpLG0PxPel008Gf+jdoBwvSfLbo6kifRG3CWC2NZ
6mxfxx3tWjKH1mXOYGUWC5Qz9F2XXIBvyqE1PG1vY3V/5Shfaro3DO38dm6hqztU+a6dWleHKHTS
NsduMVEP0mdj0SEhHbp2z/wvH0nkLFp00ZE3feXFsPF7wARyo0KG/VL0s3rasGqJam3k8hbOkh1h
Ol0lCHxAGeGtnRC2qxtgSJNGKxSffDZZAv2e46HGLdcVspPNgDEDRPk62ZFdu9Qw6bUOu6G638ol
c+dL/URnR6JU5gqodmqvpHtsaiy9SRijrueFedKWmxStae3wVsAqtBWsQu6eK9/pJnT2olzLrRTw
rfEZe813xCB8Sf4CJjsV2tKWHGUdijvLzqHEHT38513xMfrXidrQjXxOjAuaFgtdfRrOK2AvcJP4
h2vTZ4l36NlFdtaquGCb6QUbKASYs3ob228gWIyyGtQ0BfROy39sgRNDU/n1ApVDS1uo0vfkw0ZX
HS0u/1TSbpWyXUOaNnGAeXOW8MEJB0bDM1C+6dVIxdEIPlDj5smwaZDnrf6BD5AQ4+Q0WjR4/vFi
xWhXbVRos0jvN08nO61bYsQCyTUNldNgm/oqeIhXHeeExdMmV54P1nx4dt3VYOa2zFW0nrpWblcX
9hGstNhXGJMS1Oi0Goj6YCUjZ5K4g7IdLwVnhghceBlcuBcfH+NCzRSMubIBqQZrPPTcIez5VhVw
BZ1e/uYz1W6zSwYafxuFIyQMFhDqADB4U3Xw6UhI3sYUe5MbV7CLfcKLQ5MWWQ4TLdzK1XI8BmbG
hkklWG0ifbIzyDIEywfE4vOUCbeGX1ZsCEvDqxUz304PwHYKZCrvkzsdFBNUwb08TxRS9DfzpT7M
NwcTizVNfDYxz1zLzs7U8+XYIoCCcluzgxot16/rnn2sXD3TOovMCMC/1FdJxXjYcg+YJNVHwtUr
hUiZaBDEdaWlrXDa6Bi3jWQZ1NYmCWzXbEJWYuSvwxg6MrK5YMf3OZ0GDP1ziBuaPJG9aleUYJ1/
RavPUirSTFYZT7QrKaHO9rJLLIc0bzgIKIoGCG1XyyUVwftTPabbX8jA05JLjBdPquPcHun6bKCV
UHMLVgf/uiViYM90H1ndvvXl1nXTsZt2xsZxgC+PARAFDvBlR7utbx4QtK5cuq4KoK3Wq3Y2MB3b
tfrazvVjiX1inI8NxpgoDKWtB+LPtsOFHgfWeUtBhRl/P2xR+rPAVeC7m6W6XMza+CrRC2WsL2Gw
EsULKBmnu5o2ZH8rSCUYbNEis9A/glg7oEEmpUMtwfFYEqcPR87evISdlP+SCAB5jvJquRI4VIeW
CQE7zPvEk+eG9f3tlqmGceqT47aP2caKlVZjaUkCbyWMCLIrMwGNXfLIoHutWiYFCWaMRStXMP4E
/st0jbeNY1+d+V9sOzPWHJUjUOQN17esn1miwFcljj8FpJ2Wz1daRIOgNwb2TiAA4qRDTVUpVCq5
aD6caqrK/Op9wvDABvT44u2EirQ1OyEiL5VEL6PQRqvlCDz/NnNexYhAMvPmV3COqw8LjgvEfXMZ
VnEaP6GItFT2d7WVZxERP1nQ93Bh3f09ofjmRgWmljSdHw2nleNxB6msH2oMPbRQt9GqTZPRSkUv
KzVirp/BxO2dWtgHXy7Si3JgWCK6UQ08ADwLXdAPL+Loy6oqJLDpgViIwBfibMe/ox5tFnsIx14c
XyNLyTXFcRZBcNLHxVT8Ia8w1x+x4RjZ3gTbcdPE0lSACH1DYAXkXmBccPMiCVi1uzIiEQkREO3l
SpUQ9zWJHOHIggG+r6Ga0mAlbLP4aLDvlhAKv2Z1OyT76/T2oYzG3SnKWnhJW+CkfKvqTCqDq0Xk
UR7Q5jBa73cKuF2zOrIB54OAs8rhyJ7KJ/j6aAz61tpj23+O0Pa3fogHo3f9iEvdh9oQ0XMVGw67
k9dF343wEfOJlghKRVyfeov7h6YTqqvhtebXxgQozV0vGBXVditVki2559BkA/bsxb6Atyp/oxyG
ZCWRwf8jPQcGvzLk6TBevTXLtDL2+LJqvL4Rs/QsFVGszez+quTNSUWzQZpCXt4iMqfch2PfxP+N
uqFTTZRASh0qcj/0wsmAEkyruFCRLSSW6Xu9fhFpiRloSd7UJo0dOCHZFDZq3za6GX2Z8gLsT4Kn
eQvL53NUblNgRx8jdix+LlckIl4QzN8nMRhHuihql13cE2RZZMPumIH6fhbZBNRQm46Xt3s+UQbY
maBcc5FwNUHPBkY5TeFxy/kLo3nkL+DY0MdqVmliWm31yzPKWCUFNgjGj7+zDvoplaznOYGVvYfg
QQ94a1tCTKu5u1BIVs9WkoVg9T6QicTQhWC1psWu0gXIOBCc78884g2WhMzHhw0Y0siUZ8xS4Bmf
BU20d4jawYS9nCtpXYz1883tCtzprfVKDqP/DOTzhXPdVS6D01KWfbAmHUG5TgmiEkMUOwFvlk/C
j65RmBG/GQCHwodfhtkENhxccYPsDw11o60pDxmcY9lFKARTikpneSzLQPlCon50oM3/BUuXsE7k
1u2RecZusScFsC79INhw1vSaBIAvwFklEU6vdhlM0MJx7r7Zu73hpuCfu9Z/Pi9v0wwMe1g1PbEE
aiBD6UtNHK5gUbCKUWid6VAcGdHJ+uAFyaqifsPnozLvOG8UyS9KivbJn+xKuIXNVmp7M2cCREDE
SUkGN1QfBmoq2AYJWNpFwhmlQaj4Pig+dSMmsMQAN5bTwR4aqZq5kqGjZ3pE9UbZdrPMVgLp/20T
YmOo6H34e32kR9ag8J4N90M6/LCoKHhnB2kGVN2BF9l9hdB1WDvAUyDgGJrfWS+5lbdRxInCJNAl
ZxWPT+xSHeUKcwvndt16paN+J9vra+AeTCnbr6NaQuabw5kXlHgax832HSq2SZJsa2X0QhmyPX8d
bxbNhsPirQR8K2EMdbp7Rv0d7dLSGJPOBTCOrBAQJSiv146WhH6xQiYxB7xj2MnsCEV92YqBCy28
jjtHqc+/gJi++HHU+JN1eb5wxPgBjML5uYXo/XovdDvsjj5xIFEBcQnfcR54W6Aqunq+kATVI56h
Of4Fn7FzPZMBGOgIz1rJ0ct5TDDsQX3UvVkthD9Z23Uik1R62P2r2LDK5En93AvTRt5ejyEPzYX1
LZ4AzJSdXs1SsU8Eza6Ci2B79G+bsyYLej/ZSBkYenM0in9PINneExZxykh6FEmm4EsfRrpxPHSq
68j2d0VTyMldbcdcvjVQkHUCgIa+U/7drmRHafxk8JeFyp4N45Le8xSWPKel5HcKDJeQ7W5aUhCM
XIUTZ40E3ozbOLOiGZdAg/P07r/GoIIbpIH9nTUv2Sat10vvQfDF5O64PgUdcVpBA+v0VbMUeBxG
pyaalgb3alVyDKwO/GJONh1rTryTNJXPUQ486DCZdPNEfPv8BdcV+YlO7YPB4hDz4JxCgDHRIKrS
XmdihKPU0OZEtXsJJokT00ZTqGw+emQ1IXX7Mfo+NeXDn/2Htd7EMPkSWEBebWXDNmCMYFwyysCs
ooeSyPDkFs9uQUed7/sgh2OAVp6tyAfmnO40noptuhIUqvfFKBPQhFaTI3x1OF8HNnlNR4wYaWZK
TBhOe+QAheAXn+cQqd1+3QFz0/qJT4hO+dcL+eO0T8DrYGRJjL4VdORZ5TvH+IBDHsXE1t2F2Ri/
JydOqzu3cJpJpZBr3xNqz87d3oJsc+Wf1BpW8uc3VkN61mf/MljjGEmPN5Ct+86kiPQg8iWC85LC
bBnF6A3lrmj24/bWuyiruf1x0fe9z9oNYWHI1dK239FUnNg2PdZy9Z7/uHbXweySzkM6B2cdjYs7
bG8eio8iPya3UxtRqnFjX9hgszs4myvWlcW7C60+n/czBdESq6HYm++J/LI8SX9vlUU3XPi7xLZZ
IbYka0D++8R2mGc0yzWY0mhezL7TBjf6XAnJ9eIgUri5TDRPpGXVhb3qZysf8pwP2xVR6h/JxeQk
5mk8EOZXHTt0Ks4ck47PaiLHDS22E0WeC9fI3+zPYbVWHLuiVh00r7nlL+FkzM+mobs4iVPHOqoB
q5SLI5lyuokSL8afBIZKd4pcqI8b7ZiKYxCJH+XeghNWPM9aVEtiBsE5NWe06x97E+pxnix0AVI5
P36qf7F14wTqXfdiSYnST1WK9OMMApJYxwVamLpeRGi1ybms+oMKcvTfw2KGTeP4gIkAC+sypLJd
2F7sL1IVeZIry0syWjxXuRc7ug2IE8tsAr7nbTWPaBN4ORvRGwd7GNmLHmq8SSGA7zKAwXqV2cDr
OOSbJSBnbrndHWnGj/wlllo49wB5y1ItqUrSLhUufyw+mTRnXpewDxeqDlhx/f5rYd1gPD3A/sOe
Uf0Q36v5fV9vORhZEFJZ5h1I+IZGXlV/THBkHPgdVTEIuXtALy1ZkEP46OIpDq79gLZKdhhSWWGB
YJ172272sBpK5N4gOtmuLB/Iwe9cklP6/wIn5/Nn98slilc0YUyftkD1g1rwdNjBWFplbm/BeQY4
w7PcHmbao6rTTpg8DFCrfGdLven7zb+k0fpLwvvSiopfhEyKlLhlwxcKAZ+OEHGljwrlykz0Qixq
VBA/HQcBdhSGDE84uxyHH8nJUqOEDk82ueSQE282fXpxJ+05rvJMhVQsiYAVefmBjH6DRVO+22MB
vjqTtbwtOToCEzGSuLOa5acdVo9nPb2GbpkZSlUPaH6rwbEYy7w/KMcrfHtC+wZ9Pj9+sSIdK4JJ
8X3ZT7Omn74R0FQHH6UPClDy2yPnwbFMx5zhvpum0snfLLq7Cgz+bNPEkZe3TmwrOLqQSOUyBIoC
uOGU9LYYRil2GsvNszZyvPjL5wCDL6N3y4t/ceFT71FqFoY+mn0i0AP1c8y5Ir20oW6eY/eymVP5
EPM9LXSsxN0a8yQOnSaStnxYBsA9DlkbTtaIiqjCnjRrZplAQfC4xTY1jE6BFIGf9++Z/0gR0pxz
EDmoBLId0G3fBAAyUkrysnSdlTUMmpYrgek0ezYPfEKl2A8Wqjj1rs6/nmcHr+MLBxlaCGtZtuYt
YqOW3soZWuxKUF1HTvJerk9k1nP3AjsmtuV1RFwzhvCHKmw2umhg0DZdZAZeVm83bEGYKxM9YVpW
HCAcLK2r+YfcMlaYZepsDbb74l6wyX2IAETAKW9hKbxzdVx6xfHvZX2lpYyAwJHTF567hWjmTVzj
5+Gasl9IfF8IAhLFph3V6Qolg0HrUBp/vXJrgByyRHXMGFpdkEmKNJqhMv+ieBezI6NpriLbYy5/
q7jqzDC1S6Ujyw8SYsdKfihca0B83ysnMJM+uBRshoRUdSkcY5HP2ZVRTgavLOHqwrMViyWPWcJb
hwwZz5IP+ZkzvYUYf6mrxCIp1L7wmXELdfGtHdZ7dHxoN1QgdJrNDUZPZcoTryL0SoPzJuu5iVSd
K4UMm+tobSW8/zfaXBWrFOVWkloOOwxpoKcuYb1R+HQugD/had3xeMK7ll+DWDDrRWoovqU9GzRP
sALHlRwz99WcvfWaiqpOJRItaeIMymtsUj9gOpghdH7KPW+jjsla8k/kAybZAmCuYsMxEBrC/tia
lnQXiPYa8cDXL1hdoUreHrjecW7mjILHp0ehZAqA1No62YqJ8E+fo8qF32fzyA5jCkP5g2QQe7oo
ou4mZ/cqmyrgjFi//w7xsMePZNEP700x6fsqcsBIyvpDESI2NhByRSe4Hf9nUN/HPWEKTKEvPJj9
PFOFvDZPFLSMh3/eSogzwGuYXLeWq6SBdj3zQjN3+M5OYGDy0y+poObvvt8hg7UZQTTCBTHSVBUt
iSXey+G+lbCbNnTBbIDDTIlSmiR/w3wOYmtSiniVX3HiJhoUkV8BFpvgz2qh0x72BOs7olmPkfUT
ejIR2XMVi2O8+WZ/uWcECf08jLHvj5luwe+iV4AmpLDyZqo5N782Q1Ap8NCVI7SZXdR+0vKO90IY
3M4ZulyPEWDSzEDRd5EXUq7/CLVi78dpOOXkRhGUUPVLVyDt9222f+/Dm7SsmZou67VTNE/By0xi
zu0r6aGwyS8Rqu/oOvoRkqbC/qLiKFHjjKXDt4VkJkIQO0KJw1a2+CkHCssG5X4pWnNtQwAW5i6x
ou8faR3Z/nSCmit7H4unOekps0SWKIfDlGeDbPfdfhalId2zkB9UYfamKFL6VlZfyMbFGpJjnjXs
NYyY94lzb3iK7R5MtMIwNr/aV9UbOHOmA5WJwyneQRan4jHTNzlq1qqH4cTi//wzxdFTRYypyuKF
MDQEI1x51WjUKPFJ1+18DSym0j8II8SqF8iYAUJZcfiiJ8bUCSeO+swQYXbRGMU8F0D3Me8ZwwCA
+WeI/1LAnN0itHoD7bmT36auXiGCNzn+iA1xIjxy7CuKnK6A7mPc9i8Q/pHGdDPDgHPdssl/roFw
71O+zuQAGyufXorLKNx3Hh08cy7E+KxnmmSFd+RdumLmZFY20hLzB1MjICE4ateJzECfc+srVgI9
b8gxFkQE+Rb5oC/d6Sn0qtuEBgSXFQIo34CkQns8PLPjzCMf/4KnrKTkKUk8FGsKtO4VvbLujKlI
zz5LVtwDmFKWEcef305tU1I/tiCrNZ/9X7XXAgVPgXRHM67iaKhugLKd9iSTbSgpoO9Pt3t5jHiM
HxqyCEj5jfA4/Py8BD+QmLjZ9H7uv/Yfboxq3mM/WMuRUUTW2iUl61XZJiSNLjOGL14M1ov/NkD5
YvDhSaVUI1W+hapQDvT6uxyGvdVkT5S1+vq9XHKRqgUMr8gh+NAQ6BvYPvlsbqRtIinmJMWEk2nu
kNYc6EoVIPbyHXz0epU23oCF2a6CHHUq5pjrjEJo4Kyfzw3ZifY3gh5fJZ87odEvwIWF9Certvkd
MCH+eEK3u9r5M842DX3MeEc6mba48kZkzO5ox8U/pHG6Rxxi+q7eECSwKIOhiprJTGFyW9iBY6A1
+BVCavG4xtyDT05q9EEjifc+qNPJzBGA3Gq8Bnhm8o+gbKh3MH82aEwfHke11L2Q7xzbdOoGZcHO
I5YkHgjSSjxfSce5IdEqpVhJN1CclfT8R3t/rNWDezKIvnyZFNlOQFlVt2bvmy1J6VoUpqbkHR8c
2Q1NXXCmrj7zRZV2CT/qD/fUWXqDizFyUXoE6tPt32EuwOU7NS8gcNwmog7JB37wzuOwdBhbWTp8
4GVDZtdNkZP7Ai04HlC779jeYtf2LdkgFRdqgK4d24vdoieYxdVuQE43CWj8EDxkBJdeOnTq4u84
V869cz6GQgDFaYamc3VURVFqgT2hQgU92XDCcOwYxBfAyQOQCVuDafmwMpLJ33AZEfg8kn7XGH/s
wH1ezJhwQB+q1LFdd4J7vyXjIvpdU8Mvz38M+O2JxxFSqsa1I0O0N0+yCuk6lov+0HwVbDJI4AVA
vHq03O6OCle1dg0GGNxu/v3zstDaiDvy/nQ13vnROHcDIKyzGfWi8LDnsDyuxAG73AxUVlSnXmwv
tNzuh6YCO4G1zRp/hLaxqrzgOiJ8ROlZBtUSnm+hdTlzHyf1mGrMOgODJ98VWkOKmHBlcVjlsTc2
NAatRKbyWafxSmb7TMvzNWabjCC5R1BJvuSKlVdA8D+K+LLe2iqi+tKHMI5F7jEs09TLgfD4j76r
CJMY4oCO1dT98qXqfcnsLy+M1YY6QojbGAkeRQ3ewNTvZx6trPs09VNHgJUIZHywI0Z6oWwOOPEF
PrZzSrlXwzseZYqNbHN6gjkB+kI4ffb92Lmirl5hx3XMQ98bA1+m8gUAVt657lJdh8wLrQ+0VjWu
jNtMqnxGnq9OWBol3j42j1/9CDRiB85nj29YZIAirsiCTTtjH0V9JMJIpu1AgzFWeOmIQhSdODSD
ivhi1wasGr9ulxBWGBpXVEnQf3LCIpZiSxv1vbh6mR2InaodmIG0x5XUCc+EB3qJShe4K84NIjIG
SRXHPoPsXE/jljTzphUS9+2cKqJlNC5TmNjdin/FLA9DYmHfRXtpXE1tpb2+Uv7V7bJqFEe5mKxB
iDmxNBRWnpD7IucQ9uNWUOjrY8485ZeA5xS23IbgTaioY7oH319gwAxV5ll1Sb/wTaUJSJcKiRRR
IuhUpP4Biwxf75vyg54Kdbnlloweny5lqo8BrZchzWb/OEgniaWr8+wxbpXevn47BkZPBFsYw3SY
08t0EOu9Kh7drs4t8N38MkPFr2WEVIjr0ynWsG6wefjjl1mKBgrdmzaUfdEcMu2TS3YABW2mfrT2
RxmYZbXfW25xTJMYzcWV7KXnL0WqhKw/GoLWfV/NRaxz8AcxlZ6hO7cmpn4vPp/glhz/Qj47rIYg
N0PNwIYdfU4ntbnVss3ErgJA+xdg1gilj0s7T7HVn4C9rRwI0XVhXTJxtmIfu7psRQwXL0zSI1ki
mbdk+CWQpFqymiNp1ZIy+uK74QJGtuI8wTdBEH1fwdznqms+l6DuPJRcKRrHb/3wttKsx6xObntX
lm52bi+QcURWPVIikrAEpBu6uFrI2VqK0or6/J9doZ3yXYVWEr9dyMhvxbDZLZnJx72thUOHcgtL
vRCJPniLxG/yRgii/VmcLNCJRpe05sORM1A/gWEVvlO0zdIXd1ZtwRPaxY6jnbH69v4Qf0AUSP7k
Me9F4g1g2JxvQSi5TxwuKCA0HPnfX6pCZTZVaifpenUxvsZQDtC9fuGNiF3mKsBeIAOWJAr7r6aY
OTTwsau8U0H5XcCRXewgNH0CkXs+6MA3CQ88hR3RsVcLW0e7f1t/3mKkHHR1P3It8VVokkNH+5SJ
EsGYz/MXofdfrXCwdMBhHu8D/MkqmO6vWgxYNGwrvYVL7iLbFhcoK51AVIX0ELknTnCoifbMjSZ9
6pg/NnFoWxZJwt0Kgp8K+RsqdUOK3cEkY0DrVb+ESWZYjbxzszBEgyJFeK6gnHA6We82FW6WWCDs
3PTgH3jsuzrmG8nDe0MEL+hxiFAHFYt+dP54byRe20Xr0HOeyRaakCwXlen5Oh/NTfTT1V/Jr5t1
KT/tS7TOYCbL7ufZYTn9TZu048NQHNm58JmDgM734/oIXTGzSsgZln+uUX3ldTMR7hpXeZQsOaTY
zMX4QsMOV9zh6Tc4KFgACcpqguJjZouBPNiRzANEb2K58CaFy10g13dGH/aBmdrXXKBBmNW6UmG+
ej3Ir4MQYb/kMk2G0Bb3VOQzBMIqx8yT0NvlFHw9C0GSC9YzsQ9WEvRtLU+3tKJ5gFA4qUiFqLiA
Q2q8sx1Gaq9kcY2lRyyMqphNtTzpZKvHFqCMcFNgxH8dB3qNRp1QWiAOemdqncqurbO95JWmx4eE
vozQ+cHJGNtuRbGcQExm2vKwodm6DiH6N5WSoUgIqrCqEa0lqjyxuizDV+k6egWUj+fktfXVC7MO
gXe4clfxTiH22L/eZqwusMVKejr/0/X5j1mwHJFgNkGkAe4MUsRUmANj4rk05nNHJVVBMppxskmk
vzEEtCrOR0eFe8KRV0m7YY+OTzNOvR7ftvI0PvPMHgJG5l+sCxLuSQdRg4WiHJasOQvoS/FlL8mc
q1UzbnKZPH1cnLbnpJWKEI/TEKsRXjuBzuYf8+KnKFo8Ne6lMP90iW+j7bWWCifU561N3i9wSl5B
aCvENBz+FNGWTjjon79uATHnsvy2ufgqWNJUmME6eqwKd8lJp6wuVreNPPkDHiPfDZyJdY1Xpiro
/quMDddW1p6sVG05Ct1HnkQtaAwLhR4u3JZbq4H5SyDFyfiCmO2wCRlN57UFI4nzdUFyTACZJ90t
vI04vWGFnT/9zlf1VbjST5z/UE2esUvS92e0S5vT0Hi6oxtbzjrwHCUATxE4B9jEmjNFx0bch50C
rFDWICktouD5nYVrHqt0Lc2s4scLeQ6HX7u1tb8fSfeUHcJ4+oDuo/0rvBoffDUuATgXDfBTImN1
AwK/cp1WJOWVSpaJOowj5mGeBp3AfCRnscXy8Fp86p3k6dob/ARzgPN7k8iQpGR4EaDjvjekdJiK
ieD221QKzSK089dyH3jMYBdjJLrBWSlwStcLek3jUaanpvNAF7zA1ZJa/nVxD/RbDoUIp7PAl4kV
G+eoof72WAMIoaZTva7KX9hZXxqSu9g8qRstCpM083mDl5enlif5u61Q/rHHhtWwXWn5WUpscWby
hIHRblE1Oc8Dx8cjFJ5opjwam+YrvQbSGqRuPTVWq1+C4wk7VkmspiXbAyfPorbMGwzB5R3XelEQ
8FFFcvZnvyNJCF1Gq0EKgJ874rQYxX9zHwUxI0LCSs5f5YlvKI36Fsm9r9wVdXc3kDUwWgAp2sck
8ODvEimY9qo2l0C3qUjZkZccbN27KGUPm0fLpl82cvee1C5o5E+QJadF4PKDNgoXfBECSIEjdgNp
YV4szf+SC+NNOWjkXHMpSX2tz7W5XNFdiBEBIUJsUHrNY6BZ9My5Wa9BoQoWKCme+9B9P6cicePW
l++TVf/7SCZ6K64N24Q=
`protect end_protected
