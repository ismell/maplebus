`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GdkbOqEHH1/OPqsOQJgL4T8CXh1hCVqgPq7JqqsJ4KkkS08AVXAdMANNwsQPCkBLYTBp7OO2I9P6
h5RgZG4Ulg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gMBJWIaHc2sBWElvaHj9h1q/Dd6sG9O6rjxLUnXBllbrWhqyOz4E3VEcVrxfp4LznF8b+di4VTKT
IuGAUAosLEhkRr+tO+K7NsM6eO59aFggAndoIGEZUMuWaZXguP8z1S9xSKBed63Od0IZu/EDwkom
c5AWr6la2WH4+kGWfZg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4V75V8xK742Ik2kJ39rCuWV0xmc0gt2n+z2QG7fVm3iXq0JwNFZxWYmGTewTtZ6QQxcwF0b88T8
7fo+HAEU6A0/ERVEX4vdA2mg5f+yj8P084Ylo0mNWjiQPqFHdW5MqQFr00dLBLSULsji5kYB4qAV
s45qlN9YEe3p94tzQYX19O9XaCQfTsfdoND7VDlMnZvbxhzaLzoxajRRmqIyIXl4e8Aup/sTZqGO
3iBGVqYmEllA7rXlY52gItN9ZVStLZSR9Z4H4jeDcSj+j2J7pAR0GlQTTTFgzEicqJYmrmTV22y2
mUXaqJN2U1HzlUzOFJh1+rOu72tJ/fuH54HHEA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pqm1pv/HcEOhPJR49ucG0Xrc7T0Ejg779jz0pHpqnlN5qlQ/7ulfd2PeEFdcSUpxXQ3vzcwamBmC
suRYYGQFAuiTggz8yk32tMJu/Sl9ZsXFD+Pka9qUv3cDLDqPi4Kp7L2oIRvdqzSBE6zmxyS4BQ2H
QtyMBPpQMZkfgOA4zgc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lPV++dRwlGlowsWO4jLluBd7zpn87Fiv91V9Zm4SaQ5PYyWK1ryFg3vewUhmnZByzknknkMepnXP
qT8VZ5hVJ/VWZSzYTEdGCuZN66R6VpiSMBi6nOKQn3NmVujHuAEids7890JGgJ9YRmrwgOAs+mKJ
hwFz9RACZ85rX3Agba0WhKAWQCW4tV7xYOlbnGjxr6km5syu5rm6oo7B4lwEFbPkYbFCZsjbDPhw
RhMFk9dYRrYJN59qOgjq4sFQuoMKusf8GpD7sxUfBpTW1KKrWOj0FGeSmdGFLfbpOASMdRLrwTlX
tLfdjhTKnXkH76AYLs1XnInryJFJce4Oxzn9xQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30400)
`protect data_block
kW0Fp2UEdV22JTxzjem1YUt5h/q+sMN0McZcPojRN55u9MjNT4B0FbupTUqZnycxl/cbQve2kLZ4
3HCdcNe2JNW/h7ZEnTP68GMIxXJCk0LwUZB+5bLk4nazVZt+KQq4JglwXxukuVNxnRWpOJuxOdNC
gjTWgfuzfkHVrKMrQGM63zE8jyEv5BXxM16Y/IEy+2QSiHKd0yXOEQQFrESwV2gRJBStsNDhhKFD
nq5jpp0fW4F4n4BrU+vivaAdUxkf4zUiQ4bL7wZ6RWz7zEsia5F6fIhoVCPjVX4L9tmvTLbbGziZ
oz0aB3bPK8Z8oFDUoSk9uzhL74hnhjIoKOcR29MVkrxgY1qFwN2FdaqWpzsXy1VtIlOA5zm9mhi4
ru0ktKkvtEyLspvXCNF+/c6oOFKsp70L2Uq0k8O5Q9mOWzMuT7Klb8T0Rwdsyo7u2w8u73m8QQ23
uObp3qlWZACQd/wkWyiGdeC6hsW2+XnBN24ORBnSK90A1oXhLImtHQDklQcSbPaPS4c9YiG3Kjct
dor6qrGR+YjhMnGrRWHk20/6sLbquyelnvc/z01dTDjEQ5ks6S2ftXq99oj+VU6veh4KRRfyiKQ0
gTqTGj2jhDVF2fsPcfVoJFMT18TY8RHkeZQTUatQgNgBd9D2t6zGGpEPuQkSPEAP81tXkh7sj7JK
EueePzjZzn3jMBXaYVTVh9VzKgDwfKYYGrzW10GvRzkGuZkLUjNaLKCCxwGualXPoTQNitsWIA09
ayXxYLRy+QVet6K9DKgc3/sKuOQTWw7XAFJC5YgLsxYbpZixaMfpYVAT3mO5KPR0l3SbUTE0ZntY
mYQ+/Uu/zAUgZWltxz0GQmhalx1VaQ/4G/sZHWsEwGaA2FcL/giJmU8jPvRU1C6ueeAzoZTxehd3
9X/eGrYgT8lsl2mNrjyBAS8n1fsdqQRYEJLG03YFqUHNY2PFY7YvQDMCs5ptdchX2V2CqLsypMdX
pwqM6c7ZGip+sTQHzGWqs2ORTtmkE9u6WC4lh/AaCt+ekPRFnIJRxh0SANrzMkrm0S+yzW8un6mk
ISCNNcb1VaQXGF40SzVt7TNjEfutE2lfV76dTdHX3vpY2y9coB2os0CiiNwNbIGyBQ7JjvQT8K7E
uL36+7s3eU1fgAN8l/4nH9VjbmG9ERJB8b1oU9b/HFzOIt/qY9+aoBlPx44tZ8I4HybTv6jJ6XHt
NFhzxrfnxGYfoW85Np5WMQcFMfHct7n9XPne7u41KB4dFPm9KD2uRI4gmrj3+b1zFJ1KVW9ZP9sp
/uh1KGjqWzKujpyW0o/5TNP9iE5Vvg1WoA03vXLiZN0Xvjtmgj5M7nYtZ2N16/SbB/4WCb4f31WE
Nue1ePHCK4I0qcdM1fdFQFKd4mBUHVt3/36dWlfzl3oJA0IVb+LSa8NDXqIje3l/IDD1mvSGMsRn
rqgs40gbRXg8xlJZN7HXjHcxZdmv0s3FJuBZUyTriH0/dmFa25Qq0vUzhoKXj14lP+klAGlJuIui
PISRq+S6Kon/WeFtpnQmPbgT1zqdJTWIgE/FeVX20Gdnn4yqU29VscY4yf2d5HiI5DzMKBLIG79f
1/jL/2RzIvxnChckZ85saWHlVq/qo3NVkTPqoJ4jAX6B53L9Y5mhn+6blyRthip7S0kW3+84+2f1
WtVXdky3q/iHh9odC1+sqAV0GXUuwFpxSgsSh5wEXkow3Q5SFPpLhcFaWNgowneZW4R+IHHl5Q+N
8FrHLbF2h75Bvg15n+rogNVaNRxf6GN9Y40Vd6oCeA9+7UGoi+6RVUcOaJ6M9e176ulA92cjmURm
+bolvHazhksj5RZD507omUKrRzdhjB136pS8IqufRiXPl8omCDthFzYceS0p+PCLL0zKvzdjvit3
RJAAqPw2zQ6i3VAasAFshXnEs9oExQFoaYQnWskw5MhZ7TaH6AQ5fOxaqD4O/Ely/NkXHesZVLjV
zWlfsH8udP5Ky68YgaKyQYgfQivLefTKIFB5JPTWdY6H2QbDyhH7b4liFpN/irW9CNtSb6HMkbBo
u7LAYonfErAItrxyS3LXtWz3nIzDcua0AYF/9+cdLhv1zrrWA3VekP3SrOHZql6B7eBiSQz2Hnds
ffsig2muzFtTp/09uvRCvKK+4HBLy81qLDvYB0yEhgTsANXeNk2l8+tX2Sa2LLLSMaVxZHLzgo7l
3iMT0A87m0bj5STeY8vz5g9FzZbHxqixVgmkR7SbgtUtWBlZbvG9AENxGez/1o2m+EucRF9Setyq
ZEUdiMNFFeMgb3dTvcpMQdw2Chn4QAC53nsFSConl3q/HI8AYwcGjsNzZYCTO08juMtEw6VrNDfd
7inxpYdZJC3uDNECTTfuqatjHnK5lBfVBFvUvQzAs4MLcE/RqyZyUkdMxwAQEVinFGi1ENbJQwlu
6h3FjACzEcl36ar8yPW3arsT7CiVa5utJVjq4/Sl3u8MbQ1oIr9mqikOoWbEVhFzaIiFGvYMkXJa
X9UYWxzjTLyUYrwmO2+jsn0R0jjk8mqNomAxp2yW+zbted8CSnMmVzwpe3MJM74DCG0/TPXFsm1D
vXbJdq0EZ1HB7vhWGIi4CQKYt4NmhBPEXJf9A7Jg8kQ/LgSmwpZh6KOrT69q0GuRBMi7Zfn/q05m
Q+ai/LUk+jXLcHOsYdSHSmVLz8hZheTSJto/bDIC01EWVtuPHB22+Ie7ZNR1n4c8UvK/K8TAVsp4
gG8jStkjWJlmtT2DhTIfWQ31ebT+j7Bcw4P5AqddSaqF+a+8uNJ9bJ3YnOYTP6H2vFSq1J2IjqDR
1fqsENltWL3ObExXPSlYsElc/dzOeKH6pjYqedwXb+BIV0BvAf4iNgXakf14MwzTGQxeRscG9Xvl
9YinNHH3TrcW4LVYm6zHlAvw3q5ppGEIc9WzGV4vF+mM3Mv6Xg7Sd7voJGfxS8cvWHoebw3dcCQ5
EQw35HvPdqalo5jOis7GxD6rUjyvAq/s8xEZW6mAaNPEBE3KaQJn2ycDTiMX90ZudoIDsErE7cZz
qDYACUsjPxAFJ0pDY29nxP5BzbJLoyKbJY4zzmTc1xKIvYzZnBwR/Rp2HhBH1IG6gFsD1GIMOqZT
gyyuzG0Yi4pzflmI5mjOBmVAy6hb7D6WsQU2Z2ypKKLHCYy3z16Puj50yVG3XcOdYS949tM6fWQP
jyiLlxp3gnrSvH/2mO+rDeQ9l12AqQWm5IcVtFUQvKA2L4ZQct0XbcoCXsnfTsszeu8UReOCBnR6
WyMkP+WMAJUlnss5iG1k+j/SV47UUlZnJJj/+lnhU87C2M0o/w+pXs0yVMAGxmk4JO+C0uBKxWeO
E+nr6S1q80KXrJjg5rGMyEo/0dFiIlVyPxgBOxqhgWhUg2IBCP6Bm1Zh+wXPPrZRnqbgDC1su7qN
7ONQCr7sg3E9x0TAfNdzQ40WhwTJ10vb2Ox5ILslBpKpP7K4oYLSNoYw8FQHRk36WqFUcMbkrZJ2
CZBUJ1YEhEV0J8wBG3Kt1iXG722EAiwoeygg0vhrZZFwj76xZaDjlbldVvx81NXHR0dj/BNB0Y6y
0BukCe68NeqPWi9WqmrO6P43Na+8IjffXQHyRP3mHXqibM8Sk53zOaDmEOj4vofU2S77j7NBA9vl
dykEagksI7sEzfjQtedLBc7TTqLiAhQDfIz29b/MJgAfx0QD4OKPMoiQZ/TXk3XynzuiCpWwsui1
WRA9qWCMtkonajwag96gvd/4mkaezDXzCm2n9e6lj2+Abs14uZhwtCvLqAVEROHeo2dPfxu1/pzl
58DfMjc7tywdDkU3V40XivoPKJe2gMBwo55D50VpbWRke68RDt1waxOm4Vc0JdnBvNlcXryVWCmz
hZLub7fBIPmXiTcELdQNzpkcRhs6h3tgzLMMWsZbC390e9jOm1h8DqNoe9x1Si5A3O5nXd+JMp4a
MNWgqEAQJKvEoR6FBmuB8PWNDjIx/joTWoWop26bVqdNVoHtAHTCd3Qg7HWiCaSQjHBZwjMt3+al
SPR3s+RomJMuuR3Y3ZW2OfsbSJUKF2l0QgTJFTPHDLnwcr1Pk2U/OtKk5YbgZNNICFmxWeFq/mwS
5HvA5MwBkAdWz81jV7OBV3GEecqeU6+efeKs/+J2eGP0wOBRBFHKZZn5ALCsneJTOKgLFW6682WO
T2lynVH72/iRET5/GHxp0r8oVmXlrVd0RCZlxUTUxa3O65d9ow0uL85cZPD8oDrGy+KoHuFoCy6x
y8hk1RM5cntrvlXIiG/aloFxNS+LxdXoaPvGgQ1Q47XOC+sRvX1kvaZsfowNBgjCLDx1mquggacR
lqdHslIspwh+6rL5NRxkAItN2QKrNRHbcwcToSTi5CZTr1ek0VYDMCG+o42HBc6OyjdMar7MVvYA
IjjUIcY1e6J7Cvam1ud75djrEpXEUkCEOEkIJarNLFkPcCwgj8Z+rRDQG0OkCUZlPBMdIa1Cj9B4
Qt/qZZWeQ5q/ArrVOMsmAS/SPONUBivrFJdcvc4RlaoBcCPHsFxgEjvI82Mi+hojURZGuqf2FQRx
CW4rPRIYzidPiXxdQ2tj3viXCj3jurCHr9kK8V1YaD4Kg7o7302oaX+RQeew452zDCtISC92ec7W
t3PbB4IbyzIlaEh565DK/Pn+dVeQSscbKTQt8FgCMdNnnwXOXGcW7qCQXovHtQ3/OA6KFlJ70gqe
dq4m3E2DwuNfXQYKXjnpkrDegixk68DfMVL7rkDbK6MW/B44AVXXGsUC+2fBdCsjoRlR9zRixLTm
sv9iBxRcM/RGCcCEVHbt7fIw1Dwt2JTXgjwT7DoJNqytDOEHaZV6LJsggpsfrLasDM1i9C8LAV/R
nkBn1yBY+QqlsC18PSlLxQtF3H59AY74MCsXOk2xIo4qCQ82GDWwbeSY7sgOGJuWljrR/3T+5HeH
oYbxscCp4baXgwyJBdcNYMAcjQmvQdBERLouKdJ7QXAmWJk0uUAO6eGDIBp0vrRXgDL2iczFXiMr
8OtMZiQAInz5M22PB+e1SyADE9a/207Ex94FFjhRry3Aiqn87uSGzLnh1j5VML7ZPokRYs6+5kyx
H0O7/MSNa5/zMpTOwVsAGEtO83HCJK1C9vFjmu3TKMdZIrazedvrWkyMwu/DOm9ej4Gp1DPRGabb
BU/955K9EtRE9IRXummX6aEZC2J7xyAyp0Li3EWDNGgviTRdh581u1S7GkVv7OAxTtd6SLtQRZrO
uw9zfL/xOS5Fco8dN3/MOqi9xwhbBC70v4MMS+k+aTlACX/wAmJQnGAfPXy9NXsnzkrXxYi8+ZHK
PFEZ2GI1B+0YX501HSLJzOF8ge4GvCeEVZLtQfSe6vBy7KqXHxRws9PmB7HrqlHJUzzMTN3ByiTl
1GN/+Ah+ODGnsAgU90LeT/2rV1HW0wrMkZF0RTKaD7Qigly9ukHq4LMlEvvzQYI34i1Blw1uF6kq
Z32QPeiSDV/17gmKeXPaPQq7SQO34Fj6o1ikQre/hYuIvAqu8ueO4ryg4a4110tTt+vy+Yfcuu/1
tWh4Y0+vsgrc4JMYy4Gkx1XYWWSzIil9uP+n3coNDsoKdQWb+B26WuqrXQFPG8kdwoxRSA2EwNSZ
M3+d+eclYvQseWSzDR2Ze5ts6svs1Y7c2+BclOlwkhIzeAen/SLGTaz08wVkP7g+68RRtlmfD2YR
zeshstOSx4GLZzUrYqtVSnr9Jar0b42mtriCbFZgLQroD4RxbQPY01qY0HkdFGbJ42XDlV/NfZ4E
Gue769Bv9rUXs6QdCrW/UWkuVpHmW0/+JRase+lEX5ke88R7NyVzwZ68vlXCpuxso6UUTdi1zPUF
KHsJq/dcx17RYL8JQA/r+1P2DVxvEx/SBcRxvxFfsEdEQT6bKr5enlaH/M42w+aZ9sNlIrsFqYe0
/yj2Tugv32udE0z/RvvYlzRqPYNIXYD780b7msximGlRPS0kIZjduYcbu1EDescwXIRJn447o/Oa
ziCmTdhmiGhqIrWUkEdKcV9QguvntD7PrRXHHb/B58swhPRBqmR0ZSJGhkJRdRwfJbGEEtlK+e4i
9JZJ/2EP5VmQBYTEw5urUa1EDg4vV7z2Eg7i2JHf5t+VnA8rHcGZ1o0/QgeKjb6o+zz3a7gxyZGH
ZZJhi4iJcfyDmDFV/+kg301DPd7BrXDr7xBYuUZPQenItD0gwiycg/vSi6W2TZpX5lpi80/ZYdbM
E+TAIvimT+WfN/7JSYaPsTy0KKJBYeSoXbFQvaJ/2jdoFB3Q9E6NQ4wM/qQ6Wm399IVJOXwLri9r
EAMWiJkMFxZSpOjbFUuOMG/B+hvNfKK16stGNZLVKhqQolbySYCCjNzS5TU8L70SBNOnSB4+pD26
4ZI4afGCaRAgp1qgQQnFyCoS12K3/VJrmtDSogi2hYmfoRoPiP4doXyGqwrDvU+wQm6Y94B0IdCb
nBqNeD8bAInVWDy3RG6jx/EO6IsPqqVqDbKR8fmz8KFkvVTilye8UpbLiWXIcAjdPnY4XumkwXIB
21V/IMx98QDzool8o6eaoT3hwKJnWHqBB5zMkq2upQfawk9iB6ojTfLaD03gP2IZoxqjTvTiQYDA
j64FZMNgF4j43dP3SNfI9U8jUYUKIewI59f+bNypf7vxFHHw8Bs4g8ZIXapyXmH5We36xtxS8UfD
wEX+gqTXKlv0q8N33NSa22OBRyTuRDF6FSdpqqGfvRA5LayJXRIyoRdd5JyuAj1S1XahSYBFeCkT
gkS2AgK/OhujybfFdJj2jOv1CzQ3AZmMQurqsY6m74R9HCZigw9UQ+Wtjrag6wWtHXHlWTo7xWhy
LZuHo9Qq2ssXK9xFl5x+jbX8eMOufztmSpei07HdqAoHiCfz7FYPKueGWyMD47+G1GvRYGI/oMuV
mt5YhC8ar54dXdU5kLPvORVcyaG+kPvF7i9lmYnpunVimNt301dqCFsAfCrHhG38RseJRuKg5wg2
MNGEMLVHAikd42qS1rLrX95B8wuSHgHJ08U513GQc4yoWYTzqgytUEiQuMCnd3zpLaVkldpNyv2v
+SNRulS5wMORe3mUqUTTixdSsY+QdJNmKfA2Hda0TE9xsUivk5V/S42VsxF4ILymX9dIG0SpDQPo
BqxNIhL/0+ePp1cRR9TEt3Bxm9Pd3BQeaPpRos7LaIx9micWXdsk91MhZo6IxVXe1Y0I2Ruhdr2z
HJ7Y4ctcP04CZpIo4FtuA5jbbE1WQ1H5Q1G1y100vjMOd8wQBHu4kbAh/1f4u8x4dpIeSg80BmGp
4OhsBw/V64JtNg3tljH9VUiQOtlfogg53jWbB8lgbjBwLtRanUnrmytwHQ4jstAIlkIg5GPsSoGD
obbaoVWw46N8ngvPWW2vM5eyJ5QmeiS3uMUpCBQQPQpK8HQ3uNkxKRzHBAqc4DFtQrMJcttb+Crt
MnDB0WvsH+jHX2zby9z3dtxL1fyc6xyfG5TipS7QHA2QycGmBuEGgdeD45ROo+8e00V9e+VPbwdL
2deD7v7IoXrKC1+6lfNLjbMxqmfxMH5ERmqrvyuqH+NoY5zpcoTAbL+gxy+pbVBn7bcoUvoNOSM+
CPyygD0J3/mm5XfxKsureUc51xvTMa3Nxnod/3zkg7vX47Wd3KG0VBtpCgfW3muv7LNleIyaUTuB
o5wwQYuWYoZOeTejwy+Z9rD4bm/+z9ybFwoxNvO2HHisAGf6e9DuD27Ji5xoBjHvw1JXJexK1c0Y
1tL0LnZvM4+mF05sKJya9wX/zqa8YUpoHZVp8lfux589mqCjEqSyDUxC67baqKNIXM4li9YTWZd/
wQcFroLS4Jb1SmxXdEAPevq39Llx8a7ffXW3CRtPWjaMhQl5Hwu4LyU0cFDQAe+mFHmzIYuOKQB7
58RqG/+fvkXqeszflIguMCdZyCg28+7mpr5329RboVWmc2Q0AbxjK1hcQwjQ5IYQ7Nnj15qyWV6f
ipUYseVrGsbUdSFf+nobnTQ688WiPbRZ3GnSIkzQ5T9w8oadmFr/O43nc1+b93EADi5y1q+Bcvjj
q6BDgP/ce37f1IRMY1R1gxDnMqhAoE3nzkYhuTvwSo6F/VU8MNoJT14BgQhxmBSwOe5BQwa+iSFL
eKDJ6FXrAZ99/poUnaCRio1Fmp3BCgGftiauET4laVexLPrpIRXuY3sTa392UNTnsYCTd2Nsna9c
/kGCxp9/rfMxI/srBZVI5ZAcXSn+PRVjeHL5HqcojlAQ2z1PYu9jKeq/SD3Xvkhtd3OXIkGxEk7l
4+XCDceP/i+iECFFoNny02+ixFb4qlZid3FZepiZHsYeq6GCZVRkWWzFnUsVeV8DBPsxturwJU4L
ZELUzaPAxriK6vmbdXoukgAEPQD8K2x5v+o6jal8k/cR4l5ItSxdDlEAMBUXSqeN+oXWI6aVCB+G
SeTgr5Hctf2jIZDHzNO5+0O5inmahA/d5mXh8vNTzkWp7Urijp6k3rU2UHqIHU+xD6f/28+n/Kxh
oTvxtQmoEMXz/H8ZIea6nBMZLlXLzkkIX9e+m7A2iPWDnfUaol/hWT9YgzwnVh/m+Agb8y7AVv1E
n5LqlerVRrsKnF9eT/jGaBlIK9arzJQj1TJ4fjyjB5CIHHthIzZ82JZIUnmGkl21kNp3oFBAypNt
T553Uz62vAVtxEBbkbovY2ieQer91tjKgm9v4mt0M2fmW4hIKqA9obwbkAL792p9LSN4RXrHAtVk
w6CODGfv9j7Zu5jhRoKSeo1Zoyj4ov3Hm6E2mP4aaEgm46YBZL3xyP80M/zyKBY7F4fFkk2jpTTq
jnQY8R5oxSEmcZsJVSfw1Te4QBX54vj2y07jTClJVpmRU2XnYzhrHN0y75Nyywe71Ul/iJlDBJN5
qzYZmV7XVU0FQcDS6EViF0L6MYx4hvaeG/zT8vJxkkB8+Fzj7+C2GLkfgvewkXzd8/R5LMSU208b
xIaOMs4TNeJ8tCc+245PIIKIDsxL0PRfrWx6d5Z/27l0+g2FBO+SrmWpovopBCVlHkjrQBNddVjI
VZWXXRvgii/DU8f3cSvq1FNonUonZ4PKjrEw82ykA7ex0OBv8dinuQ9Quv4Pbw7jY0ClCSJB3szz
ZSzScdtAbKid8ZIfz756hzJrXECnlm1wMB5wZ2d8j31onJ6QRn5PAxGEpip1qjXB2tPEyuvUEHoL
zNJBg/jSOdzjuuNuLeYB6LOyLoQL4QaBq/Zjbpcckq8ubfRjLGDtYQAhd6dfRtQzFHa3/AwJljPv
++/OBKsV7wQcA7GYkdea8I1ssEvDWaUVszjzIhVXd4bnT61BwCKoxwuHRI0bOYc0QY9dVRp8517h
bjDgTUw8qlMOXkZ7sKuKGGZTaB3dShK+1FT/4jMCmnxDMLY5/iGjkVj3MURRbFOLqdtUjxFUen4Z
i98FYi1Av5Kku5Wk39Fhe4relZLCkjJ2FvBeSH8ZcdQPXp8vQb1If5YmKtPCXwYL2RfyHjGvZ/SH
aBJA2qtLeKyXtxVU5xkvyFtJz0DdLQo5IjM4QZyWtTPHQlkdj4qB248oamG+kNdsp3aWvzwobAnl
baohxuKTL61D1dw4QhgmLN0DS6Z+fVGAZGl6lGUQ56l0YhF8u3tUZ7Zrznb6RdtZ3SoqoHb2Oa6P
p7Rp6oxGQx9cyHgMSqk/CwF+ksYeCRAFFJdyl4BSvtTIHt+mFvdn47HVuNNv4UtgOG4H4X6P0uVp
PwHvnDAMQMZUA7RzHKMOD7njSi/aFcnGbTkj48rVa4avFEWd/jfWO0uqGMV8QG8mbMNKXrybsE85
ujwOd4efUwcZ3gyyrD8M1VYo+BEYY+KNp1VmAc14GtjT9tCTUSd3EZzMVdyQddQX32CQ85Yvpei2
NDhABXB8sW+p+cxDtGDFVJp/Cg9fZVkJW9PXhY122f0cinAjuc8lbgozs1NagYoky0oXh2e53bOS
bbi2l49xPieWqoZRL83FfKlmT9yubeQJtjFfR/JkEPRzhgN6/x2TftmrgBjTNNvoTlco1U+cLp5F
N8tuaZE2dOTEsZCad23mx028D9DstUmLohmzKrahLu7ohhzaOJXQRnzPtlMX46IDZrg9zvTYhivA
dDUKq85Ud6XVQq8ngPdLmhlVcWJNfkiq3p2RI75KmJmLmj7nr98f9t10ClSY9Djnccq1QlVZ/S9O
rWKX3dMGXhukegtA73BUt4SufwNrVXnuSGwBeTwAooAGJcXTg4t1rdlus2LEJSE0pV6ZHvjJeVq0
Abq8cZDrfkF8m/OgIyfyROLF4V053DVB0hL6+yiA9dSTW8wM3d9rnwDW4eaGrZpa7bK+hUjrDVRZ
JVXj/PMZpWvzDBy4pfeVKgTsVsWwPRr1DSbVjBmOn+ZjF8iF4WdAI4/JgR9EyHbFRyGLwPHkOflP
xSKykCmnOnQnGztIwh3u8wGBk/fPH+WZQX2MbRJcDOyxI/Bi/SzDmPTayJSgXGtGD7n0zkGat3IE
1VOil1dv0KiCi5XHdH148eMDWXJmrT6HtIcrITfVCIoyyNnDlT0sTY4xfsth9GzbV1VSKZl7TGOV
K2HeqZnts6Rbp9E644zlXK7cAOHKv48NsoUPlGURtK2lF3wBbsGDz7C6aKrq0SzNpCJeuImSiF0K
/iu8jZMWXo+N5qZcNXUpgOTk+29WAtDtoAXk2cs9Y+xAJErJc+CiY7OK/HPf5WaHoINGfi9+FiNH
1T+UDGbalxUUOfD9dRIGAAIklLexK9puKMPzK+RSe0HvSpH8fCLWZItg5UT5aFhFhK69NL/enZjx
sPB52ADyXoKrW7NmFWy/J6Wz91wMtq4LWtqG3E06xoGiTEHx6Q3f77ZiE5nM1yx3fJ28T7zTx5L/
dLSJkMGqagsUyu7YnWH1PMVbXCr4z7f3PjjxsusNq/5jfyrD/ZN8N9zhrbbfZn6oM/IAWKuXS487
O2D5Ak6Vc6cyGq0mHHGLEj2UIqa1fp9TVleRs/2/1C5Y5zr3OPte4I445K5jZyS7vd6fI2Vz5sVa
5lc4WUvjm+yxS5YCUFMOan1eS3jZwDQHV94CXDvMoCdDNFFY3YYuDbnHdnqo8fouqN7ahXQIKCqb
FpRZZwHXfi/4a3Uon1RCPSxNCQEVs+34yw+ynghkGzE5ggQSMJjNMwuVVm5eeiAtPTs8yK7MapBL
zi2seLlt/XgEPP0xwVMX8SII15bwnV/LIkylNLeHaTBh9/7gzY5Ic4/aAUqQ/g1IbDpap8+nLBqE
4Wis6lKtATsE6Ks0qqKFuyV7zgON6NZ3gpiMgcgcBCo9BMHVpS+hqRE+XbURZgf7uv/F0XxnhAF3
kkoYXkpcOE2XiFzBw3AVtMY84kvohWQNADFTORR9Jthv9pkkgcW0FakuQpqjwU3yJcYdGXTsYWq7
tTES6ivsZCOZFeChFpkcA3Lfjc3gOgZqUBBFJYQWchhVkODLN4AbnEaKXzW9KgEE893cZ345l5gn
pMPLhLB40BbSNvaUDCdUMikElCpGL8+pq+/RhzHFHhan7azElMwtW9jm7Y5WTHA+naUafCRWqpCV
OzVcZV7RbdfDbBe94UdMJd5EpMQZicQNK798KpsAI+5qYRQQ9ZmMv1aNQbnkUHU8G2JPV5wNfBDP
KHvjU8+W7UF+qjso6B9YYbT+1xsBflprv07SuD6S519OLV22HArQW/e4oBKGUZZIYNGp9fRdeeA9
vB7yXdqnou8DAv54oqRfOgJ6tIq6IpM6ZTwoHdg/YNqDdwao+FXBagwwjPzKSBgGwUue5LynulLh
uccE1OmWAGyrGfAVi6HLuP6a8eCEcAmdZz2NQqCqaC7ndZgb/6IbioPWYdBjhC3EMR74Pdx1fyfn
QrdUu+A3gfnhpsaOCrP1jRs9cppHUFPIvh/xaQlVuH3EMm+6WhZLR8u87p48pIXCYTFVtAJjArRB
+r8JzKrRhrtFxTGvCAaDpjwxtamGAncsZSQ4eCXKm+IGS86QcKXOjPbDjOTC4oJxBP2zZ5Ngiv93
+75Lydfhk0eLXb4SlOfdT9v25ATIkZD4IByAklSOx69xVTdHIwsM7Qw3hgGa6ieLD07CJQUZcjy5
9ZmSmzCD+l5TueOOVxJHWOEEB9uivhF9haByZHBaS7pGOy+YuWZC0XvPJHTGmqVQjWUAFVqWImKp
wjRCC8nZuaZKJinpUM4c/p+AWyqv56TxuVLM5BIatK8Fgbr66XrNjZC1cvseEx36TuqrmKXQGroU
kM2AgF7iKN9nTVSL8eGh1UhuFzazb6uUaYtahEHb7s/xN4qdjo7PocoPRkCDUbPABOQvKe5glLIn
+WVUVzhv4wsUaRNQxrwGazyWvbRqj2ViNnuKzn+VlhKGBEaMFhGSyCPdOrdoJ1zbFPeWvjYKb7Nc
ujKvEkK3+YNK++ohO9XwX0TPkxAF/xqUafRwlKdXTQiSV0lXMPy0YagnQq7yZpJpoYxlUCKY8rAu
VuwDjaNgeU5fNutL2HBa0u4v1f+yn1o4eBov7dKplgqjt3gyGrZGM3+at4SfOB55QAicjXnzuvAS
OonRDnIb78da8Xi10k8Dv3e/JIUF05EHXNm006QCc7X+jmXp/pgsNndKA80eQu2FFoqmMKKuhcGL
hm1+znp0cwNWGld6at/emfzjRSDlNLuGJUQTGM6413YcMiVyjd/dWlvcap943jBH+ckyN60sZ7zY
5GbCFpSrbv5RB+2UryGiRodABjRyEr3tRovzomjTfnbo7rBsEcQoUcPTjyb4p+JdaOlyla6pntRR
hmtnWMwCRn9bV6/m2mUtXCGqfpU38Dj8UZODTZ5YNdTkpKTxAUkVE/Rj7GQZ3LkkheTyCrFagROl
ciAKeEcSTwtWVHe239YgOM7T1c7PBfsIMRCSlgY2z/kfSlMvl7EFb1ovxHj0dFf1BEw0u/wbcCzo
4blY45vzVJIQj1i5xqV24m0a8ov31RMvbJeVMvqvgnIgCZjQTYzSw9V0GazF78eFNletJEWd2+fQ
sLQRemJW9KGV4+ot9sJTkKCHksxIhpf2MEAIfHFgdgSPtF5baVA6RGPbiJT8n+exAWoChiEwA/GE
PnLj6jMjuMQ0l6vZxHLHn2BxQBdIBF7UpCyKxLob1FxGk6XQlouhESFjTR3NE9XJ6qJAYsg25hk5
DBZFOhRLitmWs91eihFlOPyDr9eyLusgHtm5gIrxzshgmPw7/eCfcQ2Ats5XzQnTAgTMjA1fXo+W
A/apG2nMvSFLFkjnYEZnScz6eNGsU9nTgpn2fp8axv57gWpwH1FXyHhJIZbDpZCn6CSm+4WpZ2hk
qW0Co9MQ63pfXeg1QaRtCOaq7pnhZCJkCysgnYbUoSUnsn2G32LB0lMJcw7FKiy2iDxnOXD9Jksq
6aKZ25EU1n3d5Fb/NjpIMeQUQyzWFGkSIB+ACjVV5nCQT7nEXwlg7dgdk5kDy1n2V5g654/IUxB2
tw3DGInPbfKqxaMndwnG0boxPcs+rVlqwydVdlA7KwTRPOQjBKw3ATs0SLR3I7Id/v4QaJe4HWUr
kdNHX/A/gIQptMnKqGyoDww/n45s475jf57k6xy+03Q97ukkl915lFZ9YIoPvM2rYnsHyEl1I4HQ
Z0oY2bjjukERT4cLrnyRKgRCWYD3yjk+jc2CQ9BfPt40YfSQDasiUMOFR9daguxxqu/oSHZ05svk
2RZTKqkyXxQVG8AxXAOaMw2ejKOHOo8Es/RizHZ1+QkydSx9S4RmKmHMacA+9F/JugpkZs4N4WhV
wn/ILl2ML0Y0vsok+AwAXX3Z/s+ZXp6oMlSuCh4arxBfF7EyTtAipRl1h9putJFhaNe6sL3+qAoI
mrqjs0tiU4BwGsB+Z3o4q31//3bQT2tPVWfSZ+cbrKKCS8UDsSEskCC0MWGhTUgm/K97VTABFmlm
XzgH9oMuEqaTYpoSXMt4Z6vLQp8r6sIQg7QNhQzkuvuU744xE3qLYYNqtCIe492NDDErHLHzdW50
DQl8YGqqre3SLJMVEZhpKCCCJZOAinye58i1RSroO9n2FeaT7Wt2sMjbf+8e+i60WyEzfYaj4Umj
xnTA3H+Ro91XXJi/euRcnVDLBmbJo4a0wJ5R7UQGox6K2CwkTfr8I1KC+a2j+iv/KdGgK4tMaV0g
DLlBr+eGl6lIQ3P8tjf2uNtjhAh7IEtIU703/V9om4NFMt/ZMQpCB45b1N9JbIUou+rirxfNnVKx
yFAkB/JQA578+8d6s0KlT9gdGf8BiWxvIDGQ0cIRISye0XbXIKlAcF6Ep0pxM/pmlysEcwARqrs/
khYHOG+QRFa8wOnWTUOxRSmcpiSHJgT4nHQIfnN4bDQPvO10im7vWBuTcFxsAMDaAMPTBbMCk0HV
+yZm5W1SBbGVBcKosbT4HCSusKX1QrB7TxJhkHqA2oCpNGyF58Ejhuac29MuteZQybWwDzbg/6o8
fsB2zSdjxfh3QPpu9atcXfLoeYHge5iiR6W7S8TbLfwiGYv+BTVe39iKOP78+72rtNipvFy+cfug
Kz8ju/4GS4nVS4jkC1sMvoJuffMCpigjVvb+jCy1oXuQPwJYH92ZRYcC8QtFZVc674ruQbFox3QT
cF6WSq5oXCVXP/0GWgAPbibN9apRnxnKPbejrzvgMZti1ZVlJrKN1yZdpOQ9Ck4WoDroOcqWm0wH
A9BYxPMieJGeQvANm1/a+foNYEVbapynxu86VK/HizNnQG1lfREXXeWL8g1vZ42FLwAm0l6finGY
yEYfGsORaMMOdShJK9s9n04ssJXK79qP2wWkV7Er34lk5wY1HalM4Wc1jq/787+3peFFoP4lc/Cq
e2Zew+XbooAIfQoA9adW8egKsA+M6vY0+5flU67Nlmd1ZvLU7Qk5/zEMrnVw/o+t0u4ftohDs+zg
aNC2WeFO5W3L5Jq+0y6l/lmEpVURu6RXNpmp5IgN0nYRTDa+SaOqm450yjqttedCncR95Amk6Di9
JxS49BiiuJAY2jehFjGRm/8hDrv5G3/NYSIUWQLhrd+YeqRtzN7OYulSfDrXJo3X77qFoxrdoBAy
n6K7Ce3O4DXaCrPbMHr18U599qXgVFgxiZZD6JKgrRiJPugvNNtf+IhPlDKUbXtzXL0s1TSpnxfz
e3Xyp5Lcrft6KWa5GYqe+YMw+3tMROxQUWZEe1SHjtUUKyc79rEjV4J9GpbRqUBGPsZ2s0dF0MaC
3ImVkyK5mijQOCRNJTIEUrnz68+XC5WYu+1JC+xaIsQmS/kMdc9N7U/GstYMopUnLHyQgS17vvrv
8qBgMaUTf3ms9afX4BGKa4Nl6iS7MVb7VfNClY9AXAd2oLPev6fI7re2kSQi0ZHTc/IGAokenCrS
9DIDrklxpxlafpg7PdQPplOiBasNN/EvMc7IIpu7f9TQC8XDJIwwvMj323DmF7NhT8WMOb8Garih
DkVpfE281ui3d6Y+3gEqktJlrnrMbvL7mF5/5+Y4CoNqy7/VpyDe4sd+hX5npipF2/+w6JBDVMhj
n2Sf9vJ0Zo9GuT2RcT1G04GGrwzfitlpX2DTs0vJvmR7VNjy4pfFFyj59DglsoV8NjY7LRC+57V2
PVI57oO16Lm51fKyXqcgvPbj6l5iIR6IH1li57kuiCXSHK+n9c2dSn5tmk2DBo5bboEWsuHcXJDe
AJookfERyusjdAGSycGHueOfP0b62WoU+pkWpFM/VdPfmB/Kxli8SUy0V7LnA/SK7/q31ytLf2I8
Un1J3BshX1FgRY6HdHpIEKWGirhv5952rY6ejZg/0abocxbFH1Zg2ywW56p7EuZ+z4I5PNvA6Afo
oG5JZhE26S6aQPfiSEPk3OFIcUD5rKdOTyNukDVTm/LWfu8jXvI45/bvILN5bJXp1wrBXg0CWQRt
l3M/asffuEE1703voKfCE7m4PfqdIQvqBPfaurXcndYCIlzqXrgaECOo3eJLOqmOj2s1LvZCx/8E
2Nw1Fq3C7CYxwwme2SyvAlDKbxu6YtO2Ht6GCThacFf4VNkQnkqnbuojgsf0GS15hNBWOl3aQ62q
Dj1QzLcfCqFq/y1kYXm+dauAICipGLOpACbfy8N6ts6Mnkk7GseO7ova0yqRJ3V8aIHgBNzk9VZd
qyTINKO2uFhfL05kDVPAD1awQDfxge7x0zlGHDqXrDos0BqW6T9Ei1oQjHszPjn7FVy/WH6BwkBb
FAfcG5q0iEHsLE8oiQ4JShCoNrRF6AK7mocQeHdXSbdn9cknpwziIMBgq6cYBmK6iDzLlYnoyOHF
OwpHOmSFor0IzQpGnkslcssX9rcrAGtKIQzTJYy+Mvl6kIzyxgfHUvoiOiDLK7B3e7L0GkTWcNeN
WCv7xJteKuxQsPX7P8R9zacaN35encSOeVUgEODpI02KxZzMEiLWs6Nt7kJvtzLVRbRQUYHk1eq9
zTBY8DlwAvDkhFeWam4IMVlVWLpOPvWXBzspIMdmdHLPPVUo2FA0zaGpaSwZ15ZQBDukusTA+lqR
6v9TwFtlj4idJqyRt+H7F62bTlqzAbldAz+c8NSJ5okmKZVBiNLeacz1LBTxqiUT7si/1ePqu5E6
K+bYMtwjNpSVK1va/+grt4Net7UWn/qhstYW4T3LPZNxMSZD0Dc+8axXa7qkCelNlnZFhFqZy1u4
dxhcAWDQy7Wo6SyBCATmZn/Ncj3cfEmuLbDGVg6oNHRs5lw1vY310Bwv3FbOXPsqsoWII3Gv6E1t
ByNewB2eq8LrgABoavA3CSUoydJQHc9kgl4Lxj2zuQ9OpRvzaE3Xu8Kyo93cAqe0XyqGW+esbal5
8vvmto5wd7cdsde/7ousmn07IhqWlZZEM8/s1SrsAzf0VRVqUH0KI8TKLh+3U4BJARy6pPgiQLlo
IwcKVYUDI5ptbuQVcMyZjPW0d2sEUYC26TDzqxsownMXzwcc57+8d6YyfoX2CRPwfZj9rA/YsDlo
U9x7qtA0Q60gKeHF2/TOTdwyP+4rL4JmW25eD4lxoafrtEWEqZf3vhxu8VrCtE61nuzBO49AN+aG
4XF9uKRJsGVxSxlo7qNjM0uve5S9xw2Hn08YTij4GZQxbXkh6dhaQKWniSeVeGHMD5WyfvJryan0
IWkZ7HEP8auiGcta4S6tYMMAYQCGn2FyRs4z/OFzxKGWwK10gpyad3ck4mdRoAZX1XnmxaRBpyC+
N/BvQyjswyPGB4Pu/LzHQNHctxoRtnDFLNxgKnJCyuYofeJoJjBCo1ENLaKETBXhEXA+VJ6qokUy
WWxn3tOzOxPXUHHCCgfNl9WmjTDxEq3YmI3R0whGT59m5LGcNHt7kJxm68uWU3XA9wY07+dQT/wl
4IZSd9h9CyxjUG5whW995WG73JOnTVRPeGSPoxPLA2UN0blPX+wOY4UlSIjJYZHNKg0AZ6t+05zk
yIoWSUmgCFSz6s7zub55r2FmzWgxO9YWB2k/zViD7sD3co4ePTkGI454tu0xV4SMTf0i31BVqGti
i3qV+BwZByp52+ziJizxkBE7XKZ13IGqo8P7hxJQOkN88n9hcWX5NCn1MgTV/YYFt/u1Pt/qiekI
IwUNJsR1j5OrmuWiwzxMaez3hMzgUb+USExMc2OGKt/WDRf/JMnnWkRtvIzr+aUSeaSUCHa+LH0X
RaGjSPbEoOY8TUSfPa8KRXphxZYspieQZgagi/XRNm6vuGIHsE7SGcLlrNFdIxhP+vAW1JaFs14o
/CZ5FSq/bC6HhZ5ad2mu/IeSDDwYC37R+W/P83gxJqUOHc21KQ1C7zlzjnOeK794Jg5ewgglaHHZ
pnVxfBsvuhre49wl4mbJ7iVxO4pUTAlfL6oys8XklxHwL1YaEHMTsqpTaqO6k24pn90oXEeUExQ5
oSl6r+g9dqyXe+9KgKrVyIF7lmuvj/Q7bTzPlap0HHSInXU0Zd2V1P8Eh+fEnqlYbHiFaFVB/T8I
olhoigq2SHlDBnObSEptfwAX8Kq2QQqSqZYT/XDK5UEfg1HipREEVIE1sX7rDT4BnNXLK63wc7h9
jRV44Bqq798bNjLFG75M2d/cv8/5KcXUF7Wgt+v1VHyqi9PWpnvJ0rPn+xU/WoeJddm+vW5K+gOJ
WhbCJs/rDsbw3H853vDhsZ+MqCZ7bfRRQdV8iLREHKySezFjRg5GI4fVKBDsC5pvq5jUjc8OJvHN
Wi+xM63MO6LyzIb+78KcEGFNYUtP5S7vNpSVw1GmyaybKGI1DaasWbUDp+1M9ccVYrtq19YGVjgQ
gvYhPh6lTkorGpgaR5YE4/ZIALOgEklmLc/IswIQKTHfR3rwz3HA9JjzMDRNKnE8Vws2+SfeIuP8
tps4Wlk7gmQ8TxWSqoMXFdDZMPWozKZLnHZm9r8ZkfMZMdpDJacyYECElkO9MMOtG79LlMkZB//i
kahrg/WKcUUjfHprtL21iR98+pz7ZPDMj1NZTG1AMLIqzv+tG7q5gauhee/qakpyH2J8lwkpCxVx
fYKX8ycAyOIb6Fhm/I8EruKLyF/nt94gMIlPPQ6dQ6v2Q58XU4X6GA06beQtr25oBfkhjt0MJmTk
bsWi6m6eOKxJRWAAnFoTO86M+akmtdBVSU9G6L5lf6VMIo4JoyIm8k9aAZh8zxuu3YYDuz6Ct4ZL
dCac39qxg1ZDpgn63wI3FTs9FhopRNCCE+kAqTHiI6mmVHZadInl2lwjvf+KMezLrawKZyrTatVz
sa62C7ewDiQkUbM5Zn2c80tXxnvRlgXVCuNjiz/NrVDYW1HNd9JoQAe2Ah+B9q54l/MKuZJweHkQ
UHlb+qvyiMNhiXjlyVpfEFLacR/tTlWrsKmZSE+M11lR62bo05AdQY6in+fTbPkfkM8QUhBcFBpT
8c/KnB0iboYT5FMaR1lL4WP132RjDIgJ26UCXVE4m2gKawRYwnoDRfQ+yZZYrWWn9rTZ5AWCIe72
8rAhJPKEPj3oPSu8xDW6VgnvbYW1UTfBOgTQltmI4CmiFADDAP+Q21PEKSKfkSx0qUTUkdb3iNTh
agBd9yI2KeYmyKQOzjr6nRAIwV9HSbG57F/uiXTgpi1Q7haninkc3C8tLia/voEQCtLrtNc5u4Dz
UsmxPHXFrVEMSGofESB0fO2BVgCBPpvlRmDERvJs0esLOmex6N3L1mxje0rhDxiLI17p5SYFpJmO
a1673hgj0gUQBTnURT7pCnVIapHr8Zb+tKSV0bs0SMnUE+92qRZr6sdJe+l6yAALbL3q8ao3+3J+
Jv9dzp5dRXkLys0WwfHluA0ei4aXqUMKWgPzJ6vhe2IgHUxUxm6skyjBpiHRmeXVUYHFpYwf1Kth
k07po9YCuS0alLNR7qLfvT25DtXSZk55CI/PrQqAEeIyVY3JLvliINl1/eYG2Kz2UMNr+gT/D44n
ezlMnzyOZldggJb6dmPMb+fhtVzzSTTHXA7mx8Clx2wbBJV2bgMY6Evcg5E23CmqE6QM+kWIYrVw
T8FlGftakSOfy8JfxwMxn6u5Gt2vwDTXyZT/LLCAV73F5/q2J1Sbnogl03gzWrgaUIcVxi/tnuWw
Mz6g4VBcjZE05eqlwkyuU8BH71G0BdBjBFysNA+g4d1SeNL8ks/a8yq52IZnJXKOSKNHFkw1fSt6
owuTBicaw9hrA5cQzlBhq53IrkjQSurgHYO1T89qRbFjiTdKLlP3HbyYcpOsAiqUNVbD0gTdWSoi
HRHDUx3ocYiOVrHozrDgcEFzM7dBHUbceShKha2NL0B/60r+zqg5xjaA2NvPBV2nutk0XzTwNGCy
RdzgOQ2U3On9pyrXbDaF6jiuufACXwJ1DL57Q0cGvaZjerclOZxgbNqAP7WcVeos1NH19GesoW0O
gPt7DtJj1KjFxg2DoM8s3jSDXsNFlDOm/J74wYJqI3+NpABzk86J3AfMmMtKiHkuziniLNQLNjc6
VYBsg699HCefaPWfbYTVeH2fPpix9cMh9Rj1JZt8no9lDS7clM9J2zpTdxMQH4X5qc/kBNc+jAHa
2cyhtXN8TYn+53L13m1KLQnNQP5yBnEqY2tYOm0kcLW22yAOecGZxzUFysPgItbLSd8sybihhGEk
eLaEUmVcpgOccG4HxBruZQtyzF2E9p1UY7wNkcyz6aIbgL5fB/zdyrOT4JZXHzct27weEh02gVVk
JSDXbyw34N22EgqglGGUmFTR2ZLv58rtYqVAIlOtcsZ5jSvi5vIW1/7HoZVu7SGATyya0+9q7GLr
xQIY5g2NB2isjQtEqj4Iom1WTeYo+QFkdFAKPSKwCVexSd189NZHrKEpSwzaCnSUGiTjfdNk/H98
dCvtRuSK6Hkm0TbZgcZl8o0nOmo1CtuXNn2Z82CNfshSX9Ri2gLJdYbmTuOqN5eDAMp728DXnFz1
YLUYJMBCnHwo9I5IN+kWvEOiZEKPClrg412wppYiJrhueze1l9K6o/A82G/Vrx+vwDjHbRnz7zP6
QgIKt8Vz6dV17jcUwDA16EBbY/f0O+GDy1FcxlCKAUCDMs66YXwIllTbeHlP7wK6uGIh3W09oKww
zXem/S8ECIxTy+eivcBJM5imcedsjLveCf9hTPZTwCBAmB1k6XhXNmyuky91H2fU8IIuRoy+OgEq
UYomPMsynluG/HEuRpSqLIJW5M7VBwPwNLIBoE7J0zufo6ZQLRzLhBc0qWxPhU5cKW90I9xme5HW
7Ct/swFU1Gm4f40XkPIpIyLsIhT55FK0CwrkZaJhxsViYF0TOd2OWtWgC4YQURM2tlKvqKl/bQjL
KBxap2ZzWPWIgAEQivN1VozEiMzv2pp1dhReJwXwoEN6QNWf75RUWJy0E8hAaKtC4iFaQ8jzUmmZ
c6s5w/vgdK2i/8QDZ0H4FfEouaxWOKCkWixpNe7cczMNvZDBj8VCvpyMkw5rcaknYWANRHcHabc3
aEmxGT5WZDp9z+sNISfjaRVxG/AgeHuDzQs8ccy1VNJPuG6a/9n65h4E0/E5ClKzm46ryf56MHlJ
o8Jv2HlsnL4DZu7uhiHL5TzhNXkBO8U1Zoh3bdp3HogVNQ2tUhrDYhHIWOaKb3fPzqPZe/ObWudJ
/JxnmKatIPxEdp+db9peuQfG30P/y/oEhTWflgVuIoKc1g5DPNVbBbma7Nw06cOmme7AuANWkrPR
Q9Ztvce40GDDwtkmzXhJf0DXlssgDZrbs1N7KRW7brZhAQzuYzhGSEETcOpLtX2cgErhV239d3t7
pZx+WODKqNLwu799ZKdTC0P2CkmPfCVGzIGxu7o0oYxqWYbEsD9fu+scsKF7EI8YrrsPCT7L/gTW
Uf4K3FsNJ9FVf3CRUPvmhnggs3TEezdk7rr7vzMQ9JUQDFYDxWmFZxLtjVEy61EKkvdC3pOFYbGN
LTuh27EwE1zj7c1WycwZFpeNlniaO76thCzlyxnV3OFvwJMyWKdPjbZymE/RDoE8nlZqyUcYelsr
VW39B/oNbPhEkOf4R3xkmizXSK2bcN4BtLqA/kSaVXWX8eqYPOmMvIhKoSS86Gi4bK/3/WY3g6E8
VH0VNZdZD5wRArUT8wtgf+jLrCB5XK4cb2xmzzK30U0vDs6aItoGIPG2MIf/Ct2wPI0E1yItmD7Q
3z/jTNuvsha0N17m5QMvqDlf9X0qiDpoGAJhGDKy12mzUx6thUthWnoyxFg8MFAZ0A9+DcFx6+W3
HwKly6eAou0hVu+H65IakbwZvpHYX05dZjUKAb+EcOidWacbkbkRhlPKYquX4MEFgACU+k1FKrdg
h9u3EfHpzM4Bi1mJJDyGLmXyqwyHIABne0f3Givd0dG6SGpsqg5bI4sSFdnT5z+Uh6dYU7LFXxxm
4whLMPUmAZFqnFo/YCHEuMn/GD7hTR1PH7jZNa79h6OP9ia8T5H0HZw6ULKEVL7TFnb0lNKAVaP3
VZ6AWKwHZ7uVi2LMllPSQthWFvQ1/sMnuZv58bQ7H9sspYAoQWSP/lxrVQTXGXmOEQEPHyhkJzMf
BOxAr9BGv1yzbPHqGD09PKfLuG5ASWTXkgKVfl88ylH5D6yOEKFuphRlNSiznyypKp80/eylz6+U
xcbjk1YYEzJ8ZOupZhmGvTaQKhDcAADl/UCN04LG6pdDd5lndFs4zIv/7xxqa3ZQ41BqgJTpEQ5W
V+nu97NhH16A4rx/ij4e8LUhVfy+PKoILOrTePJd4ATII+hFRY0rYwBxnmO66uIB6BZbUCyPeTV5
mGo5cC5L2lUgAuvx38XeAAjpkE1Sso1GRrqbqKawpQLMVNC1fSq5VF+G9rtspNHjn4nJXWvBMiCe
0FfuZcJqQkdA34VA2KEKUnZYpDHxfYNqtFXRvjJKntHAxQ5qIS6fltuIUjxsMGnXhJp5vGOENPJW
t2z+v8hCe/JHiuKxDtyTXLTNRhqz2xNj8IZJ0nFDx3j5ZNwKH3RwCgETsICs6u6nj8DkYDvEJ1sH
7synNbnedl+qYh917CPtK+WHOICK0uktrXq+ACTX61ldvAa0uDvsnLZ1h2HU9Evzb4pOcKA4woKL
aCsb12mV/fKx7ZSdK7tDDsJwjNdjPl4UERJ/lBcgCFfHsbnZ6/paXDWzvVDoebHSa55xyv4Npwg+
jgy5gfE4VJrddUwAwnhJeg1JBEvS8vN84ryoacqoTuql5XfQfSuNX7KqJQ0Q/iKXZ12H0MRQe3V8
/s28ytNVflWKtc2ct7yf29uBkm4EO5RrCXDnqrvCmbb5CO0BOKnyN+A7MQcsNmu5IR2+Q1vh9rnB
7IQ7kn4WDuupani94FuDPlUz0NSoHJbpcC1bWqqnTft7yoDErbkxdxMr4WcW+YBeIF0jwetl+diS
BJ6eFqdfwrkE8ekM6hTmoUOEBI/ER1VRzOUdcranFEqZlwcKsxnTd+NSka8HV3YnNmAj1tUByEDV
cpP3Q3tZgknsdWpdH78jQlfE00vE7SPDH0PeG4a4yLz9kawN10/6vo2ZyMRqCwn/ddEz8zGc8Rf4
WH2yDWLckpQe4p1EFzkDUEAVMYxDkG63/0kN8fxWnbCfL17bJP1qQtfRkl2SOejfL5Y5sVuTxrOM
MFIExIQQoJz7DCKvG8g258iVJRt+K2MBxsIlp0se6INE6/82NBu1qoSQ+lJw0MpdwKyK6kxvlizm
GkYJ67avKne/AHsTPFmYyT6E8C73PKLyxv/oF7t+zn2CmY9AoV9YjcPZidrBt4E8M3Mbyf7VPw8/
TbjZ0MIY3EyK0xfpNlb8FZASm6EwvGXQrnmTWaKCnMhGkaxGAXeViWa+e11ieymA8EjE4GEAa1gJ
QOdFmO3Y6q4IxM60UY4cd4ZsR42ddcaZuxnjt6fJHhgF/FOyefu/t1H/aRAIEXUg/PPM9SiSTe8Q
1mSUOau/9sy8hWSir1KYGhQJ2cs9zubnqI1BbpAKux/s0QwsVHHKr6tqDLPi/NNBBXxxMGhSwVAa
HCNgaw7RbhEK+srNLjWaQt+bRcNz/yPvHe4g/PYe+/rWHxc75qE828CQ5evf5e8ZZYQ/O6oT4MN/
MoQGLFM02s1OAewlsIFgiBMCOHtKcrcmBsJioBy9jYipkmPtKiIu2WMuR/JMEtjh+IRnQg2adv4K
JnwuZyEPLbO0tPivNIZSWiIE2hbDug7DShiMaPOntm6a+yIQZXNv2ir6TV/DLSFvfDRTi8rdynkD
5Gyr8anyXsxBUx/X+WgY8r8gf3g8xOBJcO7PwValqPsvznh3G426w3Eho33gH/Hs2HVeslWCcNOg
iWukdy/1A3xcG0ecu5IBtkpbWTiCOuPFboG+WJmPRuSREqWTJPuE5qtPcfcj1ySNvnX4JEPbdSN/
oIw172DTghvEGwACAwIJohEKcMFjOhdt3YkcE0z7YmUmwKZOhfnJZP6RvrGt5mtRPZervAI8E2qz
25adNByn3TPCABtA+j6BCTrzqyjU1LdCqw6VUxgUwfGjTZUe3j2WPuYhJ2MgYOPuSzipaj6RnMze
hNr4KhGsGAf1+zjSZQ+fmyOZW9JpYI5l6oRKPNLronwm0vEp1f//0YUJFiCYMbw8XwSxOB22iyD0
79zAbaC/efFaPkfWh290sRLj5VLeTxUSRN6r+uoWh6ywywWzyGeGUPGfcL8QN6feSDhHAA57uCNf
AmHRERVpC4fjzfu/KcPnILDWN3h4e8bCAs6+qpcHz5kqr4HCd+DcwPOe+kWx1+VGCRBB0Cw+cizE
J7tt1RIjcYOb/PdYOYf0vEdfGIsbirtgiD93ABhtMX/vzzFcGzmoZT6z1dFWlrrDPx+uRRwe+uSu
5sOAn1Qb88E8gJMuYOEiE1s6ES3i8oaRnNfE29q7U4+Gv7A6f3BHYZD4T6/tXjW7Xr6z6ldTkwqm
U0I2ulI2BLd8yaaAGVBXiiRmgzE5cgTYPUCOJpI/dL7o/4OsDrDHvAQYde0kii6T3XmcoUx4ukyk
oiiz8Lx8C8gKM7/TiGJ8gzTuuJbxY9xaEk2dnr7p7DgAQC7Ydp8MkHnmK+4Vv+lqwTIuVaA+NlSr
sAOqhH8O3CTVgAOIfv7G6LEGZVJ/q5CdPiAR4Dh7LHZo2dfBrtWW2Eeh3dtJw5zA67ndoTkrx2gO
g27e2sriQ5ovJT5FFI7G00dCSL2FGpe9rDwHZjrZIzKbLO/uXFuPhlbskNhwVyVO7mnGvoomp+MF
x4cZ4+Lx0MGBncTgGyTHouWA3Ooug2nDuEVaJr7qqZBSmN5RwuwKqFjd4S930HuXME7gAwoDJbJ0
bTNm7cbQEuAx8kk0g692e5yXV5TFGOpVi4kb1WwPFTALl2Jp+p0LyO0vpbe4pRGAcIH3tanQssEF
METa1u9sa6DSjqNcdPr86QpZzLWddCsNXK0hesBRHNZJHL1dQBYu6E7iKUl+yELWmvPx7i5toRhA
RXx4DnVMT1NiIjeLeZe6NoEXyS0K1n6VOFDetVa4BgtFRo0KeX5dYAxsxVy3pcT3V2/ph0KZtU1E
by9xQ+L0d/mlJnQhbOwjX0+7f5RwteSWEhysoGJz4e2MYPp8FUvOZnENZvMwsU+ssHNvNCbIe278
Xj7L77lQIffMsSBTO/0fhCXlQb1fSXuMReP3OxFcRexloFGMSKX4T/kXgtdJTHEAlheZRSBtLeh9
h2z4UujhDcDb9PS8pyJFfC2I/9miZsxD7FIJCio0oJOQKGFHUnOgd0slQHplQRkvO7iU6s14nrK4
4N0RJPGDIRqVUGE7TFV9dV/HZGpoc4FcCD5GYmSXttbPPQMkGMEtADeTpSgtvUaU5XlXTeBr6mVZ
MtBn/jTw7RAdmoKV4XPqWu8btW3Tm7LBxbHgeBGKoYjrZ2AuhWCgKFxVBjSkq6/6qode12zdVnrU
2VXToDLwGLTzC/MQNUsZ7HzYRuVb3s7dNGIzdcZuB+ueexrRjE4RK6VTrW2tbObTIN+vE9u5KWBk
xGVBGgaIAx++g5mdavRVF3vs/cWNNjQI7KUhUvHORPRDUDmbjnXDJnnd7uwJi1KLS4eweOHYS6BF
XKqKFmx+WGxvnM598t/RSsRiI2oKRrxkJGr5Z1xRZoypsVVF24HGurftcNIofm5k2jXHUa0+300Z
Kx9+7pg3TA6QfDSjqgLLbsSz4Pejq6keXtqLWfOZNGwddIzz1MKzWIOxnQSSEg5q2sJ/y40VCtc7
kFtWFgPz//O+FXgjJhZlhiG+rIk3BNAfpWYyEYImQ0XC2ODvr4qbU+im8PmERKbwmvYAZ/mq4DyY
tlB7zmvBKhkKsn36xfsVyDTqqoBqusTEDjz5jp8O/rfE9TzNkDJYbSvcqsn96Ox+xAdO55ni/RXL
1P0SsbFMrLaw9KZukyWIx79Bip2bDe7gFciLejoF4dnRtv0Z/JJ/XV+XKvU19/OoxAZgcldYFvu7
KjyQjGOcYyiz26HGH6OHgcKqNnQLdGe0oi8dx/FT0j733MbxggwzZJbAS16gEfolwW04pKm7G4Lo
g49d9TaaaLtrrYrtpfLHGP+TsvZ/O0yO/upJtVEoz4sJlsUb8rHdR8pu8YBgCB1Li0KWKAQMO9CQ
LhYPADq6eQthUnoqXSgt2NnkjYx+xzXNED51zKMY5YmFHOBjOcoh7Xvp9ugWh1w3TOKkwEGAGBnb
lc+BCKAgy4fuHY4S+4WATvWCsxO6Jmupy2l3hUS9v4zFyRNl0fZxvzfgCBcxxvSErMAwCzt/ng5o
2dvgl6Uj1FknERCS3CQMbDzScoS1x9CpbHM9XxTO9whtx03r7+pBbO2cpJPeo/t/gl6UB5XPNTSh
3IN478iR05APL4Oi0Gk60d/t+s+FAscjoLchpoqLJXHf/60jCCeHS6VP5sp3l4KonFBFWPgn2ilV
/++oTNrXbWxGgfJsrLCDmRQNUAL2yOVokcYAdTvYnJfH4MGIN1e+Eps+Jt3HZp+/Xe4olgv4CvV6
cUprhCYSK/vRyY013YMlzyFza0/9jtQviZKBSFRSelPPT6UlJRSZhTrcUwsnNU4Kt7MQqTEovAW6
uNCZ9idERdgaH0GR8CCvl7idKyqflKsphV8EfyA+msXMclVbTyds+1SNb7axyqLXsIhTXPlkCCS5
qMkXRCSWuDrakbNc9qI8rpe8pRqVYQ8lUsvGWMfaXONPsshXNk2O4mIp10EY1kfdyc7BiaGu7Daa
ixbfB33tH81yPUHqLCG1RmZ7ELNRK10lmj1IJfwM3oofk64PlXm0ebURavxWndQaySB1IalqYrBn
W3413SiAvqP57xgtKURQL9CEEoHuUGSE8xC67Gy0SESXcIPc0YlZr0If6CkSl9fVZCHFpFbmfEkm
LBVYpslzdKx3lt3nb60MGdz6s8aRopOLe6dPuvT11aab+NG6oYFS3ep6Q6jMUKGG1G4RyMqNs8tX
QRrl3PjPkkfJ77ng+UOcMHWWaMDvkfgbXz1jH/db+kIX0vc7ULft2UUFQPLAKJoV/mcIQ0Xn2Biy
sgsJkrA57alJyu09NSbGEsPYDT2wdTNRB4I59tmVjH7qhAa80ibIFrG4rQDVEIp002JH3VQk0glt
PAD0FbAjWv09FDtpxC3F88yO1HJk70yXvlBAaByEVCo4n0U0m3OvzbvCiviZQZFB+J2Z8K2CtXAX
Qy8MtpLYN0C047y8x07BrDRT+pqqtRFIoVT351TtIn5+FzxAAyqzJRaa28VtUfms8q/tmQ8xVkcr
nOMTSJHpNtuLQOmqAaBJ06zKWbh3EyjxtTh/P8Kipznb+lf4x0QRruw2NOtg2gVj0r/dY8CuAQZF
BjewfEJaiRVBHaYs6s+FA/AgzZdQX8hh8ECZ9qynlVGsspKwUrQMBdPktxIjB+b2niCZWd3fD7W4
7fi+8M4GN/VmU8HSxvNdHKEmOWFkC3+sDh/bn9+V7yeZYn3X47qx1ilb6YcrlNLtLrrzMV9/rZXP
gIduxZ2+x9sm800qB7ZawfBeyDmpaFnhUEJfDF3Yg5b+NLWWZE6QngGReinfg3ap8NXeHbrxEj7K
jOvxdNlhoDJxSvHIdWFn2gwrcYJ5Tkuz4uQVqieLvPVKv8cfg/YxNvB7DAXJ6xZCE+8EqGEbWpKP
t5uWhKLvaUhecF8umF2F5dPRI9Ldtb7sIzPlfB6NyjGSx1uKNcKitaolikbSU/jvWsSRq4ci32RE
J5I2+/0VWSUvRn64vsoOlyNSXzp5nRfjhG3M105Sk3lP7Gj9zuof0j938Mvm43H+sqQLic372kwF
DL/KGpHFow1F4PIHr2RL1Bm7U7Aw+udGI9Fxx2V/EkQR+P9O/qEve8PjiSG8FTz8PKW8PdnQnsoZ
Dp+mCgLWkKFuHmezTyUCRVsNI4AiOxCHhEWhobi+Wnktz2p1hVbCjJEoCNk5uohRw5ygq6rV2HAW
/6cTJbyg19oCSHuoGNHHdSE91FxcC5NHNw9CpfBrKVFXaJh0n/XuyAPoT5+lDBE09kf0Vv5GPV5l
2PjuFq93ze/KgWHde9YJFMgwkgqFdsHkV6lLpdYHKaVvS1+QnZpYcucjFshbgEQL0l6SKx/s6VJ9
Bv327j6DaD6eDDv1RwAyPKZpIz3cxELUcVLvgJyzAEFtFDRXaSKX5XnhRsB6KccWy0wYlvaroZnz
3xeOOmlZwRp7ACZPoOxtTi5qD7fRxsP6Veij/gax/KcYETo8wcVeSDD8cavoAa+8nxZsSRqcoJ6G
qVZHgIPCxE5sZQNEjDn1Yq004HabZ/M81D0c7yJzMzoit4mhcgf/ygHXOKyTrkjYjkIa4uGL2Kx3
bsyxNF5KMFUZpBOyrl/IUEI+llLQM1rf7v6S1s5AofbjV5HbaLvUte+sW9i3wz1tlopvzLOI1BvZ
Vkusguwfm6KC5x12UvLcN1kGdmZm87j4dnlqx6/I/BR5Tnl5F9f529yFWHiGbM+2JzpezpQkRXTt
+6gmNqrf8rcZzkNaI05U1fdL+pnVI4VjFhW5hXfsNnSFqs/X3nlT1UrZSQU3s+LPbY9lgTvKHDNf
zd6g0tIlUgwxkuTnR6yxh0MU3l+5ii8D9PMyTeXWkC1WILa7bWOSJTExh4B0gvt8V74cc3FRl1l8
UqC0X63sGMuAPFHKIy8cUO7b1kU7RKGUgsnIY2KuIDuvZFa2iHK27YvNhNSjFdVOZsWXE+2vOc+7
jKuGL0dCn77vmxKpaiv8Usk0oP1VfCPUeaUKYvj1QS7tgTM6q3EUhLlGEnmsiFGo/sVTjdpnIrca
YPRiDDS4sR424ac8DVmLKYHkm4U+4+NzdTBcSvSCvPpePddE2jhSuP+XdNvFwUHGEfYvJzmyFz/V
2X6CNsAPkG6aqbO48//2hwmMsRDb8Cyq5HKg5oqOVzML1Ampd3CVZJQ72MLdj6S5sg3tw8s8prLa
+wiDjfGE/AscWRtK87JIWJgOgKgp3sWDpXH1ZsITdTdYcR9h/djllFf7+8Es4ZGaHjNrvT7hTfKy
yZ4gdiY4Ns00zz3B441XmY/NkoJ78aAbkTVfZaVFMP2VYOfP+DFSpJtUE2z0uDwuASc8dxL50Or7
/IziqPQzpalswnQPVe9IvcvbNOamKoJ0uo0yzFlWcTgBZBsLunXv5KKMQ9ix8ikT1C18ip0gcYMv
TvnmeJAO50OObHn4t5f3ecjzMJgH6JuEQeJuHLL2TTgBo3nYDRPq9Kn40SZw9mtlxlM6j1NBqvaW
RxOI16QaNyxUGA/lSXj1fyur4DdfSPekDXs0EqCzMJweF30T6demzZzJYDCcqGaxCkGYT+kyg95F
Q3u0GWoC+ZE2wb+8VRCczMJsxtI1MUWmu8PIm8+LqMWioJDWv3D2w73kIAiJWulwheGO7Gf8HWjk
b4wFhKt6Dw3pBO4hFW3vWBQ76JtlkKuDd6h0MwxWtAAZrTH1FZPGIjJqmmU+c83PMwE0fjP7Q1q+
t4wy2YK2l3+822NQqW+5Y9Gz810l8Qpj5PIIVJcPZ//wT58Vr6pUWG35HytyDbznapRDxkdI5Fau
Qtgby8tOonQvxRisNf5U48VC47OMxZ28r4ZuchV4HRRiafYeWfV4dMbzDmWMycKFWGo4qjJDEr/6
iRbXGUcigHLJYKrrRuisIr+1YS1CcaxYuzVjmXh28pvOylVqaqLvOnWTvqUERk3Wlusy4OZhpvuf
pDeWv+nbvjtnciaQJzmLRxT+mJzoIh26kNBG+gLCPh9NksPAi8bilII7qkwI3jZqrDCN7PQ/LWve
CC/EYwjwoLanA1kg7zfYIHWrNorVEFkK7TpDpvOi8rzApbBuonFpJ+xDhzBmvM897AcyUav3eu+h
LayL+zIgQPQ+/6bcYMpW6jOGzmJwhNyl4okojzZ4yRsx5ChuCRh6MtluLAW+HAUSxv72Kq6aFm/I
qvx3QjeHnryT+QtP8g9Nzy6q9WpnHbK5Se9EuEYOfscmzUTd2RPEjHKdHdL83bAn7lzz0c/CBC5L
zl3a8ihk3t713N6jDz9sSqcrbjEB1LI8z6OhMVuPAvGYBjgYUwDABP20fBdj/9C405WRsrBoMwPp
BAWe660hhQ0ADAj+DaP7W8U7vOJ+nflCXRlK5gBYUH/g2cbsjGUflY/5gyD8h39FhQJWgogq8Hs7
Hd198Zu+P6NTkE2Px9/LghCtaIn+OiEdPUTVpVq95RzO3slveDt7OxbqgTYuP7pxD3pgLoaG777T
HwP9zUjJqI1OiWQ/G0c8SGAl8zhnFnYpS5NBNIdWWjvUD6q9mv0xXt5SmIFoCYpA7jjjmzA/pnnI
4mpGdCy+Ca4Yf6Aq4Eh2ViZPqIEHxRmGPUP6EHJmbLNmfRzGTby5q3G+gnQD1AapHzzPSuK2254I
JtZ8SNyIdmXkLMwj3eRhVtUy8qm9nH42HPP8DfZ6baji6qFMhCCOOeBJhvft1IuSfQrwvWa9yPQ8
M9Qi+fXqsFc6vDh58vvZ3QBLiwrVffRotAtIyEcpFleAW/yrPD5xV6sNhKY/wTZXTy87Uia67DGd
TlEJjQNqhF9nCO4nBd3P74OsqUUxzogIf9ItAil0fIzZk2lXyfBa1eZqsHiplZAQ0QXq0QyYFHfF
yCOTKQm2F8yJF1WqOuE18JW9zCJNrVCbGhCFkAJEP07O+NU22LUR8QqINA79HEXXoG5V8DiZKhej
+P1leXC3Aa2fWN76UdqQEp5VcBseIWxa9+mJN1scZeKP5t2YtFy/PZtHjG6zbqStI0Zn0M8TcKuw
WG3Hlh5Wx8qaEYuI3RfIJBquDy0cZoDLqot4rB3uyP+eguVdP6ExREhqfFAKrZSZ4iorrBFa+maj
I/GmQsCEAX/v9kmg+f2eYiSv7Jwfr/X3A1Ma6epTbYJFahBna+PokU9FybqpWDw9NT7r2QkzsBHI
Izrqc8nMfQaee72BJEiaAzi3nNhnRlZEFxFf1uPbdHHdvmUmcjwPuAGrgkvPc7XStkOdTG8Q5QR1
7vfGem+iNfcFr5cxqm/29sG6KX6ib16LeQNANCbZYLP87O64KBzwlglqLcb+Yz/nj0fmLEoH6K4m
x6pPT/IlGcpHRXz20qYOQtFiOwxbY1QwlSnWx6s8SUtX08Q+zPWUWgWs/o+FYQqQr38mTzJ3gT3K
dsMymGSbMq4W1BcBTzwta7fX5cG8tvsYW/2N6fQf+OGgMNuK60emiOhHE4SBZjBSSlu8Q3qyecYV
Hodqq4vX1GOgTVMAIIFt1yVWVgkQ0KPSkmnUQnWZTQI2BuewHdPyf3kvLQy4TC3hAy6J1Ad1BX+1
6SLsFWHsUadMBACj9RDi4tj37RSxdQF40GOd2n9iev+CIDjqgAsC+4TcQapMTVqLxS4udUXuMflW
ZcMK7Hl+FnTgBj298M/jFHxORjoBkeN3Yw075fkIBm+wuTZkfgOYTdM3TWQOadoiUKQA+js065yO
BKMD3jltPYT6n1Iv9uLT8tmjkXzHAP2h+D2yd5z5iOU0LMIHpG6yMH5lVuSMsHBZyT37GoDJM2YR
bfjOguUubsWj7rFSO0WCe3lS34YKqi9/HXtFOcyjZHuilS/waIqN1xGJV4COm0JLA2wlq34/TNUI
lheNvQDUC/5MhfbPWAq4FU+6aTwLFBxa3RH033jgDk1LPmdkKbEsVEH4T7mxmcLfbOcTx1Mfgdbu
1pJVLe/u6irbuN9cczbFvPAcOB0FT0rBL2bhp9M6d0Zvr8wtG5mv4mgjcu6JFvPlIvg+ZhQQcxs9
uWKU/KGiVCqNUV5AzIYFiqLriu8MZSNURgnzdgMxLw2RUYWCVbqgwsdTkf8m5uIwu14VO9wnDnf/
cgcQ1VPfBNpSa8Y0jRt1ynkllDePWERnZv+wc/8O/XidfFeXbMqAyVyesO4iprvNF1aFlru5XyPR
j9Z/0Zes4iPZKuWrTk/uNfDy5RYoohiFtXjSmsGX1cyz8QFQ0MZCZ4hN7PTIqNzajpmKOVfROh7f
3ppxxx0C999ZEQiWzgsWfQBj15OtZuScwb8Dc6A9YUVuxC6uqlW/2d11I41vBuuDvGXuHxRp8ibu
JQjlpk85SGysn7W/tv/512eZqnwr5ZPDn5lhZa08Y7gDdISzHowfa/fwT+JsBqOOxa8vbWkapggX
iFc0HhLGCKN3qZGF21nbuy+1iGt4NYmfMTZCU/xXEjaxTlvXEhA//fJxmWPvl0epX5LSHWGhZ27j
/h5z9dTqVd/oyqE8pj2yS+wREasj/m9nG9nYAMwIDMCqCR5EM+BppMJD/KuWFP9hEIB9R1VJBRa4
c3D7uKhnLEeefzxjhNtRcdhJxbSuF8Wv9WimZ8PiPWFjtqNkuTEhRdNVQ7jMHuLMyLu6JZlrn/19
MvpzJFB/rxIKBX++8dXHaxODIPzk10EqfwPn1T6L6DbQey7PxTlfdIkQJTgqjj3xSta8YOHt3nR7
tEIyTMl9zNFt0qRPyk2pu6mA4UFg/mAc8C/rNBSbVBENnL8pLGERAYdoWHNwzbp488EHZzCaWz33
f+sP1UK+ywj4jJijuMkTR62NICMmscwQcCrYUVqMZbV+aKp72IcxtqQzNJqx9HhKbTbXWXRtOxPM
uTeQlGdStUHwZFZium0PZqGy+4h830PptQhRBEQpQqbmES9tsPZleNeYh9TWWyMrlDKxlkCk3Yx+
JPjgtPAPMQyFKJ8naWvj5DEEd+MKTAO8tTlzCtVoJSb2SIX0V9r+khrC2yLiBMZ95UyKMqNhm1Kf
WKSITvtgojQCRa2T59kq0UhDYpkVWA1xoYogCP6gYN8l/U0tj//lWQj7gsJrjXjXKa3bLLtCfl+Y
OP6aIwtzRCvl51Jv3Nr5nBwCgwjs51ZuvF9iB7CXlngoRbDdulhVWTpqXKTGl/Wx7ACTTPlcraaq
q+KAp+tIG+nNt04KUU+TYNgeTzudjb7m3f3mB9ZNNmomgPiRAHkLlNMj1VmM1wu5cURDxQWXUzAJ
8CNqCcrCcfL/v1+eJmAKfQDt/Hj1Rt9gl1peTssmMi4tEe8qVU5jfXnTu2wLIPuA/NOFBeXZv7HD
bx5vTZ/nUn/oWAim/ne1yTeO/kR7VNCMzpBy6wb32EPJXGWxfkD7jwhVtn6WC4mAPt+126t+yZnL
SKi5OBDCCk9JoX5lW6jLlwsdiSnJMAVQYj5giR+Jvl9xS2E5gWzfwakDrbJPbUtet+a7whbPKJvp
hhFwcWbR3s9qHlUOZH4I/n5Zobi+AeCad9sPvNXLESLYD/wFzsoggKHdEPn/YCDr1JtOrLs5SOSs
LGHMqw1FW45SIcZIoyf4743T/avkV9/SnMGdy1ri++B+R1CmDsskJcV+rXaosEqpg+SAYmki8aMo
7Z/9UYSDGjSpQd3QJe5/NfGCyPPa6yz79eYjmsEkHOoCMCfkfp9FI+8h0sOfuvKr0AKmqJyRrsZY
QCvCOLAJ9E9HwDbGss/8LavqxVitEaImdjVA4aiCFbjKCzXyHIKeZ9No+S6/VcnixkA6GJEfebWp
n2XiYkZePYTygn66JDuja9AOJSu4D03tMk3jbzRDoWYR6vvpqW8BVwomPX/2HK41DKm9xkvq/0RP
PnK504tLdre8hbyWC0hbjaV4UYmA2waqaRSEV157ilG7ftkIuvIq7sEeu8BxZji3ZAbcvw+uhsYw
7j24O0xL4kJx++4bpwrgwhwWqPvQ7NXM0YN7MGHzMLiuyhZ0aW9L5LjCJxpAPy/PI3OvTfai9rgb
bubvRpFO0mg7nXDxBjy54yU/iYE/IVuf6zyU2wnzB5jEeHP/9dBKwIcwTBAvaVS+9ZvCcFYNeQJf
jw572YMOFs4TntL6LFZp9PUxra4fPQyRmG1gy8YAAS1Pqu9+1MG72gYBIDIPBPNqMsRgxfVGRWcN
AO+bkSXEBmU+KUb5wTg7etzQmvj95pQhEtdwdr4dj81Xl+twC5/XzcqZGszQ0Z1zIvUDVI59fgib
uQv4c/mL/ea0RHp8sorPm+u+I9o6DKQ6nw1n9f7LW/7fbcEh7Rh0hYnt/U3Qss0lzUzpySg+VQ55
WVhbIBzX+me9sny6JWBCWe/UMvgEYWJ+zxAdP1kpj8m1rbU3lDDNQlWjESaD0aewKJY0ZwUnfobA
EWnJurQne72ToNrQos23UcKOTlxDzwhkX4ooWgpkY4bulT31FUp2TlijKBSNjkKre/p/MWujnFzY
m7igGbvSW/d96B/Uk/Z5VVLHB33M+mBxJ0LH40fASwNkjWrTgeSMo5lIngsS/Lfv/UOaAmlXfRYs
DymTKXvEWhkDutqoG1bXGspW6h5T+DgQ/mUr3gPI9MFGIhnA4UfQpOfow/BSYMUcd7yc7zMirGRq
pcuLxJcht5bDOtAL8tHFkWk0FZ4CzmFbgIobTLX+WBuTLHyR8MCGWzDhqCAdaicUbcfD9hW6rlfu
PKqPITZkwpcSs7vogIhGRyHKlw9y6rIRx9Dxlli7L22M4vdJO/lbWOfhVSpuAJ6lEFDvXZBGGmQA
lhFnMMJh7+AVIsZTmFrPKHzgG2MbtY33FWxK4zJ6PaowXK7UmP7qEPLAiXmr5hD/0ReADRdSj3pj
PPK4s5GsLT2sXqSJoclrYw9fUOmgQvORFk+SZKlPeNt0JccODMe9/RQvi88CJFX+mYy22NTtVuf7
EvDXasvWhh4qgYudGrCiBrHhD192xvTYnnIkhiGK3u3tyURG5yzt5/0VfJmizMvw8YqiA5JZhGdK
7fGAvOzvzXbeiiOHNln25UvdKkKKadHsNm+cG799Knj/g45PvVqcNVRHdk6kpAUJ0d1yDCknJ/sI
CyhBfM/7CY7kLWhP/JZFdVLUbq0bwItfdsr0sM1cy+IRywCSMfWbDQQ+ZELrBW8jVnr6/q/THDJl
uFhS+p9aWlmiQ0MQ76OsTHcJ2FTFuvVApnrWO6Jy8cV3M9tZorWHhy1uREXQCAsViiW3sq/Caoen
eVfv06POfl9XX+GM3GHhhfMqqHRfdoqpUxqwtaJJXkj1Uqb43lu40L28y3E4rfzcAB57pB6u+lOT
iPgUdBq3+d/QcbN+mOrJUEwzhx8ladaryOsXgF8wGP8an4kfyYAubxEwY54pIU2eNHvyF88Vk7Jh
YV0OcOTr8zqB5K2ySVz1rDKbZMm6MbVcR17aZuaPZWspRj+5hvtBKdlnPZkBHqupQdLjMsHiYkHM
N0LmlcNg19oZs8F1KsakNrueLT1NYs7PNm1Lra581ZlWRsWhcMR71s26VW34NSDZ38shhkmo+5wV
kvvyUfac1OFYbD5bMn4G7w+D2d9iLNlSgt5qB1zFqaZsRsCAEOPxPHcFWbPWZ9G0KFZbc9Xaco1q
vKaDIqjQ6okLqWtMwWl7XFPx+AuZ6EM4fXWHs6CQXR8WYG0uBQSkIVmSxplu7sIl2jsOKnktOyrD
V4aUakU7ebnAkVejluy4LURQqYD+Xgp6EMofxqa/GwKpos3dxQ2N3hJiRrzn8bPtVSyr9iPL8R+8
wdrzZ/C7r5dWR+lY235UZk9dx8wFei7sPc9FbOOMGC6y8oRN5a5uApKvv1bRXmVkxl4nZ9jBw7xT
MnWfrjINgXH0CcVax8RXNQJNsALL78bLr9Of0Sx5vdt6HlG8Umb01J0eVh7czh/VawzsLo86OyZT
khlnAicjIUY7k5DK/lDEj4bhrjJk3RMc2Cp2w0idv4I5Yk0GO1ClaYW4Zm75S9GpzsPrDB7tBDFC
yk2eUsEcpq2nypHAbh0LWK44MbStXIemoXbegUvmOllMGBFMPwD6gXUmygOAxMqOSljLj3jZkLMJ
nYJ7T6usg/tI9sfhP56evGl6PjGYYXCAZA4zhA9ebX/u0P9AviVcx3ucnklaykFXRfLzuNxQ7Tc6
JxlHdoqcC+hNRohy/3ZJURxP9n0Tp9Yv18ohIZmd/V6d1xPNRvQoSebFvd08F06bo7OUFkOEHWeT
EQCVd2kVrBKoT0VPqOERx92HG5MQGmM+2Sp2SzNQ/fzxxdTPtKfDDJwRCDOIfon+TF6nYMQw1TSC
/amOX7e1epfeL543E3dtiPH6mWWV8QAR0s8koX+jld4DB6W/k6HmZIX4/iqdN3cIVTRt/jagyN4N
JyFh39ZOPtE89rmW3gUYIK/wwvbgM7KdLdhODxQWsdrkRcYO6VRp+nNBLH1bE081SY8iCErc/rBd
//iq8nkqdX29LpAjHQ8gEw3z6zQQ3eTNGPnbGwTUt98ZJInaSpUS/t8j6DcEkmKQCXT/mWI1pGqv
j++Q5myerwmwcKEZK1/lz3YpZfGDwR6zwuFsuqDk8GzheUdjvluOIVSUudqCV1z3nFbGE3OGq4r1
V41fOY+m3JkE5UWOOMqvXpECDsVwzrSuSXU+NdvNPiOY+1wt3LeWYVfYEoauwc/SntqG+oOFP1gg
jTpzhWAffH0P7kyK/F+TeqBZj8Isass7Sl6qhZhBeTfK5V877E2PnS2xiFgX7fuCrpgkXRZweG5V
z0qN8lIZfIppRHgwpL4B6ZewisUJtd3mPE3kMMEQC5T1D/DXfjqfqwpfIKkIw11O9PY+zqExrYL2
24SFgc9jDsXBzeWW6N+VLmVsN6epYA7ekCAUaCFiSUHHw+4YxeNI30k0SbyhUWixGVfMZtb16mYk
PJIqeHWzecqncnjn+6Hkp6eBm7daiyG2bxgccrR01rsHDSAfAgDGIZAcvM+R1hoRtTN/zI9rJXH3
eagVKbNGPk+lNIQTYmwycoUxSDV5wrPzJNjKVaqgT4G5802YaFANelfnw5AN/1beLj2/3DlDwB/U
4VX/HfUzhEnVCH2hRZm2jTgiBvtvfKRgE7FOTv2zW2Bkabi5BK0j9b7Y30rlG0tihsa89or4CfrG
T+SRtUS/hwVTaHz4F5Ud2r4FpP1JjKDm9hwaMCN0qhasOEcOAJpL7VGML/aD1D5f5GrZgRBAV4P+
vgfZyr05MaKbBxuuKbJji1ad1w+M3IeysYbvbXFqwBGL5w0UWBhz1YzGfNxaTYXIiana5CptYiy1
vL1enWAlgUZZm0CmY2WvLZ0H+VdHBMGr0ThKI/JtfTWx01SzhBUAnIIYgTklU4wlOQfEDXNc0Jv7
8rlSCWoBsDTHtycvAK+LWLr4XVLdL25unHGiCAtIDccX6NkVe93ZXO2y2+JmN6cvsd6+Qebn/CSY
IlSPoZ5BDsmjiIDL7NP0bi8x4cpZWtlVtBw7Ax7S3CvaPFpS13tX4jC65FUVgk94JJs0P3e6HHO6
hV5w+cwKp5AHb+YFmRYdBF84+i6ceKtBqpak8QiT4WQk5rW8r1W+kzK8JrkilA/1D2yE9mn5Z8CM
0WDFeYdbe8XbkB068ZjxkirfEZf+qhUbTPsE2g6zgi20MpOtyXzecu9iQFEAvwtsNEsh4i/2vRdM
9w1AP9s9tBqcIQZa0cbETyitpE+z4MUXvYCo6//7CjAL262nN3Ef9oPea1WijxkhXP+7kMuFtzUN
Lwp9PZU0A/QzlRJqnsubdJWHsIKf5E37E5GfqRv3l4WJwFCzyxlYMvFHiu3JA+Zzw5uKJVLpoLlk
S/IF3quaM5rDjGp7tJShAbWplvW9JMUKetOkX47AY/bo9m40aLp/ISHWIuYEWxk1b62WsT5Z/kPL
RN3PLXrdEyu5lXT3A7Dj5u5Kwn6GgzIZ0x1z/Cu0uulinFZGmn7pRBILJlnumvFoyK1IdRsXej7+
eGUSFAZ6Gj4h0iKqMIqHUPnib29CkPy6OHwi7ItZCAD2n/Vs7McRB7jeGLuNb7IakNF6FNA6xVJ3
P9+N4ozOYzkIXUhcSL/BNSx0NNGmZXnaHCsEP5OufPCPf93cH+HJKCuz0GJJsfCv4WlbUCWCqq+W
1U7xLNUSuvmZ6NjO63f9eGP7q8WSKQGFRgmHU+FMb7yT1+sxwPWuY7E7cICFgdFYFcCh6rZgwaKx
aDsajYVQflNrpfq665HoT/yVKdSQNR0WvZAZ3SfsGgylPHPMQHn//bGe/jy2lMZtLd4S60uJbE1y
BofhIzLnY6lZINVzEGMY9ELcjlbk+6cy3z/xNI6sPfRIdDnfsUD0vmP9AK8SlpNQxksQGh4tXeBN
O35vUCUTcMmtQdxQe+3pYHhAs4HRBZHMPhn7wZl3TawAzj7V+MR2E04X1DCN1qUqcUySZWhUAz1+
rYNSfXOBKIzdUkdkQd/xyKVuOVy7OnIEn5GaNRkp6M1GJlC4X+nyLepAG9wKXsP3nHJgiuDkY6gu
VDynJAb380Y5dAdYIau5QVpUlD/RrgL3pHTlb2KZwsmMAkQ95Z9HSZeWnHVrIOJnmBE0J0t4K7/3
jWlnByUEQegpKCMCd6h8uVrAdDnAT0fjDrpUotiYxxWxugX/H69XrToghx7ydp3nWtz/QsFYwSQF
rGOjskJMua5kyyU4wj/OtTpXkUvHPHsygnWf2MoP9HCUpnzpX49/PpzqnRVPA1AIWdyB+fwGkm+u
3ApW3fEIQW9aDL42YeEe0ffvTj1+7MTibXDLQ+i8toDL/HwCzPjMLsyaM/gK4ZDZqlz/d5KfN/Q9
XdO/Y/Bg1lDyQdx2KHN4nrXy/hpf9G8qo7QXnXh5dGNiPhBi7LAOWOd36ArscR9JiSnLhgkC/fCJ
y74vyH3d2qtHNYM9hk5e+Ox1178Y0Clc9eSTRckqKuo0x9QepdMzmoMcb28mhc0JUvAVD9znF3Fx
I7GBGIeB5MqM05NXXBX27CONldJZL0dsF2dBTQnkjjLOIbJGS3gTYFXh+waHNyF6m2FXjYm1GdTW
FFDyXK94QHPeZ/uuZ2tjQxFbfowveXRknOEQaLYz1M4weiuuPEs9xqHF5MQDfJI+uHCNWZQ+ibNg
nO0J2FJewtHPyINh0++UIenPZ37hLbRPbqgyB9nUboN27okZP6Ytwl5Pm8im3OUvW8nyX0pYntZE
xiyMX8MO5i6omrKoRb7Pe2aiLqtrpDvNS7BshmJI3WJn13po7/bUnyP6leyP9JdWO6+fvdcmPNzf
H2AQrJ+fN2GPAdC0qUj6FIbIWRfT1g4MH/93dmFsFeYJhGhlZq4J7gmOjK2jplqCB45uhgn79UoL
Gj7NNic/10KXAGxFxWC09cuwmNJHpTLVakRWfdxQ+iLBZDgCiiL/YYsbgz2oPLlX97aHVXuDWjgR
5C0U4p+Wf1Ps36DkjtPXCYZg9YUUvz9LssAGuWvDJBKyPW2cOz5b9EPSJ8itY41V9AaQIvzT8RFz
Bh7DaVMSloLsYDFlrCoe6Mz8f0noBHk3Y5ufvj6HYluCGI5HecFVEOv7j8pXANMcjjkV7Uc5XjSy
ucfKOjm4F9WROLvSBgB/lKV8vJt9SEuMH1KuHdl3izUfBF7Ya0L1a1yQkapAzWFXW6HV2VVmEr36
NDrDpk3boAbUmx5luLhsv7DQ3TGnFL5oVNMKKjxIlfTrZPZNtK9YbOhr0Q6YGBpH1NVPgoOist8K
jFBof52VHaQk0CT2cF/DQ8hDd7mz3L8xE3p3zbCxSgMIpZH51cIMghNrDcSpfDikUBvToxGj9M5H
1ZNbIyeONtbix6yApIK4FHEVHClnhEvFZUz75BtSuOhJyr3xCiHdR/7s16WarHxH8FiHEE2Bg66j
HcNr8xV8L/dGNoj7CXcY0+7cVsBPBOA5uOw/D81ImGzUodKFW+TQ2lbk9gjimO32kcqJ8R6IHnwC
kqaLRZHox7uYDgncNRU4V2cnqUgajmNISMEY5gY2EHnPwcD9ZNHAPjW223KAOD184GDfRYLTkoeB
lCyvStIXPD1u6tI7SUl35zj8iho+CwAz0Ep9y4g9GvEbZPIZb8ue6Y0RpqibiJQF6DBYx4heyhn6
bhcB4i/7Zh/NcKiOhMb+IN+x/zKl8OcVuy4CuANpZruFGCFWfugTNUnt1bD9t+oq1xm/OGAtdfd0
7xk9QbsA9dwuZmKHReOFo5ZOHjN4PX+GlbTzIN0PDbmkqSmjq1g4R80ttOu77huCPv0K8pTuXB4e
TOTmVInpLsB1Fu9ZmFXh5DuS6onhFs9OMCVNJLdNV7Kn9sPm2cWcg3IRq8RgCUxU644WWA/j9JPo
VNwHsxFNNMCm7S9z1UfN2lhpF4azvzKtmfC6HA+Y2GU6mBlcW1fumNuPsQnmV6QryvN14tUknekH
NkdLFl7XLTbeGzjNWYA7CYdwt8C+UhEqu8LqK9St/jraGqcN1e7mcnk/x7f0u6OCowWV7NMu6rMu
iniCsUaJHNzz8umO1QT2H2ZQrJvf8jV25EstV4poepH11gPfyUG0bIcJr0pzXWVd640K/XFbJByI
geyEcOir9G7ipikGPbn6BA6EQPjqpyRo5FLRKsNQ1KFyS2ALlriJjjr0Y3pAf4/6dvE1BK81/Zlp
GW/cm9q2n9a8DP9BIaBclerYj0W0OSt/OlXw7CM/o1vPYU5NfJPe6FJIToFWlX4ED+zKXa/ngWph
wXuoQGjgTxZ1HRCpiaOX8KLlWGYt/jCUaBdnDLZE0NIIPhSJb0YYnBLvnTxtMPNtaKNu3S5etQzv
KV+vdqfkbdR+pA2M2xd/Fdkw466hR9p5Hd+UUkZ2RLGlsyEYFGtAMvvvCVIHAux9D6XhPTxSjG2V
9yLGWRo8p0//1EkAzPpxW3kA5kROKNfwzUq9lr6zAdbE374i32WNGas4AW2fqiEpZShVKXOoN3O2
nCvUuNevSe6RTxtI6SQjQy2K7Q==
`protect end_protected
