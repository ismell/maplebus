`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B1s3mbO/MjGG8pKFImjEd054kGpu6RMOzIfZCWlOh22dWrdNQvZL3YdTqs2+SlcJCN3T6tsLepum
phBwKO7DKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HCfZfAp4nhmEeoik0mrKMJnndg4CI4HVy+gfeagBhZV3JCotSgs9QDaZo78Mg87b5tlloDsjOHah
LHmSpaHLn5JHplK89fJbv4sAQiNdCs7jRJFVS9Zqoxl8fyCLisBSSFK2HErZ/NS0n5Uav8fEPbbJ
71aXWJz5i9f38OggX2Q=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DsZgDclwgmJh9xYyv5I16RbwwNNfnQoHUU58W4MT22vpsHxUxcWRu8jNVKJsgyZ9yyrUVPAbz9mo
7ihn9KAka/UtCcwgAWR/t0XTIEyv2fT13eNL+j8+1CwlKP2Afl4l3k+vQUNBteZL8KHNfdrO8DaV
OZrzGvWswDTCnU7eXg8Xv6ElaQQOorVeo0dyrVxnffjc8GESovw+e976D8qFkgLClrU+hNTAdMWl
ISLN11PDRgFi//7c1hKOSQcg6Zkg/wLxhMbmlC4SbYr/IX6EetP7JXgRnx907tcdZmQYGo+bJErp
+P97Sbjyjews9KuY/vmr1iVMv7wX2x7EZ9sNiQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qxQamstdMFwbx++wvtBzPPHaNCWs7fO52RtqqyG1kwnVWHq1E4TgqxfsUih5e8jsmAEwqn6/faiF
bS800SR/dRgir+jvY0AuICEFLbaIH2ldiQQpNXhmGqqLPGltAnb+zF+kj3g68R7KloeiUGBCSJOa
jQFt0Ia8jUhuXwEDcf0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
phH0vTdQAvcUl9GmLkoOis+aUM/ycGf2jBlEKLjhD76Xe3APy7ihxHfAWUp9WoOKtGZyhekvci9u
AJRGkah+x1z3yPAwZF51SjNRPtmfwSV2T0bBUpDcW7epujoD9qib7Qcsek56SpyXPB5Ljr3KN/xC
7oA2B5mwEB+n74p4qovhOAjWpKMo/b/K/hboTWxaSk8lx7FFWVECa2MN21XmfgYeKu38OQwDM9nc
ekNISttvYdUWGwaOPit89xp4XYZBNYYEKvvpm/3VXtrQMSjW404082z7nqKe3Nfjq56qdUKyFE3O
kA2cXu/I6a238nmHtuOIm2ELii7slHZ32vJPtg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
9l1Z/nTLLxuHKydlVGmmv87RFwSOTrUbu1lqSEZAWb+30PGsv7WdzzwJHsbCMrHJW/DR7MnXkUj2
DuPW320EyyC1sWJkAPGGDePMcRzipOl6Z7EH/pV9rdMCyFm5JBBmS6fZC6dEWFEzArzlL8sr3rK6
wo0qOUWsW+xktoTnqFWAXZtyw2FUOKA5uaGzuqn/e108Mo1Dqi2ItStlM15FDlCABJQlhiz/3GRH
YCUCXkhRvaPanxkXL279keXL3PyRY9leDJU9Y/EBTBJnulFj30D8/QHiVrNbdDwLNa34/vDSE+oF
m0fAx3/u5Kd7cfsW+t9DRddpXirzb9KDwAE1g/IoH8sQCns4sXhfm4dUTNU1Qn7EH54hWfQVm4X3
7jKXM3oNKEoL4ljNIYi4y07Je+KSm+W0n6qwIlIEDjyqHpHhopsSl4iYHnOBfhmlOUXFHIXSuSju
e+ACJZJeVfql6kxvf/s7UuDFnACEdi5q3YNXGaag2ArGf4DLLJBzHbjrixgCt5TPAsN41r0RyFb6
gxoHNLFUHs+KK19Sqdz1FvExWOILAlFv+MC8BgjA0DueOmwGMoLbRqvDBWrEoFDqol6mhq4nufqy
tLy44dNgU/88j13GC6YWTy1oztEkDeTWXSHkdYbhaHOuU8xmJSa8xJndNUmB1wuAgfwEckKl6ggE
qJFLCF2DAqe3gkylBVew9sw4i4QXadrrdcMKrJFM6CL7oJgbh8wCGAt+V1Ogl8Tq1crcH9HwJEEl
qmISeE5LRhIyxxlEtSD8OBV3ll/GLylC6uBdtEl13IW1SvHZYrL13sTSnlaZKRCtxmtqMUswcZYh
wXtfzJ94DT7+2haVjm3ui/JqW1Hjwt6BG8UKZ+Zc7ucFNW9K+u1tHEx7KYXFxF2Sc5if48iYTKQ+
KWRZ/U2IiXFhLIcphUf01wmebO3vUOY1cN+VHvFT2mBmTkqfCP0XNXbbp9Kcj59CXhVcG+kiDWtR
YuQwV9zdzXvZbvzF3tL8v8YSOhE8UkOavpb9PqX92njB0w9p20LKmtH2sktOn62Ab4Ab2I7N2oBe
04VOiuuda8irro+rpj/BkB0EoBjcMjPRJOcSEPlpRgdFUO2y1lurpocggql7lXJv0BGtDZZEtGV9
vrqB75PepXv+10UkWE2lCEkmFQPashaQLWIPkg/xqF96J7lyaAAzNdgv71oZsevSUVS3u2ItjUDJ
8v2OINDXYYtCekCJczzNZmmhi9wLJDmfuGAR36EO21wHd2upo2rxcqhrEPIzhdwrpDltLGGFoyuw
D03yT6yKBrL9nwTJxVWSmHCuJg2sK6rEdXgKKZHnnctLZCo4skc9pzE/iJsSE9hdWTZpb6mI4miq
z59GoMrbVsqQleTIgOd4qqlPSJb1OWaHtav1ypno7moys3KrMQYmqWWHiuhaIQ1PcEiyyxj188Zv
lBolzd2nzFc4lfO4nmXQoVKk+PixNwLjieWVQHk1zhgp369HGNbo8rhgfl3g+TtZwUMW+4W8pr04
zpV3dZlK6ofCrUYIUTI5SouQj2I1CoJ0LgHRO5JrbEkuGp517CWM8Dxeb5YBuyTand0AHU0P0/MX
+4uFIFXces42u5hXy7S+573dzSuIY0OiFUDf5a+f4ZvpsmREZnNKKWXZLI6UYabgdpqsNQ2O3T8V
Hs2TXXqO5wkpYYpYYyseqYUAzly9ia1h0Whix2ZfYeUYAmndUc3xxBdD7a0bxELuvbNLhLc+DAfu
2N3KvyuaU5qqvggwikrhfwmuNnk067LHW9EAN8+oPc9Uh6L1w9GN11ERytvH+OifIt4Bk5xXZmG7
a1H7Qp4tmk+79arNeAQD6WM6s/xxNfLt7DzZnsjJFLLoGZ5z/sRI/dz11eTLUetkrKPh04LID7qK
5QHw2VsIw5RSWCW9vJJY97ZFx1xj72+pqAyBkyHYqf5Aub6JmbXJ8CuqRpOKmdE3r2C6voTrY18M
mXxEqmP8saNm6f7XzHNccklExMfxUm+a0f6vt+qY9jmzjl33pPCvMkZItu4U1y/6Hw1etAhXf/yM
QuV3Ho0n29hzSG8h5h7V3nezE0UsW2jTzWVCTRjJ3xNQQtQCA0M0bei0yllq3K5mnqK8O5o8nWAb
wM7TPGUzQfB7kKGOCxfo2cAvX78R5RAq2MOqCxpix2+on1+2cqoneW1X9CsLfXfhOdbC4vyX/6+D
XXz5l/EClb7LSPnIun+CCvC+gLKpPWJHfnCpzoZQE/t67GDWe1WIPDELgzBWICoJv9M4SYE4iXep
TPwQCxdC/q3mj3LW8R2wIRnLAOZoJlBWrEQKKvsOAnZjTCRhaWwJHI+qgGxGHWdIfqI65fbD/KAF
hpRC9UZRxqYnU08lc9HGpS0xil4bRS4znIwn0YlzViW9W1vs6AR3SsMnhXlEUj9Xf/VddtVVIvlv
96HXXqkJ5CxU9DM261LHzxOA/psGx45C8Ia2IDRKQLFB4OLuoK7pkjwSe/N9KuPjzCYYyNLf7uzO
9zpwBMu06ElFeHSppMA4slSmi+p2StIWMeJTdecXYc6B+y9wCBaQ+U1voj/NqMwCe1zeCaRU3OlW
A05I9IyzS9vW7yUfgSY+xVN9nASIcZ/lUiGyCam+0TOolCEK4HdsKIxi9lZvTpdmND/MkPmozZPl
p9WWV5iozTWNLi5RoFpnPRD3NL8tEiF2v/B9MIAPhJrSXw7K+ZXLtaIrL/BELLB9d1Sw4V8RfP8U
FIzf3pLgepb/jwfFNojFO15BL4piL+HIX+fGcdfNh3KjGQWoBI65muyi7hGXA8h/F20l5vkCVmkz
/yakCxPpLO+xSgEKhsR40Qxt3Yo8u6nBTtN6qveOVqTHbA2eEhcTKfe9wGUeL5hdmLmbDftDAUw2
DQV1aNzFcFuog+e7JSy+k+ibQb2D1iTR1xqB0QWL1P4LcyKPyeMw0lIB3UFdY35etk8Ghkc+NHYP
BD6ePnYryFauJnL6GGkVfB6f9xtkqH3/rF9/x3zIGt1YG1L8dxJF6jN8K3hwZDjizMjxKl/xoolk
Ea/e6fZBpqFUtfHdQMT1uY/525MWtXq7s0EXVR+fXlTmV+DYIQvdu+zlilD6fwN+Fyns3riBjgyh
AR65wZd2OC9QLXeKMIjqkgSHZfEGAuktslojPGsElkGRJ9v351ZKF/WCIKSqqbMD9bbFQGb1KzVS
kuQAFoD0p2v5jHdnVJdm2+XEZiPmHnEpjGRRdAjHzuqP4tfqcW0qzgIwzO+cTNtjiFALkLkFfkzH
UbAK71HVVH0MDJ8MzprWzONQzQA/2ChedF2WA+FwMBVfRJGoExoNWOyCQ7KMGFM3/B+/oHEIITjV
IC18LFehNuYzjRXiejOfBIuo9rulDdnxvC4EaEmXvjmKT3uWba59th06mIyUBkv8CKbLUo2kY0L/
dPM+h5IGSzbIGlmqhCVoTCHJgJcsVhW8iak5bXZtee+hUYpxrvzd7g85mvfC66zHGVdMPhVyAEKo
iv36PO/0FoBtDoSSB9rAGXdScsky3+Lpy2mMsFTXB9JvdMSTJx6yM6p4WubuWzHSWahzhU0OgYCG
hKgeORq+gsScaeYuVKuQ1mqeALSFpbtdrk8dC6sdaJUwZYvTN66Z+lDUCwibvrxKChM9vvLstTdD
rq4vIzSyK1ulbrgttHtPcHUaoXOdemqGBcYLQF7vx24EkcKw60sZco5PbfsDclLKPCLYVpLzsQ67
/MQv8Wm1ASz6uStnjXRlKB8YLKUR6Pjelp0KHauYRDY+0wVfqS9GqfzeukEIbvxO+eekSuWacTWF
RD7bv49hRtxp8J50KK1OWmJ88YGxMDhvHHPDbr5lNa+P1Gib1qLONb7PRVykXGV64RVixejkEapF
WJWXICcgfJTxXB6tchVeP1emoDDzwzMltkI4/6LnXEaFEU7T98xmlYC7eVTtvZ+8fxNlF5FvPg1E
78kGBRTLhZLUvzbze8qMQJ7zMZiy73xvt6lfcaw1YafO6L4LvwS+QIigkxX6PCRz1rbe1BB8V5ce
Z5n5kZaHfuy1FUcu1SxCtauBSdt7nU13C6cU0BvI9yrsZeehrkGILCjSwVPwnlNVoc6HEQULojZ/
jZoy+AZ/dBLJcsX/OSVm9h+VNxay3C2c3CL+6EOybxv8VSbdiNDJ4GGRD5bhMdGK0d3xuG6xp0iR
oJdXLjcqvY5ortMwhpa3axqQgGSjhlaaDxh5kvwXNpfM96c9nR7Kdh8FTxyGIkZmbL1yeRlRIrLa
752ThKwnXkumbG+xqfiakOsJL9ZDJi12AINjkSiYjTE9Kgz5wzdjBVz+jubhsilsHQ9RLZYqwa7K
swec4f7hOnVm7JSLCxwO3G9uuMVJfPPdDnTA0rYcUjZHp5fTh4faB+09r4rhvJwln9rQrfPD+kV9
UBGEirGZK8g8R8/ZZRVqzpjnh4RTWWtX3vD9e5cspfzOWnlzq6WMskN7prHCLbVGRZmdMPrisfDv
x6jCq3XuEFmutHimoIj5JGaFNZyOpUllofBa8fG3WXNiJMczkOgTsxp8YWUeXWymIdDbiCVxL9ip
kHsafuJmaTtPENnRv1puiWfzzMraf92JiA1X9eftPVznqZXsTlZX2ZD3nM+qbzxjxFg3i3Ub8STu
pEHBrq9BVbr+L+riDF2w1cyV9v5HZuK6+zMSrRH8lBRXiBjg50Fq2m9DEzPaKEYaLW87v7J8s5dK
43GfOCqeI819CVKQJV8XUkU0/kB2G0NMp/g64rGAkIq5aeoP3PhodeKj6wmo8PSDbJz84yA45cOB
UfiueCG2JBNpBwERwKKY+Dc+qrswXQ6z42NJvyuobpTeRvyZJYiPUHD27YefIzZwn1ps4btOG78/
BhK87ZrIDmWuWfjPf6u85csKP/UQ2A2g69ZwbpXuPdGvYWxMub9AX37wS2jQCuJ4dqqQVbcWlY/p
J7vQw6ativmIyXl/sA5lBPEo9LuSnWijnWSu0T+3hyd9kKoM1PZNgRiUWM/+5XglbLttLu8+xZLP
6G2pCpeaHrDW9+YFifcy1YrbD6ze7Eug0Y4079XHcnm9MuBE+C0eWAen+v21rTCGhMLmss5XgyIx
SFCkj9BlUdBs8i6QrwwVGSKJdMZa5O9Ekz1jzgQ3knOdoN46/qlXkbEK4wnKIkfoaFDESW3KTuYc
sxeRBhqdWP+jO44LWEZzaOReJjSIpUPQJrUrgPtsfHa+i4upKn0rhG6Iqjhwo8cE2qXiNYbCeCXa
uFrW3WIaWb5QrKDeDBszc8Yywo+3qdYwddd6V7wlqB6VcNfi6JbRbNLocqsdNPaukxVPSOqrQCT6
KCsXadTB+e2a9HXm8ums7cIITbg8c/CLHMbYsDEs5ZCwhmxCinyF7lBsf0dTLUjI3SHZHWQJEJIg
BWsk/fIbxbjzMpp9Q1Coi8kwBS14RsNE8w1Muwu2gxlhr2WONpMGYo+KwmJP70FBxcyHHLxzECua
FDWLKxhGxIWSDQc1WVy3cn24ITu7gQTRIN0Uxc7D2ojHg2R4s6M3q+KTVFMDFdYETmcOncfdspAn
FAiHljBvk1/tvZYqbB4zsATTxu83bVTcsULWoSp5/DQmyGwagUYrm/k7MBP8cfgX1yl54sdxR+4H
NdZ4R0Qr7i5ZRW5ryulx7JBd4h7CX/zuy+pwK0gEyd/7vPWpzzhdS4+bZu4E/cTVbGTMGm+bdApH
/v0DoF3bBU3ZLBYEqd1mNLSMfEKp9wwI+ID6M+o/5Gm2bYNQ8N5x/KlOyK19KipMhuNjxoxgwo+y
zcyW4Z7td+Jg+Pc3rseEnQH4r0to3f9GeOXcDpYMRnEAFj6XEIB6sjY9EA2V/9SKA/GF0CkJC1/z
HiZgJDsvUD5UdRdAD64xA9tRwT7/Zv4P1DB7/6gGAx5pGVa7oFPnmXQdJ7Il3kEVle12W+XUpNiN
klWJLntg2PGt9yImH/0THZ9/iZjzPEO+HCEHcjM7fcD283goBfYnN7o26zpmMzxNVacK/42igKCF
lzP8w8Kkum4owlRcq1vvuntqqCy9dlaMx/cHp13hCYeWZ5BPF+T0swd2Othh+YQDF6EK6rarTwtO
hikNk08s7o45VyhB3tYAfp31OUPpoGVVDuwmgEooTcpqWWm0A5/lkmBcUaM6x13qdSuf8/z90nbi
rli7da3gVbjPi7WjSm9EiM4I2NRWEbCQHOn4DEXSQLbpwrIV72pDVonSg4IdzRXJJMP8b91+WrJZ
+TcyZ/WkDc98kVPUDAnY8rz5tYWxIZRtapdBNW38hvWxWnomTztV2GxITXHQmhe0ibTz0XIFgvBA
V7wjjfz2Rz3k8MratiYUzV/ag03jX/n/kOLNkaume5eV9y5kNDBCt51MO47wv4uFprRLvT2kG6Nv
texevZBHudxC3P+BzRmTyXvgEN8RbGs4dx/eFUGlIFw7s78LrE80FpUrVXGILXA9gyGIjQ7wnZGv
+jgxaJ5GXYU0Z8cpW5bjijQ/za2WmzmvI3/NgaEVHxAnN7ylJ0vKFWQJWP13OHTrdoCb7Xwc8GAc
JcyB/hoUf2JDKEkMkfcVMOTetMk8bLEiEFUQOlBiqqkqUFbDvRyxs3uxcGVw5UhT4Rgcr9Yfc2nC
FES8mEgu018xSxOq08V34Ee/iq9imK1XXHbgdtl7ViWvMM1UoN8dlvrBHcpljQGcMGeQsH2A3QSu
Wi/IG/CdV2bRiB7EywluOSugN4QPFYuKjf1EHIalr4O3km7Vf4WNW1Ng10QLJarKGvSbUYNRrnBv
4N5VY/c6KObwUIG0mGfG2wb7F4Cqc1EHtOMNu82csdgog/EapmgrD0X+xYe0JrT3tlyrGhkAAA00
hrl2sozuDt1w90OytvzC7fssiwBl19c6rHlDlfGIElO97d2LoBzy9RREXT3oamDTKD7kYwD+z/0u
+NOqQ9bwYH8kYbQETzs4iXkcqZ78g5IflUj1HhNLA4qUHPQ5eHGqXCpdnMKAdVIcW75ELn5tf2M4
Qg5L9zPsREh/UqM1tp+sfOKYADMoWd8piyVNejU0yIpqV9bkPmlHhF6j2T+z1kWexUrgHJA6j6eT
ZMQQIukC/fPjxilBlVV+JCvCuAwG4JLUpAt9Gp24DCNYFd+DC7TGHWCHT4/ZVVwHlaC+RKtw68w9
Dgy0DEeSDia6I1H52BH6DLsKPHk68GGNVv92vV1kmnAhj7RxLmdP5lF2yrl7njJwPmIhx22rpNYa
CRDpZFknmLhLihEz/WC1DJrHc9h7SGz4syKVBEin+wVSpS2yPwTaIzFmJBcz43wBPL7be5fJuP0X
TUby5CpUA0Q5fSDwCKlHWOQAu+fCp/QQbKz4HzR0QuJbYBXaJwpbCOW7u2D6gsmR2Uxt/EQMAn4I
mr2yv5O/dKZY5P132xDabXSJi0TVbsbUqCstKk06C4CVfzZTqy7tgtiNqL+CW3Nnfm8fxiiZgco2
FPsqkf0NiP8LtGDfkczg4ziLe7AcqVGZ+OCbdmA0n/V0VuuHBd07fBDBcWBBANGZHa3GtPRtB8rQ
zaQr2yP/d9bxCEoMSMml4U4FlygrAgo5VeAQG3b0jQPru06R3QOR/A52leYDXll/IbpsvefixnCF
F79qgIX/8/7UuvK/S676ZzilxCvcPMZGQddlFAT/CLu3ttUgtanhOtd0dJVbqHFdkbA+EBmxAFg9
hU61AJLViN3vReGn0rV2F8BO/wvCdzVVKO3m0NkEUW6A5csAg0NNuzZZpuRndyU6NXaf6FskslUX
ZUId/s5bqDltXsr8nb9ZhaF/YX8XzcBB+KGpjrLfbtfm9c5UpHX+XGXfIV/6uXy63oafKJb3qSl5
VJnX+Wv1VLnPZtkZa/w53YI1C+Q1wX+wUTR6iN+9HWN8dIETlA1sEY166Y3ZVsY/BoxRLQFA/9dB
9DMSv8tOcNToe2FfkrbV7xAVgEZi7ItgpxY1fjUR+E1p7nKMz8o4VWKpAmxyXed+loKpYmzxhfP8
i8Sx88SVr7bXI777MyrebUAs2anF9Q2kVRMeOV8L3arMrZNAsNmWVYhq8ZcmvHsc3eset0Q/I5mx
HJp6Wetrk5XXdPMr/+xLQqMrSDhW6oHw4WzHAItGRuxUdac4WD0l1v8BZwwY1ePphQMEhAOOlyy7
/RN1DGkjpr5lPRsbEXcbiFLui+d4Oa9Sle19dK5bLNZ721VarHDpsaAEz9WJfd0Bs4hQMzu4/1A/
z1g8ari5we0WtktvtBvsSn5mOazCuiG4Fes7Ul/7QEcLpUflVr4A/qZXJfKIgm92EK/iH1bl6RkA
BvbMPpVjEDt5AZS2UzduO63AV3xTshf6Bw+zsOwXSPYY+PumDLLzObdQPSutk/RLrUKtm0LNzjB2
k0LYpVcJ+AZ1Af+tgHQHhDBtV4fn6E+/2oElUV3cjLNGYta0EHButpm2q2glblXEWMi+xK55T3n/
ucpBmNiKo0vK6nrxpVrl4EAHnhKQmp+g0T1zrd15qC/357lxUkMqtrn6zBAEe4VYJ6/DSuSRPDkq
6woKq/mzQ9d9ZtqsecUwJ8QidNsMHR3soQqnxsUVetm7d86+VicHXVEr7ywzVyVT/PZFkEoHSnPv
AI/ZT2uhd7orCC8pdmteQ1FVz3zjFjhfdyM12vAbzqoabhSyU//TU8bedVEkuhAB8X5O4Ki6rbdM
XfusiQ7R2H1E2PdMmUImPnFKMqR33rZ8IcnoWdWV8aSRDwGbuoyPjVkwliCW13EWCUjGFHSjml3v
ZAON4L78I6gi9s14mc5LLon4j+oBqveCo1woqKg350/I/IT7BxSU9e08M3glHNMrnJOue2lkDMNq
X9Vs9SK4MJgd0JAjm2ElE3/CbGcOkBx+5xjd56PAwGccAFHOsLj1UrcpsqZq15YkXuOFZ3b4q3MV
IuDxjrK9D3tcU0Y8tIMWKaAH2+CFllFukKsppACgAy6NBhj3nGySkgiAT9zRgWWhmSsIp151ocwH
DknpErO252nvPUEMp1nQuyo9vCPHgY82O99XrNpOY7azYwTpuPJSOeCE2+rpKvIsTBsOZ+LU0fH4
0VZ/K7xl5Qx3eHRxaku6tNPoNAPxZPSnljgXmeTu+wnuUOPpIYDbBdo15wZESyeAL9SPTBn/uigR
fzPVGadOkqjxWvfomwnDdrm50jnVy6z5t8wjQknVC3frZosxPfO+63F0O5vJQrRHb6ThNkyvDybm
7VThgQUeIx5aSO4B7QnXl9uBk24ktNLzr8hdJs9UR+MJKT2yRcMVpa4KEzuPXCd1tWEI9SO7Z603
o3lhre+oW2VzGnS72FncILRy+e8HWiA70vkP4hp49RQixUSJVgqnYKava44+I9EdIDD6jDRISACr
AZEAClT7YpucSxAPv8Eo2XdN4BtwUjCJSw/zlruJ5rWkatS6a0WcDmxrUhocDqyv7BLPYSgX2flZ
rh8ZdNo0BjHHTBozrMoKAaflwQN7OtlrkAZSXpNGlb6gY0RRh59wGxkqAgvTbYB9wa9VL7/zf0ly
7yEBpdYQZGS3sffYbJxZo2jeJ9oRS/asf9e4epkf4t/IyN619egd4S4CuWanaTVcVFKa4g7QkGMA
iHVfEON89hEdLo9n963f9y1aU6vZMbYkfiLmt6EIyorWED4NdZnAA53of9vH9vXk6mLSly+xqSAL
tp/RAluURGCf2pEV61caHNb2U7/X3aGlCOZj6VYQmuDr4+r4Wa15Gwrt+nxEiw4oXLhf32Nf8ER3
tYDFh+W8jiVfKnJ8WSFQfotqtaolmKuk1GH8neSjmjr9/c/aFl+ck//T4wfVsCoTQbebUxwxWeVh
BLuEmkdTr1eZMBSIIZksXFgu9wjguuxISg49BsH+GIKHNgZeX8xiww4OYWSswtpQ8yh14NMy6ZqX
wX84l/YNhlcXJ1glhrU53a2ObUlsU4FMgy0RPsxu41QKAt5nuovPMZbaZH8vYu9jZoamdKH6eadh
mUNmpMyuWeYmUhOurCVFIJ0n0MZZyUJMzFxUxqlLqxblAETXO3M68HWpYoLPZiW0xR+Z5gzBfiRI
/J88HD6eO9RX8YqEW7zYFLN+BBi+L/91rLvFMPOe7f/M6cc1Fk2p2tlooNX9cRqWjw6YfWJXzZI9
gcAN6Rt4n3TDGOyH7CqlaV4d/JBmZ703n7WLmA1KarS0UrpL4dbJQ37Jqz81lDM4+RhYsYoAPRMx
e3nh3DZfKtAoQrsChKweq3ww3T4Lgh1clGnuFsusrA7KfgD5m+kc38CAsZ1j+8dpU5tmt8xJ1p4A
EpFgS50oOgy/AYz9iYrl4hEPIz7kniO7+2Qd5jB2Uo9VIWeAQea6as3Q7ng8v4SNaSdEyJWA6Pp6
lPw3TSErecrkAZaA4TplS+07OHNz/Zo4fHydHmEmigMMXbvxhb1zINNPgOI0QJnukSBw4RBhiLNJ
Pr0IEFw1QCoEmjXy0XlG1BKSFZbD+5IB8NKWnPJZkFoWoTAvnk0QCj+HP3VA7zR/nC0FeDBBYNUH
yCFAigTliIqhDrgdD9LECgXtpBuxKvZPINADmXzFd9g+eiebMXgFRd8rvnEWx16aQ5vMgzAd2dCK
11Mk3h6/9/mSpuCqlkY4BSoEIGf7XgNVGQ/6HTNQo5K/7zUGLg1rAHMhNFj79MDIugSJQMogE1MP
c06Lja7YgPa71/tn4THmMVRhej/8jA3P8SZz0pYZ2NSJumseKeKm+7JC+tkpqw3KlUp4SefTjKHD
GrDIIEoTWxBc+Sh4+HwW86f41Ffs1beTU3UKtY0SUEhkFLlrYNGaRS8jEnwOq73+u5g1TWYaRxvw
s2N0VnoVhk5u5I/fBVcu3DUTAR8uZr1bzLSvGf3N36V3dfYVgBXJ7EZqxrUgnExVtmjtX7nPeXXr
VyNJAZQbSLF/ufc7QfvdRgvReez/Avbi7j0UPps4RUnjnV9I3J8Dh5bJwMPqoRZuB/4jXo3S/nlr
letFRf98FrIvB0IqgDl4J1QPjl4XgJUGPUlMaBS8QxsGXNXzfhbaZUow++83pfqo/OQnZUKyu4IU
LviyyM79cvf6zAXB7hZfqqzkHrCMFonWSeCzbbq5qLdZDwFiCU6Yhxr95yeVrEsKIeqNxS4Daswq
VaKopT4s/G8FK7n/clgIL49pjidCX7UFLnvtHX0Vi2Z+X//4nLoidKmC32opyTl8jhrUDF8jikjC
TnnnAbr3tKgiq9fnTyWyDhCVgScryDHPdKMJbfg+57xomMkE51MWs83QrGTT7569Q5xHxKH3+G5U
TVGMq79egzgoMX8jrQ5cT3NtKRyFYrbQK+wDzClFdkudml67omP0Wh2sh058OxKMiBkWXnsl1Dcj
T8oNW2WytD9rmrfkzpyDpRtDcgLK3DcGiosn2tf2SUFGQ+Uby08urUVkI5vrlmqEV2pMA2FnqSGH
cIvVDbbHtrT4OYuPYvly/BEo1p5NgYK/piPdHOk/btDis1S94SFz9iOZBCyVRrFWIrB1ywQkisjz
Kz9JGjKngRMOzgKyM0sbPAG+gJe9bRWO/KEOwl1Efw3QhlpVNb15D0osi6INohfBz2IKFktm98zA
vL9T+z9wK/EfYPh7NJoFaclAmmNvNLMeOwh58eudzV5SvxiaBAwinhE/jQqs6PGoEf6PBq3M5KPE
F8DWgD4mBHC6INGw8zt2X+3SenmRFznn7N/ivQnd11pwfVZydnw5SFVkxk82Venx93oxhU+2AB6G
L20qcqAOP8afGRcV7OGqsnkDRHtAZEmyJXxMgLZ9mk7DY6ZSpY9cmwTWxPMkrU1SvoAtrrlZJ8pQ
NI+LUkEuaezWYnjraMBUfCITKC9LAw2OsumHVgx07igXQW2ywOsk8S1fAHPJ+sznDjIThCvOxzRb
qymbb6yvMrzIg4aeEvHpmBV20yO6epPLPONtgpC7fX+F5IAcLhn3yJN/PnCoz4+aQEk4C1wMdChv
KgLwQO8Te87WqMgSCQC3m1VvqsGfbOVqPs2/v5Av3LD1LZQX3w8Mpj64k2jQ/EoUsKCXvSosf+FW
SOHZZ/aQa0BBhBJqZ0mQ3AOd69FdmX5PGJQ8hFeqRmMF/mC62RM7crpij4cef9nrypx0M4FNgqLF
QbMnx+bC+m/omO064Qg41FVHJos6aKcMTM1VoMElFdVB08mjgf56wJRA6zjLvRH9Mu1K6Spr0ZnC
jYz2ChrXly1U5Ja1HeGzT4hwLttQP51X4BQkymKCGMrcOFbIiZ9Zqnq/s+XZ7kbRgVTesZFzmzWu
D6D84EP/CPryqPI9jlnZDJpaJ5TOiVvuqzJSUi6fWnrLWm7UG99GJRHr0qtTWBxNQnmOe/V52WZ3
nNu246yM3xvLG6HQjsDs3GpVaR7MQbSAmaSyrLB/h3RNHTs2EJlpaaAP+bEqoc1acV4EhgZRtL7T
K7SEcdNa8mzaZb61s+gb6n/QVnbN5Ys1xWF/ep69hPCy1DsvHGqh5S4FGBEReVEGtx8ehp9bEz4e
jvwc+vaHXTMdyK1YcVMhMNiVXxi+27ebnQp8EyhxcV+stfQ9DPV7hZNvpeQBucjOMmcpye2WJCWF
RWPq2M3QrO2M4GTs3iJw6dwXibkGBAEF3QB1beKoVOxx0YoigDNt8glTWTzssc1IUTptDzt56xRt
Ni6egSShlhH1A1jjey/6yw/adGt0Z1rfc4RfNitwwUAz1WCmmLUbsLlmFcqI9552zKombmWx4WJc
0nBcHH4HtduBTPk9/sO4NPRtJx0OqAgRPiQZXLljbF1CK6THdQirl8IMLRsixV+gNTwGZVTaj/xD
lPEPLSVd3ZtyQeODuA+EsXWIah5jMsLxsqjcEg7pW+ym8pESFEjdaB2LJXK43sRUZaD4o1hNasSV
lEUQdifrv4qvB18IWDx+RSCJ6tGMNckb13+JIT9AkjnTWYYQLnqfpwFfC/2bB3fkCjo6O/FHxI7W
uQ7VLRfykTUzChMNeydeCZq6LDDAVscdcJFORp9LiZFf/zuOcEFupbLvZ9dXFdxStEeTuC0gtwRh
COBZbySLTKevs0pKa3IURMDClEOofVPkRwj85Ew5l2Rr7NUMc6sM4y3GyUzsCtq7qILWrw+Mmdng
OYNxwxbaQwTWM1S/B4jXD7W5RIosDkeQMOvyBZXAvOuZ3R1BMy9dr2UfVYVb5bTlbhzhlpLabmNw
32+TTUnd0iMcFaqVJqAfWZB6ILeRQSt/7HUZHXTgm10iNKdQntSszlX8S9Y2197Wnjn0IiBkvho8
ht3If5S2DH68rCPDdIf4/Rqo4y2gOuqNcO+UH3TdiC+oZLw0X4lw2MyvazdIZvOf4qHGrpwckVH7
4d8IaHoW5u3K9qicOXeNnDLSuoIdxduItiDnt9tLwCLqQwNSZrAGIZP0pOf7TwwTY3J6C6G05NqV
XUu62nyWD82PFhlNMKEeLKkTmohlS1L8YUoNgT4QAH2MHC9w/bZZB9iqrk1Yx8BLnomVI2xE5ux2
itXsv1HJsJxttq/6wPd8acvYaxAa9BrhM0J4ocDnOPTjLFAB1tldAsachBPaZqmGiu7FV4f707vl
TIDOXx8yZbx6MVY4/Le6vnHOs/TqgDnaTYPvVKymr9kvx9MXGxpzNGyLvWo3P9xDEwGepbYnpC/0
BVv2rKoYIL9Kfpjm5UxsjupA6wCDuFqvgNERrVly1tLgZgk4Lgr78gmFOy/1XLRbJuZfFmtWylqj
xRNT2vKxNc9/sSk3Tycp3DyqBsj5xWyVjnzICiPFgas++hcsApNlUiquFJ9gZnjgRayn+q61j3H1
b5r4cYT592SdR6YEIMs7FMej8n1/6+9rWExLQm0xUyIBZWb22+IblDLsQyxS+hDYaWYiXamuJZnA
2WnxRpWI+ZKN6YVmDr36GOiI9pHS81NPQKQ4/VLpfHAmg2MrN9ZPHj9Bvjw3UZ4s6VkYF8D3A2Tp
no1KAkzORzksPMCMpz9DsMG3bK684tp0CkQF13i3xcpJP0wpKrzqaOKOCr9k2A2JCvoOF/KI3OxU
7vD2STV0yD4UFgs7XhRAVU8y8Z6K5yGsofvC3xHHyTZ0ZhHdzEkwMikk4c0JbLXbIHaMpOQuyHFa
faxAKTC1QH1nXFJqm94SsMMLAEsFkvSRreQfJGZSp4sWQEpnewayBK1sTL7s2dJQ4Paem/0Pz+mV
TgAVuJhk7/JzBQCwZF+U0C6Q0gOg7ByDkU3jC6K+sa6cyZx0znXIB+BlVaTRChaOt+J9JE6C26n9
E/hsB9sB/yFWIm7GPpuhFtOO6CJcT2tO12ufCmrstIHuuoMTbYoCnnXM4AxYleWu0v/UZzC0/IPd
jCPI1nj1jckHPbNCRu0saIP2lbkQ4LwMEOBwx1tJf73oHR97I6Y/cj+rTmR60twAgWXVb5SDYr8w
qTetGWwY7OqqViOCQqoNOVeHIAAgDBIWZ2a1+dwfqb5DcvyuZCBD0BvgHVtPHJfLq7G6Fw0bKpLj
8+6O5dVxsDElq34n61Y77W7sI4NSMZRBPJQd/1J97s/Dm8BuWb88uXO2LrPlDhhtlRhISSe384Z9
GnaXdPTQhhryx8t3X+gAxHHeiFrlnNEcoPun+WLiyzHX+gu/f6C7pedqzSsMm/J97YjNuqGPKx7W
0JkohtBPBnmm0TyR/xJA4zAUG/990xdG6NnEX6NlwOWkDF6KLjzZ98LBEPP9dp2SBQr9rsv2ZdnA
zNt8xSksgkfBbdy/1q9wiE6LN2HGnwPgq3eHkFrKhIyrlH+13Tw75XIBoAZfNFpLT6aCDo4mviFq
//w09qf3SW1e7CKzySzZX79gIFuFjTcsIIMdwriwdK5s9R0/9uT+tgFjb1f7YyPZ5Az+QzlsQjOr
fx0TdA9RJJVaxycCIhXSz5Bnizg8shuLsQT5fmdjzbtu3f81LYFfcNw0ooEbdjgTTJWQxH7sA8OQ
Fr73syyZzivJiT7XfnbPMRNH7tyCbkxwba2og1LfhPgaEX9gZOyyxEG+0EpzeBaQmXU7WSYemzG3
E3eeh+dwQtjuRirChQ3w2TLdZt2VFljemgQV0Yf6WoZMjVnYJ7uAicasjrEHDREDrsqUTKM/A3Ei
incTo3IK6+kw4qp0K4AErj/Kd2vFwyahqeiP0uX6JR9RsV/lqS9WlUJdTleGI2FxQ20xuWZ+Jajk
BX3Pxuv2rIB4V5obP1BoKAKx86qtSO8yNvwai/caXRqtaM8u6iHJ2kXvOErofYI5A/4RjjUzQ+9a
gJeGrcYHsSHEZTFaH3F86FT4w4N+zrMCYy7kt2P5fojBjc/0qlqSE6m+e7uLDhT7lKKJE+qq4Mme
Qiq+FksijnzUqOQbDqjG2ZIZw7Dl0PVItJoRd1s9qGlvYx2D5P/yNdYY0kSOLgTLjCHXD7iQLJ4M
jetg3GLo4RYgOFiJS97YXvTS2pK/wp8zIf5K/9LJnRbRgQqBPVI+dNuyoPvwpGl18lCa3Tl9/Ujg
nABNES+kkwXnH0fmhISLjO0YLkuzUR0EpQGh9MraCta0WrWzvlBPTAX3Mdr4Ld/Bge4gHLlSPFjx
slitPEoSVOi/SEvY7kwkeAGNCLk1zGgXOQyFl+M5upGLVdXpJ1DVEsYCwmtJcws3UEzHuwqs1o1g
PqUvSXH1ZJGOGsV3YNbd5WBZcfEHgzQPH3FO4+xIn+tNP3YhwC+lh1i1CvozE/R88x5GkYhkSDvo
AkmxKG7fDyHMJ/V65kCqWGZxdznoYtND3xwvFXGPgeE5+fafENuUux+6sEnrMPQyJqqbWtRXIt0O
kaXERX8Mh0oYw1I3hYDUgghNlb1T4axdrPldgxau/7JnXa+P357JYZsT71HDj9SsMnQ2mQVqVewJ
qiyqrtH8B4r2eaNLuge/pZtjbhaTN0ZRoLm2D9+1bOQ=
`protect end_protected
