`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
isrHiAxWVRJAlvHNm7GjJHAxGt0pyvtoxxv5t0Wd6WB40cmMDqHcfYDGYlRmbGHugOVsmu7z94BV
Auhxq2Oopw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LfGKz8fHsYhrbAXeSgdX7Lp+9ocoAXBoY4EV95aQjceOUd9zgdFemn1D7cm37K1fF6MBnPxU+1AP
aaozaItnzT2wxD2H5kGzPn+OmTnoTh2MtnqxILq2A9lQTia94KFlty14W0EXM4uIBmobMY9ken3X
dyVbR9QtzLt49+JbXA0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QSNOHEeeuUeqpji7ip+lMNxlARVuzEUc1G0iEzT+ysTlR4XmsIueBaX4wI204pG9pp+VcDVn2Lz+
T/wnCVoCDdUsF7GcP9LLytmEX6M82+LfPvevGX7uw/qMAJ+kpR+P+RqArfg9kerVKBClVMJB/TQP
h2FGRIXFuqKZbH2AajbHA3a7wlkfkiOSsAg30PRvuCoJ/unw5X/Fag11j6PNTTrrijtuFN73JNyb
5kOC6tKyZtoafGyO1Wa/36HO6r/82r+ll7826V+FzmYGjc1MHD4miPT8OQhGqd8dU+Qpe4VZF+J+
mMz/IA+9yJp+9K6m6chI8mivkv/eF9AsT53saA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mebZ5+XGavNib0tp8857kJ2AQvUURTal6lOC2EqBJ7vXqi+hVSpgqZRUeltrJlIthAvWQ8FgqPqF
ivCcoPFtP4OhL5E0Z1AYLM7+nD2+6zwjnHW0aFb325QmOVjLVMygQMWoIbjoKCeX/MYlB8V/tbzB
MmIVCJ1HfBLthyBvS/k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e3f6LzPvgF3mbYxynCmrVOfzDIctiZTHRtxeohww7Sq52zZcIggfkubbw3DzRxzKZla2HPNH4Wbt
egBQpYQwzhFPmLK98gpt8oA8jvC3ypM8SlvAT5gjy7+WMuwfqW6D1WxmJ2tKx0ArN0kF6soS3xdd
dtSmkMPKh76J4oTMIKku1vkgPbLCDgD1XsVAg7adQVo2n9CuQGvD+2ILrnkzneyf+xkMdEbcabAr
VDxZjRuGh8lLgBn3LLP3VbGhM6QBB8SM42+MlpGn0/56QcbmtnqhJrTJBTFalKfy3xmxs0MbyOwz
L9EumFR18SOY023UwTeSl9pSy8GTFEeyFAK4Tw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 80800)
`protect data_block
xp++znWXFMFd6ijegZNckFOno9DgDMDjQJqV1sUu+r9AFS1J0bcdCRvq1Cj3k7LEMjzs9o2KfiAL
1QfXjlpY43Vo3oDXNcBWpvqcDXYH/NdJsONG6cjWu/qzyCBXycz/4VaCCgx+Ia4c1lGZFMKIjj85
4jtVGF0hsKeDOmgpcQXZNdTBrhuwq9bV4kc20fxquhH6ub3lEFxzcBA8DwaT51NhbCZk13eie/jo
1eoemBxS9USX0J/bVAHzVlU2xPSa9sSAP7iuRgwPhRrtBD2Br6sO66CAc545sD7l3ccCVu7U+Y4+
rzJY5lwc7Z7HqAoI6KaCcclqBUW2+U6pfdTsqMK7xeSnjeZjZ/GPmjvEUMnYBBGrqYEIDuFbdnE9
UqMbzM0S8BkbuYeUSiZmaFkO9+CUWRB0+2s7K6GAQG6KAhbFubcQrb0OYJKnt2GIo646ft3e21Po
P4ihK5uUC1Nh6kfprVmdRIbYZMFepNMJyC98gmC0sRuRWbg+G6lXzlIzoQOJZVTaHKduHxHkBDeu
5Sm5E2ij+/aSry24QBHW4ALGiB3uwyKP2aeiN/bdRiQ8njrRR+KkiJ/9PmNGq13shy2YKgN/eCuY
FfDxixtofZuONMMqgNFaAPFmORnpSNgd6dVKilMv6PxIUPFj9Qs4AUaQd8K3nV4yNniAtlyqrr/g
1HSbxJa52I9cgSZPBeqxZ56DhwAcolrtSOKU01x59vcxV8SBr4S9AXMqJnIaDAL1gsLBMklwLS12
cZ824xPfXN5MlNu22m8PZMOH2ee23eqjREllHPy2zuhAhl/rxRnSvPMaT+G+1ADtBXz4jc9ViGkF
0hcjGfT6Q2YSqiAF3FKck7/nBDdEwY7+CwpGFopE0gxJzvr9K0z40+yDO29SsaumeRBVwVZxOuRd
5nH6iCZnzwUxO3r2ChpvH8rxbWG/gXZ2wMfSq4COJNS+ocKCWcTIAFOMX6oqldNliW8mpv/3wICk
gnaYhFO8E1IKqyZmU83gnRLM5Juv/3k24jyMm93DzanklWqyfac4eMp/Te6LBNUoacHyTdW7k2Ef
9JyNbftA9aO7Bs0Vw15d6GHAhS056RHcvwZ4VOi/vi1J1JqY/1TA/HSMUaTxVmDo4h5eg6p+K4VF
cot/6Zsb0xpWdtS9jMfZiQe52vc9krAyJiVdG5KkeyFnlYOcgww4VGo9V8qX9KrAiOwZwTYIL5ya
qsdO8jJEMm13d/O5QLR/EIDRL+T2oJxpNkLfAkoeKV5qo852DbFnpwEfNu7u86qzi+O/KAX56jOx
mjMwEjf3l8W3ZYPlTkb5LcoTLBCqHC+KBL80ieE3LkBHh1Mvtirrr2YeCgV7Ik/SmCBvRte/scEP
3Dx0bbXfz6yjxMFUPWtz2xGmNGRArraGBNrjFgbfZVKgbJx7TQD45c246ZkZC7ba9si9/qjaURJU
1IXxM9z+kntzXOPIqjNuVVyx0mHossgASNFi+32EPucPiw2RACG7i0MMk5vglxPENFpM+AbrEp+c
wvQtjZCMKajoW7x0/ZxmSmdF00bfDVa+2afbvzUDKBLKE+QC+mtJel2wH8ayZ3H2Z88ho2FXFcft
OqMm8F25tSUBqPOv4VVKgjTZYKaQusudzXRRL50R8vSxJe991Ps68qUXkwHkVKNAPUV762ZAB0qC
dKeedxMsFQjGpSL+sH1iH9IJpWyf7Cb5vZuyugyqgrtSXC8aEt+HQy1dKbBRcxCy6UAFPFheLV11
EnYZMm+aq8NNL/QQL8n6KG+iAi+x5JqoJOgvf7TQWJvFvO3462EfJzYlDyFfnrVilVsJiAEOivhq
ABiPk9W+21BqI7nLpNCtgOCCeTr/BoUcFDqvS5uelAihUpB24hZdr1decAx0kqds0HRFUJIXIfYq
ctTTsqKXst+nvFE47i3JAkGRyb9d5ll/XqYJ6g3PSekrvVmL5dU4LqlVN/IvEyPXnoAbQAaM3fVe
HqhkJzAC63N2GJErb6tYPSzERkRyTiMvCJAPIlHniGsM0f5vZcfAgST8qGzAfkOw1BP97/eZS3r6
V/Vjzyhy4EepLKVPBowPqBCRJSCcoD99hRD/LyuMfPH04zLdJf8Oby4fPGTfILKMxnzDFQkprdpn
6HROJw+wW25QLS1ySbHIM96Ydam0eo81uqssRNMEuehxuzpqw8PY4d3D1sE7BDxJzGG/T1C5LOtA
/T9Qshz6sDCQ6f109e07GZNt+hVSeVQ+fy5H5+49ZE06Pmgkf/wn1++jCvJIdR73L+S0GobAAldI
FMLlfmCSmKqOd4/M0Y75+hDpfZFjIfbCe6nElkdJP4VcBC6U4Vt3RVnaMXXHs/kptlaij80mlKhn
hjph8ri63ZhyZGg/IovB1c2TS8OErii4QNJyCRLKyBNSQEIgM/w3q6mG35bLa+iaw3Z5K5IoKmhX
EEs/JOESNUs3Xty5li06rKsnTTSGAySp07rz1R5ZZ4ix9SR/rrvQmTks5TvQ2BOjwDEwXeD5HmTr
x2aG1nBgBPSmZZx8tHFfhj5FGRw750QS54Qxepaf6A/iAHlp8FkRFENnMuYeU/QJRE8jNKa0IBx2
zkMyP5FUvTrG8lvBWvD6H5z9sU3v1nFvSEZuchDrg3qhVDBg1o1enN1raslEu9kSHoAX8dFc64nF
3USU1GilupTqXNZUv0jTFqcgMyDZV/jCLQUDOCBgLvwkrwlJY8bOKz5hnuO6MLOViHk6xLprfJm/
lOyQ1sVi4yoIZd3PqDoEy+iQ3Py25h60Hr4SoYH/Y6+0jQSe5OiK9JfscDZFyCm09sbjEv/+YCdy
rp4Si4SdhPVBQwVCmZK3LRKpufWDKVem34MgOQJpuZ4RDIMvYbVpYZM9uTKS5xLF0Ti4OsctPI2m
Jr15foCnP6TfFdbnVy2AsC4Yb38weo2mbnxq9MHdNjqpi+a2nQsl3JcDSOl6CJ2Sf1Kmi71yQ+A+
ncV7VSZ6xffeOa/FigrDjfV3cK1wEyr3FPNX+S0W1pDC8DZTgNNl9p1ha6sh5jrxBNmirz/4trFz
HJGYjZcm0XBymlcA8b/k96N3dbPStlLHUN2ooxekIaLFhcwzGwZ5lg8Q4ikBHApZi9R6/MjlYY8m
sCcFnyCdGfsTUODqNg+iGZQctbtStNNhX0TtBq/5Nk0Cihc2mDnZSgmDKgFXtRjMSdLQO4RftNuP
RoV/V7JWltOxC9Dui/LA1bVAP95wPzCHpWhOzDJ9mUW99Sro/PP9IoyVMSgm9osPIJ8ggKnWZR7U
Br3dbyRwNyZUKVvGs1Ig2lFxw+AJpVjl4cgT5R6wb7/iZtyoSqw9YDjzStVzQJEY00dTCHlnUDmi
tuQUkpZIKT3cJeIngQm00CKjLEXvpNvgpdi+233PqMBszRsjwl6r1mRF3JY6awkPTXnanFdsQaHt
mNPdUks3+OXkEfG63VRZ8Eop/3QCcwAH0123/NY+atXoxwhrIfhoYYBAtl1pEmQhlPm+q28gXz+/
BtDRoJ0+PurINffk6AgJrKaxRcrDN6Dto0UhsLuPb2JvbCrhQpvSGd6j8lrwMsbA0xsXd5T/zLMk
y7wtOJ201KwEW/awAktsCffstXKzwAjVC/qyAG9GWVQ0lGPSRSbTXXUo7u8TEseCCvtYQz+y5Rkg
IkqpR9kK+zdlRlN3B4s0HTLZIk/VlQ42YQco+STgkQSyAHce3NamHJVybaJ1WsaeRc5X53uVXKLA
4cIKXyotaTkVbjA8yNrAczAAr2wqcqlcaesLSEVkxEQaNFwO35Jq9PVwQdh6SEvNF//ilWIo9shc
vBeta8dL4z3s+uQmDlIYU2i2xbLhUcxuYNmDrZyJoIIg1QNq73Dpk1QeVEFo7T4YvzBBXDoY+4nU
thhHVa/XVwWdp3IX9x9VVi/Mge/JSD2tPOV42gb5F/N4n70NMtSTsXjYM5LNPYPCUqKwbFZAPaXx
CoOcG2vtVdVPJHbfIMU8FcxEHZzdlz46/DVonOlR5dIY4YTmrFY60tAzpgbbjpKij1ur6IOs52qz
CLi9yWriJUtolKOelguCw6ggGSekOuu7eQLXxlutMLLpyhoutXKp//Yp549I0nqpmw6oZZGnYkd5
3ejr8QPxzLsBYXyL21aeefO0b3maleqehkdcyQeeKj/enlNAf9NHO0sonab/dpUZ6+wdPMN4l+sb
Gb4rGus+1gjI6gt8niT5wA6xNYlxRPLW5eDdOhOUTuCh213PEMChVJOszMrapKIUEsdEzvxPhFfE
0IDY1anJzAr2CEK2TrwSeSOBWK3ksXulh84z9TkbVZbDUgCLP2el520rMNYB/0OaRt13nu+Ojmhs
GOMdmhLR+K28AvGRiTnVh896OLr3DsWf05wV9CNBoPvFek1SfxB9p4/sGTJMutVrSKW///G9J8QP
ItNXLIN1A+nQ3qQCwwdWULMBDFY9jwF1msnP6HJ+chnqKeIYf1SZqzMhDUiKvvkWSsG/aouwzU0W
wuGzc92mkjWEJUkwp3CvFfsyf+NRLZLNLvddQUwhrWZI+HvEthjpHsG86f4/vWn5VACGuo1iVC/8
r3G94AW9ZjGlkJuiHeIa0D81XnbO7w1xmHO5BK7BE84gPf2vkHFk7oAeFTZlbCafEejxh2jbEUO5
gF7Eo9XSMk/F+xWdKIIVT1YeZPpNI7mF+EME5xyGNNkG0mNoZmxAFya9cbonOSdnKyoNCid4eRL7
zR0vTBFo2b3mmwIVc8Wk7QpT5AxTGBbvUD3jU5NG88CAC+KJyJPjBPbqk/1dJb6ssCWVG3T4NVCg
v8/T1aHFNzacFwe73IkYwDXOr4fdYDz6png2x+zGNU1lWkrXtLVV5/xjjVMXIjBK1DL5f8ukr4Nq
LM+Eal9ONYHH9ySC8X2ZA+R6El7zwOr9zDuA1S/L6xzZU/OVowtujqW9MZ5q9MQf9mK0DY3VttE7
Ors6fi0WzfHdkf7TxiBfIBGitS3ws3YneCBVjAE9xIsi31WkkSCLIg67C8KqSznNhDgrQljr10qY
UpfhPfckQ4e0sBuKMuXvG8lfcu9uUkhbYt+RxrYBFHzYqSDwATCpJiRnEVRBhOwz3Y1sKhxT3L5v
mLb5slh5/CdxI+VxBBOesn65ulVN6fvnHtOe7erjmEc+zYiBBYvhipg2YqwSJ9XJcevnJUBA2/Wl
caFCjBJkc/zuNfT2nHXtzam+GbxPyDtW8kap67ENaPIyyKkVYx2f5rgriBjzKRoQuLG6Onka18DM
uREz48OrxrNfRvooDyqfmaKZzdS3+t7VmTv8jTZ4XCs/4mmzwA7c1R1osPRB/RylG6DJCeYU44fQ
dAABbIKI7fu1X2jHHRQOz5wy7N2Yd0EmOZPZaKLtmIGaPTLTcXCZZR1QGbxC/6arNEx4HyVv5L/X
5cqEzXeAe51bO9QPC9jjlm9NRD/IdBldskoinnwWBUM7+ts0NebAr9GJH6umUA/OVLSxyo5Sa0Gd
bESofDbOxhycEKEZejvhHLPJHBh7ndx4I5AZyMt/gEFRcXW49+AjZUg4r+b4/01FIJhVAjgKnzp/
Dua63tNQ7A/5DU87XYKqB/Z4PmCB1B+DZbJvihm40cNKZ8pihqr/V48rGOQS64cAUCNIlY+dLSIZ
Uw7wgC74BkSCr+zGwq8DTwefqQiMtLtsEtvNbJN9xcouj34V/C9A3zUdpa/90+RUWRdzw047XMni
TYMjXXo+gLBKobvJmGo8ydJFxnt6ayR4/DCE+16+SINQn1YG77QVg7txHn2Yyxj9a0O29r+/iUXa
r5q8SHmAjHSL8Rn50LxzaC/ReBdSOaDOIgw4N09/cDpb7z2xsp7hq42OOIoJs+C54SgPh6cUFz+6
RVQSwLj0twaITwn7sQFzPwlspfvud5HYKTUuxv5HsfrA0/yE2PTLv1irV5uMuzzwViriBsiPQt0j
HKzVxvDwDvdXJghrkY2SHa3xmCJKpO/rkdPkNxKmiMGqtEIuEGHxqdcpHZYEgphE0SY4W6wnUpY/
GyAEkKR3kuu1RtA2MOwNsSWHDDwjEuKBiO2bXud/x3XcscDn1bglzxJL+GWtiPHtKw+YB/a4gpvS
0AsCVhJ1l19awaHjjlh/to2F5Ajr/cAC3YOFXM0qrVu6H3mPKf4rpUDqbh1PeRjPzibbyOtv9EPm
fyixzCtDS4l99ITQQ9NHQvsQs8f+evqz47+n5Hp0BZcORhJ/ZhoeoAnfNndWXUHpHjb1rDRFPTn6
SI84/e1m9K93dR1BB4LychzZZ81bsP2WFVfFt1cD3GhF90b9xZiOaUVyBw5iAjg+tigUfw139siZ
JRjQzLh7g3AVwS00ZTvH98VYcLiV6se+owWS79xnL/68zem0dk3rbvPZujtoPMZKkmbqUZoNRbPT
05jv8mPq4rW/0QwyUQf9TfLdhi576aVs2RxIzs9nnyEGTQRaNHS4Cv2otlW1CRl9yx4tA1qRRyXw
IvugUDuxhMi2C90HDf6ERGiL1wxBe+0u9LKageGxMS8pQXYbdypbVNDyT86UrlbXZ51e8wPKPy/Q
+7qMIOCKrZhHq8sOyNZOpsShRNItFbypmUecG6P5m4dE4di6Fq3okrcE/aw/q8D5U6oM75EMdt6v
dlJ02P64MdpMZHV07JEkVUbxFpzY9v8llmVH/1JyKFH1EsVwvkvU7vCtSRQSH/K7Vq6dZONamdvX
BpXUtbGmSbh0Q5zlqjrJWzcV9Rq/JKTtvUhsDxBSS2sF/9e17avhvuvZr8T7LGoeYOdTFQqPuiAw
YPQlBfYLgHIvOZcAWXx7q23vZZCJgGIry4mWFavugvylLXzVOYdAiXFPrw9lwvInOnxdzBqw0RdM
OU4m2G+X2hrL0aC0/YkyUtSOI+oxf0WOX/X03bdV8hgYQ/PnOT0ubH04bsZ9ZuGo2EKk/B/E7v99
kWIQtUJ5TLAuRYE/kVgiv37XKkWJ2mqNLMAmYPFp6XSeZENfKIG2cEAPwu+qwYFTGo8h/FhafPe6
ERgncUp0hhKnRvPT0C5Ky77H5ieikI4p0Xgaul/qSz8tVfgdR8lEs6kLIvWjooGcaoGKfJlNdIhb
Wuoj3ydHqIvTd23pwMnd8F6f4Zz2olDH70ZoREZjfj0JoCJ5jtvIXgkU3C5TDOYrLOsAZTpwy778
+tcWBEHm5zK0l9SYWhxldAPQuXb8NZwdy+ZPkdow60wSGJlvdRbeD6aaa/ffZ4tn7VthkXJSReHF
wbFNmrdiiNOpEp8LJWuevsNCc8na2ccdIYMK/EGtDSn6CwTIVF2rX2hiRBnlN6BOM3XXyy6IQkL1
f96BJYgRCExsYhzc3aoPcBYDTrvy3K9Bgjw+gx9wunLqvxXCcXPLTPdn4Eka663PQstIdHQac1L1
eWg5bZPeYMbQ0oLU956LRS3VeT4/GdNRy1S7T4A5w9qD8nCSOEKCm5vUEAAG8D7i9tqFzhaeoUKz
Q8I2G3woNUYXSdpi67IUhiHIkbfMkoz67UXtZGEDAtgM0ohbKBB3O0xepUCinu4jSRXmF12+8haO
JdtTxn4IuqG5q5BzAnL1My+IsynE3P5Y/yd6/OeCf3z4s8qQyif0DumUGuLnyD6jCAaifZ9maLyn
eswn4FlQlpVIekPBBJEkB/pRCctBwIJuWqvUzl8Ms/SW/592R5TCYUo653aFuGVT7IcBP+qeZs6G
k8p/wxAlqaFSvMVSoHafxbGVc6wNDzZGo8LcL92rWchjWRpcFHXc5T6O+lRStuq9av97ZbI4FOJn
E4Rc3sB5VISZUpoGGet6i2SgH28OzIlRJLxTPpkyM2b9yjAxstpimL0pqD/EJlrIpZe6cbHCjHQ9
hiJXYKT4/Z591bXHZAl/5wu/rqIOc0IhbyM4SDQ63/wSkBFGF4AGme4P9OtbhlSF3Pj+hIXtwPTq
CdonLjsQfFtLGsEjLr2vjKyvvi5/bb+IJnuyXviTJONbvFuQzmusAnz29++1drA9TcxNVaJdcJiT
U9SvJ/AxHpP0S7bdwb5a4SmZC8+jo07SPnGHgUyCU6Uz6CLJVmll4oQmxoEqRODW3T+6Ai9wm/4Q
38jSPXRMYkYh76VeKdUpk2k5wPGrGQ7o+8Gq4NNh4/EttZjg/Hdasr2vFPwYQQDKssYESWhgB7fq
828+iw5ZUB7NHtXz3W+S3WK1ZHSjv62ufarIDQaJJ1IPXptmckunoNZR6UZEGR/eU9psHfx51S5V
CqRE/n5wDP6wOEN1l4z3hzQV8jmVoG0CAk2ofZVefsDmi6gxdJ7L1AGE67waIgqUX9jqr3aLaH9J
vQmtcgKXE5GTPNCjSaPpszAToSEDeMKBidLyXQPWoU3DONkDbD5yM5VVW+VLHRVN/IDbvhW6A/j/
KMRHz2ZJ5GTdI+Kd9YRJQSZ5b8pknWksHaJmFOPgWNLNuMEZ8Tpzmvmtqt2U+9EtU/GL2tMNpXe6
2pV97ZkC5KGT793s4qJNPmEVVoLoO1HETXkvUnDyaxAe9OVah7TU2QS3ZPBWi40pPsIgmfRD4zW6
uY5Ae7JeacLCiSvkGazFpHc5abdDHPtA/YzSyR2Z5vJvgn/dpdgRCFPAisq1GIIJV0c4WKnEpdns
H8BlSXowQpf+P1KOkQARS+hyIV2PqHcsdVu4a2lrSfcmhzcpDm8FmdUOUlQNYICy3JBse4CyO7tE
KBNXnPeStoJBO+tyWWUMhfMYW2ycIyzJ0HUgvUqwNG4DuWNFCuvjFVSNdnv9sw9Sq5mXTTkOgtUC
egT9nbaOuZT21oFDHUqAG9G6Qu5VE8zXB4MRHsC6nZHvl8F2XOb8lPAHGPDkWhlZQX4eqSjtuXHz
Zk0Scs7OUVcgkLqAsy4/z5cEeHppgS44ZMour+B0GZWlDNDvJs2oup4vIZNabe/563o6ge7iynGg
xG3XawuULSzDQa/9fTX7MfEt6Tni9eR6SSiX5IoqLW/8JsOAWvySO87vxxQnbhntysG7S/9ZsUCv
6CSBTHS2Coc6tQmTzdTFww62XZLbJUNtgjBU36LqSXS/FVsO7WMI/i1U6ZlJ11B9JZAW7QXYa6ET
U/tLEKVNdp320EitDIaPxH4xh54KeSjmh4ziGQM9aMO4OtYNwi37rsUtYR5RNig44bJcjPpZpPat
y/wuzJRCNu80wCxng29Ru+obQeDy8wf8uZoyaXhGcMr6Q0Qff+2Cls/khzg9pYFYxFBTvaUOwmBC
6uF1ISmJoK6oDGMjUQ7Maw3P63v7qW0hYkVR13tZ2uUOMSwTrGdJa+bNMcc8pfLfFbqN08PuT+RP
Fn7JvFEdaSlPuHmgu/N+yS7JW23XXX2XG8h7fsW9dAc1ovQChoj0u726Gz4KuFqE/o677qTYWlEZ
2x9jIf8IW2kQ4fB8E5mW0ZDQyS2IC+p0dSTNTGTmlCDHaYrNK19X6by92WRRmKJhtxJKU1lZnRoQ
Zd/ggi/vadqpAoHHOFZwonKRig1GxksLo5TvGsCX4lX+kMjk1E8OhIlm1cu43feWmKYqDsxIBowt
cbSAaT2ioUwgSUG79DKQVuHXgaBPRbyH0cvPvooyJRxaoHeq5f/bqz5PadMeAFVMPxGlsbSsE22Z
zj8DMzonS3eL+Qk+sot241qEkm80KzHur2qGP2icB4OS9/o5AKk9VPj0bmAN9TGAG7tUMXtn221u
SEPlx6Qw5kHrY7kk0/AhcgvF0Myj+K3TM4JgTJiQC3V3uEdDvCHiZRgIshfDciGBqHpy1AolT1UB
2knrydxWZvpfy443WVYA1J8nZe25sYxnyY98yLfgBkr82gJu4R2cdcxIQ1d8GSHpEMIW0UyTozOm
ekGY1+we6GoezCHig9GyUqkAwaMuvwmCYaQwI/HEidubPfsAy/m4VM/PbR0j/BXk6mLs+hiX72Rs
sX8GfJPq/hQsNFw+6L+WNgjGurF2BVBBsC7TRNo+c4KfGjrJVaJn+2eDgmUCOY2ar+G6Xqlw8BFt
sVVC0o/AXRmXKa3p9WPffdudF3j8UkC8Tclt3edRXtR/HcIvdvBpVw/vpNaSoCVfZXGxVI5KBlJc
XIbWd7WXbBtSa77hoJTtZ6glbvAk9c8qg2OPUr19+q+ihX26gP7o+hUcNMolaXcD3j0t59kPVJIY
it2JlhXhXxbWcZrbrWbuGI/cft0j7f/9FN5XivpD9QWzizZU1EnakzbMdWobCu3x2Uj5aXNwtXT8
oKXbpptXAo1n7ql1VyLCezFN0wnzi8fF2zxqOkDHayVcOexs1LTchjtNXUfMs+4TCw1iKyuhWNip
8yuoNlJlUasHomkmZUFRekywawZM1Ogvy9EKZBiIHqci7E9dV9efifF0mVTeVVz9Kvyv1rlJce61
huQhToOJlHHxBOLabaxGWK6ILCTJy8qw+MZZG3Q82/KIXYzjXUEcxxRd4jNw6JH1cHobZTRxA9tA
QSbKfz/ByeAR9qf3aWzI0ePV7khBBJwJJ86g0w8yD0MOVYEJMxagsxNeft+tphrfRMYGto/UdK5K
UuZH2QZyaYUDS+wG5s9tn8xh6ezBlw6PecdN1uXaEW8ltZ6iCqKp5GWjPwRK7wDejoGb9P47HdFa
Nj7fiWAEo7rDDyj5ydnXVxFlRw3P/gTnxzgJpnB8xzxJ7jo+LhOsU9O/RoAfuz37eKSKPo+t4dF4
xRaU5U+PBU07hLaRa2OW97njSn/Nzrmv8uAZD5mN1eeR+gzpi/0bdhvhpuk9ANViDCVr6YwiQeQg
yp+p2n2JrZz7oYPA4r2PFc66cWcr29b19t2bBTGpuDySJ2Gadjg4NtIixzYDV/GLkZENIpUuRt3/
NeyJIU1YSxIB8HBaLR7gT4o1T4tpe1vAeDhpmbOsYBuBLJ39fEhFHoZW+pxj+aGBV9dCE5DFXCRS
U6smIz2PysnUGxZWqLsZAqM0dojoRWX7SFaEdfVeU03rNAVcDxDRdYXxEc926U3IwWX9CE8a4Jmk
lrlI9Av9OJ+EyJm2t3glbKW4LejkUds1zPDFjsIJXk2B+JOcekrjuDoHiQpwd3hf+48tAu6gHeRR
6FkJFdjgvu+z2owEgG+rPjj9csON1/oE1yhBt5QbGH/dgwIU4j5ZqDTzKzNwmgeFAV3BSm4ECMsy
szzn19hymII6ljL/zVkFzUVz5l4nYXNhWVP8nYyBKGZa6q8sQkpH/TwNwNu72s04H7oBjXvbBZfx
TwGtx17cZCprT3BFOg555U9clgTgv0rJgr0AK3yon9Mv3I3r+meSxGZbBBdv4HixgzSTqNMLOlVL
VDPHkKKLHqzqtoBKXNn4N5PyT7hhhV0pqeiWo7xcexEnLoyiGwszo0H7JfYo9LOwUKx+b3q41a79
TucJKKI3DNApnV87EhRTLB5TmatvaQRphHUIl+NHBOKQ0Yoe/Hxo8fH6K0wnQA3upzZTMMIbtn9N
fYqyVmQzpHLDHUptc9xp2T+LRqowQSAb1/4IAv2bEo31BAl/f9hFo4kwXE5atIuQqs85tnKabBNd
MMFk5pHNtDC7nXzKfIYtfuxSYxIa4nR4v4Y4Z7kF+rmImxVxXRUoo7O8fNAVmECXz+AdHT3dqi50
Yt/S1jReYd9JfElj9hKC+0WybqCzz4BO3YeUZyCe4gZFH7H57OUg9cYFXrqvEkZPzQ0oWWfCxvKk
LqKODLjZmFjKjhhOJN4si59qIw0DifOPVoNVE+7ckIje6/OW1l71+0EdPqzuxjeomKmZHcWfeNcr
yBc/yX3YcS1ArmxN7xJHBB00sB/eB0GoW2gjMuPijCsGMy01R5PPpFFxV5PZFKD4uOg0P5g6RHUC
zQWnVJY04RjRbaT5B0ObBvPccyVGyHw+8J0oUwy4MqFPfuf1+JfnrLj3UKM4OIv8GAsOgwn1mcGA
O2smy22YbTUnqbYpkstp7Wq58mqvVe+Gg5ZX+G6xv6YyBlRFekJggzkQ7mGWk5j8fLiDc+d1opwb
UCPmiy64XCSNstvYzZaeRnoX9g24rMVE8wbNJgrkAOHlPKTS9L6L016UmKg0k6x7aQGJaR8CXS1L
MQjbdy7Mlhnsw8h2vq81D1Stj/U72vi/p1Cdr/COT+i6TTWfGMUZbAaupbdF2Cbx3h+AmOPT51Y6
WHqQNGIdbbBOhX5rHZI2OiMb5aihR77KQlzr672oSA1ckY6tWkL9mGL9l/LKa7j5AQUteNbNADHC
ciOs09zNdPB1gtr8NDvTT+7/sxpRKFTIMmR2DZNpwffSq6Z75OJqiBZsOzzn4Hxe0gGry1kGgtrO
OQD+FGzfU7VGi65j7OmKFmMtYwe9ZZBrwHVesJClkr00lusgmP0xiFIrepvK+ygSETSVCU1JiWCa
6S2RPlqsctnwsWH5z1bhxN5/BA3H76z4N2ynlNJXL2usI++PZaiFQOu1CrBOGXlWnAxo1kttGL7l
ayePPVeVgUFBfFSSTZSgUn284C1illL2kiqcKcibXgfuLmTQPUvJcwpSbQxlbB7Gw+0aY1OQfDJs
HTbV4LZ/Hf0WBsYlJmOV9/mBWNQNk161WoyJVp/V5Q7VqrSdy8TPvA1qo1v4G9YYP2jUVsUfS0sj
sk0IIkW0GdVX4mJqHiyE/rspXzazUqbsPMw/k53B82SSgJf8FoU0lSw9S8svGlwbk2qioL7kxkUM
eN9KRRbBjl5zAG++Cw1tEUIy+uiVfIYVYyal/7sBLuNigdq9f9nIrn7Wim5yzPIsRLngbpUkxLU7
GA2J/m4GG2niIRuKdLPfwbW+qCszZQGKHNXMTRzk7wNmsY7UkA9ErHdFqOj3FcUw/ebQ0yNVPbva
SEdYou9GGRyzsuprq5FTlT5Jj5hwf+H7YQB8U7MOSeO8Q2Y/oR3+KqDaMZWYmye5PyYOhv+RCylD
IOwaNrzXRiPcQsosXwWNkhNQ9PGmGyCWNSZrL+rl7V+DKxMBp3nNFbWeOkVBoWnwMXJEIaQDxKdF
Pynd3uh8uQGas44XVARqgoJWc9EYcfxpuxvS1Rs6Nta0I83+0hGDahceezVDD5150Xwax8BNXtbQ
vix27ZUmhROKk9S5W1NzMZc0AFmbhPTkHmd5m9wYXSk+Zoh2bgXun8OgihYIKaLSP/LPafLm5mmh
qsgbNYnEflC1X+xw0QLA7X7nQrEnmWci1poqBViQLCBOrSTkzv9yQWC2PrNdgjGzzKPBotoioEw/
u5CmE064eORvy2kyhiP1YOLtlIUCD7ahX9Z15RsxaiRkIMfX5gZ7mkrRZidlujGb4cu2+wGFHv8a
DyN5jb2qHn67Orb4mqKx038smiCUxF1tHLavZUL2xPRnWYIW8NBTT5q0R3RZD1+xYy+0liKmUu/3
1RIC6njz/23zA6/3ZJz2HNsnGcWNyVlTZZk//OMwUdjbn8lvUVrwxXhmHYu1ePAztdg3PDbOKfsn
KolzDG+9Q+VflkuIOB0GlCm6IPr0Dc27JFQpzkeDJk9sGOFEeMSeetpgK4RIhdyO+vZIA5COhXe+
6s8x2uPAl5CUzDA1SDxScwT2g41J1LgAa6F9jmUENeTdpj/GuroPt0RD7MD1rH1cC7viSXLOykIe
xDJ9YYzFE3D5LSOFXFJ7IpwrEQdKnvx4YJq/QjuyjbuB15Yv3KiirppCuI9WzZVhffph1DHix3XJ
XBrzwSavxnuEI1+VUhvD2SzkEW5VCc3XDaTbbcSr7KSL3lUECyhVPFSwzQYhYmLWnHtWUnF1N+2J
byc1sL4dyc1lOb3Zm5yR4VxOuIOdPzf/+7RLkgWDdZfppQl9zePPsVKIXuiowlyFMuCsgR+fikYl
6NAJhJk65lWjwQL93rfeA9BxQM2uSxWXp52F2Pbb00ImRkJFJmLoRHd08VowbIWwG8iPJtz3+rH1
q0YbLWYyW3SSgHpNUDopC4SddsRQ1IkAU+UGGFiWEYAnyo8nmd34f6JguJ6j9zUkRt4dDvC5KVZ5
ZLVKLzn/chZR6G4bvd6rQIaSfptVtyeFsRJTtzUz5q36cIidHPBmF49n5dUN0Kouqd9OrcviG1M9
eQz5ID3h8HeIe57omuFUyLIYf9DAFF8vMPHJkEe6KOZ2apv9uZjNKiG+gP8c803unD3yKmQCPgiA
v2I7iVn4wGLGinrin77ZpmdBQ2ONWXEUS5r2PIx/3Z+Xq4JxyLEbkdRpK8THpvqx22WR3raynpUn
MGdjWvqQuPfOzRTccvRVkHaGqY2SuriP8j1fGqAoLYKExnixQJjz4+MYz8XcAGuwa/NOaxHuXIKW
yMTHUAyRCEvR1i9/9v0wnVQzF2iI9DZHrcRjNhqpgym1hbSO/XTD5bfgkTB5UY36S5BoGuwwyiBt
IP1h7kxw0/1dRLc1uWxD9cQKwoP1gBAp4/pqhyRi6LDfmJAt4vfETsFi4U7glwNP+aT8v3r/eu0l
R96aqjz1TBT+oi2Feb80rbckXnnFql6Kjfil/vbQYoc1KTJNS0hM1QENPunUp7Daez2bbuOKHLTE
O0l/KmRbaLC6tQJKH2i3YaoP5kYt34cVDZMjt0sv6wTx8NKmslizeTHgR9scMyIIbOt+HqIEVZFM
PygFafwRf9AML190DtlKKIranXnl9NTKTwiYcfFh7m34iPMUYLIQpCM+8KLKXAXga07/RGwEBkkm
uBQ9zWC+nUAsNn5UOjq4rYhuSpfxwRoULC+EWrza1SSvcWm3Fo6mgXZAGnrwEGmZ90Tv6KXHurGB
DrkmkHace7h8wn8h5m/c3KuBr3K6sgSW161qIzgWS9xm2Qt0K37yPUd8PUAp+m4i3zurQ/WCO8U/
e78gOy+AD+G0GgP3NksbfpCs6vMl9Oj6/h2S43uNtD/KejbHtExnEAZ2urwOcj2lY1gAb/IRgqB8
H+k4IbpJzLq8W6CqBd88P/Vo/9C3wDE8M56tpsqpFo5VuJwrQhBYUPt/AG1LNM37cNM0Xlks3jhq
dsF6k8VYz8OKPoOsphrBbMi+7l6WYu/UIZzBg3yaTUd89/Dq0B2Nc5gm6ewojDgzoJT1WBEm3gyN
W33TV1Gxm+VfAPvadrIv1N/8g1QlN2/JgX1JC9jaBlppLWUrUo1Om767LZei45qTvHSMVbdnXrwr
wZJX45TcUIfi4CmFL8cB2E3xCSoO2HDhhG/2wCM8JI+frfLra9CVBWct2E0YRxCLOkn3FODTcuRS
MKHLEeuQtJ7kbTeDzYdyaOb2Jzc56DkAX+eL4jqdraQ5qlG/A1ONp0glkfI4zLl1V0Pdd5vJYW3M
NJ6awdjUcLuul1gipt44SmZTbDlAVx8Edq8VfVomuNDnxdE6ljRylPV4+NDljxCUUEjEB7hnr8Sm
bN+qKhGWISV0RqdBMk/TSmyqcoXODJ1uoRpXX9SlY8H36XI7UNh8wqvU7TY7sqqZC5xv1B07MPEA
Kep3FcrSWQTZeeES8ndNhhmHmB+v0uoJHMGY1MSwmFU1sp1ZAO8x9AmOpA2SYHhvFdUzjTXRvCEc
xLVwxtoSG7Q+MNMU5X3Z/LQj5EgVAJ89xV+KyMkO1lI9o8p7NkgQvz+IuBNc9bb3Hfu7vcsFR77n
/a+UuN74VkN7YCdhjT1XJWtdOY+lsFbvdAbVAqdJe4kLMfRV+gquREbyhqDr1/Zh5leD81ctoHFV
fQXmT7AH+oM6xZMZ2aBPg2mJ+VH6oiUKqgdt483g7inHxjFqbn/VwJHFpeUXGeUpuA+1XXzayvOl
WN1B/gzSnIDgJ5RC6gpeupFtOL7kiy+wLMVXRTBHksojfvDnRwT9moRzPGzCBotS5IRaWMjvnhTJ
wEyPYaZUfxbE1YyKvtuRknR7W9MsX53qlEJybRbTuoQGTqenAW+OJlM/stNwZsJTxaoV/G52HBy2
C+/UyJRLBtEEL2z0fSOY8gLSQxgh2UTQLVa4iEPnrJuFpDpYfe2WMwxfshz7jgV2iM/+Nwk/ua5B
QiD/KVBuZj1rRKhUAasoFgWhUgbpuxfhfMGc887CCJT4N/w5Ib/C+txa1ww+9EdHK/YUf0CCzvV9
Gge7432grZwYULyPbHJ8y/KAQKQklrY8BjxzgFI3mMXsrc+gRqsSO1TIBEpXU1dBvINrhoZEtt8a
KTmh+1ML+NOQDLivTARDzGjA6xbiIlOSV8mC8p1cjZUCYkYS1+826CSa+HFdW5vobanfXN/EwVPn
S7+HtBnjNlNM1JGFIcDBfAd9MSpcjHxByRKifASFWdBmlo10fGEgkoX+khE4zYTyWhPFfWaCZhew
RvBpAh2F1PsiaXms9Al2nDEwYeIL+f5x8/iRt/1ofQPEaaC1Sx7DvoFwNgYWAAtn548TVqUHfl3v
hpMNoeA6FZuhosiNgCVTi255Pioe7oLpwSs6lSPOvJGbEguZZXRRcs87b5cV21jjnOL/Yp+nfT7w
7eUiC0OPdcaP4kubIjYdCb8kByrWaiJb/9ubDvXoTY/JztnhUU4dnHdwkLbV/KwkkiajdtXKqDPR
kjImY+N+7OE8lZeYsfchs6DWVyuEDKI0GAjDDR5sRdPWyu+wMrCW84TgI7/OGhuBY7qZ6/23DKuF
+pgHyjjeGWkUl9m23ZOITOFaCoGYm1FZln+UakRY0zMdJ1+LPQ4fajetwTdT8I/CADZyl163/mTs
uOITtdQcKWNMUE/qhVghuKyvcjjxk2+eGRipoVXwRmqtZfRgPNU+YLwoWxQwdco/4R8jrzEYE5NW
yyC+f5SZbAcepvzsxJAkm+kZYgAHx3F267U/h2uKsirdnO7JIwahzdyF0OvNn9c58+xvhmgJos1i
1jmkPWxMjBYCnMb5Dkm3GqGgGsLZhEdWi8/bP3Q5VwXJrRTJwzAmg99LW6wd5IyciiXnuwewxIrh
Npt81x2jqZexRb0jMVBvvNB0x4sPrNieQYEHbYBBS0xqQs4LG5gGobPUSD6SSsCQ5ofGbkxze0Ue
V0/ALVzE11OSBdSMqQtsEzr8qQBbHRluEtbGG5RE4Y/H5rzTOloyPP3INBKJHmFFBuX4W3OMIE9M
OcFkCmWtm52mK/h44vIaHNinLG4Eas6W0MaaxV8ShUMxu4+I4as4UvbXs8qOl/KFHdD+Nc9tbkbD
Vp9jU05CuVCakiZUZYSxNf5EYOH0V5CP5f6PhN3686P8UmeoBJKDvpN+uZijDC7xavJ9hBx1Ud07
TgtiFf8ZRRvDlfBVn6pAuyLXEEBCQwjS3gQ6W+YSRPiyEKbusW1neMtpOwkweFRZmPP3audyOnMH
j7ILLwN35n3EEC0/Fs7I5y6gDN46hBLNCVBpCQzzg+jzAA7MwoUdXdqYwvrnyo79hU+pHGgUkYFZ
S76v6KUgqbtBWiU9pOmHWYUSPnXYaHYY0eURZNm27axTdo9vQzJ5r9A1sryRW6PJ/HkGwGAIsqet
PdG9xGKu0kbx0wL/RbV9btbmrwdcrl2xusmit73nqRVOZ56M5fp9vkX/WVSvX5oWenwzGHkgMX+j
cXrjkaVoBCKAFmA+oeKOZwbGSpMJaDxxsIn3/6Ra+VHwAhZ/ZY5cjuLwVzki1MP7Sp32xVNqzI6q
RzRpgJRGn1Niq1PXMh6z4K/iFeotDzFJ325s61dUjXu+BeWChYRlwgzc6RdVjouKBMYY1Z7Ut/VA
545nw6m24H5FNy7ZbBtctnSzvASnrRNhuATQhRsor/pfYkZzlwsCvqBWvAG+DqbDdP3PzjXwG2YF
qAA+L3IrHearOskrNwA5fEYKSYxTPPML1AICbeAet9PaJRvwnO+w9WNeqlQcFMdII/kXgJ6hNAsp
TvsiGXX/WeBGtLrreR055RdAWpAr49r1xSLrH/xzwT9vQ69SFbsv8dq92NoEDJBdXq4Mb1P+DUzi
TQmLjrOcNsAr9STcEXs0x15Vd4a/zjpQXypTQcUlLowyYFMFKOKstxsFhAkROkhqXEmWlNoPm6BY
Hn2Zrrwf/V+HC65kqsJvyZ+bEJU358ft9TMMBGW+3iSRtrGIbUQWKbTcbhM0CNa+920fDPQMB5sY
C9dUL3cq6fHP8zaIYyVMMF/95TxUPGMx2FAOZL7BMCH2Xvxw027Ntl3Fmz99oHCgwwagUW38M2pB
G4rZwl51QcbNFeUTtixEIqcHWKfw7R3Q9lGbBjPL0AxzC16buPRdPYW4tw0DBC8YnPXRRLN721HD
AYiwkpfhU/gOfA4zmIOU3Xw3bDBiUXazbeTZQdTPhTPclnl4wifzQQR6gSDm2pZ1VzMU1Pa6LA1Q
jy8r9AY/Ld0M9+TZTXfPxDqFDfJ50VAj3m+B0nlBOKtZs4kIIDTfUf2DkLcCx3NkzFYT238iJQLL
FktV0dg/EdXGY/utU69KLQTIyQ2Al4cJD1LtQQ7kDZJ8PCH5//JzQnjlpNIglzY4A2At45MyicU5
gVzR0o5upsJLB24Is7t9Jd+IpD9qzVFqaJYBnY25BJSDE8kUILf5f0eIfcsuo6UdUSX/gD1YXdmu
KLPJgK2+AJfgk3dUyGZwFL02VgcEAa6FSI7AHR3TVPzovuA3XJtk9WoOHgN1EShgR5PXFyiTCRe6
OdE6ueYvUdTYGDokCIcBJsIFgQr+5j+3RCeYHf87nsc5uTPlrTwaBnMSTtSdxonSetgF7415GQME
FJvX86kHHZ4Rp9KUAMrSmA2gdD2jEc2MREpbJtDeRTeOHrXx/bm9SQ4ZLk/4qXNm1wi1chabHo2J
O8WeEHq3H53yq7T5T9XPf0ZIBbZ3Pjy8hZAABsNVmPHbuHe2/1jbI1FSbEBhO34IiPrhgE07LgoE
jjDF2jCUTF0ziFZlGOjGiKixGG99pcPlUZ5EZw/U5cR1kirlFtyq1JGJ0VvEsZZOhAzsxbJ6P4/e
uhfSbb2gcI2Oed2NYXzj2BcuNqZat4ZD5fNyQzDdc9cEax8r2AgVNuO8wLl3UAGJGwjzUAJ/aawD
MiVAkYafXZBI9Eawwl9VGAxgQ2oxsmiLgEWaGnb+R805XMVTFxDbQdC24V4JZSGw+tdHXUwiKR+J
ALaMx1PsyXx7nGNLxoaYvEo+S9fBXehv0/qyoiJhPOlN0LRkoC/qM5DUsKvOxwLbCeD/ykBJGwDQ
tfBe14AQQjFrDlGG3LlUBBEyajVdvS0Kh19xK/JSOdG2Lsf4lcPo1jotJgiaCsNJ49IFf8wK1XoB
OCbyP8pG6uKNwUYk2jadyQolBlnqtLewEu3X0VjPZfmSbyP2zUozEMnx21pU3ahHcW/H2V0p/xUg
gXVouTqOJBqV4QmKVqdpais8exsErR4qoN3XhAfoJC3znQ01cNKQZ8qQJbTpLgVIKh14UyLoczDT
LFtWinPqgBNfP+3V5DvWX0bOngAzb49ayCBrUayz/T7ghbwJSjVDAWA7YHccZPML2FWSQusH5KrM
GJglUZJH7vx0L4/gQUVZMSckx+e7VfD63LWB+l3kaSlrAFzs4oLLPa3X5jaDjd9rPBC8jCPTfpsF
70Ri86iRPpUzPmuUTCeVyDWkBH4QG+DHTruxFOyNR504pc+uEvy2TrakSwJU5kAYHPCxd/HZr6f/
n2SM3TBjvomhJZy8HsmNure+lmueFvzeEdQmaVqCqZ8dWjXXQ6cZaMujweL0Tmztxdl6hD5eeX2v
cLDNMGEn0w/RhhPf40Q7GJJz2Hdv6kd15/bCetGMJsOGqUkAkBQdMvw4WFB3tzGYGOQ9LNZ9gupx
wI1VBxXdnGf3xntO4jidS2TyBtXJvYqAud/0n3SW9knvF0/M89EfU57+tMcM/aAfDYgK3CwNzikj
+7eq0JM63lQOFEmZDoUDvKGyIuDUnrcWaW+jY/r3Jz6txk+aVtAlRuS5KOUdlgq9nomDgliugWwi
Zrh+K8tpUMnfFC77H/cRJKJ3PIc4dgAaf7vW88VqzThsVFR13NC3GUAI68jGBejRMIznc08GO0YR
bkomFJLPUONkjpMcCCCInN9wXUzmhyqq2MvOk/VTfmvoZpMM4d7Wd1OMw7VJjqICx7F0ivrlSZQh
dTxRFSfvwdEL6AHEZOHXEBYbOuoCYr7pi+UQFUZiw0cTaXrg23OzvCXt2EDfy7krjXUT8d9km4MU
opyNDNk1pii6/ZqMtHqXkVAjDlmaJf9555DOpiaSN/HjSPUypfUbSRz4SYyK7OcXOjmqH7Uz4VHJ
6J0Lu66UoJIOH/8VTnU/Cuao9WBuDBKj0vUjc2rEggKGn+qo3P06bbhAFffvJIEiJGWm9T6bplOx
8B0DC9ZuoQsKGLiMcE7crRp4g3JJFi4Ayu//3330/cg6vsB7f6pNa+Is7f9fWsVDSlDFSDWnyOY1
YTmQ5cBpZNIrwYlWVPn81SXy5rW4vT0voC+mbQH6T3OSqFKqugZZlHrKMUdNtS3CgSDhx7zpvqTP
BiWzEg5su3BvCeyGaTnsnBrV1KlxNoTakYm7/9z1dZUKxz038i8Iit5bghvnlCM3KlZjDGzLW0Vv
C6ssmEVa+UXBv26zq7F7D0sqD/XhkfJmRr5HaAh8LfUcbaoHo30DAVIkkTq22/JUeaW4wkxOaNjL
XMkSjC1wqg0zukLl6TC6mSvkLf/tmKG+5rLkOKuRO3hPTxnaqElDbQKGXH4uzF+fkiVyCd04b0p6
8cuj0bD0FDwvusfFfWkC0zr/BeJvy83zut4Zp2KOVPcgKIe6nokFIbrr2VFQPSMADom8t9XX0EDn
CFGSeJZW3Cv2pMiK3lfIHcuLCGkw7WghW+ASxQ0W0uzhkiabQBQhzO4CE9EJ6U9dC8StALASeHlR
G1GDd8sbkpNZxpyi1CNdrDvyPJqwpCiQgdYSd4hPE06oO+lEl22O0EaIqo6AG/rJBKhr+ngR5oyJ
VP4vMgTC0xv9oP51cRAv+T8jTGHpJhbVSR98kDtQZmVP89LIFyKpurEn8qBTVBv87E+5DlSt/aC3
Ds2Xj0xi3Uj0QResptNPsWLoeu4iHa7Nn6UUPhd1bTO46ppVP9s5HosI9VK6C3vn9mFCDhbmwS0G
3ds8nIPDnLhAnNZ91lrWA1NnetphCBBejPFl8YVuxPz+unYfKt8GyWLJb+eYfKtupC/su5EbV2Jy
ZufZ5Dy7r9cMm+Oo0jwBfPaoIyBfZkmr7PY9QXqoTIaMeai9BYXkjtmPA9ygomgMQ1ssvNcu3/AY
hh3P5sPgfV0/UqUXnoxIrEZuAJl4YQPd8G4YNwVCQl46Ll4eRkpc/QDA7gzHdqGKlRJGw4H0Zl2p
Jcnop7jcdju8uGIl1Pd4hNJRbeVTA4PAnyrMnAkuaadaTdz9guym6UuYP8I34kW66Vgg5ATVM6Lu
W/Bx38GARbL85YFoVhwmwRXb4aBnxw8+cWiTG9sJzgLU89mtK76A5t1P0qOBkKBeNyuU8udXGipR
Nr5sBcVn3woodnkEVtrQRN2pWRbg5vLyX7iiSHV1FrGDbAehNpB+gPTY6hYOH5y02R6lV1BTEA9v
VgWou8w0AZ2ZWEuN13V8nyg8bdvHs9VpQQeTvMH9BHCHW4HIwaIKZeoJ23k6s1yoecCofQbNlD7r
/eWcDr/bMwubx5yJhvWPRoe0QrmBtDgdRHn1u+tyvN5VB+M+rnH7JnnvDRa5XtlkrS9+2HbwCXXC
LJptFEoumjqsxTm/iRE02pttrLO1GFtzCHHOwkFLOFkVwOwhXnU+5oIGCKpka+DqmrQDecd1DZEr
A2PEQ5r2P46FOXVh1us9GaoLt0JUhN4HpziNubfe5Hg51M3Rl2To7efmgXB2DPuroeVcCcsNhSiU
RGRvArGDYFeQTe0x3y6Ve8ZhDNudp0gBtcmu1xJ476vBVlcPpuckcp7QRJIBAC/Aw/C1jryH46C2
XlkdKV0joos7xgnrzB8AkultE2Qk6V0QO86S7k/2oIGWuQ9+j06rNme5thYvRSHjnLDnYGzxxiCh
F8K68iz5+Raob4EeAaKJdLmM8+KbOoLwUyukYrrG6RiUtfFLruheOrDoYs3wpRntDZ6ztvF/VGyt
5KWteo6HwbfSKAyDwYWXUhUhGFMEU8pV5YLSlFhfmX4wKFeWGHmmNlXN/2gw80wZC/g/HWFKFMX0
llHmqjtLOPb3chvdY61AlYonPqRG5mJLfDRXkBEtakg5vVPEcSeVZpX10zQfZIP+XAJYMLIwrfL9
6nJpUfj9VHhvr78LGQ64ijCW4dQgbnF5sa1yA50s9OQqv5gKmJi1R9ijsy3exqvcIPPai5izasN0
pCm5xaf2kPUtr0JJgFOu4CW8TOzXyQyE59dNXUyrDM0dt2/nZvtK68kppW1l6PmJH7JKD+jggtgJ
RPgjFrEDMgFPEwbbrGLep+GLP0cndYlXScnPAc0CK9roLrTyvXT9uXD5Zv+cIV2Xc8n/Xna99LfY
qq5xWfAqyrbYkUYv6TO8FkeItxgMKDDa52E+PM/F52fJwsSMX/rAcdwmNkzkairDdrCgX83jYGCl
3WNk4wZcVLMWAxX5T7XSHOFsjtxZOdTphyB7C1eazWgL+0eq070vXkFHmGLY4uK6B9hspwJkwaw4
uV25pPN5+8WHQ4rlsdi05BDvOu4wSjbECalrs0gXzjwk06FXkOZtRkGloxO8UJwOFGhc8cGHFvTO
4q+nvTmwpBGaMt6eO48kA+HZMQQ2XGFlSeKXxutUShdKzshm5RDyMnI4XPc4BaSylx3cipn1Aw0S
uZwtnAc1T5gv0U9EZhR6hMPMSn3px/AfeaPdpTMQZ5qMLmknWTbtm3ZTQ+MnkbgsNT3CkGTilFhA
QHP3IjfJBbVkY1xYvAA48cuAMYk/dScNk/EA/awhIrF0ICh5yIvKPW8SwIZbtmCaSvA37fjsLMar
a56vmvhL+/PKsrEeZ58trdF8eL0+Po6KMcfay1fcNpbrVkzm/OWyS0hgIgbck8LUbbxO3C1+QeVp
5+LnzbZZD5iNlybla1xfyIc/zhhDiFa+mALUWVqtv2rZ3Xf/OEwebBrYn8e/yauU0jSCL0FJp1tH
SkYWxieiIwGknIG4+KidPJ6JV2Thxqi2vQS9sepH9vLqECniLzlT1zaJdOrzpcdMmYcoPFJapVHM
/rgSTxyTfdP5DPfJ4WGP/tGL5aaupTjY9sTEDSo9Jl/Xslb0qIOeaZVkCXMthXjPDCESLrEIWXL6
/7V217vJwZiV3C9KxOEPwU24iajf0qHNgQs+cZFwdLA6dleuR1UjFEsDbiHUY3wzbJY9XqRxoB8S
3RcHCz9M8nyXUb0vvM6jlOt1mHQMMst+Iv1FT5O3KsN+ZmNq7CxspoYfsz4FvPV/U5Gz8zsOutce
apN0+Wj5jGGaTmQWg6VrVtA741MXOBpinvqUm/rUo+2VlD+5A6LxZcjOw+a6F+WwGNYumG5q11BP
pNPobZibtd2HM3AFZ4QyrjHGSGnXPJQwRcudtHxs5G90hCQUlUQkL4anUCGvlX8Ru6e70cnyfVJN
0X9pIx7JFKtMWzO1GA94Y82fPG1E+itmtHCZrMgIqN/4ncex2X6f+puAvSpQNx2/zjMLoNJAZNlN
Rk+C/t/aAMlOYQ5xfKkXrFT9gKnnVKApiRKuKuUhNWw/+Vw0egCL+j6ULNm6Eq8Lo/HTSbE2BHOt
Okd1yfbenO1b3kvPI6RowCyZ/THakTs8C3oe7OEiTIiiBt5HISvi8/PgdCqogYVdntG7OznvgQmT
tMuif8Q1jZj6oCk6aa17BNVm+p+sAMQU/jBhsSGwA9EwqR0mVbkEwy/zsBMekEdMXCLhTDrOysdh
B4gBtnqqlH3TthAXojNvwZw1XYjw51oHuPJpVoA5znBFBfG7fZdvlQITzswKyp/sahj62BIofY1J
Gm9GTPkwGJaN0KKAnVJsHuDGYxypmhdQSswQSJXlBzE7b9tJlR7o44W5lcSxQv8RmD9tS7C64Ie2
TuJtOzL9WHy5+AbfRFm6e0d0WkpuA2Z6EKCaKx/qBlXkAjtr4kgDbX8EsK7OUtY5dz+WTVn+SHRc
LFPBz3QuOsPIboqznJtHE4eV/rlM1yTJ+4rtX7f+EgSeLRZ2mnrlcmT7rAoVlMGR60nVWytkGP8x
3NnqX+H3nMs5dxMGtyXy08CKhY6QtGNgRsGoQWeK9AUGXsIWQ1ypHsNCJH7JfjqB6ZWfUii2VPGv
xVSrM4hZMeqZ10acYxG4ECUBQCcBfhd2BsB7ygYCOe8d9k4mmuJAUN3a9yWxQe8Fy9zDcKuU97sW
lCPF2yfcnhi9FZHl3SxyCLhOpl+HqmffITmVZATK1A3CwT48Ly6B44hP36IkZ1BV/+2uQYLqn8U6
XYkQzzkIoTDC57R7QXKxstKITsmM3FO049H3pzAz9DbgX7e2os9xT89R/O7p+yNeYuJvHxS1mCqC
MEV7BcoyaWlAVd4+X7PGFaWcxF4Ne79mEubysQDUh1QLf494bFyWATwuYyNTLWhVeXAMqq4qSfA5
nJPDM2qho2+lmf+Nyz4ce4UrChEcYUQI37fNtlNaSgsZyAvbuUeOJCYT2WCFaVF8fxRLCZNHvsi0
M1mkPsJ6aD2NAUvQqFMZzL/WauQKdhXymEOGYYkKan8Ls0iauf7Tvu37Uc82MSVOp8csZfYCpTNc
5aU1Gg/mW4ZAPkz8+jPpzeTQpoGU/MY8Pa2ce49l7Gbf0x+wkwbJzFtd6O+xwRH0s7GzXq0Kb+Ee
wWr4uU+diSHp9CzTXmfTEOAY9U/HtZd1GrKxfSC5gHA1xYWSyUTu0HQ6fMdtITRuybMrMeHrb7Xx
KMo6GqznLJx0MfLrW8n1G32mv+NktVzy/UrzcXgSsv3LfoSedlPWoCyQYwXp7ikmaEV0FwfL6Yi+
2izUpyVLCIr9+JuBnMKtSiclcskV7htGE8rB234EWFHLo9RrsUiwoaSBlcAKAYTSbAHxkCjZICtl
yemZGfzLFUkEq6zhTt6Yz9qcMP3/eRTZ1Bc5aORGUafTOTRmn2xD5hDZZfVq17xYlmnqhY95xKlU
6roLiQJR9KAfrsqzVGUJfmtm5EiyOq4QnlsbOd/BGocEgTyIOu/rbAgbKFjUGKP9y5lo6r9RTINK
QF6bRoEskyDCjREJ90vI7XkSxml3UHLRxIIvc+mky4jH2CVcavS8zPhIvz+ubHKr2N94hxOGJHCT
0O0DL+DzUEO/R9CwdAPnL5P2r9f9+raL+2KadPy8YbHwwbQe+Z9uC4eJrXBoeu9XlBIR76ZFu1jG
bZGd9SmaqUuNuI+7xMFO7JuB19h7QYwdElA2+u3FhUTvhvVGte0kfSt+4vTSpR5LU+WtE9TZu0Ci
CvTja6GkhUQMqn4A2AR4H8UBGMO/d3LCZPt3JmTPk2FSwgM9//94Vz8XzGJrpIWao+e7nGGrsP9x
y1qcBXEOoHQgOIV4TAiug0qkYKEj81330oOP1faMiz0M1GtHvhcD0KIBopM10IRjesEc30u6SoZr
wWT/EfKLCGBGq8TfkxUFhNrHUYEe4PB30qhfnevADtQk0iKVRBWHS6aGtcnr47B3cqP/dkCqEEbn
lM94y/u5rWL7e9LdC8cTVeDtIacUxwG/y2NbweMFPanzujdWIE/XBtE71LkKpX//M6j2YYBEsVC4
yURgxbtzzWpXUB7g9i1fdaVsIHR2TcEZSO0ib3m1l4g5/dhQqe8JVj2aqvvAh5PFQ9K3BYgoYQpE
zP2rcgULjzZ2TaZxXkOIkiqxRM9XOn7FpBkh/L4zkiF2o3CGIyWSqr/PH+VRtu/8crMhJhxasHyV
uMlOS2uwRdXm8pWhKJPGR7/2EVNqWikWuMHyRuJWNXyrnhanRvUG03086C7mrPlxp52CbY8II09p
V9arofUIBBSbUUsLXL8yIQfXCgUxYm06a+m9bLVNYBnU3Hvk6o98pfkykSc/bsMmHd0jpZTN++lc
jhn6kMXpFHgoAQf761fYMlH5ivGDrjbsyjElyLn2e8LMbgSCXG4uM0zCgMjEV/EnM76jqe5P27mJ
9i8rYENxBrizmkRo4NaQBdtgjmfSLI3p1ic0Yju52GZ0VVDMi9N5BKfjY5kOGFdazT7Bt7Wqy1n/
s8dQKxdQ2dkjInDYtomsQzlY7NLQlLe8YGbnZlJjYo6+9BpQ2WlnQC+nZT80miICVl+FUMYhE8GM
8p57NoO+6204ce8dKVU6drhMV5HHqtsa/dtsEFx8u+3g7djnv5h3NGM70RYCWRK2EjqpxRjOTxSK
BCa17sYhCpI8oOM/hR5t+YUWFb4S9Yih/s5Om59R7hm6gvrEQknzrSVSP5dBrwUoS1ou/Mc3iqve
V1yVKK+mWaDaqX4jJQpAkBWa8cR7cgmTVzg7jChRc6Nmr734rTaCF51TUh0jDK6D83cYPkWOI/e8
b+dfTTSK/Zu6m1osgTRLQohFDzaBwbiN5medh1Z+1aGxDv1MA6RGrDvAkJKHM2nmI3eDf9uWcvUf
aYcAdmxEfNsJnUy+jB4D/inxQZ/IxtL+P4C5F8G198ZJd/YhW38JyDEkwww+CACoICtl0T4Gih1H
MhcX8GpwmPJ3ypPeJxdMzDztGcTvwC8qkrwvzZGKLbp90l970PMrRvftImhNA8AKrSrRdg3X0jPk
Gljh0OyZizE+CDC4xbBYd90wSkfjIXeDRMvGzX59pPKGkW9+0VXeibqPHmdRyg4v5Vthk0bFoSyM
S3fhc25IQY0sjijYbJ4pHuQ3RW7RbHxVn+ALkd/qBPRRT9XsW0XEB+atPSiii5YcbfwZtn9K0V61
BlGQggf/E1NRgFn5+RCC7H/YZ7mRu3ApaGK0I7PwwDaqHCQWdyJQXg+YazW2+192SCOtKv5uRHlc
MMtMpbF/68ABNukg7zOk4Fr72EA6kYxQmd87MfnmoBioGUEJrAoK3MtWmQy4P3ruNdsQ6A3ORvXm
g0gr4YDoWPUERols6RcKnGCQXUkMj5Khalv86FyN0N+6H/6ehGXpxNDPJYSYPh8owyFJ+dgW1Z55
e608btkZUAS6pjaUN7iWH2UgpR7R3YXr7ZZcbwtf66SpxK4CDR5NBV3zBgYFHQU+L5Wm4FbHBFZH
sunLRR7Djsu/rM3sOLdrpptE7m0jzW0BYlcZb1DDwVoFMUkfdv5HsPEgY/lO/UEeFtbDddlF9F1V
9d2nkiBc77LGINwJXeGhr7DiCvKmhljtIiRzO+odSRT0cx82D3BkYDdAIRexxa585utUcOd38D7u
NeXLRFiqcPbOxlPIAZldcNoczfqHm3t1g4SPS9lP+u9YhFeQ3X+uoFKNlmq3+6VgLvd8/hOAyNLS
EkQu2tVcDzg+rIAhgB8uiBEPGLizRIi9GexcUQ/1cgiSgbZjIsDj3SYOgeuOScbzLAdYfMddhBTp
YxlmcWwQ0m0HwDX69HfdtlHFSCpq+iLMfH/ozD6AHwo/QI2eY4PVPLsgWC7Lurd0YpB7YQfmb8Ym
lOkLmdivt3rMn3+aOsZG/lUXOxB15oDEgTgtmNGqe/SlSWae6/vbTYqz+Cy0jSqB7YfLTYX8fO/l
ks3cgR6vd6PIvM8pR8yypB0moCl/SyDrnbTKFTRHbrSSNWT/1txS7LtZOQCCejBPtRbcZOLjq+DW
ntMw2sGlh4Ahcawx8M7eMMgicZbOZimFbmhtTVi3F5zpo+f9Z3lxBckaSpc/zgCnEqt+dH7dOlcQ
kpHW8okFYhgWVX1LqUKc8rrmMpKoOlKAtAruwfFYYtmKOjF00ILetHkWmXyTCJRSnGaLhl6rjMwM
Y2COpzLvw3g4fWoDOrc4p2mQ0WBD0aPeVYzYkBzBqWxKe8RG5UeHEekZt0+rmqymgHwgtki1AInr
3mCJB055QAFyrCcDvuB2mPdt+UDfZbEnJYoTQ8Kx9S5OQGhSzceaQ2QH6H+d0ylwhY5xPdtR4/XZ
ZQUizC2Q56UNOqPzu8FBT1NcYAlPiyda8gCM0mBTDPbbd/6bNaHYwEvTobCviDGDhxTDyhX45a2+
wTGn8j2QVI8xRIzZnt/5D6Qn0LijZyiTNJsEE4JRgOHLTMVbUARANcDxiuJ70j9KJ1jMQbD8xkO6
kX2rarqXVqhJ1Y6pT3tYHXFHC0gX3hWNSTcMvPnHgjS8FctT1qsVte4J2rUdueJ2litdJwOpFOsx
ibBPGZbad1P/GkKiC7lK1nzWqgAak30h+dzqOvH82am9R1uC58V7L8VWIPtlb7PzquoueWAmE10u
X1iZxVIBt2hmryeGhxVDLxFdCeMXPJJK8jdY+Xc4xB+SCyKZc977dn8OBelUlbtM+qnjhyPRBxYf
cv7jplLzZDEDVlUNpZJJT+LVYTzNNiWMi2+Of/XaDbe4Saafgk9dSTbIIeGsv9a+JTqtdSGkHjLH
nG6Z3trLV2/8EH+IjX8LqzkPIE3682j2gBqVj6dLM+1uDKLQjaB8uHKuOYZgiFEzTYmqcXcy1+35
qnS2pMX/w5cWxSBTJzao8Vo5G3Y57h9Zf4XeL1JkfrDaO38ZRNxzBhKVdi0LTEB3n+BIHZYJnS2C
Y49zCQTYzIQF1OKowQ0HoFQH1209MS7wGPm3A/DFKA2WOa1ABJi+rGMhZJU2h1R2AlFh06e6WSQP
VtGc1JzJ/VK3JcEBvMhGIYVIndUOurKP5hSepgviM1yB0wRzVQ5ESJvJufCzPmMFgdJVH1bs9jcC
vfNzjMokZh07ifsMzEswpUHUFFAzoOeqhhiv6iFGJMt5ZTANla/BeFB4yNOtfE4/zTeb8qrQEc0E
Pii41SfXHjiDxhm0ZhIN6/usO/5jZEhg1r+Y8ZqPHxmHwDvyyJWiRmUVq8H9HhC45PVa9BbVZS6Z
Y7rQA7a1ZOC3hMoqXGoO2INmAoRVtyTYlefzdZQjw0uyquStgkP35LLAbnrww3zXC/ZQqf5ytGXq
IlRjrIkAH2BSYMrWWfkWcI/7migLrXmGXFrIdoRMVNoE1wdYXd2x2KiQcQCecgzXmTvfroCdWW0b
sepy6tJF/oETd7M8QKpT2128lIkOjgLbBbc9vWMDVoqrIN+qKml8A1bD0/hNu3urTPT2OOjnty7Y
6qdRTG0QdRbjsabuhvyGVNzcmoil3Odl/cx4DrHXSilqbAtm4LLBaHo1rIz3JJ+4s3ivuSS/Ceyq
bPJ1MGL/OgL8kt8JLScrpe7oGyBxxGbxTMJV3rAr5bNAgsdHTIPZdI/R2zaHtIuGWApaGB4IF9y+
eLrQNXkySem6swyc0i4uR2UNbiyx8s8CqZ8/ewRt6ou6tK8FwtM1HXU8jTQAANPCio/cZZzPnHLC
eUykiCY/NtyBly/6AgdIAEM6HyF5MV37JZ/NthSqDB3LfwrVER3EiQRz8ILnnqs+V16s0WuMaFAn
tGJkU9TSXnT39Cc7iZa1tNsUqLC5toQTQWnWciWEC6M9ZNpRM8I8o9ilF6e15WfBCpQu8qMkByQk
2Yr0aOgVJGdNCed+u/jKXZxwZ1UOchH2JatwX4jEx7UG7FgiL1lsz6xgzWqKsdgZ7fVLBxfMZgXw
mwswA5czyrsnwaY6n4Z1IyNrBwB1nh20bHDGlrVMi6dZfkzHD8QEg817oGEaCQkgX+hCYAH0He/z
vZPer+u+dqvDF0ReZ81gSezhEdTSfCa9OKsJSHytujtEPzof2z9OmE6mAj+lfFl5BC6mTcgytgZB
HwGBKEMjkuqP0HBYwie/k7beGG595j8WOBKMbjebIJfPU0HeNeNC25n9nDKGzDW7MLI+AqftcvwN
Oev53IzIE4cZRHw1WwiQvcW3SZGTxWpO1hoFAsWZg1E5stNepAFe1IocxNTvYRAJ1ocQQzqF9wt+
XhZs1z4tW23APKe16t1N1yPEEaT4/f6/f+0NT53sPUm+u78VHFdp0y5+OP3KJSAPKH5MZzcA5mtK
seT+xa0QnHTw8Mw7vbi2QIqCuID323QVAi2gO6r3tkwPhH/wQ915t1SeM2m5ClgNlRr8nlWXPHJg
u7rgI/HCFNKPNnSKIXWlHTzRjzaV5Y8LSOAQSgbSyydrNjEkWIJfIwJGQ6HcdGvzaP8YjyvfTUA4
Jrj05ZTR0D0VUjXaRXFb7uZ3ZnbxqQEWcOsGbPC9HRMymcFcZVSDO9o3+e/Yvq5RRa9WqgLCePeQ
sunJ8nYQxReUslw52khJwhm4fwJPrF8gPlSwTwWYyF6qW2yUPNpgJZO5VVe2oyV6g1OTD/bSyPWy
mFUHnUgHzP4X7iACLZEJ2i2mgxKS4SAgAQgnrhzLLp4uyXYjVyW1tvDN0T2lGXjhPlM7MUwl9yg0
aI/mXv+skXSV2MJFr3xgYbv0JZK9RwaQ72WI/E7r7wNY+P+yRHVjt/xDz0gZdvQDATd+ZOGSYrVv
pm70dZcZa+HLDSruHTc/cwe1ZOP9WmsnIxEWLCupqkxRwd6JW2TKLRPMcHgjvMCPbplya61dyVGi
LeNSSmPbpqPFyO8HqbYUSwp7qSoJHdDeHLV92L5ayypIw1e9G0k/S/9TcXbY605WTSQFAKqpYm/X
htM2cdiqHPg6U6NQMwEQ7MSFt+YuimCSI19KJh+vWgRir9TNLDP5T7SXpCnGLWUNOSGlpaPvhYa7
OmzdB7VkigA5WBHa6Dsju0lJn6xGVF6u55RZxQDs1/eEqai7SZUfpFcn2a2lge4oCduMGx3xfUAf
QQriCn9jJS92cDcfwpMNLxi14hS67ua0c9/sbUg/53JFP/nrEFc5VIKRtA0OatJ2PIaZPj0xw3N3
WM4H16I8IgsxUN+jLbAAZl4J1KS/B50AurEDVdyD7/1deqX818DtEJS2KVMoDWV0A0pd5SL5Lhcd
T4uaBq224d+71MLWjG9Zb4Kec0fZ0idpKTyvFF7nT742v88R/mmQ19FXrE/ijNrAC7y1AhXe6Mxv
TR4Fndavv85QxLJrkNAu94K3uLtaRmvH1COy1RgC/laLV2/wYfgbct+FzKUmdBIQA1ci6DCYtbgE
VjJuL607LS8Yj1H0w+qnvkSHIfgZKxFT2Vjm5iUQaavo+lRP5DMUbcNuuxudX1i7DZIC/eRvzNzv
MjVHZyf7iYzfEioWeF7fd5Ce4AcFJdLTs/oBDWTUGc2Mh+rd4tgFTUST7Skjv7l3zuLK9C8zIDQ4
HhCkTlVcbrxNI9K2kveBeBm5BG9HlyE2/z/Ry6MtwoSkcAHg6pLLTBuhdWNA8wG3+/3CWcjgkWEB
dkklFIrRTwu0uz2HPy5wfxBX+RycMyie9g+ObD9xH6WL1wF9wKJZy/SMjSOh8oY/aXCTa5Rr7bD7
OxqDD7gt8dykFRxwy/fBTY8TpR+nvWNhBpd7DcahzyQh6qRBLJ5nDH+myf0MJJT0Dcj9HVLj3/M5
wTqNVbttrRuQV+NSt5GsmARwivNcnbxtblj+pZHj8cwepOyYEJznHRDDEGd6GMJG1R5+AbU99AvR
U9jUEoB4XAN9skGkTF99xH9xSJBlsE4q9SeezzitHp8z2co5Qnkk/e3Z5B0C7Gq58qa5Ni2vja8z
KRCmL6ou2r0ZsCe9ljsZvjzmEYzH8wKOCbPkryaNfTw99niyVvUc+s1mZyLQMuFN8A4IZm8xHjgt
KbU//IcXEO5utir6aigdLhK6+oNs/O90pgD1+Qck299TU9ISBjUIhC8pAQfUr8Y+mGYDc4dpTyQ7
leHxzr30zAwikgPcO/MoQPIMbP2jnBfxdKI1/qmW2GPm9KCy5ZRDsBDyupeGWdpNbch/0EY6s5s+
E/KEYunLLeaBdiokslGUBeodaD8iu6b2M2RV6YaMVvj2xzrKl9CNz1pisUiWxjPmmBVIzRsYk6hX
7/Ju7wGgiZJUxqmYmi4e8a/gqNXrWn/Vm9FtJDvUxSPZ/57kzifZ725dMXjnJcSR7K+aEwKJa5Cl
z9pI3f8l6JfHvnwX82AvVeBEGxylTHvr3aRfN4c1mOqJYTJqzX2tFlEmXQS9xC1IY7M7BmOHEuM5
eUZb+BBqyJoOscFqtS2wcEifd0le4fujbr2jTERh20t+p/QHoHodkJUBupkEtG/hmvELkKPKsLmv
dFjNkDdoP/FEBvCpGQ48VIa8qyVyL9rVQBsDxwFsYhlE8A8gA1iSRP0pYZ9BuSp5AZAxMWUNcSeS
fIflXJIinJHHM4H39cYUKL7GLfv1/4+d4w1KD9j1vPHn6PmCZGANw1KL2kZncaPUdu8ZKCgC0mkw
6duwAVD9Kj9eKyIL9763Fz1mjgftPPwRxn6g1N8BVvuKccqIPC3qeI8QjWJoNVs8D/vl2lhldhD1
KtK8w3OEOnRa33wr4T60vKchrx615UBRcqBxRaPkFSk8FP4ZkhkSa8o038NQDGdZqOmSNikTqviu
l6CPbIQ7JicNif22ggWB+qYABgReMGMi26wCdit66m3YjdpFUncOpv2GJn8T69ui6kAEQWmPeupP
PF961yJYTinQdN1aEkHU91r12Bm2I84acCuZbEKA7J448VBl2N5RK/WMag3gFrgr2i9341qgDb1z
KctZpG9plOM678T9PQOgAEwl1XAlqHaRt/SH/KBY1H8JGw4OmOi1taI6+Z5kZ/t+hs/0LbD+wPt1
6Eycq/uuL2q1kSmmGIcyEsDekhQmjCcFVHjj4nMPQlqYyTwh5ojecAoexRPT1OtncZ4IEpTgGtg1
x016MpXFq0kPvENy+/OaUCpi4OE4Vmp+dquF0uvSyV67HEhr348krdZDmSez4Tw+6MuwXpoqaFXK
XHNtw1sGaku7h/N5mC4j+PzV4gB9PCI5ZIcqPzqVQfhbbaPgX1H5svguQRShqUsQHvRL9pz7N4LY
fOZcAhoc70DIyeYMQdy/jz1eLQhv2WSVZ0C5n6dUxFzqAfzSSDrfkPqFNI97MLLGI4prHRECxm+a
3fF2ZCJaSdcVRHYMF39VsVPRiRSKIZDqoZHAqP/nR6Bbdx6Y0zf91CYq/x2S3fQ02vHNQkSUDqqf
dlxGZnU2ZYIq/6VxgEsVrktekHKIiX26vlyNVXHSe1FXZZVCktWosgCIg4ONXgoVPDCI/4mI7oEr
VicnLblnKmF7qea2bsRViR9Dh1RKxOAKo1Ro6GwQpArzcBnFRskGwHV/xbZ/XhINMPljLRLawsmI
ieoqnKlYtbd5WaO/g9I+R3A9Iru5MnCAsPQ86fGDCYUN0orzAx9qPUFZsiL+Py+aCp0svEDrsrKR
opPRFKR3qev9RUWddGXe7T01WQDr/tBPyfc9ZJKQwO+4VfaaVOJlg6Kh5MYKa0hQJaLiOEs62eFI
uFuYow0xseOhzRUQexeMwn8fW2stdndgLoeRKeC/3OpWbTaYfR9UHNkvHJnm/GY44e0yShs7jdbU
IBDNjflNtB4T35URQtUlq8iM20Hc6GG0meibiifI/B9WqlKKh5uF4X5ZAoc1xiu306q4xhS2KeK1
XON7wCsYZMYMqTPDGvPtwqhvBstTbMYuRWNzTzWG9+4+cK+KEj4o+XmJ8i91M5MHIlvBTPIpzr+Z
gwQNw9BNHEuKogPtPA8LPw7lE5N6ADK9zKgK4hziKBEpoX14xfDnxG4bWXw0JJz86qp6mkfiMwq0
VJwjsRJ2cb+IxWvwB8846q5c1oL28jlq1VCn9Eg4HDw7OADHLe2eeKZilRDiCp7paC5mYt4p0cVA
mY+mXZ+JTXybx0TyggDddSsYu76+t4huZ2+ulUHHU+yAtA8VhooKxhrkZ1/GlWoo5LmYvfpYnhYA
4oO70l/1Ox+66v8ah1/K5swiDC/yia3LynBtWOjutM0udNe1ryOdBDTPseg6gSUyzTb0gIV1IIW5
9MAwuz1Su7ahSM8NIOnWbWmA5KHAi27Vsmriuu5rAVtR7+/46eqcZmpnEqJhCYKLMFr/yqnEQ6c6
W1RVrzDz6mPeLV6VP40zM6iLtKlL9iGE+VfhbzIpYVxWno/tUGJ2wn6QIRB9PouSycEbXazNDZHZ
s+VFjP/poJSNONshk5f+kK5gDEagrXJ9xSnNKFaOuHopMqg4g9BM48VVPGrfvxv+54ka/HHoPI6g
fw6KBAtOpoNjPcbmshyO8a2l4SnzGFbDz0UwnzBmB9VQez4Rz7/0wM3JISNDItI9R25aSyqRHj9c
ui83J2ea9MP9GpYb+j+z1A9hSxUipIlpQrN2QQhRySlPhPGmOgY80ghbXwAj7lgupyP4Vrh4wtgA
B7sizm0d98PSiQHWupEmNK8uuk6xHfX1PI1/O7oP/gmMLfvJsBezg/rlZAAdyoW3w7WNTylVW7yl
hlDoM/bNybEC/dQvVd/3UBOM9ApLCOptaDY/rg0iZ/2lUh2M0bwaWsoAoOGMAa/kFJBlTbqPvDuv
SNSa/HMacVHwMl8kY1ZGqolv2A2rN3IF7ePN6MkATcj2t4eWZjYr5BsFuBorOsYo+5C7hT7xI2nI
J5+tkFVohVZCDyB6TYL8UzHDPNBBMncJvYmdoLu0qbNGBCk9dqHonFi+8sYU9+iy5D+WGN7mTA0i
hoaFgim40E0qfOQmb16cn89dseBOVGVhwAJLp11JNf753DYI9Fn73jUmGanCYp/OuOVAQ1IYbliZ
I8gBhJyje5GjSZJqvZv1NMDa1uRg72GSLTlkeZ+QPh50WgK9yh6PW2EAHPW8L2v+ObTOkHmMO3fo
tjp67cEkmkjnA6qiydXkIcXez0AFlM/y6bLl13g4nxkD0lHhaoJzaVbSzmOybXWi1lf+oLTMNeTJ
Obv8qfXO8CBd/u6QYHGgoO/C0jUNJ6Ib2nnsEOum6BqvwyfU/A3wnZ0OlnqcYrVmVKy3RlFsVe8j
bzVSo2D79etL0uzRAZ78B8Y4E8qHzdz+7l/px7RyQ1x1w4u9QvMi5ORZkg0XypWLBuYwNT96TnRF
YclKUvqKvrxWyRjvJglqPOknIb61l/Ly5DmLCQUNEyp6e/ACVCP2ZP7fzNyCw60fUkOuAdPC9m+j
1QVCH98TmtdK6MVlnlsEO9ZuozqPt1N4zqHv1rhGKSJ7WrEyprMiJjkEmc2yKdjPFDa86YJim6qO
p1YP2+zltpXmhRrGKTWuVeNRR5ytDdvPWdqo8b9HC+4oMgqDC0DddFbEGN+D4/xA+IPT5+Jd3PtC
cnfW9XrB9D00a+bOYf8pbs7oZ7LYu6wPaDLSPg2hCUuTBtp721ZlA1ZIIqgIQ69xgNCiXG+lCfo8
wUoeVEYHsTEYMSRiTIc2t93Z8ho/QkWe+62/3SW3lSy9ejaSTMzIj+ujYjJWeGBzNeY/4mK+2hvc
O8NKvuvo4K5VWeVqtRMF6+N94ywKZ179j6ehEkQBPOBHYNnfm1zAhd31w4MtqqOuhlHNhH43fchK
UFQGyYQb8sVEP7oxxEC7YLiqSEQhustu0j/2kv2t4UEbRD3GdPwqACB6HXwvZcwP15ORTEADJKiK
ZYEEHdR+gAW/Td9KgrQAm7J/Mh/W9+ep0KLcOKHgHnuZGbmfFoPL531OLMokpVK+/LWcwbqufLNO
+P6u4fLB/lZ47x95qVD66S0q5Vmhvb0AEfKtAw2j44qvOMOFT34lnko7nC2Iy9jdwbd8kJxgGyhh
GRLxIHQvawXvGVH/x0sQYogjSkg7vem7/zfUumUWc5fMxZFoA4tWJIWoqBRIwYApwxQiHoJ4/nlb
iF/UhkOqOjgwIsVr75HvwY8ODSPT5guK0VruhHqDXPMYjoxZeOZvs06IhcUE2j0n1iHzYX/S3w93
+4TumXCJVWJNT2wzERzP6sF0KwaYKWaYYe+MMG7A1LCLQnW+uHtpsAarx/ad8U1GoE3Fau37xFyJ
cf4DrwbW0b4HAL7B7XUpax6GIPjFNqGOeMdKGzIwEUiRUaBOXsRrnJwC3DlfPWyt5wVjljW5XwW3
DXY98IGuaV1TApcocQFR5j4SJN6gP3uSkdPVNrNXLGaIrWQTv/mCWk4I8cFF0nlk9koRHAczkUuF
l/RtN1fs3rLWOTh/MvfCH0yvEkZ6iOPqf7zhONeneMrrOojqTb/d2HWSjitYG6CrIS1lPf5bRaIT
DwKb9kGvUpV1oVJD/TjqjkKMTGX9aGbemIJL9hrGEjWQcLvYk75P4OS9dDGyB+Gd/zwyO+0naU2H
dnWXTNICMiw8j4wCBuY77q4KDeLhYGlw8618Blla1+XFSTY27NIiJTq4LSwjw2WAEUNPYKEtXN/k
THDCfIamW7Ju5RUS0X7sJoFwoBxd55hf8jJEd1KCj2suX8RpcEpabcqeVzmXPWvUqi/IcpYCsz2Z
cOROreaC6kJPtHjrr+0D+pj7LARpzVSVzDSVM43feLvPXTyWCWFpV1udfNHFr9ELne/F+E0yHoVc
7UShjpjKBd28Uw1brUcxoby1FwVH6dXJhTztSa2IZevvtKWjOU/QdqrkdXe21talGHaQticgqANP
XSfcnTseIgZx0x9uQ0Lhz73V10Qc85IYtch87uASuCdX1DabQ7lHBFyUwPDZmEaJSegbA01+WKPC
8q51BxS4lJpTV3VdvIr4TAaBILvPgVjJVdTsv3M9enjNlGLDN8zQ0ROt3kYoV5Ybh6g1sMfkNfBJ
WdteDOy8Ocao/SSfjwFwZc+6OH2uOPvOLiFoyBxG0EcowqH99GqQuP4oJj012ORGGIWkj9kNXbbd
9iCy2b2jOEHhOcCtqkMHMjDg0JEmibmos2a+19RwfOUCDsm3dbXEwAbd6b9LbjSkwjXiJuttT3j5
VFne9lGo9w5K8CQiasqBwm0Yn5r0iwSxOjTOZ+yBt84s5/dkEOMz5Noy7YDf/m6xUewD4bPWQNBV
oecxyYC9Mdn8p8ehhkWXKFr7e1a6z0bT2qHT9NFwnlqjM6wFZEMoHifIvZgMtbh8hzpXuWMWA3DJ
6zO/QT5r+dSBtMQ2yz8HZSTp9/ayho8bNfbfTR7Ao5/FCTWqfsbxQvRpJO54jW0yPu26blHg9m2B
jm0NpMFxtxQz+NO2IlKloiKxBQcb2UnKi+ahn46vU4Bv8wLEk6Ix3qGQ2g64ZAhbYPna0Ildbf1X
hPk/ldASict6aFZlRsm5xC/cqL5cA6vUopAjTQJc2yf/yXGBAuaUUlap1PFBAhrejiQTYulwr0Gr
ioVNVKmlOeMaopQubBtUe+or5zCa47ZFFdJkVVkfb1ULAI/c12cfBh8wCxxQYbl7WL1M3MiQTVSA
/NxDDWS/Qmi/hCA/+3+TEovw06cEl/7VuxgJMX+xMWLbGjxveNjtLjwIMDJfyEp2yMfvGyC+gOL7
Z6QvukNJmzzco665f4GsZuTVQm8CN6zPe2ojlKvfVSh9src3ytxRphsTLWEV+emgNvx+xakmZKOb
v+ZAByk2mHfBcX9xd5Ws32GP7rBDcwY8lH6hb5wnIBXwg3cT6XBOslw+PMUXnX7ENxxanOrsaZE6
w609NUwcKKPNKmLR7wt858ix6Y9aRFMcLGR1vWEIAJ3hx/M5NSm2f0a+HJm6HUg1iBvE+N9zSUs+
ab8mnEsKRtgtkeervQI6+xFBlUMkAsuX7OSTVOCTQdxsW3ds429FFfmS6fgJJOms94+lIoIaolIL
pGt7vtf1L6sfBGfc0FVIoeaKYpXv4Ctde0tro3ZAcMQLdQQVHbc05+fiKvf9Md333BYjpyP6zjs+
XZNkz4NovSiFgb94lo0Z2PExg5fM5s2UPQK+fRgGkY+X3kaNN4MY1ELyLV5i2HlHsXzLG7pNDUGb
x6FlYVKLrwDcPBTn8tPF8RiDqIdWaB4ndf9Uqe4OLQkaZVvtuu8rJejhtpnAwoUWRFSXK5ShGYtx
SYDfOhiovJwhHTlH7X/eLxWbtEemZ2/wQYryFb4uyR33F8h5+0k3xF8s84Kt1/OEjRYvo80FLqIG
5j1UDhAK0PC/4feG1aOe5DC/V0UgbO8fpqEkW+UMOPaxNPjgk88YfUjl1GsDIRO4Nn7iBl2HWJ/d
ApqrHkz0zlP6zCJvP6CPH1/EJhgxJzBH7x0erqZMUqJ+nuWjv9+jvgvKUxpre+iERM5VuFkFe+Ui
ZtDWb3Agwsn3jgaGMNxUiJ5B5aYCbaErwcv9wb5y50HzcMIVj2obcwm1fjQtxhIBhCaAur41FRpr
SCJ7r3mRUa7YXub6flc76A5fDirwMnojXERpfjf88z22itxpZwKoCG+lOAhkF1X1nw7dOKqHCdDI
JNoRq0BUjSgVWjaJ3ztJYYIMLS6DujIu+zJYQoY7AqA3C+gcJ+5KSDgoMqb3dTvsjSKm+Wt6u4tF
aGbeBKKXO8rnZZ1nT9got3xftECb7rx2BMD5Q08wLkMKaBEv0RRewtGlKNUBpiXpV5pNUkHq/m7H
F/ZObms9lrczOdcDIb81gPTzAwdIMf/FVNUVU4JX/fltJZT9bOC4gZ/uO7Htn+vr4ETZbCuwq/dU
ZnvzddmZFLxjIKhDRfrlKR+YHb/CKPaSYHCd0047PLPTkfPMLEbR+3VLnvnLLSQqG4QUcm7pO4Wx
1f4KlMEmdNURPnmRzuEldoGsMhq+xsi4dhvaP7rWpQZoZe/L0552H/SGaqOllYNr5c5pC9z405WL
3cvpBJjP/mcTltBgYd1xrdXv7VFKaGyB3shSl8JpGp2LEmYulJd4wqfzqWinNycwUrXY7PDzKkT9
TtO3cfk2aNVzJmV9urFDV/NGNoamAbJklVL1jjZmNcUNLhsny622JEymXJt1RITPn+N3rTktwZOa
LuKyjWNElk3fv8W04uyeNMv54nV72OPDOoupzLSHuqMOhQEi5bRXx5SAUx6UraZK0wZVrxuHF3EZ
y/9Hsmvq9ONf4hyZXTZFS1YQCvRdIebSpNjRwJIVeCAwF3CVQrjJCez/6mkCjrwT+aF/qEjIKKk/
luSsl4NOruQFQky5gIFBJs8Q/74DG381VxkWm6FGNLNead28DoYR4BNG1fv6jLPfEqk/b1JBqvSx
JRtM/NnFLVk2/r6Ssp3svfzZhcn3/rQ8+fFO1zvH9vGa2XgbGTfyetfRu+UqGcVZk+Gy+S79+RL2
V5Fx9zLpwSdF99HI5U+Um7ptj/CHs+7zwFdIFtoLIG3PD5alChh9V7gdTfm5XSqXac/LcyT0dCvU
xjxYvL/jgcAswbH0HIkmzltAXMBbJDNjmeDSZVGtowdNML2TVBTu9EBjPaSgd/YkHhc2RZ4lXE3Q
xn0sxs+SEVDSDukMuMH61Tym2F8e/RTTbWfo1hO9y1jkT3tWEqhFdy9UfZ3X/vg/Xz7ONg5k8w+b
uDFtSu4PHMSEnjvIoxv6e2KiijbWkDzkb6gB4Wip6WNBW3o9zeuKjnY2vFjb1xM4sY6kpas+jGLD
Jr5a9PLvmm5r9SKGQssztXttITTAQ1IXTM4BaekwI2P0MjDjqfZdZFGGar3/uxzPx6FFkIaZWYEz
GRX5fjJKurn0fuM7JKCCFMgBlN9GSY+5EXhmBpukvZw8HOTF9YapwtCKztfJt90JDzeylvfsOyg1
Gqn0oJ5n5xaz2cP6QPyFEFNdf6cgNdRTtwukE8ILZ7Eca3KnPoUp57sU/H+xQBQSnU7hwxO6NDHS
NbKT4chRxsIBu47kbwqrm5uZ/DaLlwnSHaGPp3Qpjz4OjKNUSGjR9vjyurFF9AgqexjU+C6OObT1
7JqkfgcpppBlxNlB/ud9E12g6EHUzU9fPY8pPPiX5rGZ3plzUU7yglAgnubhReL7s0pm16tPzbOS
I9L7Z7dktyDg4H9m9xInujOGhccduMVTFstRrs/BCjwFR2RiXFYKWQw1LjoPGIVB6rrVH2PDBXeV
89h+9ny2BEF9g5zCzRPd2X5kYgqONgcwWvJPX0mLy6AhNFatQiDFwGgYa9BbZNddcKq7n4KAw+wM
PNh9q4z4GkM88uPsD9i9AGo9SeURmEGGiUpjXtg95Rl588tOURO985/IshQOCuBMJcVVh3oGBOse
w6YGUILPkvzGqUExOV9CdpUTAARUHNKVaP2FDzUHNMI8mZ2AZgUifY0QGjuBWNk5P9oYcktnq98x
jbZ1nklisMTQ1VzGlupXTcCx7MidRiIayj42bgIip3qLupbSbmSKFJNEqlv1HPKIDlSzztN4JW9T
NvvJxtWI1eD9ogZQbIx9l0sWXRDMEhavSn9+EJlEmY/kE3W0HFIbJb/RHIsNbqPOQourDoelANQ+
roXv2heXGg/2YOOT0RiEOl8Rc3rpqTbSiVoCsvy3v7I6+F8sdPsQ78BNu+vjjbsGjQF7exiNZcoD
DhGLN8shYC2vuQa3T0aOhkGL+LoMrcdqZTdRfByVv/EB/dDnx2nVcSfuoA3IZs3JTeuQs8CvjSv/
075tSr4OkLne+2WzbE2hOtum2ki9Y2XX0w2sdCrb9F+sIRaHUAxWrP/71OBiG524wchKSSPjJl9f
IYm+8rfT3rDvZ2xLM/btv8SG8wsnh6MinvO3o7Y1/75FHb39mvkleBKjXL7eLVntut9r5Ya1BkRn
kmEnBVNcN7lXtC/PdW0jfsqqTgsT9w0DpomXffGgl04CvaSVFY56J9wXa2dNCBxDDcjSwKr3e1Xl
J+c/Il29esXGONluy6btiltBNRg68w2oLOfIs8mL64fWJ5deCA+WkFV6tjLGcNHHcBVoj1SZIpHj
ojWdpDY9iAF4y8FyckcTE73+4UH0DRFXyHofeIPmu7DDXidW0xrYs7VvHe/6eKlIJKtRQhxDOxdU
uiUwvbPbDKLMMdpa8hNePKbz366WFXpaM+Zr4/CCBinIuNKu89zu6cRuirsRj55mqdtP4WMIpUPG
srWgSDbOyBs9SMiEeLwjxROQaYTy4/Ni/sOB+cUL5iE8i+d7xO2mZxNQFHBhDDSX3UTLKBUWc8uE
+ftzmeNRjGJqhL9YGAwwKx23S9CF/8D1vJdfjYdFOBySNE8eC8Byf7fnpDcSahRTQOY5stwfBwiC
fQHlI9b9DtlnEdGu+o6bXp0ox12nXv/Smf5AZuoi1HGjONyaAlIv5WM5jGPkfbUa6qyeiQX4OLV+
HNv2hZjmk5hnYjjbnkmoIeZeOAWp9p8iLdpEu4WGkdmbDdZDhE4mjtxvQ0486Vz8rz6xh3ZBpsWW
Xs5VFMMj2j/7XQTOLE0F2f1RPWIm852pA1Vm4KrbracTz3TFhv4lLwWTx7jknk/8zbay8DhsY+vz
/gThzViI9phh1qd8uJCpwtrgSF43yUEi8nQj0OST/hGweb3ccX7XsETcVVQRRCiXG1r6rm1MidbZ
k6fkRKFv/fVx1qaz4VehM0c4eqkRwqMydz1zlrWblyTamJrITF7/eQRJNH2c3zbZn/gDBO6/5TTD
/IZYIJNRgtKPGb3pK4G9yu780dGs7p3Isy1QnIGt1dwI0FP+YX4PX0PW+8VYcZABm6lwUXZFb1om
j9THBl/aoNK4RAcvabz/bbyocNoiFKfdNwAujQQNeRlSMpWfeLv9ZCWaTPYO44vegQDPVGHTQeCa
l1Lbs2ZOkyv3vQv4Bfl7uvK1K5cVYP+6unVLtlC/zFlCsuAn1L+cHXS30JwLMEAjp2+WDuz4HMSg
rIA5CdrjzodCuHYgXKs3m/5XDtR+FTWWbINpSvMYWgd1lBc3VmwJkQAlWggtxLAs8jx2BOw+CWUE
SbKTtucUhkLKVgP5RBPWKGpExf/nKywijuxYJ4VwOc/rfOQ86oUK1slEoPUY4LibfWcUg+i1uGdB
GYh+Z60pyaaaAkYONFO/P/io/yCCjfvKr1eszAcOWssSG47ZeM1/AuIRU95P8WDFtyHexpzrAcjL
beWlQxPDaGFyhmKMhlYs7ciK6fBdtjqUXGkqR+W01cWY4ACKk6J/B++cNsNHW5PXiaclRdtQ3UTz
IfcwyZ/iUsOuvguIbosU759+oGEzYz+rw5mtCl1Tgr5pEEyEb1qu5fy82KrdRKTzpWLEeOb2Kzal
GJu4GZi2VK6KmbZcrlqSBBUTF77sLAzH4WJdH07itZLL7AM+6UWp8kH2tK1IUD9WhOydj9gaz171
gQ2S4WWp4UbNghAP5pFCVQeGBD/KniwWiAo1wFyXJsfhRgjUbRB1MtwlTG1JGue4aYtrpb87j6Io
jLn7/jbaTiYyzGW6U6AgnzARlKGfDjsZUNs0PcfH2M3CXXabtpXu9hGIAkbBqVEyvh5zWCt98bs3
zU3PpptU9skkIemahKchijeJXFFYnvfzQ4AaCAUDdYGx0OAMTSWRgdLfH2i1tAnqW6I+CtK8wsPk
Coj6pTeQyiOCqFYC56HSdyPo/kSxdStc41zrAyBGttC/REMcxqKC8rAheb1id2PlgPSmhTEE/hcI
xlBfJIY8e+f1xDlNonlbaKysEAS2Y68wAXshnDFBTgbjI2Wd4qv74XlfmZu9eZ6JsMNzMKE6hsFa
cSMPeLBmq3tFSQT6m8ucIGn4/RWdQliXULfOwojzvCP77OMLOIwkk2k+iF2wMr5l1MS4U+X7qCLX
l+fV5VWdGoi3SKNFj5u2DNZKO+TpE7OEnWx2b2Znv66IpDXp8zRtO40u+epyDtIfiB9KJyznKRNb
v7WTgcP9LUrGbB/SHtxutg7773HU8nfHt17IxuwAXrAYuUE5lzW8St/ixt508QBpTR4gpM5phWvx
kC650xmLWhK1rdeREpJxxfsXiu2/MjVgC2cYldeajKsIv/kmdS6UXNUG29sUXG3xuvxPGDwDW2Cw
ebKHc9kt785CRNFu8o6ApAZQXFmwNGM2NNdykciCcegj12AmP31GRM/EyYVYqCXqsZq2gZpUJUQS
/+8+92SgFTThId+6NFNW26pY0tI2/9wdwYKZQ/I7UtpxPBYJLyAxzZWsQur2PoIfmGKR9+0hbVBa
rtPKi18rhnj6klUkZF+orx1mH/IdcWyLutW2qwnwPRqWVmb+Ub0l3u2T4/kpAE5elsfO5udS7SsH
52F5A4IkrLdQef2Gd9CXpkZ1zWbb8uYn48nGxAkzvsgxCIygrwhD/WK5lSoK4M1dlt/LpTlK5fwF
nDDnqaxlYSuFmcI3F3hSyu73ke3ZyuVr653g9eOnHJD4imYSfWhoU+jwKwr/urpN/JIKpFbdqNH6
4YiQYwGBSzianP2jj1yE+Kxb3TsgMTxfsVlrDNlZmqcDxzXjc3hMMZenOvwmA6rA3H2kjLO69Kx0
FA42GEZwGvwXZA+YRhtE7ve/81oWjJ8SwgG/yqz0wNWEAvARJUvlYS0GB1FfKvjSI/V2ydhEjmHq
HGYa2QYXaDO5tuCMBhB0AQ6YJna+Iq/ZQiStLuqOAlrC+uN+3dTKorurfj3gCb+DK8utc3jXzUUL
CHyAl9/OybSTN1Bo2KIRT9N1rYTnCDWZgqSqI1wzkhX1nRoe1JWtkP0RgYO/fHHZ2xcIunAzIN8A
JBiRgFmUB/HvacKsBaF/O5DJBV3J5+ULMEGrRGHUodHAIw6aJxun9X6EgrHLNVfQ1OCdgVd12oCd
K9Ore8ipMDedQYfcMD/1nHLdCcIJiNxp3i31v0BC+8ENgKXKCxJeJ3b5ITfSnju7GfOgJtp3hHSS
EMDGhjw4uFMuiXuJigQfZWZ+iUKNyMdnNR89+IxLuqWbgTe8aEUc5DTIPwxbsejrQlGieWp4TgRL
HyDUqP8KlLBiIXVT8ixU6QXKbSijvrC/JONdP+OLcxJ2QFH9yRLL5WuZVhHxcv578W4ClwO9bB6c
v/G8Cpqy8YuNlDAZ/UsS58F4tQ7YXM6+jV0Nolet1zjGTU6ps7fkxdA07Bfr6iJ9UmjyYZrrntoE
F6suA44WImv+xxbAxZMc5Ql2pwG77pOEAioInm6fdvvVapiMC+MXigi7FIv1Z6mywkWxm+vivb6f
CPgKIkQ7O4PJk6sUpRoJDlVwiJkG9MZLSMUusMBOwd30TSIVFOV2xD3/42sUGZiG8kZNqXoJjHEg
QosYZVa13Inf5v2AwhZ0N1X3s7BDsioftYh2mDX6kDAaqWYO1GEYzxu4O9BpKBDgY7qliSjQlHjI
/V6gE4Gc4kbTEWQIF2nFQv02Drnp0atLedjbIv4E0GA3eb/j5Il4k2eLYUPqC3FVz4uZkcSpmume
sVMiM2PYaW3p5GXWZbAw/xA0Bqx878+GsvxBgUczw8F+VZMaJDw+elut+VShUUaGNHvZEg8d0JCs
mEDsflwu3RnV1R54TYh1X6KcrP0mcfuaymgSZluHcmHdBC2igp7YORLr0rCugr6bWEZ0fAoIdSGe
Kw2AefhXzadqc5LfIPUvbfXTEzvuFWAKFzUzNBNNi63X/gp3XjvySVXYJq5b284LmaF9kHRttTWK
C0M1DF6vvbCNe4k/psHE1zei6oV8SY9ft8lFTgB9DkUxYhYpXcFMSObHzNKJgw/s8TQOQPRYyAT3
UEYFNGLhedn0v6bglAKV24F03abm0I4h062F4wKsDOHVkxnHer6zXzv72y9NZs9WZgn1UAvmzUwb
H13H0qtMVh8BVi6hkGPqvI6PLNXinwAcAHdsinyQ0NYRGGorW2xyRGBDBm5i5kKguR/XADbF1axD
2Z9TxPhR2U/6owQ2NqhhU6+lcFkMcKo3itDnhkerX91ga/TaBGqkFz9zE/nR7VMPHA5gafWFdSPu
AhzwLSdSI0dtU+q55TRzDeNB5E7yNA3fjB9CZzyaTI6wGgw9jNovu9PJO0O814/DG4j3J/w0DCAG
9mdPk8FRFfXSCvYUmERx9DlAffm3v5L7hBJLOXMmKXonB2rgNWx21M6RvFay85iYfqcb+26Zl6Oh
OgIZz/SZMMhkgNoHP+glLC/Cmjyrl1a8crJrM8T8kusJ8ATbjMgVqFyY2hk3TT62F1LryDHfd+j8
E0IClYrBfytN7vTieLPSIcL99qAaT7Tj3aceQQ4fmICIQ+oAZvxm9tDhE0WvMvirKMhsB7huFm56
/zlP0hc2Samo4FXVgwdqPa/3tnbAwUogB9ke79CDvXj9pJL1fDxWDL2FMDI2zl8pBFZK9k9sGh10
CjWklrsjVhu8R4RnD9SjDbTcNwkrMouVdyb9oH1ifCePz3wPmQsvmNmjb72CUF0Otn0m98V74O1d
uBHO0O0Z2APbCvG3blu4NLgG/vfMNrykSQLXG0cxX0I3yuCOTbVLBPq/ths2gXjDhUx7J0hPuIXp
SubwC8Gk/gMXV+FavkZusk8/ssZbK5ocsjrlukh3KHzfqT8ogXMimLAVhNtfA534zKr/0EJCPYHo
D5wCGJ0FiFMbaOW2FxxhZyzf+zaC9a3YCcnX6XkCDgiTk28gqlFkby2AoImqr5wYndogNa5Mfzvp
z4s0cDdTtXvBIBg41ND8aU4iW6JdZGzZWjduBEDy82sW/eC646kMya4zOeXmi3SsA2t+MzltZwMh
vFe5tw14W7u+ak+zbU5MnTZayZi0WrkdtvBGV/ts4uxBhqYnalcRpiyu2W9X3OWbX4oFr0z3almH
7MciRh7t+W/u7+q8w4+bZ3+vMSlnPNI+o2lNky2zZpd+c+ECxkj4Mzehxo+KL7NHC9exDy4gmlZS
NeGq90HXW99l+c6axZhdISOsTomCSPxKCU0jf8XwhGPXkifYzWxeWIP4FvpjhMC+1U0vLXKCwdmv
pTb+ywedSgQCFRpr64wW1miM3VVviTCPF0a41GTcMDhv9+CFbhAloFXsL57b0snhAJxBTE+d7IfM
ksogj6l+SMlJaUrZyGb1iyP5AWODpuhS1Cu6L7LXpjBS8jh1Kt7wtCZ1Y4DaTo870MwK9l5gaOJs
xKFcEZSUiVio1DRn+Pro5W1q6MSy13QkvZHqWDF4jP4xJDYXOnH2wzwMPnVJqTXgUUrJ5HbgYp0C
hXU58kP8NIkEbdQXDlvu+DIWUL4yCpma5ZWcfDPqwGnztn+XyNaS1tiKzSU2yletjnZZ7gDQi0PE
r0zcakjtDXEUYY4QrvuJsBDqGM54h+eWrertyA7AwqTdGU8pfvawf0ZgBj8KGp1nvYCpKXwKeoJ8
umiIsiFpYRkNAE134CJegqMZuP16W9xzh+QY3lo/GvgweS0e6X9eIrs0476iCr8hwsv/qdxqf/9z
0a7jtaACK9T2r446EGjOsMQaylxQd+g9we8R36b/ZzapSxIoeVnBFSI8CjagUyGmgU4cnLOull2z
yg/YsTlI/4mj2/xz//3DeVojvCOYAWs3CoB/WNRQHVdAmCwy2V/3oywF96ZcikIuZWUrDa/APZXS
vwNrmHZ8kpMas2LxrPAQpTO1P0Ibmkii838Wz+4BdmNJmSCPkQl4rHfdjLXEALMs7oPJfBEy10iM
x+BTtvkzCRr3kej41qQBuhdhOtbSACdMHaM4i41pxwKLJ6BqSahTOCArEW1aHAh5DpDd5Cf31rME
Wv0BtFW0q5HXMfQDjywQeL4rocDt72RimIcFsRw9lS7DoTAwksDcB14u0ng0SHUxHYUyzlIzRKqR
GlZzbtiYPgPM2fXNhET0j9dA8pwdfBgpYprMeytFKtvut5QrOHWOKDOv+tAFiWGCKBi2kVrrEJJI
yCFVy7LN3yvyGdLGatOWHA/IoMUL8MiYtmKYFMFY7up959Os/2M1i1qc7BmEzkTcCzY1RTxSJ/JQ
oFn7GUAYHBSjGTdeucBBsTZXPZbXQqCVVXGH1ms7TPw/NmdjAgoMQhlI7CQIRAtIiE5QTJFyCr3J
nN3H8ziEY7/ImPHfcGVqP9ra21BtqnzSXYsy8+cuC3gVhrS99w5nn8ZszbZwefbPtQKuEx7BJ6kH
euRb6VJzuslmiN98gNuTAUYjQI3MEmegzX2McA3Z/ZEDiBSrW3STTHo2I8/84bKIhDBiwyydwCeY
8J/CjPXqM1chX2S7V+AoMGzib9SY/ArSKf9IB0opuKRhEBDUySsiYwksOvtz+XSfEXw9WIkm6pf3
ey5qTu7Ka9CdQa/WGwQa4uuJ0jJKIqkWkeiwmziKh52fnH0FdHPk5aT7c1lsknYjtPeQ/5QHCwOH
P5btQjG3mkahROuRtKtHa2S4y6XibbPa23zepYEfis3rtln0DoEyF61iSgAiIgJN2OaGfdpkoB4o
lfLqvtFU0Y+BPDGdRIemW9mb8Zge3ZFWlAw0DH9x7hDLjyOcnT6qUJO5QgpIMapob+TdkoESAG9a
V9mZiPxG535l4Pg/KFI2bgH4mY9MTaUqpbHj7+ZEhCxLJ1giV4dFVA/D7QjMKedcQ/XXsNqZEMJb
dwOhzbeOMFDHZX8MupiPlm2CcBH11cFtG59WZ9OdE2EJVVgqqcBc6/6wbcyNyEmspSuN0UEHCQ8S
dnE3joQAW40y0YO3AeBkuaoDCWx4GPLlxLJHKcE4u+0AUdXvNp3sYUgqp+Yob/urlUJ19vA929kt
tTGmrP+J4NS4Ion8+TSh6rNFj1vRnLDIEUuKvx0K7nHQubOT54ysklLPgXalEa2Y4k2MJLq+WSNB
qhluwmjGUGAOQ+jmQT9W4ceRQ19ivfGWJCqsb/B6ezlRUetGryJ/MZ3RMH0YWkY+72TReZqh+lik
DJwibqmK0qxLcy0CxQSscad/1fGBOjTzuBI3T9A8R4adfFx7+ZLCmhXTa9pnQurkD1EdjpL5lyXO
ptnAzKCiJ+RXlomZ8W8HHSgmDZrZmvVSXJ5E9d9YZanPJQntCRSqzJdsanKxFXU69e5zzhjZn2dX
NXPV4oEpFqeabkLiVcltCtI7CmavBPRVAtzlqebBmjlQd2bDxSRtJPRdNf2bJ/4W+fNXlh9Rs2y9
N4/m+XQjeGmdkmv4drtqPqNvuaTg6As5Ut3GSdauJ2OyrLlqPtcFRnu/IRKwzvtYqPn4PJhkiIUH
joxFTyx26Ez5d2t85Dq+KHXG//kfhvV9IM1u44CRrbe4F21k/huI+KPE/uPrvSkp7mya707QNqN8
o+jGv+Y9HP43O8AM7O8ksrdnUfw6mIEkmrVJVni05J+Cp1M/o4xxnc90AQ8e4ZUPVdW7vQfMKqpv
KUB5gnLDxsnBiAyjUETK640mTGkGX7rINbALEi4tnRyMOOvBGUicJrFwHEO/S9boXaVCXCSqzqG3
lY972PFx81EOi7GS7o5kELj2qSloE/VF1CQSBfMCK+kFQCmCoYOJ59JdIlmx04MspHQO1045CZM4
eyhyWbICnkoXK71KyWHWiUEcHSWmohL5fyPVxzu0g30eCVMibA/CV1V6EE94fcmiXj2GZAo7Aeqk
IEpJeT8vvQlUDG4sDlXw4nLwDmiG6mT4nrwKs/BMEcLkbLKP/ivGJd5hsTQZovtXm+oPk33uNtGT
bZqaGKfjWCfNUcY7membRM6Jf+Dnsf7ivwU9Ahsb87HvPU4bucN1Gan/5cDBdpwtH1jYUv9L/4Sl
YAbxZ+qDBl42YkixtJHkNrCUN6EgXHbElDfTyuC/d/MJO3VmDVc15G1gNMYZcltLcFNI02gxG7K7
lc8lbLkOk/k4/ZKAoimBWDCnUi822CxovPLMMNUudkD4+Q9S/39eYHtsLhB/ekRWeBAh6jaDtiji
iEb8QTS0qdV9aBR4dmfmzNRs291OaDfYRgv725pRGh0M9Ox80aMYFtOxW+VNeZp9rdUsAaBJRoQx
ctQF63privdRhc9/O9HY/1kF8Ju9PiMeVQh/ftNA64Y7bry/pV28s0hnUbt9C5WKWuHWgDQiNdEW
Dpd9FTOtItmGmcaBOTrd4nDYp00GNQ7FnT7ejsJvS01GIksjPohPF789zF53JDNWhM58RkxmE6wt
ly9jzrKPpmKD+gZxeaPcEwvTHDvj2TvNlTis8m7DPkuyT9HTRE81qIR+byjgEDfihxhqimNVFXR7
g/iO7oWIA6T/zXYrpnKVdqMYFm8uvQnwR3hJ8/E0lWaTIOfSOCtdSyAb++xIpXNmfPcoIrbX34hG
qwkm4JhJoeVwaJOxSbKCDbJbTGNC3NBfQtMz6YuhxUExuO1Eb+U9VjPiAwEGGr+p7rwsDorXMsFC
hSEqCcRa4LiDsykSFFdCReNtNnbY7dMQtowYRqW/UQVQAj9pb3cUpvZJa+1l2nor9gKs3wdvwUfY
W/UsiDksKYxUtKbRYgjUSIk/V0DGvPZ52tjPPzyWwHhP11nAN5gk0mfX4KcC8biXE1ggkr2Tqsgb
JdPt2u5APUePy4/jFv6rzjKXImifvnJ3W7BAVawS/I3KmVbMzNHXciG5D4lRehLTkNJFoKv6C9Fk
BTn+W2j0eCZaxBxMNEKJuJM+39DiViMBP6b9G2IUoIotYi/w1xlBFuhugMNKK+JceYaxRksKWWTc
hi9fcRApNQF9doB00vQulck9fRTG7HGdNOHV17WBhX+K0Wy6lh+D1MFkqeIzmJv247MlQbRIB+WY
KiSKUMakWXsTXoFBGN8lqo7iwPTY7Lp4Jkas/YhyGJvGoXsGq2LxKj+WLnaisnvVbwclRBt++5Ea
uZ9rvE6jWsxyaDXSc5kw5Id2CFo60/DuL06EvQiDVp0gelhprB36wf04diLtaGqo+XYYluvnzmWq
NMP7gvEgFnRpneuE3TJxiKSJeS9DIekA/YTEXdV+lwA9VmJg3vxquDQu7QXVMyL3Y9NkmJ1gGsh1
MQZoKLJf4JGB6xqF2wsOqYPbX9Yk3ao7LNlOgbiy1NxMvmBydI7nPDDc5FBVICxIEuR4oPyOiaOh
3Zgho30R/eyuOb4Ef762J8FHvO7efJGbHs/a1+UipXR1v2tVU3RdI0qknUI5femyos4nWF0G10/I
2WFr4kdRCFBsa4mL0mqh+3yWd6Vob36yOtFCRrDrLDY2XUhK5FByrGuh8XLrRxGleWMmogM4BzCn
whFe6V6PZST/L5YjLkn2zQ0Q6LMvtVJ6fEoyPnMyM4R9YfYIfH7zIk0sVoMVp/rcCJr4789q9C6y
50A4sfiJzFoGF5ll5NtbWAj66YCnWllUbSc/CZcHJE68je2U3PazxpmaNHHc+sj+7zjrwc9Lg6IJ
uxp6RhHAyLUYSqZkA8HXUjq2y/68wSmzs71LycxDQLyjuuAgtWESFFTmtci7CO6/1y9JkK0vFtTe
EuZk4ks0flBSEM66C8hNMTFh3nGn1EN/nvguFevl3CfNBB3WNBc3vX38pbV/Sxt0vkJEc9Tk+KPL
bCf0A9YzxHWQLxcSLa88EmiNX78v33hPzWAeLI5v9TZAsfpMHrj6NJv9OY0uEN8yBaVI/0LWOzB6
rzx0IFiLWuIg9LFZA6y2djjYadm/OPQDpShqXE89sgFv5D9vSKr1Mo6O6T+9mT0A4xJJAX192pOt
N0gBPBGytK0jlsFFgS8K+8eFzE5r6j3pYYl6VT+uI3wLwe9d4tsy6VTkThAtMLmQxqSvggqE1NJV
0cp+56P/JJOZi7cpHtuKimNTfRTTVCESNahbLAYhpjqWKgwDZhz1C4yRyPS47WuhLJfLyXHBNmlD
PiaMssmgaNkPYbqjlDJkkNiUE6Bj2z7BBaG3/eotCJsp8gjE/YQ8V9HdJN4DunAULSP1SEviFKO+
J1N5sdam7vmNCmV/rx1YIRTpFBXks+XyjwdduchIDnDUE5OI04nJotHTlulXsLoyj/Sqcbs290zr
sUcHIi2jCTl87e0W/7QafvvXyWAah2JGWOZoK54VL8bqSwO8YnhJhnzRfnWWpOfyznkKDPdmghyE
PG4IVYax9Jfw3f7vJxEpvHXa3BRty0nJMycWTTWclPOx6D14OboPv9bW3n29uNaGCTl59R3VLyCM
7FILteXQ6bXWIn1/3mI8+uO7fhxnKzF9NCHklEcgzFj9lj8sPzFlmXvfVNOFRe7DrV6yu+WeDZCE
jETPY6Pn7UrGfPFKK1LXIEUKzfbb33B5wD7M0OXqK0Ws6aFWN5wPJXCb9rZtSovVrTEyUMOhsJ9P
Iwfv55wDGIQ2CbmL3vk9AXJB77ZLcDzIBJJtFMxeiiWMRe0SpMIfkTLR/0OSz0yeM4E7H3nd1Imd
TWdcLGxo2a2t36WhHtu7xwtD61rw+qLVM24aowNL9AkutAE76l99NWfnZ7BIn+CHLTvzxb4oHlJx
R5UUwgaojx6YP7kePxUOELx5LF5djyi6Nxs2Ga3hTu2Yr1zBq6kr4uxw1XGeBS+inkcLUtPWDc2H
O1gLtgS0nsguBcqIC4O7jrg1aQgeIdcBnRgfgyd8w9fGxzRAlq8/BUPppWWqPm3fBNjp6XSlFXOv
VvW9azUcfcg0VLV0ucp+lnKbOVsiLxKMH88yZbvJRS93FM0eyy8LDcCIHhYHlkzKgv7j0+Z4Ykln
lpmigrK4yBNnY9/AZzVL449OJDWLs9/mZBbLnDn28iRdvcETKpjq61B3GI0y9hD9w8M78/IH5YZR
5g1SdGYq9KBrNGQAP1Bu5nAzU86yaj3h4GK8VQxPXAN3pslV/8pCZZtZonsU3mQF5oC68A7lBiN5
igJJCNKvCc9vwSfmnRq2nMMFvs/VnmgTHsNndXmCykeYBK//Z29M7nGDoGe5agyOg2uta1/uMUoM
zpXufOpDrgBFff/W7IMq4dO5sgiy/oNvfmAByj/ZUH5abmMBLVPyeGW8hR9XBQ6YWGwuSqLNmpWq
YzzqW9+RtpIOwDTEFYcPgKBntkBrTiSXzNHTR5dVT5bKRaq8cWw7XH3g8g7lvF+OYaqhugE6XNzb
OuBlt94MtIGCW2qKzvkJKd/3h+toBDNiyo+kupqqCIZGghTECI/h2BceWq0sjuxoyqxmWWSvAXZF
i8atHF1nrNawEL1hcpEfm5XWs0dCLCaXTk/0Z6GdIoHt91YCH7dwFbV7ogr+CwpLfaPVNgwzME2t
w8TJ0AqvkFGKPt6v+Bv7k8rh0A8vRF9vZxBD8xapV1dAOFbWws5J/fE6DuSjzCiXH/EXKl4XMGhp
Fc6Lo8DVwMX4ZSmTqKj7Utt0A+d/QlRkj+pQyoFPrX8e0gcdUNG50CQXdyNZHxQaWyIdvlM6eWD5
85YcDe7YhWieFBaU959qVnWiIQ8yr1IxFGiJVosme49y1OUtFoLdIuZ9/bbU1M2AYOtTOmWvydL+
eowYQE7lNv+kmEBj13MKFXT6RGFNnoYjF7t8ojEHvScSBadf5S1v6yXXIdTjOjDQwtslHN/ywb4Y
hJ1nHAlhn/X/m3tGlDVeyOGfBdaWAdWwPZD90uROg9rZsA1uN37QCYhQJKVWAp5vcyGoJDcWiL6V
wlm9cJ6OgMqOY5h9OrQqEW3V7EmWs3gb2/dccvUSWdbIVWxMw/FH6+ES2T1MZiJx61i5So7eoaBd
Sm9PAIHbX4B4oL6GvizLBlTYT0ViflpMASAgsqnA4jysgMIMadN75URvJNkwsStPuU9tbMGgvwIs
nqwFDFyIrJ+tHTnVFLpLNtHmEZsPIAJX1+OWvsCbJ1ngxbTdBkx2H514hFdH98oxzhB+3HavvrdD
7ZtFdoz9fxCaZPtehHVDuWoFfVVCoUlX9QTMyxwVv4ThkqEIw8VWyZiGL5oZ1sFSYdTMirVMXnAB
atNB58ZjZXGYt19qfyxXBzpWmLBdUy54aVQw7t0FJK3z9Kt+9io6Wj0q0YtTGSNtbidkiDsJC/vu
JkbLcOsI9sGbEB+uZo3kncWPMHD2On6rfA78HGej1TXUyON2NfK2k3GRnBHPfrpxXjxCozT3nhtH
t9gC2OeAcbG25Z7bXGvPR2XPuV8PNHaalUFM2O2GNHHi2UAhsRY53H7tl/e4lhACVephTyQochKe
KD74XQpJqyfxFRXeAhoxyVR+zzsWtQGr2pWtAHcfv9HgcKLPrMKOI8wXSlV6o2bLhjGKH1uzf9Kp
eD15niOV+z10+P3tkd4EJR4YWewL384mVt/w+tBKiiTIwdsZmNyPgrMow6UvHxALlFSIUwNiIA41
lMp94Y+TxlUvvGiGhoizvE7HRQJez2xzh4KRrZVzOdx5mUpCfscVslOyiGyRK7Lrpbmlhe6lo4Yu
c6hBRIpR20kTWIKCcbmXD9qgW05kpeVrNhWeLhc4z8xVZQjUW4Ndsz3bfvOaBNUR/D4rBlYc1jXT
9CBJDtGohm5qOysLFABkGz46RXmI5hgxSY2cKb0mZT6YNpjsbKf8e3+tlgCL5kx4UEkjaMCSePkR
FC8bbs1b9YJMr+A5rk2UsVNLNAu/nU5n7cz8NxJe/2oAbZh5j48STGAdG63dia6uHhlPUddEuHyV
cR6ncGQiKgnxKcLlgCohYRn+WCnK1CvpR4f1nZ46tIEYHQPrDJ38rekFnJ1W/5cf/lR7JOvRS36i
v/BJaoorDmQbWRaKRxI3+vKHBM0piOzhlS8QyhVn4I95shZhO+0BST1g8gKWaS4Z/nelgUuxx+U5
t3pEZYfHOqbFwmuhMxdQRIBIRkVBIOTDJakqVOIk0XqeqPX8BNBuobPH1GQBJQPprEmPx8u+/1iU
tHnY0q9VuJaf2zxqifqaNFvbWG972JKp7t+nlMpXyUZ1UAWRDTrwA1mM9QxeiwfJMGmPe4DpruHG
q74JLYErK4TaXpHKwn+g7JtJujrCLuxAASbHbqdvh9iykjLQJbAt4HVaKt0sw+gShkYImu/ZV500
sEIeyhKSTzvFMWjqtENCraOqnWZ7pMTWHfFEDB15/1qrKJ0X6teMSGKJBtfhKCTw9g7R0MaUnliw
luZzIP1zVTxSxgLvOe+hUkTi1YTvQDf060NMN7ueBQNhIGcuAa/HpIlFVT/yXJIYJFVeWFoOh5Vh
0Na7QaJFPvqKT8UP5fQghCP9EaWabETTplxeWfLRGDvTReB5QCkBe0TtbvG1m8Ss0EUrcoFH6aGT
upJd+KWt2LhmLYhWWWFSdidELBOLTUfsIWhdk2nkfzlmys2TfjaqgTUSEALBB7ilNgYw5n4QDFnv
cEHjTcVZ7Kbrevfe7qzir58rksURh464aQ8zRcLNgAh8hnbQUR3GBp3pH1PmeTZ8yjT+XhWQEIAQ
+vCdhSEtfxUGfs5A2WQdXpPDAtjiOU5esS8PJdNzndX5MS9mR2d2v4Gb6XwhRNfiCwk9MVsZtDrm
b9jyLOkWR6k1IJSxaue0ESBK932WCqkzsn+DJPkFTeq/rEAuWTfglK08LFOjWD2A7PE1cKR9V7Gs
GWLAPiwHCHB79ZSNtjqNXcZ/T3TaePIPD/4IAdBPkFfAFV+xsDLbcJo5+eC9mycsBhkz4FN0Qbkp
H4aNfV8Q6Gckwg2cjaItWd7HIYoQFL8IgraTS9ZFajltyM3vZ4R7FQ6osV6QzI4hJZDFHdGCyz8S
uzZotLAx+7APz8ePdEU2ssKI1FoUrXYhkRUu8Ko/OD9szT703OJKYyMI2Ught58mYIk8WTnWu9c6
nQLSBj3oI50YyM2yP7gDe3Cxjk/12gRkV/G8X0BYQZoxoX2sFz63XO3yXgmcUDD9mmDvJVuKtwDE
4HvNceiQQU2MYqIx6HRrkmGviKW69ZF4oZh/x0zSzUTNdSzKbaHjQpM3RmbiXSu7vYrMGaTLV4zF
chj0NF/CGbQg/j4RTVj9aSAiRJZmxs3BPzzs5Uhtqa++ETO81n9mPPqWlI+nriFW7mxWOlsGr4zj
98ljviVNYXdAjHcYHPRs/NI8MHDXE2TflDcywxf6kJ1m+NtqotL5h3dInOXvTVJ2jsqyEq0HooQ6
WS24lUfLq1TRMjRR8jKmLxQO+iAtnQjDZt0mCI3swJl56I/Tb5EdqowFFA6OHr/NVMjbh1GPeG0P
2ik7h8iI27ivfntTXzcJSEF95B22v8fY/uHV7ilFVkbYyiglCLaojJNtZAKkRMWAAKIV1wt5pn09
1Hj9evg8cBCviCOuJz11FVJWxPBsnll1mukfsWeteCbXF+g+4h0ShsWVGX4yiH203R8hW49YzRXk
J7jdL2j1NESJBPjjXzF2tQU2Z93NAoHomnEgEml8br02M94Av6bDegdTwbnpHDyFOUQ7b1dCrjpS
GK1bqusb7z/4OROLrD1JC0Y08Bdy7CuC1h499wg5YvI222ZiNPjA0OrxmXm4Y+VjJLnGYsru58m/
uflqNQrDiJJieOWEk/Y8nLX2tf1gKQ8Kj5e5lZztOaYn7zbNETJqZeZeQer0Z6MkhhllOtb+2NGj
ZqRpdG17VpPcv5N7p0kkzPPIWRC+MuScpGOi0s6CZZWkji7rMSlObQJi/VvEElSR3OGjICTKoWDR
vHidrlp7Nv6Gz+G2FgdR5GBOUp59R03HdrG7kAmeDpUgN/FqyHwdFuhWUofYvewxEppNitjVQEPW
sGXbQIuWdfhDT907twBfpvqZ+egHA4DCViHPjEs5B0XRP+WVKxvAysea/sVKFNL33fn/gEPkKXxZ
3Tfm4ENJSp8cV2DaKfrhKhQUovK4AmX5EtxkdlnHuvcf112bHqn8FNk/8FIyKtAGi+O9ZFmKx55b
7GGpHZYazpKd0sadh8kUGleUUPldF7bWozdavqNmLKmdV1X1yM55q7umHVN/2nplvAF/mODN24lf
YQ3QHJl8wR3Fvv1YyZMTvFpBPUOq44ZKEQPEdRPB/WZ6k72eWSzU3+DzGGQPYKrbv4azVLLgWX0M
hSy1mtwLkgm9wQkz4cze4cK1cbXGhI7qk/D5Is2uZ1rgdcbiiAlOnTI9C6YcrWlMnXvGIMz8wOfx
W3gFGu4xaQkogprcj1BkAwF3/TERYrc/hk8eNh4lg+u7yWp+1tIJL6y7tHvDxi9LBZFnpw5ZqmuI
52BVj7gft0fOUYNy0cm/hBTkOj4v2n5WheI5nmf92bTi3o6hGKPm+Yjp/Pkve6LSCTBEUbW99grm
Wzo8DL+pXAbPQ37Mw/AP3KtPqKcMURAprnDDTMexHa79pnK+Rrf25VfMymSWKzt89gA4CIMrgQTi
geGHrtsmzRXyDbWgIwqf2PQC6GA/FpEAk3leWzMBhrpmQA5hUUtnfRGC3fqdsDA/wCIphbFsFssP
G6iGibL29PXJLxhDVL/2BK5zW9rqg08ocAhPLqq2joVTRFn5xnPHJ6L5oMkAIT4vuv+ZcZLGGsXE
m23S2tNkduCg4ykfQU9Fa46RnBJB/uF7nrQTEnFNPNcN237l3YPb775lyjROBdB+MpO7D3vNaUU4
qWn8nsQJS61IBHX5QRABRjPZHMRsoGBRdqW3Sjm2FMWr7VEs8F4vGQ9Q9gCIjbMA3ZLRaQwdHJR3
+eSk6sbpCoOWIFe+yTPRoNp0L0myUDgMFQ+pRdp4KyqIpPOhcbXcvKOGt/andxfk15LY7FHRpiE3
7R2HPfF2GsCYLRyjPPptCn58LyY/zjnfdGtjxv21J4I2zXs03U3qiACZgln8c2FH8J7OLOHQHaNg
1KC7jAZHA3nVeXPOkT2IyZy8JdWBbeK5s/uGg5Izzd3q2V2/wYWwt+NrKN3TtVdSsANTugCzv4M4
RM5rH9vdcc+gtdSnwvFr0rlmj3PkGS3Cm7I2VRN++1x5qy85LXsdL1wuQZJJXfJxC92O5wCSK8xn
paNlVvY6ua7tyBuE7NXqSx1qMUDH+2o6O8LsILM86pCPdto1/JYpXNylfeuItYRiGPR8mOLMC3dI
MboAd3sRS4Eei4YyI+20DiK4G+8vqW9DnT+VShtlfOWAdldxKfjbPbFqQ4M8wYK6eYiVDRHwY4eD
vrHfaqJXEVoK6wy+/0iQWPyzbUTFEpdaRojRk9GhcKQXWCQEGaaDsXL1KwchPk6Uz7cm+4Sz4t8S
gWyWuGEBPUAUdVs8MAk6yvrNsPEmzQRkT7GSFSiG/cDDI/TpMEJU+rM4yWvytMoISkMPcVYWVZqy
rngXjf/Gftv6oxHZlueecvwSJixRroq6Zq1yE0REBIhMIL6OGaW902hDeV1OzncQSHihAr+gg/gW
5PFsI1Sjb+qqMNoAWS6Y63zTWQrf9vDzFbLYsaueDlkeBJpKxAP5exPygr0ayp+yuMzZL5TGY3fL
tJqsK2ACLfB2h1PN6AppAnrh+OZrklXwlyoMqvSmQCrJj0WyDz9pMTv204/fAaKPTuIn/r/lBDNV
yMi4A0KSXWUkYyfprP8rkYZovjJxwRSGl1bQJmaBuWvbPFS68XrpisrPPFmZsNDR3vtgjhlL0qfk
jEnSfxfCDmHA2tCgvUPIchctqZf2N3pyXQCFoiZUpnmAtEihwnQ/ysR8YmEwMcpEQ7TODjCBagsD
vzzqj6BtMioe2DUspWlcinepeROrJKmxihJ7lnfm7eQ6vDzAyV5uOi0h43Ie8xGhQvdKCWdmT7KY
Q7YlUpjN7UNe6iEVfei78u+AuYQjJrQQEsA6VJS24yjUUf1SUBd+HBLnDF/pczzXIJpHhlJ32Y9I
9+f3rmzYxfXIBVYtDgvVvg1vu/eAwhSmXqgH04L0RqAuI1RwLI+HS0Emq8+gsepunEVERsXyj8eB
faIpwhLzFqSvU9YxnW3y3cICW5ExqO3Ctn3trZwWtz1ibbqUIrwVOi59aKL7J+C6CCt6dhOQm4Tg
VBElzlE8G81LzBqoa9CEmTAC7hUsO9BZN9PHhanSovbVqznfb2M7cIItBpt0TEFTHkEymaYW4Ftz
IcPCanvWxdnodGuSMlee0CDEVl4T3qjkbEuj6F3PmNqcMXfDeOTTLOL1QbNZW6n3ocHpKWp924qu
dHCktWokYCKapcSaV57krWGEJou4cJcjNZLl/lFN/CleaRwFCvFY8CRKwmhhYGZ4far1p46zyxCk
s3D4ef6u83scuWtlDtngps5pDG5QpvZyAFTdOJ63OnAqWj25gH25rjdQZP73jP5ySyWvfUbLc0TM
meiNDW+E/PAVjk4/peHrDaCw3+ggbHpmFuIgtncYLaeTPlA93ufFrtEuXonsskMt5Y7ITXnbz1LT
ZH81j7wyF31x8CmDNiZQ4c5AMu4GvWjk9R7TRkrZCTjIO98w11+x7S9frmMKHYZxTnfrs7unWr5d
xblE3JsqNj00fsmX6FCnag/ERB5SQlsC3ANj5d9n+emfSUsmkgyzMgOEY0nAMgUdqByZhACGfjc3
Fp0J0jW3fEK9iWOUA/f6JMFfIzbNf/I7B9c+GU8lqdCAizlTduJlUgXgDoiBxiv2XQpLu+AzjH3+
iNtnsJj75LFRgiUCrwW0IigWMh3+PdqnLaIsppswJeM993y1pBJKzJOFtOBW+wpK562AL6XIGhye
onqt81BI4PsXM6ZzO4tOCee3O8VbbFqlhzVF+T7VVl96gu3L+rQLJtLKcYws7mx383Rz0t3Xvudc
oTgsiCTn2CuN575+aF9aD/8s9dvD1skoYIYOo5JM0mpikU+Rir+dy8BhRz85x3aOVDT5ARObI9E5
RhT2hoYHrYmoKn109IOk3H5qX5oVaIIKsXy2xVXSHpNcP6hQM/vw0GdcGNkNo8vonnwcJ86TeDZU
IQWOYEVmLTpZ6zoFpGWi4vay5ajOvil1jiaoOuXprSkb8NNrOseVZUgm519wlKb6QdGNfaLKj1xH
/EwMqELvr/lLuhwdSHSIsL48zl6APtLhTOa07ZFxldkTc6L/vvF38V4PKoQjfv2oTooA1hOOZVYE
F7lHFd/xmx5VhQAanlJAexyGk1wnfFDo2vFEHINTeI+RRaQvt+1d6QUnJcQ5U6QwoRhhdLGI6fSg
D9haYwkY1BdH7roHPv/UwhbskAkJV22C88yrA0XYx//gSf/W87GLLRicrcsjYUmjHqNLzdiO9KRC
vHaDZB7grkVYrt2MfAQ11IKlO3DYb+UeNaQYHDR9EOMli3KYE1ErvpIuw/wo//rAS/s3GSmYPFrN
7eV/dHcBbtgoFxekVZrCokx6Up7g2MzrW5bKZtB7RdEatu7UqYSuSG9BSyJ8RycqmAREThBrtEJ7
a/yMkZE80sRqat40/10Jrf7HtC+cfCDlix9LD4bFpsOMNR2RXTnlpS0o4Y9yt+b8bqVsXsF+nLZf
SmXcwOx7Qz2G5Tz0l3xeAJQdSaZxidDvs4c+BqYiaYbOBaUAMjDnMlTMKyn7UAwOPfZL86mRJPgJ
Bf3X280pZSwHTW9M7atk/+xuL03NBCPFmKmAQbPZYMAlRUablLQNCbEHuicK7C5vUNU4IqHn+flO
pRNDI7eXt64BP67ZqrZMJuyXT9mu6utAt8M+4Iu5Qp9uE+HQIDTgQ1IwPT8cUgfR+7HkWzkzvd4w
gfEeZsWJt0BXp7ibBar+FG2YK72/4nDwMVnwUI/ic11LPeaWNOTLfcIFwvoXd95sFWBPrAWhaxzT
dcdCwngh/wP/EFxoTvssBxgqbtWE+AKLpEt4G74yVLqwZrFP9j66I32bJcv3eS3RCfru6iQbHArc
65gFF7mDxeFdgtIoZ7yE8sqCLypfDxV0o94Mhr99LujflBQo+XD28qZ54L3km9xe8wstCJdp6N4L
fUW1YHUNYr9ZJxz/2M4x0e395/YSyOVA1HLax5wH5AzYY2zZZOFCvFoVBAl/mUB89XI3r0d77NAP
SWQFLIL+I5HaHvVG80hQ82rLKjVzzwa1SUEeNA8oYK0OykEnFlv5oEb87Q3RtW7VcwnQ20j1/Xa/
JdzcyuZAWggP0rQz7E3BvyK1iO5R5L4MuwFCssSzXmpL9fPp9gGT+53RqtS3aCD9ji8sben1DomK
Fi+xB57CHZFOnOqSWwG6iaV/96XVhY0Y1URScK8fWYUBcYL8OM/iwX9Yfti2PnWro0stNtgHD0PA
+NkVPOBJrQBY6/wt8j4IsKOcAB0va6t3eNI1fdSV+/YPIuQiBoqdPHBU/f8ztmjukQ456SVzmvbH
j8w6i5jS56kluEg0H7FX0ObeDjVYZGff7p7BMG2dg2lugVv9QgwCd84hzacrWq9LHDM10YIMktyh
rAfMk3mw1LNPrNZHvSvjhkEa7CI2JZzxK7q+AT9wG3961LIvx6MDwc8S9StKzn7n1B30ZIUlIpRj
KGO7RGUWj0EqiVxjkVIMWTSNDhUUF6eMqAUp5ZuyaZQga+PKGh7QPlg+XWwVyJ/mhmdNK1lQu96B
HDRGC6wNCaKs95/85njSqgJwf4C66SmOL/t1b0iy2gB+15+KKkrloTvNoWT2AY7qJLqMAPQk6yuz
uN0CxUxFtrrBSzv4qUOq/YUVoXl8NOBGdrtl9DUhTQKAIdjlMwuYrqjmfBjAzg0lPqF1eEvco9fu
S/0eGakxBGZ3xLNjUpcWPi2J0e9lgg3O1pJkZRHVS2+L6ea+ozg8YCNmXf95aNS7ZxPimoFOH5JQ
Zxby8rRyzsWBsR70urLyvLtdhk4n1QvEMmIqfXHxeyO9k0ANChndzlSsDSaJ4kXz4yl9I2CkrcVE
YZOWE7d1xsYTVoaru0sDVy2BwZSehtMZKrsfDCP71N1vt4AmRCi3WBD/h1QCb8G5k6pPwHEIdNQd
zlvAryo3ej0p0rBolMrTH2xy4sqC4HrJkR86XLtmi2UeZjN1dP6OmE4H8UT0LCXW70sSoEMB4jkK
4ztRc6tqSl5Umks3ApPWXoSVxYWCh4R4tZKA5CkXa2TQWX4Wx1KRrvPOYRIutMTlJm/52++npmpP
QtGsTvnhoKqGf5kgGfJTFj8PJpghDvmPaR0N5VqkOfN8krIFs8Zh4x4NSkLs6JQc2mgZMx+nWyvj
WgmNj8756NSrE3uf7+qDM8OUfqpUY40iYx+RdHZfJ755qle+1o5IZXMgbtLdhcF1pGs8JW3iUluL
EZLVRRcJ9//qGKWdwLNC/QhUwQZpgkmV9keo8YVpZJbH+IYYL4ZGNbt/gdx0rjLVFvNGfvZ3ACtU
jzRTELnNw1+BT1zkj0G/vypVL7/o8hUqTO+vHrXkR7qxcNb/ReMa1E3jXK3MI4VUY00st3ukoAnH
XRrecIotqUbGXWQod2f1wzFVzTidB+H4DYhjGgqAJLgTBUZZ0HYUGCDo+T/KF3SfrFezBqaWT0dt
J/hbZXLSe7THCW2hN/dgf8JtfxJdOOxtnmyBpLz2X2M9NBXMnXZbzAEjJxw2apJi2FtkBgPWhLxp
5IE1zAOsWM9GMk5RR+aD9JOMsvV/sXCzL9fO8l854rKpIqIwFhyNvv5PxbQA90CJvDtHecsrZ43S
ghU/dryJd1+c1A+IHJNyax7IjODihF+MyL9cYSq7zcRopdGXezV0xL6nikKH9PEWJz9KvPyPonsY
b+93e9//oCCi+/eafCmA72jxA1fgBNc/8lglp25raUn+Ko074Xbw5nX1UFENHYLIPj8F5eFp4Gxy
2ZmM+Kt9ys424V7XXuaGN+HiZWD4GYQmN2UxsTO0kKPNp5zG+WvoXMGr38qK2ROf7e1nJfjOVmCt
Te1seEQVpYoDJfjZq6Vx+uDI0ParwpmrZNeUCN8yxrjLb1ViG4RbxLlcuWvg22aCgPtYxxvWUkCO
WJTcjYVwkfLbxXdqBgzO73SEYPJzWQWni/yxWDUtEYA71vmIegW09JfegNFgXdc1yzJeGcNj7Vn8
sVz5HNkl1cpwYBBdWKbv6AQUUkDYEWNL1J4gMScierspRJDwfuIeA4a7RYLiobdVp9PF45Tp3LNW
pV0s1D7v/mVzfadtBe/vvEe0dRkglzXFSTrbsMNK6G56Ef+0ARZ/n+9/CYJ7mHd3JkoAsrGBm1wE
zKnxcVV4ag+pEl2f9GwautTb2sg1X/kZ5lq/YN0L1iKHoxh41RY1ak2H+4F9LdCk1jeXPcBSmuQL
eqiiX2CoF2fgEQJmz2EGm8lFRaoAU6ZZMajcpNenyvJdt43yttv067RFMt3tL5/gcrmq69n4ZoDX
4dSgPQV/5njL0BDQnM5boqH2NMlfTZzRr2lUrPsSZfYNDcTtUjfxqeDKQ4jKdzqs+I/ANI8bAWoG
9mTXqqDtCdCJCgjgaijGJfiQ7YLT2yvf0GK2+5Vi7J0a9aMwkbxzdmt+cKJVSXP1H4CEzBZHXx+R
XieYFG9A7EwHWib2r+wzvgHt3umC5kf56qdXCG9BoZJuCyiCll9a6WmKcPZcS8Tdng/7Tt2YfjZz
ET2xd2Qog5ENa16fK33rPQKGOT+S4lW/ThezKAbpgtx5QkMVHNVQ8TdMGTlq3qoPSzrRASjnVgDU
N0gMTFQaSmB6xORIOGRxcs7RpZCH1iTkyquYnLmfCzYijI6ryQw5IGqKHo4YR/DasbWQYKUCNSS2
B3uRK74ZoCoYxL+r1UXKbwW4AW5KlVHMelby2BsPjkKOQNuxOBfrwIIlRmWkMtJ26zg6nizxlMEp
SziUVCjcgEojVG4yvoUxxoIpkHjuyuOEZcBx1KMn1m1CVFWxNtC7X+Uef3O8/Z3bvxr+bq86w167
Q6T1i4Jf9kBCAB3E8b4Kg/A0DqRh3DbFX6Ez2vdn8eh4p6Ucs3u0phBQY3HZcdwrFw2m1qpcqam/
q/rJyN5oQ4WPKIj6o1hukDkwjUD3XJRSZQurqWKGsxX0QVhPHstxJz2ZO5xzllV4yUG3KNkhCA1z
5j/QzgWjDyq8F7qJI9kxzADZ+jkW39FMOz+SkEymkVm16752fI4B90axGXtU4YnKgbh924NXQgaY
nlWqwQhBC/qEVFPMFYm46F3IAFHF6hLiy6T3qyck3ucZMSq4jqazN7S+8gkTVX9+oWT3Hsqg90fu
8LfUwFYvLYkTwNjBSbkmHBlyh+q8RSlQGulqZiERTwB/1Kl3Cf7GRkssVmWvttAMIYLO6KXlqFPs
A56FUYWPSOBzab2OyaFHdpjp1JDlwhLFoE3OWKbZg/sQxA9R84zcfOHpPLoL/cboJj3CqRCo8QUB
BtquaE8+wBL2UO6zhoQLTrsi8Y1xet/dc9bYTTYyPepm9JsbUiDpk1PP7wyxIKZVQKdikkXj3Vdi
tAurXJbOyVcZCijmBh3ZkEJADKvfzLpNjfrAFYM0P9hRDERgh+37Hbm/gEnL+H4BSW/0bjIB/Ou+
4j4boonHn83MBX4j5OnfZHIX7Rfk9/GdATHgkqfyWcsSM0bwqSvEpvXue7EoHzRxM7E6Pgow6/mF
Y50S/BSrAKL0TgsqMFu++ObvEBP9JqzCZbbi1Nzmjr7K1Q0pmMzdcnDu5mPiBimS3d2FtKaiI2Z3
/p9GeEj4FYiWfXnNoeXAdPqi601ykBkZBCz+puGDKN1L0jLRI7VbOf0+6FcY3j+/onVc+KNHnzr1
qfNt4IaB067QSVyo8dk4yK1LMYF/nKb4aHo2Eypz4acQ5Q7e/emCiyMBDieIt+DSOJXy7hyOGxNE
n9W777hgSrSYWjcUzSAs+EkrQZJtQSHEjh6/e9rplHlkUD96XqQToXGDUrS3kxEdziA7x8JhwEF8
eTHSamTU8QbzU3DyOBuuNDhp3XWxi6IEA6Gz7nd2gzAj4vDWJWK4jFWyWpOLT0ppG+zKNi5QbPXL
/wNmmxrQ1GqX+nRlAAaUkcvNzeG/yDTxiMbBq45w0DPAeGPNc0h6JgMtPKx101gn8QLQhiajIyxV
d0+5D3ymc2NmlO7cqewwaHi29o9qMEOWjnXSxJvz3CMIZut6uVjko3eyOpHhNziDhtQ6CMWrX6EE
HhGlNr/lu1Z879j08tJMLtDzDK286oM4Ubog9EAcYSSFfbZy6ZaZ2uUbKK9Wm4DSSKpo8aQMqTQT
sU8Da04EyUbU7DSbpKNyWMoDPc2rDCD8g7NgxF8/z6myZojimIPhgr92YuWtWrpngMNilu9qqkTg
huBG7fdqQj7Pjw9Bo/BOOvOP15ZWfLnsRYoqF6RrxU5VNrpFcmJKQOnHoqKCKZ80Ji0rvXeUdKg4
FQfH1POpAzETtpWl1c92s+Jw8YkVomy+W8+c3I3hV3rytMvoyICvBlGLC49nGsCGySuLPAYcRMcV
uHEATi14CVWtGCkyEptIRIFU0kc0sJGopBz6w0X7Brjn8OU/PSRVIErWch1TmfZ/Vwi9e1HqDi8c
tjtNmz4h4yKN7sdMoOQ9v2Tq0iz43F9Zg+2PraeS57VLx68pryur7ElfEo3oAmOY3j5AnU/P/AHe
krfDxY4Qi6JM8yCpBIYVd2lT+kl/BW8YKuGJ40vU4x2Wy4bm9xXs/gUO/xLZ1Yf0XbUZE2PiyXQm
3sno2oENo0UbH5tjfWzDqRiSHVERA3wQWplGUK+mmAQmwP6nRv3/gEF9RP8YwiQHdsOq+Eug1dXd
vx6AdoT4NEB9q6eBKvN0NkuTF/JQ7QjWd/5If99qZGxvLrrETgYBBYcBI29hzd20V/PNvoAaPy2C
NaFcdJBCA2qmeABxkkMD5xcr7p1zvUfjmR+MJXE+wyvWRS4etJQPbZHpLqwdrhOK3jQgZIMWjVuh
TTV8gXWOl1Wciok587ru8/MjTb1gZtNudKWU1ZhnBD9rkh9GW9uox0ncyJue2hujMSecKstwlF6M
ehhZcviV4yq+bvMSOYRk/83msSTsjFxbQXvOyLDJA1wg2V7K3zNViqPEgX57YHAp7cIsZv6K3M/7
zyJ9SAuvYIltzBVVpeGcAiPg68LRedBhv0t9aCKPngYkmmXbShA63YJRkBgGPPH5jZV7fc2MDqXC
CR/PsX5Sji04dFBqcVT/2wS4d11bIw85Tvwse92U7mmVSj9RimaBEJBQwxu36yDFdU+BM7oo8/Re
vmS9NzRWramaxLWC4+b+pQf6ftLIX5L6iTc5AiPmAGR5fjOngPPa+VouBpqd+XQ6i8LErtOQaKZC
bwnjDsMJQqXp2npScy4A3lGVpH9CQQNUm2Osw3NLg4izhr0e+ORvPOxnELScznwOe6eI+lB5SW2t
imAEvkzGE1KOdLKnarsN0bIQZgFRhGnf1I94GOnhg2iiy2hx2FhCMLnXwdZl07cvMZ/3fcvMrwOW
A4JiJMc8T49WOZXQGQzT0fnReD9JYrzYCSB/ds8Xt/jLy6MqLxZ/FmAXtsPsU5UJYvEDgD5CR96x
Qqypq52nghFarLKO84VfH5hkEQIwopd+KX6NQqqOW6rBcv0Ak1FNQXQzX+8x4nrZTQf+/HtTFePg
V7z0roiRUUTISwA1PPUwSUxH+lCHruS7MzyG+EEKCA9LnwrmfV29U2iFhBiIs7oaN4LNGZT6W1Gn
LI8LLnwmqyemZ86SKWXLd3urdR+ZiSqJ4HxnPPTbxiAngDIEYNNhuwPgXktyufGPn5r2rIkMl6Hr
Ze5XdFQCVRfnghdCrfygCvvReJY/Yqy+tWd6cJeCmQ+sXzzJTQiMEtxvzCM9QbGrPnYTU0ZwXYTE
dsbxAlx8OHM7Tq3BXgcdNzGgpE5CPb6rC8Sxc/Vlp/SunE/8fgS+pJXz3LRXpmtcu3XBHUm3AIFD
AM8+lllWxuPqNGKvjY6/qo+MUpdW7+MGCngfwz7D9Ay8uPGeCKqPVWqJmXKS9gtKbjX8+epg4pwv
K1pSXx15DNUrwj9yIblve3/khU2e/wxlQQ5CowmLrrjnOVOdUMTov2yHYuETd2k8ug1U+/flfXoj
0ZPbTaW69By03RmkMICBkXzAzvtFY2ZIe0QBH3CoVJQcE5RkZ2U7tAAWCE78LNgnpvruSiSt6m8Z
lT9X6/IInqEB1ztao5FiLw1kdQGctEbkHxRrvmXAcV5tmVRVy7uNWaUcyiUEnTIcqLw4TK5DVnK6
Jz2AytLhxSPZISQd5Yv8thLqBM5WGGhVXTPuUWoTyo9a4fu97CCG50gzKAUEbBjq3ff8utFNBapu
J/zdyzHtkVF2hvS4q5agbrcUp2go7Xou6ZqV0EMWQym1asB9RIgZNmfaXTpboXvJpSHj9H+e0WYN
kyZdAJ1J53E/3cwpVT2Nw4HGi7rD+pSEsdto5Q3tNBKc/CfoHvetTA7e94r+gmnt+sszUymMJitZ
dywaTCpq47/aWqPahecutpyHMnLlzvZUMk9WtPN7A+iL2eBRvMdDXhTKQRj/a9Vm+3hEVuZdhbiq
KWf3BbVw3rYJZ+yw45ZhE3q3eDurIyL/1UZ1u2K7z6rW1jYSBG+7UhLTP8i97B1p0J+3eIfX4Ez9
Loqf7RtvSOwvoSKOAOzsvlmFUmyYLwvDIPeEtKVdhvTGlZn8h1Bine+AKc+C143UElWDavd9fdQe
6Gl547lR9JP8XWs4Jkd6qwStJaWgTcPw/+hAbEuJKr16fz8t6djvnkIiF5owWgGl2+Y6ErMTALAj
SwUJcP/QaYgB9D2l5BrLdkD3gXW9Ajif7rsTNn8o791K96JVcllgl2n3etO6Rwxlh1GdQEGOSsWh
KbRL2rapbujQreCTxXGI75D3zyWdlsoKvpz4TyROsB9Yrfm0A1vxiT8GNfgfgSHa0hbzL4OflT4f
t6JFxdaNt57DJ4W4MC4yp4RFVHJ0taXnlpxO+p9Xft7mmbIAsCcpCpJWk84hoHqayXCVj7XTwz9w
ZXLhW6hwd+OocDtjrqedUPXFRIpq3xRb1dAEyp9AC/o+3b25nRF3R9heIfLgrYUBCfoCIFK7a/Wi
CnUm8qixr6xsNk7H07SeXjBiUFrn1Y6KS8PB8k3aIph45h3xKDIrwE1wg9JCLIW2KUKLRvu/Pqpk
RnHMq3NIUzJk3szP7xxy11SkgvZpWBcrPujRDUHpNZBPAIyRQ5pMFSajPkhiSasygNJndFiWHmMR
DGgiHv2N5ZiQF21G4P3iaqA3UENlu4wNFJmIgEysBrIdhZFxbhz+uHqZPbEkRwDMsr5DaTyKgknl
VtC0gNXdf320Mr7F2ACFsPQKmK7RWnDSO7VXM1OSszFdhnW968RhhLNSKiv6thaig+SRhaR9PMrG
rV9Aso/UGB3rFbQsCw0OFrDaU2sBwH1ttqOLxjRMtXsUakJ/pdY94IcceGfLJu6OUSIPGQ9Vxwcy
zcnp+x3Ps7XbN4ciM5ImowT/J/DPV0j2Kbiz1aSXOMLImINzZ23eqRX3CpwqyB9Wx03vf3FWpnJI
UtAh+7us/PKkzNhVC2gE+Y8x+78DjtxSz2x0tKV66eniFOQO6oQT3s3LuYy/H94etyomPBmt6XJg
MutQiLeWJUUILgwZhlFtVwiXXln18nWP5UyaO/Dc+QU/qNcQW81r0f/SZZH2h2rJGyrIpR4c0XQ7
XJEHu1JZW4+A93J9GGVRBBqW505eEgjMgXN57pSj34RAxckod4SDTf2jHCyENVIxzpPQgSqqREqU
d5z8QdpbL4UeZYn2TwUbytP2TeBeo9aLbXun8g65tH6JaXbPnHXhdf2pAEwDqB5Dpm0FlKnEvzpy
4O0fkZ0FLmEwzwLllUtbUktiP8wuKl/8+ap0dFXPIEdpAfTsT57kPtM6+vQVdtj5xlGkbacaePBm
SNO+LGme4m52ioG7jek8/kGgf2VKOddhMZ609wQLby82O+u7MHmalc3LJNyMs1pomAcfRLDnuIOq
85WxjfH3IKQBJwPEoknQI4irLEtRxmf2pA4ioLxDjt6NXpicIbIcKOPRmOSk34jUuXuXEs7UCVZL
92DI8SIVNUA5bWvbYC1s4MCDqjHBbzlL3F+m2955gNlpd98Aqsj5vx1BBvlwoPD0l2ZI7EaFnWQQ
Sxuu7WsvGxrp98NwOpjxu+7aWDsJtJVKI6J6XQ7ugr7kw4roY7RX4XdgUR/5yhus71N07RQ+99B2
ExwVsd56zerzXfTbHtNYlqcXVjNR7oeiPycaUk1rXJi4ZJ6F6Ejh+ywin6sY23Lf5uUPFRiP37wv
pqtQNo0veF1BAQGMNGRL8+k/7Nyb3hSveYjq+Qy4uezygq5oCoZUn/ZanPb1QR9USVjUGVdRSoFb
QQK6SrRmjmjp+JmO8ZhwnHEjYnDyDYbVuY4JIrR6Vtbya1+Kay51NjX/xjANmsWGCdPU2HTvg8sZ
B7GIMJzNh4uGVPbnE9IuHzQrgVy02LaUXPW8izD2wm1YRGCVT6BgoCu5/+p9sc6xcnDa4G4n93my
NVDgqHumN7whauL4II8icowd6Ihu5xT+X1Xl5JmoYTDIH8XVBh0DSdVR5eQCTVkOsqP1XBWKQqbc
8pvjYfxtjBAG2lja/UF1udSNAPFPEjCGgiBJ9LMb4YJ8p1IE6nZf/DUQKvGk3qud+LRu7k+uNHB3
BCbiD8sl0KSbeEBLVayvK8+rWcrq8OOyFGpFcm5hiAW5SCHHrSrkHtbkwkYAvK0N5s/W/5u3ZjKv
Df/PA40TUaFNCKC5YSbN6sgkeaSiGD3XFfwQRq7KeLz7OecqMv5iOQBmiHOLoBzdTCbFH0VJyUMk
KnYl2DBOhchTKTtgmu+wuEoC6afLRET7QcYk7kyGMBW3dffYTL2cpRT2VRRa4fhVb2JU3eB3FUvX
FcSHL9V53AlCCA3Ob5svBdZOOStwgcubMZwjMIUi820OMlmTxbtafYSUUm073RbIUa9h7N7AG/Xu
umYZ8MYr658W10YhTMJHHUnBAC2drjBR4vTG23hzBMxCrAb2TCHurgHyxl9PxqXKWCxSoNoE4yTU
aCcDGGQULAQZThRorcuO8dgMgGjdjAvFAEggeAigHVqu7NjpxENlhIUO0nK221DbSMsAIUKqXpbi
KHGrHy4zsOdVLfR1MPDRWIASe3khH543Jsz1RcziBPY/7aoxgGqSu0qtvRMpsvv/sC1o+gFzig16
D7+imW/Ty2OAG6zGVCSMNRez8rkATIWMXh7xq+4RDILOBHysJ0r1FfTnZ31v0uxTFbtbvjljkIqC
xznHqjbn1KnqgLRXLc8/IYevje5deuERkORSuTDEbHUBQPPODciBmYCx3U2eVEyNKovRnyA2e0/f
Q+zMRogNhVjmDN4+2FNpFJTnnboQIAu0mDiVj7k++aR7Sqfh9gnAetx2CT5IE25PcdiWa191lebz
LTqdxLRoSxOm3EVy5iKS4c+xJlFROpnzNGyzewezD1u/Q2dNoQJ6Yi+dCO91jXn6KHhfYJTWWQZO
wcjRtyhz3BG4OS76bpPqrTk01yj+Zc4CAp2eWyFgG0BsPOmDHkxyK46buSF7KYlBRNrocQx3Nwyj
m5FZXWc3iBfqLR78FNYYnqsy4uPeinptyj1UPXNanol/fqLOV5Vt+qnOtIl6d0m5XgAJtcYrUtjj
7onL/P25rmAf31YMtcJ4L4suSBexIT2jQjhUhacyAeiXEqVKQcvn11JDtgADRWBVN8CFWOs/dgkz
gmrc70N6k9/kUmdD61TDjnDR8kMoINGJngq7zoi1wImcp0VvAC3UYEagsHulqCK+vbUnhhkHUKNP
C514dNf/WBYo6uxSkvcH96a1rRsQtekSR/F+APf5oG6DVcviKhbk2eiUghwJeiSZjDuKG5VZtyuu
Now1VdEEEaXT/x2Devd/gLm9oLSwTaln1S4fEE5ydu2kENWGoL3F4kpnX+/BiEOSiuOyak/JINDU
W35welxhHqqDvGjela4wDZyDGUCOphCvgsmTWG9W+2X3tRnyHf1+wKClT9/z081ZeYYdK21/ZhR6
hvJAuMbGOtcr/PWAglwd/rbOr8Nmfp9D0HfBsmaxLbjK9j8KSRlOn1cv/BZIcCioJzlGLitjlkgg
UN5QmILQiQTdWZJxj5sfDSJo2wcj1XRIEhRdnhZUm5Z6Qrl1cyZX6z9Vd0dehYj38kD6ZHrCaDgS
bFUgLjIvbzZ8zR9kwX30G5YI3gNGtqFTlwv9XPpYGeqaYbTr5YXUTrtnLXOkLtR2t9YOrpN50kp7
ZlA+ep+yfj/ACdL8q3tdHuuS2+u+zfVYYYlcKPs/bCEXxnTMpfQK+6DXWiwIxHcr6aR9VLPx0r+/
/Z/uzRjbWFwpLpALfA2KbcLyBRiu3bL66JyKXu8Qvl+sRgG8WmGPMhaJVMmSNuzmD49x07rk5ovM
bXMeskmB5DRMum/YfimXXtv/+iQcnqKSzCsQUfaRRSQwie9dF54N7hqh/8gnSXYj6Lsdjs5CFkSq
SO9gpUmyiMzyiEdSg6EyHor0T5fHLa6N9ToBby7rTNcWc967L9Ix6FD/nv2eFWelhTf0qZ5J9xQ9
DrIeLbOic3xT6UTxHF0l24sHQ4OY34nNMe4DwRyi3uhMalqVURAinLMWMGLB3ZRmHVRO1ZDnC1+T
tKXgvRFbB4KNVKgwL3eLijIzVmRFoU71RILGWKTbX7tcUVc1d5y72mTWcSnus+MJaw5pCIZ3Oc2K
rVV0bKpk/vtxkftUK80zRjkQLmCVFLbznktgoH9wg19MZwMee2LFrKfdfIm6xzOXWyxmIOdjfg5z
/TlF8DdgjkRDj3kIcTOYZ0Lz30bvnhzl0eupfg+7/cg1z/7hffiB+Gw/Qv28GAoiFH301IXfFHYk
ZuXY6cq7b+R8QgovA53AGFYYAlSssRxYO8QYvvL681lXHB5XCToTvbo2gg6Oys20jZWnIcESTAtC
LDD0RnNOiLSpEwESNZU/6qxpA10Htf/j1UbVP4pNN2M3e8zfCCJqhKZOC/6JXuqn6IQ9Aib1C40p
hMlsA7H03y5DloK8jyZTKU6eQ8lOpjc7P3ilhQ/ik+4+bTTRHAnUyijmmaP5euOom1PNubOMvBC+
rdOcI2uiuEBIld4uPm5BO/TlkeTmXl6vhAeQJc66wKxA7OlbjyodIA8obyCxbO7+iWeMAibjzdoO
FaCeJEKfbxJdl3FezMpJ+/UGgOiOLgwz99D5dvgraXM30Gm/6386HVL7irnhe3M+qA4hrgcC8s/j
rPFoNo9T5Ns/93m4qnLWT4/KpeXEwEru87XnUI74qAzKwTZUlbP83NcLDzgXTxuVP4uzZyA1SLwU
KkS2BDwC5qB7APnwp7SYpagw8HhvTCFSozMkmcPEB2N7xQSf9N4l9BG/Lfzb0hpb4UDvysNtPCtV
FBMWIovSeHJu6UwTQ9PPO/8bdRM3NHXlOM/tOum/9sXXyW/b9jwP0na6vnKX8yVc9QRt85995nHj
itkfkr0ylnH9IfmPH47ZIKeWteiTo1nRLXVOK9/WJCpNJqGd6gb0ESzzRp2JUeRJ9AF/onYp4PzX
I8sbqsQcDi1mPfaYQCmk7kpKrcy7gsNB6icifdaFz0a7/2fGPNiQvw49CNZNVJrwps4M4/k18OEX
OW+ijXSGUDDyCCa4d+byT5RIoowJJStVhjeKX+zPutr0yA8lNMlHldkxTC7MYYVYYh1fmSk9NoJX
jqOfH8rJXVkgcxuj4mhp3KU7FPN1zZ5Zt8z34v3zSPf8LdCjE3Dt7cjlkdITW5Sj6vrqNlUk6gqz
thY2RLqQYyj/CGvPChGGCVcdCklEAQco6XmFV3bL0SCd8rOK7btrFh7a1Dvo/ds+0iAgtwc7LCga
8crSvC1w+xFXhF+zUJQGTGID0g94/eWZxEDp339eTJ9z3U5aMbROJq3zy7bslDCAFQren/CmGw1h
8PHf6rc4hhKWAVxyU8w5eGTXGMs1ovrBwrW8ViAYQZUyFpCzfdDDLYyr2kOM1fVD1jGPcaL/qlAT
CttYOECZyJ2CEjDmNOFX3B3I/JXYHv/nX1tHsP8mMedukGUpmizpvrVJdguoVBGJQh5gZt6+qKeA
o412dUs7aVAnDCRcovdjtB2ogTS7gleTPQrNlhLc3enkLGblQFgq8pMQwB6fkvrbqzpaLEcx8wwk
izFodXMPowXIeOe+tpWQbhTYsQyDAlwza4ApgXPKxQjmNrAsgm7TFW/bV/Ht7zjN8xXjYLiaQfBb
5Zj11/IoDJQ9m47DJOxo3XprzbqYNyIcAaqnwYW62J+/foHAcJvhJTSsO4D1NBwMaxwdFZoNjTCv
ikqliD/pp4GwoWTz0eaGNfK83IZNWLrW1dlM+MG14Jq2kB7uyOHDbu4puwilBm4WCw/cPPjcLt0/
HiP2yUXb5mL4k5EVFIZsC1CnleW6hk3XxQJ0uVnHL18sh4KMNxbvc0xxnm3WMmJWeCbRNv1H9/z6
6s8HtLiywMPp1heTAdRenzY32VxKtynzZUaIcQcQdCgbE6dSvTllEYuOLRrsze3jmP3YO8yB8NEc
BlBOQb8+3LL5LVUSD0vLwFbXZhjY/SIZoVqAWsjPhuPYrUHP8vQPwdYlBxS9eK9519yf+RQqWRz8
Y1U2+EZ6QN8Ev+gFx23DJ9j4TRZql6daCF0XTcbxeDEgQsWus4EqEZu1zgshaPw9MUrKjpsVoIwf
0A/eHlsPk8A/xxxahZwK7J6coE/1KAstKBYePlwidXU3SLpS44m2lqBX0dffvkeAnHstGyoy1nPb
ZKSIpA3+LAqru95U81Iq8supIz/V43t5c+H6YU05baMGiWpchcDUku0TKon/m9pdwh1ixtWkX2Bo
Iw1sMFdqfq+76+FJyR0pmQAog0BUlqD54nUcGWLOndI/R7Xc5/MIo5T8tWZ2OaVNX1NrkeeFgYIQ
G8Blsw8xOJkEq9YobBI5J50gWm0ET5wAx//uSLhNcGgbx+edxKKRCHlbKvKR4jxboU8M1dZo9hSb
4EiUd+qOpO+lO8AW+DN79WJN2X+cIc6pna7jRKpu3aj8C+0HnL6+RT1zAGmJBeCQS8hyoJYSHu8R
Kj3qIksfuBMEK4/9EQ1NjKR4e0ICtA7GQNmBWZ3vf4p8Dyu2prqM7A1c50ZrsByNrn3EDbgVnDwt
7Pl/Jnf0nKMfcMHLPEP9XO5KrU7pSEsYEA1v6H1pCIRsE+8FPJF9K6fnvToffGSjC8i5EM6pn26+
a/ym4ebenBSe27SggKsAmlsSI4KpNLPjIihQ5NofPsuGwfjCCeRAJ1Tx3cLKhyZyg/sriZzlnDum
F2yrATBiWM/m9Tt7B26+94f3JqGZl/2sd6g8BYLxua89TAKZwD0jPtfGQ05U246P97M5sYs47nwu
WdJ+lGrcQOdLoFRVYd+mdJBcKeHhT4nbhtGXLuBN7y5lrCBsJpXpOCvCNBGSVTraQncGbQ3aXazZ
OrZteWyM+yAonwxQFp2GIEbS44fPrsTFgjI0k27URSYz3P6TETj7T81NQp9rHWC1yWiXhKc7jmye
W5odsM/r9xoq6w0wfv5iLWCQP7fnFxCxJQcTnFyeN0jahgCgqlod/df8MCg8SVlqm6K1yPc8XfuZ
iL87ymW4gGNO8nCmOZh0JZn7kimwr7DBv9Qvgh6AserJ0LEB+gCcp9qlopo7kMlQ4wgN6ZxrCcdq
7qK/xaPJrRv8qZkEj/B/dL+Jggo2/1AqIUWnfmeEeHX93/uq0/qKnkG6R6mGrUCDY/gcnvAyOw9T
QiU54IsFmTgFkh2v9XMLaUS2rl9YXouDRVo0AZj1/3ORMQ2uEklDxeb7fmKW9yDNqjG4AGBne1nf
vVb6mwZeshmQPvaF/to35PAcXKtOuDxy99EFhHdvsFcphip9/q4E0MKVz+SmEqmeymOvoAOTcC6q
BOHqu3dR+p3atjrDqU9vbfJ+TWBaSpn2KiusMGf7B3kbjyB5v5T1SoLXOhLLqBrkSDTaKlVy1O/7
I4RkwnvldnwpE8z2lB0zfwjoiDCdXuidpoZB1Zwx1EZlRoukPXAavN+kddTZ1n/rE6H1HLQXBrp5
6iI4J1yR7kknw7U/Z8GL7rf7p7v4/vRaZziOdadGi0pvur3n5kHbvDyk3ecFvxiMycNQG3/VTB13
aA8q707H0W2Yo0EhhCnQcQ5GBibjWkKyDCSMkUOwymi10UrkXBgEy3qWyYuBxDuCnLGamUAapsLX
zt9ugVyw2JHD3u/oofB3rAD+NDhbGaoyrG+RPVuL7nxf8lqH0pot9ecG3VupJshrdj5iRDhs69aN
gnHVyZZlNUN5JIfsdDTeQNPjQ5eePJ4jPxN3Wu+BvHkEb3SyMAadJy2WeDuFfLnk1LOqL8eXQqg8
o5zrMOPPel7xDGMU+HsYYB+LDQpRIGoCirsJIAXVqBfgKsslzHai2D7NOtNVg8SvWJNv9hxZJlnA
6t3ZjZf0SITyftqxN1m7NJDWGS+5ukdsmud1S6s1TbKcl3uWFm+8KV1PeqNeHV9xiApB94sTyLnV
CBTFVc458NoMRGU0rEojiPGfSm5NZrlkQxGZ7NXboXnV4OMWd0PHG+YBzIgUYg1lCc1pRacbiNn4
NYalD3ybadNgMGIw9Qyh753bzkpKk4sVr61t/KA/6FQ6kv95YGcv7XabzXcdCX2J7dpdALyn79Xi
8TPQQX3QZNPbsyaUGW5JH4EOUZ6bYwjlNafJjh1hkH0h3xULbtvCPj9bZJqBpUvoOpPhmrdJZunE
aKa9UeMyaov4A4CKNRZTiJKxfohu8WQcyF48Tsr4pRCqFpMwJKCpBifgMj0NQ7GLG6NaoolMeCu5
qy1SLfMOvyFP8Ck04S/yunD2hb6uOyb/CGAvBJ7TSqqx2f7Ocrr4UV7RoqyDuh0wAJKelm07+P8I
hKRxeTSb+RYMzouDmdGLuOSgei9bw6K/vC64ZYXpzIEWvgEOpeOb6K6fOazENffiGKdjudYbarim
v7hSU78OALX15lfFR8kb1XGNIWNnJl+GAm5DF3/ONwsI2/UnLJfE6beTP1LSJ5E66SIfFVzYP3e3
dmtoPpE8qsZFBDpF8b17Zb4dEF9O2A2QUtM+a6ZIMv3BArwy/1gE3L/csuNHvZhJH2GQuZFRt6aE
8LRNDaWL4YW8NWBG5Ak/MX5Oppf7cwKestSPSdqt+sufDoGEkO93LY9707KnRVNVL2SOWPWh1nCj
dHr9ihVechPzEN5VXL6mUiS9X7cYXWr8pfclRt+UEcDDo2PEao5nCrZlOagSX3wsQ0tD4KAulpWW
Phn7nL/0SIQke0RLVSwiM+/143ldT8a7HDEQwZI5jtmszFz+nHhOgpcJcAlpVTwP+9N4+hvfE4fZ
Gao8XLd8sSL9a6g9JoMoYIIu9QSqEmPwPEi6lKwytb26GAVPA3TmLeZ/sFDkNeNHWdFmA4nSoVY0
Q21W7wOH37E7eq9RnMwP8O+BWOJHmS2AMG8IlGDT+Vx7AXvrlCSBJ7HM4r6n+MuLu+tj8bHEoti7
Aku/PHYFysUmmPxB6I2zOL6rtUmBgQJZ7RJo0wvuV7XN1Gk6zOxt/EsbUgvTihx3/sn3cxpLZfv8
nvrxc8aXwWdNtRDxPTUZxR+pTndH5WfY8A1XvOLsH2jVvyVHaqIzTQhHrNH9BwS70VTQyKsCmGLe
0QvetzYVu1HE3+GFcyPrWuZjLGnKAKZx39t0Zzfg8XDhSoyyLUIgJ2DDHWfdZ1JH8oWNNfK9bMIM
65L88UmwhZLfQ7rejaT+Mu1I89Nwiqt3e8frVf44cyGned7NfmJe/N1LAsYQX55rIQ4mIfPsZYUW
eUiSwBDTQ+/UdfjFHMNFvHG7RUSzcZx+f4KKXGs5QXSC4noX9D8b6Z8TvZbZgcgeG4efyyFCNSpf
DTqaq+vF5ZmnMFc9wnVGsCfBcZk6708S1PqbFAJC6Mz6yJZThKmDA8hZxa+gVKCapL33MElecrEZ
2y2LRTurRtXIjL24+dccS2lZKp2njStaMPz5Y0T4wi7pZTv/U8y/sxaY+hpysq3VZJn+hihyYNXi
ZVizGzoND6D2kCKaFI+/N6+WHkDb+AwzA2xnx4O+C02rTP2UaCk31hqEEYSamOmk1g7DcjfWn9fo
nXbevZ8S80V7Ad43BhJq3I4hEDPJPF6oo7CM/oh9eEO5Wqg57vx/MxsWkQPvRL61dB2hNm0QeZei
zEYrBy+46KG/0Kf46bu7DtvWQVeJHUa9+fHDR8J+tmrN3RNnBzz+EkV6d3ikb47qIsCG1RP6ySe/
5zmunWMR/xJsaaRqm6NQC5LnKQyE+V0uvtpwK1cbQ+f1Nd4mPN1DOXb9RCnafJJ21YAm7CmD6jR9
Z1BvBsJkC7s6p7OynMkqydvyzr5JLOFKswC/SmP3k4JVOaw8m+BUymy6N1/qiWsSdodzT+5aRSSW
3oZOqUKcO7L2DjIN/DhjpuHHBE0yfDSes6NoWK+UBpgH9DEuD95jQZjU/AT7HACE2MMkb3SGjh+Z
2bhGw9TvtaHrT8ImuCv/7ieupHP/vJY9UAXBgzYi+E+aQsSNI+GU/c9u06SdoEZ11uFmOhJplSX7
6iTxPZWXmLPz++usleJiQZ8sbY+ofZ3Y4yE0YTpTuUTRHw9Z/6RBZq+9s753Up9D/+C26nqJ1HYf
AaU4aEDGgvC3R3VBHupfcWO+Ab1tLm+aFW/LcrQVt9JfFH5ydlnXsJ2pqhtqAGiDHUFtxWNy+V5q
mxrQYsSFlFdFcd+8YSJkb2zTE0rBHcHOZVKYFvZFMnZxSbjsu5sf30wrQEdmJHqyU6Sqy+viMEy5
K4EDAJcNb+LhrFqPqz55iqmDWgOR0XlUUcacYHzqYD0xBrGiolNXbgT90c7h+wOTeOnnsXjCvp/+
8XAgKLnwnJ/zBNo5CIGvcCYAlGxhuVa+3/FN/NNslToOv5zeNGRg0tnatNMNFxbcPanhFlt5r6iF
R5IWLYiAYSg0ZdqCC+n4hs5a4WAOPckGg90CGqYuLuDQToUhwuFw/fIKVZi3Bb/KM+j4t9uhpuwg
ms5EPFgnIlwdldb086drtPKvgtovc2mcaaQFnaY/QU0+lwGoyNpZNaaktLrxMkChS+pu96QmQ+uO
eFiwNryunh9LTUlgt98BQXamvpQSiPCdVnqU4/EqeFMBz8NtBP8XsXneYlK7IWFY1UTyl84sdtHv
KObrp6XlvMizG611M6nUX2LO7OZk02q26YmfTSEEXSEGb4zwTYqLW+/42yYAYRW4zGVZ6O3JIR4o
Dtbo3FXgNM4brJ43I60R6c8pRj2DTMNh5g6etyrE+yaAo5ET1Eh3DUNik1gYklideoO4FfHJonMR
wRvMt71kek9opToPqaeqJy21/FUU/aFu5XqFICXNWiwrxXqJ8nOrptUlLkchHtx3viB5n61GMtaf
t6a82sVgZn6AUh+IqjbBfudl0m81DzSHXxIl4n1iPJzHlNYeui0zjY1+QrSAehLLsDX/YxG64U/p
98n6qYGw+xwS7+C24LH3hVgUivRsU4+DHEK7bQ09q++4A2REEgb8TM+Pgqhte2SIXmzY1prAFnz7
vI5S4AHJJlitzME+EchSu4NcSeke/LKrAAYlvuJPKnHQ3FYI1SKhd2OWILTlvRlBpm6RQHSHw+pg
vRYfsdVSfqQ1GXgBxNfzRt+Sfe9lAifJi2CjeGMK96QQCW3IOj+FDKUEPjWwnFUxGRGbt3PL2/oR
6uBLY9rdqcQbqbUviG06pF3X9xHpsLejlCLwo4lcjOCVFMFunGrExs8F8sW79M++mkatUVQl/Liq
H2X6lu4dglGC7Cv3gdRyQZMsCA9+oU4Rzy8Ql0KStHC+PtuwHLXGUsW17svCau3I0nQSqYJzVh2v
2jyZo/wHI1nobnMrWOYpfyCGLpCOtHoG1hsNd9cttspzuQl5cMsnExHpnuvgUVFp6fsMmEazehlO
YFZAoavIZUjwasm3i54D4Wd/IDg12FwgAEgaTr1g09ypstfh/vS9FazUvBM3/6QR7JAelitO8mgX
4Aa5SOWzzBitq2yjaxFmyrfoBG6wUDux7bxwIVlJKQ04V3HjEXZ9VMZXBOkVxmvs0YpcxlnGD+kK
CcUcV+ibya9kXrztpOGuRnJDvACLfY8mYLxWE/PnwLSw3C+X6Q6xxCVFOCbPYp6jSmjWtVTxRPcC
sdWfm5GKdWQly5M/VJLAA5Ykkthpq6sj83G0HuME1X0Rpk+l15EXR4O+HrwhHLqcVfvQVz1mhpIp
hVQVCg16V76IKY+mUoOMYRBLDTAUmzwn3DgUQepG6Fo5HdMAqL3Pbtng0/1Xm6Mv+1lZa6VceyaV
T4OnEu7J4GjbIhypYRc5r/rmBpfi9wsHREQK8JY1h0sQB5wB2UROM/aVt7TBg5tzAoFsH03VtG2C
PLdsSv4Q2D6QWQbWfZj3UIiDRwfVuwlJNUV0sqMrogxb41ELKjlNk0fyUPEYLWNbIJXZF8LL/Bsc
V6/qrtcw/2DIpcyvPKdWh79HvEC4dEzYnoQ2SjWwLbWLajK33uPrtPFmQjf+Rnxviw/qTLxbt7r2
p88GT8tYaC/xDVcfkgwkCKSM71vsh7Qx/CiJyt8jJL884t87n98+Qin238PMgI/cVVFWJAXRz6Qe
5RNxMgYWiUs7qVeDBbudsKOHmWSKVgAkWuE9WgNdy0XZp2vS5C9lx64grS8sjLlETWzbK9Tivm0S
uU+HG2CkevUD0kSAhzJj6ObMEC/tDZ2xYo0RUi2SVUcpHPWizJnGVDJboU91seVbQCLlWGSM7nTg
jNu/f3PFdYsT8JYtr+OFirE5e9SQPqvrzxY+uyRGPcfEG0n/h0/kvd6dpEpi5sVBp+BLaVPjYFhs
kfT8230sG9M26aHJpwU3mb3q6ukg7a1WucGN9xgPFcv5dmPcp0p/EuyVJei8DUyuqJr2HUr/iTnp
PhyMdBy7EEZf+jbQOJNPCowKKtq6TaYNsiO4zV4xgXU1BaxhoTOQzFBaAYaWsf0pLzH/TVi3D5XG
vmnYWvxqNo+fBKRyC9RtI21oQ3i4oAey7YDh8pUc0A8hlAssHNQLPxf+h8+pmQW2ja3KfroNHHXO
sI8/5R0MngI3QeUiCCCmimzR8+uoFu0xTqbaEZ5GjhkTIHOLweks9ZhJtAwFeyurtX/1FC+giZF3
DZ6VFNTLGn8xHDSAy6GtVX+U+mtrIrOdN9edlbkF6fKGak6Ao95N6SV58FBjdCx00d9vcdySTLRr
ycsJJLFImLRD0CkVO7ywJra0MdOvKjOJ16yOQUggXJzqKe1Syc0KNFWmsnEq6lRnz7hHVgjTPuZ9
Mrtxg5F+pTcYH2nzWWk3+JNbGRrbGCrYW16UkTKywm2zEnAF4kKr06dC+Mv7ag2puJt1RP1LgD/b
nfb4+835PSSUgxYEzzkXtRwdG8TpOdBKfUUi51XNVyQZ+t9pYvGtrdu7pPdue2dYNhQABXMeayAW
w949wgCI+upqkY1cdtjQRmttcYafMIiWVCfpqcMzJINqJ//3asyVQspcz+bLLtuh8g2VPLnGSqHS
pJ9EXE7x8K8tj/cd2QlMUrS1ZH/z2gHyYdu/do22Fgvj1woT5g0ck3YDedJRriqumAwcZkw4c4A/
/9YyPjydO7I4MAKvrIg4PGLDCyDOzTq1h6/xdBHIDNexXUspI7UfY3HLqzcvBcHMzlSkUBjiHB0F
XrvWguBVK+vUvwOKnF2DGajzJEc7RzaaV6le4PsEOkzn8xU6DnfAhsy7iOEutqLdZPZw9rkutt8j
IRlaMmOZCoMeEfILHuuaGVCyB35pMveCuL48tgE0PAMhgEsJYvMJ3REKaTlno4UVGv8Y4xhyXBkK
H4VAaRD1PWH3n7XyLKmrVeScdHFrm3PSukEqu7TLVYS0Fn2yeprUbsBG7c+2/ZMcQdnsO5IIIzU3
rB5jbyGPXkMim99Phdk5n2sDOKmTOwTKYG/b0jgb7t4XL09RyPSU1fcURzzobqETzJsXQg+j7Q+p
Dygcet9h6mTL5hMwu274WMArkbH/H+etuulCDfy24SmYsSpThZe/kB95ml5XbhPEscdZBTnQ7aNN
1eCpfW/0X1VGDJItKMYsr+PFORPrbrJ4S2BiKVj/0DCW5fvAtGJKn4z4x4gtgF9YB7AKVE/oOOKv
Wmb42PmshgrzJYqV7+hMQY+pc5wAtOwACa5suCyGHM/LamrqwJnu0s+ljSTLbhsoM/vMCobuubIv
xx/aEBFV7FOq3PRFgirGSlkNhoPWSHWuAa1eN1ZWruX7fN+O8PMpBzpTi1rUr9sfh3A1L5HQsmdT
9IW0QkkwyLHUKEVQShyhvPM5ariwYn8L8/6D3PsPzuxkv5N3jJe7YE0VBEQhjimKQycB0bdOSMFB
clNXHrlqzcU3JCfc4Jp0cDllz0SAsi8UY2OtdluqHFnc3fG/psHE8OiAifwDkavf+xFQ17mP1arO
0QPlp/XdFQ1qGuXhX6KZRkgEWaPi7n2eVbYn8hv5cqy9fefIietla4Pc2wKeLhFNW2tG+IgmH33e
CfVXdwSX/fLYeNT5tlDllFokJllTdq0vs9vne1etd3m8Ozvt2sjL17ZqYHI1umMNcwOYMCSriq/6
6GX8gFx5G7mRtPTT1A5rI4N8oIYpnwDJjWIWep1lA9gHrrrzkU9tNPo0SZPXQpQI5tMCdE/yqson
T8eJzumKGzpQ2xE3lMpWxxNUNJzOQhwvwpYKpijHdXIwY29NmNuue9NSo+kuAgfK9+jeMXWtWfts
aVq81zognSZWCTQ0uTQXfjWwelFBahrlPQsd7IJcj3BLO+99ZN3Nc2dd6FF0AnJaqlHMSeuFyvw2
x06bMhGYSUVT5P1/lQpTrYsQWvJWSVf3YtKdDXYqrHN5tkv7Vwcg09rrtUXXb89TzHB71WDtd1wa
05IMRPkhgdTd/1ePHv/A5rE4l8yikXJ9rRp+rw1GCIo6JKbZ7gbd8bJXVhRnRxNlhlCs/Mlkj21h
ytIsjx1rhxLG7ZD7OGyZ6llXf/joV5Pkc/0MtyFiPjXu1FVwNZRvjcQjaDnBDFWYUeCTfFqg1sse
o3jxC3T2P2gbAS+orIpefDhbziL8J7UK8HFjLtPrVounIYXXm0g1w6y0ZBllKxPPCObfCV2mUz4M
t4wLfYGOAaoq6Zs1NkXAJCp83F25UUZbpjMom2Hq39MDMmNpOAUHPIEJYzOyWWNSFwkLRuO6/W4j
+wqJYEl5PVQgFO/En7O5MlrOmRUt5fAH91eHgU2j7VW3TnPYTYFh10Ru9cbBBPGIQ6y0uMpjUEJ8
sN7HnxgTIG8vF96DPpt0rWu5FCFdSWGzfKMWI0WV1zRq+tIdFNHVJkFhZb12Q0lKxbp1LHxv9CFs
SPa3BFurTdjuofs/U0Nx8e4QvHy5+/o6/ZySgORyRVC+qAArBHwuVHDIklNoIeg/+Un50KhQ7Clw
dKZ8V93PFpOTrU7I+zczy0pAvMiYEVmhp/AAkorW/dDgDgsgHk5AVWXtDrpkXnRQdIIxwEKJMTVr
ggmUcMefhsfNRybsAypMfsTP733ToPPmPV6Tz9BNazDYchvSJfdKlXtuy9aBGwuobQ41RwRiwkM8
F7zTtybWi0spneiV/U7uBeY9F9+6dNaJOjzoucILhU/xKqNHkyJ2lyWTKZegNC3+AcHZgv7ugnUp
yc3qm5OJRvfb1WCUrG1X0BEgwwkNAx/2zpJNrFC0PjHJm2NCKH5hXxz+nH2A+arJl7HiSKwkXdDK
Fm5UlovjzqIooCshbeMtfUfpW5FkeZv+8OlK9NZMyFfS3kR8I4vZxbdXSKbq0YgAAmKL3LTP5MM+
XfB7F7Y+zXSJVHNrR7HUxphrBDRhlsmcxAY581kBE6uA0MkSg/T1dw8zYCyGIKP0SCIDcYBPHS9g
nVYjwfGnvzXfHwcG9dt/Qz3pUk7Rc3zZCD/K/mNrukQc/S7Pt7SRi9IcPecdhtqBs2x0A77tTBp8
lHBmvmqDXu6LXkFNu8gVHkBlnGLJL4KPbdZiq3EdKMN1D8voTb/bOnFvGy1EJ6QqMB2EuslF/JOp
RceIxlwLToZ5K7AMXUJYR1/9YMhcNqm5TKDfBlQyTfvNUxI2EwfAILPRd4SAjKLoFsKRao27UalD
Ci3HBdzTkbXMJYQSpk9u7lmCbTTkT+s4sn7nTAcg1Z+08eoXXWovf/CfXVNRLvazvoNl5W05ysB/
xkrv7i2e9ORxnJgXBsO2W78AeXdg9RQ/EVd1fzUc9k2bmxJiKoQBdl2ULcVZbHQHx/MD9C4B72t0
tig8Uh1G1y0bTsnHQS/5878ZJO8sYSQsip1yi7ytWLrHhr2OyWztilfITjyeOL9Pm2hidF015g/Y
/pA+Y0dxdW6XJCYdqcqE2Pya9LlGAigSb7FSiRBK9xPkqPSFfNYYghVefvVeaMz2BWGhQEhcVCTL
MksDF6MT6cp0x8xqc5xwQXjaPHBgiER2T4JA6TnG2lFVSkk1aZXeCtuhCLNxbHn0JxATxMetYN1f
OTfx3wcQoNtESwzNnChVV8S2PyeX+rqxXKMSb40j8iJlN5cAP7tt994Bvp72MEoZItLhnIX6IN4O
RqTiW9pLu8lRBIy+p3CfEAM25rY4z5nfLG1hQLJ9co4P0z+/v7iHv09g4bS1N884mJolArJCKvjA
Klh5osmAHNhi03xQF02AACztb2YUpBe0W5tNlauIH8y2l7D6V4RBHKI7VwmCYhn8udtY3uux1YCC
MDJ3egDUmR5pkqOqDVbgdv7aw/LshjIU+xoqsyOTYWJAM3wwaHmXe16Q1+n+8LnKh56VElYudRxT
GassmdXJ6FKJB5F6UqY/AO1ZDl299NkkIhNumKozaLpRBW+ZiONsoQ8dSlAMxrI6ylReqCGXEc/W
zr7n6WanzCRtR+MKLAs5qRTUuN0+1S66RdWIS1jqtS/PIjfq2b6U1oitBwTL08WN8KUsh3CJzMK0
NmfjFthIyVLt6I2KSMENmAbMmWbAaX6hMVY7OKNgKJTwNjde8UeSni5Sne1nfPUdqLcflay7c7+5
gNRuOAwDNWINfy9BRlgkqh/+xFMPPn7/TuJKYv7gVeP1Z73IJ2DBdG1VAN46miBQAj45X7Qas43C
KfVcN+qPL+/HC+iRL7f/+WCucBn6Y0+3/c+4hX3FkcQGBRa8WMCw1veYje9kC91aGLfikkb8xSNd
D+sVuntxyIECdUNuke3J+Z4t3CpIiGnYXiGgTATnsvizeQ+8xJHGJVVnYfjnFS+aYriX7OPtWBTL
REcP0YHQ+JccJDPkotOAT3l5BVYk/zTy6CzkTh6Y771HTJTvIla7I6Qvuqu8yrohYQ6TgTBz05gK
heVU4PdXCJTwmDKnQS9TH/AfDYtGM5aCcMaB89i/ZP7wF2avgATmcB9c4Wh5LRhomFLzybgxlwWL
CO6rGcTQfzP+LRafpuisPoSAMypue2TJWVvHOqD5drqfucPkQ0Hdhh6LH3S1bcu+W0mfFT/ca4N/
ItMFs5JBrjSkGP7oXu6n+H6B5nv1Ys5/S6jz10yp14a62Wr/kmbV2c/9XrKyuKXk+aPYIMeXkqH3
oEtee3FtwR2KNHA3XECp/jrLm9OBxL+Srj8XnIgzUj2cCHBS2+bnuAqoKon9yf8zExLZkb+wJn42
T76Mvodm0e5tEA4bUg0YI+DSwbkvUSZqTD/hmuRIDGBAtrlDGxi7e7s+Gdol/PkHrNiKZfyvJI7f
/bMexmuhj/t3IkzaiAfcJflyYzMooJRmVpG5pxSSTSZ/7TEXyxXawTvfBlSKz9gXCfLD6YxOT3GU
Gup7+2ZWK3DS7RpyzDyKrLbmXS5FtIsuFG6qRz4s7tFeThR1NcqiXdkIntQR+YachDhrpG8N3lif
y5OckImqzi6tIG+IdOEo2/L2kuj9u9zpL+/xyx8JBtxG8/6yY3OcRzK9uc7y32bvhRaghfAJXFmc
4EH2LEiTm/+x+0JCk/6vb0md74roNv+JyJZPvkfMUYND1Bku+z2/QQsf0Sr8g+iTz1PZ0t6CLsIV
ogBb1jqKt3nRE4e3j4yPGdVQQomgfViVOEifQ2D5MDctPK7oK0xEK3h/2JtELn3MTg+RHaDt0rAD
N2ndvJl7RCWVfzKnsX5aLSWzwq8cAd5+eweHgTw/Bazq2J6vPJiADynBEiO5tfH3O4g7ZUj8v94c
368GH3lBn4sTbmaXOLrpk7z8ZO36iBHhL555KeQGKAsVbekNTyqn28oYYNlC3dRqkoGyvHRx8Lxo
kKWeKTRAogf17kOZt0dRC+fWTH4AZCiiByWvm7PA9v2LLCfVGMw8yDLTOTe1nGEuF4LL0ihShjFc
Ul+JX0E0Cud1lf/PPe4uuhKQnQYQJ8raOtsEC6lv5dwsCGFEVzfnFXtRd1HwXtiaTDTfDHe7Pa02
QNBMlER7jfxj9kcfSAZGcXFqQ/C9u+cGvJesSLDmRoi7gmAoPUhaE71AdegvlfTU5ErGglgOleRX
K1SC3P4EJwcvyF+6uvGABdaQlKyyxiAtqzYhqzJznWb1qSEznZlupYzZIMV4tvYcdtBzp+e3sKCy
qMBQovDTvx015odOE3xKV+xT12MnSjsYnsEz7rZ9vhnx224Hp0bpdojE5LImC2c+X+fkoJ5cLjTC
fMx7bRoYgzGsXU8ZbFSIXAP8KxoVvbDPwrdBCptYtFqyEWvPDIsM53r+K6LhT3ivCivi2pRzzU8o
5lztnRgGmU155xQKAZqTFUD5yNvdOK+6QtRlxo2IV13hQcCStvtB5tQYZ0BPxgONUL6t8V/sUs1s
RsWR1FPVFKMBm21/LtiKz6reWYNYgitmn3G0amCtIA/Y+lXRuXM/326KsQoeRU+Q/fxEnLef5YOh
FqPbetBCpO1j4w8xH88ZfjqMzvXxg7jYuRynva0og1EF9Y3QMrMcg6Cx9d7lDS7SYkDV4YgESRcn
S/m7R2A9qDXTDz4qhrPISsj5SWlcD8aCHKFveXL//NrKWkjb9r2tsVGZSzFFcf+DbAPTV60KStLN
Xs3mb/doM7eN9rLG0qOdEvzWeTnRUxnb1qQ/aIHOOA4H1f8mcqHGbkQD/8ipYGYfECzfM/IvN9W3
esMA6GPmbwHI+UrW5vBtqWAvlqaPdWjKUWODHnh/70H+bQFh6J9djLCif2FfmqeCGz8TwRjHNLWi
Jd0fdY7YA6fLzxHSrq0EIwskk/KOUdCIaB9A+fyy3sjsaOHiu/ORVQZMZdpgUSSa1tu6+0caMBoc
UIM9hR31Bqu3a+Ak6NyDYK809+wf64aLJgG/vYdz+TdZtvM9RgSvv9qXO+YlEqhMLN7Nuaooc7v7
UeapYpy//fkV0BuE3hTsEZBUTgEcIbhlEhWHtj7//mJZPgfXk8el5bzbZGOf5iafwKaqTl8mTcg1
t0q4GdbFizNrQdwQYK4DCcAccreyQx3kAxUAm6no8MWeXge8JfESjrPO5UAiIzcMxDx7srsDSPIO
Er1kRTBOWzVwVqljW56Tb0IGNhvQm3B4R5KyudMBYU7WXXrhyO349aMXENlHZ9GRmsry8FDnpDIB
kyYyU35Q0e7f0e7SXzWWlQqIAwdrtpp7OYivRXX3eSC/P4pjtkmLdx1lTybQxeFUyuivNltLMKc7
qWDxo6nacNURtHbyP64mywx+WiKDtC1fYafyStX69i/d5/VX/U+QYN3Hn1/IlL0QdfszEKvpyAhr
Z1bNhybvs1a6zMitK4GEYy8ZhuDb4Urjpej+88iJcZbjkNhpOe+q5wWpw52adMCp5yyG9dMtbWKG
atUmOWTeIB2mDKNQzxDOuwPt7AshZ+rviC+jxn6c1lnx4npgRMVG8KsjLc8a5RDLNVuC6QP/PUND
OeORmiF3xDasGtwG4OeMebvbSc9FjvyrpnbllqKZyER4SdzDGOXItliABuj2bAmVcqYep5DDwUmP
qUnkrKykEvw7nmYIlzbaHEoqSfMlhllxJEE0T/nIBuz9BlvuR/6D04CpSOxy2R5BpFVtM+yLwWi5
R6T1nLpPuD91+/fWIGDUYelNxZ5555RUY0/3TLvNIrT+thOqphGrlVta9gXfHKGUrT+Z/hS5FLmw
dvKdXG1foLZzbeaHZED36PLxZ5YszMCyN9RQbFTHQMSeAI6yuIQPbdoWKxn6guAViy+bB3ip0HPL
3QmL/pGd370lrLz1po7lCRZesHLrxLIgy5MFtykQayh6Wf3V5haVNNIUupv3lM6gCrY3iAgq/Czf
MUbh/Nsxid9mUjmRMAhiuEPrid6dnR+mA1xa86udF4Tn+ScIY0GAdl4RXlOyubOfa/dOhoFWeUAf
TTvaj3aFBGNvk98mgIkwvrvZBWrYI1ir6+o8yO91eZPoqZDUn6vu0URIxdtjLuuuWmCC6GKScTrH
alIgWxBowkj7h3q/djPM74L92liVnegv2KbjmxPpFVK4BX8jB5SEyh3v+XFDmfoWcg1Rq3w0g1HM
PHXxCOOT9/pbKXMZWJX9Vghf3NEfpmnV/SK0qs0oIk01YBz4n6uHhk1Xo/Ge3vaE/OWCQQ/R6E3e
LYXwPg1gyWikZx/XNM+Ue4PVOGTuW0TIKj+VjQLWomwS78Q/NgYhY2XXkmxZlYyqUwwY1e1DEXqW
qSHjEfToMyvaQY6q0jMGNg270gm+EY8Mhsv8lEs/4UJmSQrKuAePGEFGPLlZwx6xJQAVAG+bCdHX
Fvyrk1iZFzOwchgghVvaSdX3vMSSl6FDQgsqJHQk9iXKVO7+6GUANIVgvnI5+eAGxjgaLO0ngmb+
lwRw9lQ+Jj+wTOY2XCowrlPlGmkbOh0z8b2Guw1yHf0jOiJOehHZ9tWuOJ+x4DIt/rgH0c/kOMCN
C72rGk+PlkxNaIy4sQ7G5B/5e3xuWyOAIMYKaIkJe1PvzDs2ZSHJeVSEu/kDJm/7Ka7wg5UMMPiw
CQeP2PLxWIPlktiUSb1uCjslEl0pCjB0yGE2vi6mg1/P5dIAvleo9bAvCO3AjId9VX3C0UghO+zO
YZYkemTZLIXoy2T7YfdQ3/z6q/AAQkictohE6CDB3Krl/znKvDhsC8Nw5F7J/cfKTBfPo8sCdS8l
0L7qPCRUJ+KfMtfBtSktCeySV+bkhVprvXN3DHgMWesv3iXg6qfGctURmNCya6qrTvPX4B0nQERN
Vslq2wtZvqv0jmVB9fy8g7OyLX1Kkwy64t83ec59iG7BMmfmvNqDsr95LAUD66KcC9pgEuhD9b1b
GP89KWv39FTUlrl/2LFRAUfeju5TWKh/yTQvIKOygN5X4fHXGPI9Wt0zBhxwqAIKbVBYwqDCRYT+
16Sl36vb3EpIzE6gQtY7QX18E43G0fP7VFPk029dOXmEqW09D30/03j4zqwsMGu1+uEb6ourO9AK
Y7EWQL3K4oVfobwTX9jPj52pvyCA09T4WPL5/Qu+aIayi3Ns0Y0cNJK+L3RhzuJ+UU59MAtTomPh
t99/+s5Wz/hGUd+wDi8m1bDCcc8eHQmy77c47Oq7gP7ll3/wSwqAVBQdjMCWQaUM546c4aM6crex
xZnTO4kGb7BM3QtJB4jOLX2K9MAqQkX32VdtETI+jJbeti0XBhbfIrqj7nCHwq7cx0wUt8tus9vk
z8AUy12Ix2Up3eWgMV1xxDnioI6UswYogyhTZjWnNR7mb4M7VmZiq1cDECsT3Z+nUAZaDEzqvqBT
DZs9Du1NDyylzV5pr6m7hntvE6EboyUFaQLziHurmZ5gUcEMJEI8p1k0L5BGfktDwv3K4EUqkkuR
T3Kb6nnmCYiLiPsNmn5bMGTPurdmr9d+zxBljPDZx2yG0uPmVQJwO6FrZu9rpXr7ZE4J1zCIbW5x
5NnO2EjQKkctihO0+4MBT9w29Va2TveGVbCqNqPVqYE1SahLqh9w//lbFwraCOCbmnARs8VQ97GX
Ft9QVS6D2+GjnRKb9cZp0clss1XJzdhUUgLp4U43kImuSaJRkvg+B6gS008s9gpBwAgGG+4wJx8D
uR4ujQpzI7YFKIALM3JqPYgujfM+TEvTZTKiskF/8Qty/RmXZVGWvbFSHO932WFTMqim4bXKkyqQ
vasePFYiB1JhLxoJVKYDUEe1BtnzrzAxEy157Z80djybfz4XPS7laq8Ro2gALBAbR8tX2XHsi2j7
d13sSH1NfD0UsaXGcXNsrHw0QzqHcu8WAT0EcEQe322DcIxoqhrKSn4psH6Oz60SXLrbZDV7zt15
Qh2bm6IOKZLgH2BdjmyR8XiNjH/8EHFVwTJ/KyDtVXbvCiide0Id7G8tRdlhD2r1lK3QX24Q1a8z
+/akoZ44RSSMLUWTW84hsDZZvbmoH3dCT2daFqMa/FS0yTTxBcAKfYpJLA9cJBg/BlBGLN0Ns1df
Ze1LpWfTNmd5kSdf+MkPcPn4+AXGUvuetJIfki9bhKh7GkJqHtML18nS8Vh0uE6z3p/1kJwfZCSg
haooi08dof+njo473a9b4hr0r5WC/5wAE3v+GzkNKPPAUyWgttqU7dTmItzJKL5dtTqhjJ8RxOAi
8hxkZYsdOdfPpUnmN0teMgKrgSXCYWRv3OQ5hCUIQSzMRT/ZUE48AKC1LBw8M3ii00p+GB74Yi0D
8jZkv/ZQzcr5HrTU3SBfclXfybUhUw4hnWBxSDMY1n03rvwPKpl7rw+ijlmpBPG1QpmujcVu4VYJ
TQs4qDqP69pUrAlPQ+wviK8CFjdx9IKYt0dbrrgeR95k1e7o/Qfs8Ox5+PMdqUJjV/tjv4qurPHC
LUsE1Kf6wfq3urtmMIfT1W0thzkPXO/D+eiYMeRVLMfVVi1bUB8Da5AKC0gGXJcnvG95Kvef9VTx
4ivLYa0MaJ08THe6b1dpEl9rs+VuV0XaqdzrEVWes8cOv5pRQYnY1m1HKfNwmrp6DmiONCMMys+9
HM6wuJVXwk502P/UFYQNYYrxIDfqMQC24edt2SoLesKQo83XwrgR9uq8803SgSaJU8qWCO73X1Gg
nZAIlm9/PP7/+JhUyiL6auSd1vCknLT1Dy6wvaigWf+yC+BdDiSwtpDbGg5viLILcskd6xQv4rzQ
/3rMXjldBcgIupatcg/t9b5J4Sp9/aclA/dVUvjFbFvCmhdYr2emdcSfx42pJOpLjkai9A29gykT
S/Ugj2lEbXKT/htqnXGUSSaq/mYZHWoShnet3xTHZE5eI7TaPfIKkl+L6BwmwMsnsrYbJJ7gNdSi
j6jl56vLVgH2O3WJ4LblU0RQHElSJby7u0ologgwsEyfZrDx2zaYK7TodbN3VdZOn3ibC7VPmVjI
yKWaw+T+R6aO0gLOPyK9F7rZvHvNQW8OeL9M5RHhVLcAcuoDffjCK287ZNe14PDNG8VgG2uSn15V
oBYvDmPk08qvWIpuQzc5WmpzA5dS1JijVwlL6ejeO4Afu5vsGtuRV/SdUvQqM0Eu68SJTmzlBRMc
bAipVEZNpnIPsg1Eagh5sXmk5XjhjYj1lg0wAl+vt6UefADYb9OVOlFu8Oxz0DyEQCAxLo6BPnIU
WVn3BPj6iTLF6EuOSYAtsxmu/EDLBAHyawSNy5j1UfN6xhkyXk1dMWjVDn/RlKcYZYJqFJq+EFEJ
S6eN4XLKeV0YOPqDPiPIvcm7bU1v9+95PQc294DDPG7MB7OK5ATF+xi0kwUDpl4081smX6MnJ0Q2
NIOjHraq1LJCN0WOwkvtSi8vp+0FR9avjxHlU/RYty4RtQ1Alvt0GRsBzafhu683IlTulJoLWxOZ
EUFQvrKqp0xCN/hexE20LUP1cNAsS4/ugau6Yr1/4oc3qgJw5rh59wQXXpyA/mOUaDh7yxK7LE2a
oAhbO1zXCKCaranwGMdH4uboXnMBppc+HHBE9lbvwib+UZhzzCokQ96Om+qXyFuAeJ8Rj2HhP0i6
c8icfDhsQY0ZwMDwMYMPKGlgDW/UQoPt6P26kPlCklJVx9cO5oyCytcG0j+MR1zWOlQJ7GUZbXFE
iM0ASwUIUklfFYuY2c8UALLEGnZg2jePBJdEo/lWO/FAUU1fvD78zp7/EBsZ3ua3CH9GljS52juH
VWyGRWEg1CuOQF5DIAMK0cIK7E6I2i9j9ZKUU1LY6xFY7iRPbxIsAQNY3kJPqUoKJVZsgpg2tM37
n74iioT9VjlCQkLmBy26ScWRok2F0p459ph0rpBZHZSjCGAm4hYdZ7DsNYYO4dTn9SEYhBMGCYx9
KWCu9LelxHsXFg8jGIqHw1TK5JVJb8/38bGa7zZHDUgv9TirweKkFEge3UzRvO74w9hi83S930cg
pVY0Bhy3bFc7Fk1BExwB0OCMAARYRtkho95ZFU4lCzpn2+BWPxsZxNBglj3LqARl+O2ZRf4PDb4z
G2LYtAMStV5N4sAMCFluBMzq7WGWYjRfPPSf2FWlqDR8uR7QxqcyRoOpvtVLC9u/2/egTXgc3NY5
zzXoaznVFwg8pjMLyR2QDst93oZDwZxdnkONwgvdTf76u0YnRaswoGPP3Ivk5+9Y+AM5qn5a4dUB
153MAkk4FJG+TqkqqqKnC4rNeP4Mw0KGs3INIvnl2EcBls0On2Mm4EBZKz2/YqEDiVo0TrxBcSM9
j2L3NM1NUKyq8927CSIOn4K7rEZD17KGKMYB5TQl9kBlRb8I2AlXg+h32Yad33Ibf/e/NSBtSFev
sAEKZO8USbFj+qLI0zm/FImM4YV1fG+cXWppmDnzVnUdtz2eUmrkrUHAszFVunVXbKsPbTf+Wl16
ELITwJfC7TyWTZ85uHehkHu7bnqfki7UqFS94yPkmzGLk/X54ZX3TEoJb+Wlkq/JvcN7/HOsJe37
KHQu6x/DxR3Cgnt+F59gM/29kC5wC/ZtXDD+BlOZ63Ihp4SPepQhjD9urYG0RYyLzmqdCGxKnpMZ
UyoTLC7ekF2fOvuyjFExYWLZ4qmGJqcBVfhXpHSTJUrbSS6QzdVGmq/AnAGsuKxZDu+YwoAJszJ5
TXJ8gWofQHumhil8t+2LK/PS4M5E7xPOgq7/s15bk1dAIDPsYHLMSlsOGeZ5EbHigE2Ro4+EuQzO
V76pQ3ibv+jpSzfKRmIcdTXFxv9gzlamdpoffGsQT+AWE6xKl4wJzKnYEi6AduayKmF2zrDr2pxc
OClXtEomFSbHgbc1mwUq0unuJmNnnXRaysrpdqcV9YvNL18RJ3iapEPfs1QDQUkRGBKtCAAMo8Ur
Q92rhe0PeJoLnW65zOzh0GDiKcRaEWA6AZ8zPMXvRNU7KzXX7xmOgJ/kIfp9KD1aLKVzLDDcHrqA
C2IfsT1qoAQhh+XUqYrBVE4jxQPhuZBxve0ebrVU3+iZBhdP8Cdq2K1k1TgCZ6RhHnutWOIjxDRs
HFOpNJ3JjpkYD538w05k5TJepx0EoLNMpnxtefn4cuWzXrSiGNb78tM40I76c0ekXi1+LlD10QZQ
M1VKMiUIxwDTVC/a9lnJJ2BSZcci53W1rkEshNX7XDG6ZPnej5Sw8Dx782uoKi0VuQF5G6UOoKtY
TCpx6RRM2KP4PASNiO7VfE7sau5eeg3x/dznNKp+NaN4uL+iuP9MVoq7CF6phZSpOFsZN/85qe4V
3UBoU9bk7m3voG/6+/jmcNDbXJC2gCbF9ogGNkJ3unA+c7cTbXyK/83kR0IB/FJaAq5eKyvQziOy
q5xCCaHedTOI1Zx9vrk/0BwgoF7YphFvbvGZm0glTPwB1ojqM+Jvzb1ROLRzm+h7IWNpmiQ0DnUz
35lDWzp7PFwyZxEFwFm0fq+tJ1eIi2t1iVWcAswJf1YlG5kGSFv88UiCemRf5YdpLWIMJ0Ruc/G0
J9jaAs6Dp6eSiB34m+6QoIc7vDZ8HEb8WS3WxO2GTYSmmJEOxAM4tPLXwBEBPPq0H8ITQ3idZYi5
6pD2U450EoRdx1kGygDKpVGbm3KVVdY0rXsNKwy8+DmsJ41WzSLgvqDS3UEdP2KkATIR9I1PcMC/
eHMcPmwIqwXEvRrIW15znFDy6ex9r3jFhm6R+OlMB/93dSN/0gna1lG3qbMQTv3AOZi8Vj7i+6d1
tlzZKWcKOq4fe9UBxu2i0zBwsm7V7Sk6cZETvXP9/qsOH3OjZDmZ08bQpo6XA32leVaMILDDrW/L
Zu/FT3bkNt0pHMSkWE09k2KydPTe4EgAUf65rShDfGoLQzUoq7SiVsF6rUWmD2LNv9bmNfI3EttI
9sa21Tb7d9FcDDiKnFMlBYmJTYXn+nBYp0FEmF5OtGprBG6CqEkKlw/OLYuDpBhEtwfbtoBsTulf
EkhUahANuCf4rLeUo3y/KEU/KxcFVw8E7E3DWm5Wr/m/Ue/sjNXya56oj7EaWGI3fC50FPKudRTz
mCkpR0KVOWM8RhKQ0u8+3/X2HhTGu/G1nJlhZJeyZ/nS0br/IAyRYpNoLOzafRznERqwz0OqcnKB
Uo/hf7EiG357bZOG/FdXY9LxZ+4EbCXj29aIqFB6wB+RwJnodbX0GpHL/erVX0O+t2JQ9xu5x0+S
kQNOd2pzW94wFFx6e2rR6LEp2z4pgLKM8MCrw53JeTg6MqOPJ0hw8BIS/Bc2MS/PNg8XzXCwqPMx
NMxqMlBIy4jfw2B4OYEy9jNSnjyski4erOWswoZqYbhMBRQsJVvlBo5HeCpDp2z6gnfZ8cZjAfm1
WS6tbuXpM9mo5Rsdh0AMTfJixRgbQE4q0quUZRwdnQrjY0x3lzbHKJAi9gzTotRfdCdgwa5Lzojx
fM0CC/Wm0b0OdjfZoRqtM4Lu9HghorICZSEQZnBWHNrSDWSVG0iz2Rx+y0Q7etgRjhcGNLcmL6i0
a7LXkupG9npIH2MB0171DgJLSFYH8Aw75J1mTT0j3Ren8/afjmheQOlse/G9wC/daRpsBg08XxmK
NWAtRY/qC8MBDpqVRdSCYq5smYPYuTkL2FVXJwGgAGkUYOTGWCdit0qsY92SCINYIKVLznGwV7nZ
PC7SIp91lxuUi2I175+0hdN+JndaIff+tkDEWu5aBSrbXCjsqgWnIX0k1noRTB1erWMTvZeuucxN
Pa9WgHyldG0rRM5MzsKZvvIZdX1pBHAT5YNHu+bngK2U2xcLD6uPnYSN4tzxGbw6MRj86Mi8FhX8
ZuHrd4vwsnoX5bFcl1iiZq8amiNwqqPCetQatRyYEPP3XhD8OosTqkOr5YxCbgvya2yzgUmflzxM
IR3YSFfPCogzU97I655aDY11uppNblEJWN4Ei6lnwcoOwEkew7hbcQANKNLH29RXtrMxX2gEtPx+
odW34jLQT1TcEAmp9sSzmWd8HtB8PA9+0rNKPdHJ5X6wLefL6GnY0rZ5MVjAOpOCV4dcvzlr1svl
hDH99gztREzbhWivGom0k2DOyDIg9ZY+sfzyj6zFXovfkYhPNLyNdBWaPmYlpNzpFjoTqnir/+85
Iw+4Cj3MNPnVOZyTRjfVqQq5xtDd1SjGtdAJizwXhsZ+pkssENIMthaVdYVpH+t5YiWeMmGRvCrh
hxWkIhyDtMGKXyvcFVFplgmMgEDNU6FIOUfsTXpwOwpFXImcl67p/Tn1aYQlnc/5roih1BQqF8L5
b3fKjyiSRXUk6Xf62rUpyfRd0K7RUAxL3LRh458C+YLplnzvN2Y3VptSg5v6MV1XIsuDnBmFHlmV
pxo6nIDZ4enmiBaH0GVoNT6aTrfP3NjuiCz83gsv5Rs/tlQiP7xEHuU5VXhWNuN5Vu4G0Kr7i+yu
TbBHj1ERtZZO7F4zCL2bThcnNC+d3EKs7q53BqKQa8fMNr+d7lR+By4ta6319lttzzZoaxCVgPRs
PRQhYr92TxDQQ0KNSTjl7EVnm/0GtM/dBBBsRZ8FbWuYOTukQcwPNwfn7b6GQ/q+4E+ZCeEcimXf
34qEuWUxARPM2o04ESHChEA/NsJy/GSWRIDKcCApOqVFLNfJuC0DHbyf3orSIZVtjsl0WidwLYeP
Q5p933oLuccB1xRNetLHHSg9Q5nsOWZrCrPiZ0+2oBqvzOhEMTHc/giZ3JsCOA9aPhDC/kW4CgoV
s/a8n7PdN2Kio+Q3hTZaSi/Nf23D5HZ1IB8Xid263iGW0q36/P5sZFxaPJSy99d/GjWr+n86k2Xn
Gpg6MeUXp46gSdV2uBPelZvD2wv3KEE+gBKowi3dYAjHGvTqCCYODWYhLU/fPo7+ismYWXxia91F
JS1A85719RaEoMLsc3GLvnPmLoWvnBfqRLXGgGyL7F7oa5OfoTTBh6furlHNanXe1z9AbCO5/rBi
bm9v99qPSyjKTM7b6jM7bOwSVLvC7+pFGQ+p21u5O3EyMLdhgVabX4feKJSPnKBjtH/PoT9HMVq3
3X7mBtc4DADvMANGpkcDQY/Qg/YNAnAXhDi62BoWCkcoQykfuh1m6P3f6ozkV8bZ31Zm0AK40865
MAtJaTZdE4LAxo6wMYMaFk9si+jWgo8F5tPP32GsbGvafr1B7di6Q0dje6Qvkc/7PQw/TRsCZORD
xJfRxZ4okJzNEP1TpqaLoCID/h6LKA3IMXTtew3YJBB/MrXsLKr11GztxMr+DisZjUyttm17fNhC
2a59equYZUYicdU41oz+Pag9b2/x5brTW6aZTSIhLG8nOBU0wBHbWhJpsgJ81MiVDw/YsCkYE00q
yW2tjsPEVOgKHIe2Y3GinhhYp4sXxf3iTsdJgF5z+wrL6WuQBcZRuIBFZNwwfCo+ENCfNAYcNU+K
ONReZFjwJaJeptBJttDA2T+kQmRqYsrPFfwRi7pHrF+pjVVGeH+ZTKq/3ro4aqdv4+P8nKKUfB0u
Fn/R+lhVJ3Fm1O7fbMUPTKBG7+s4wRVC1QjCrxDFmzsw6KA6s7HiuoN3MP3jjG7xDFGtw75lShlz
62HrF+Oydvi+gurAzyPtWwKNuwvDiBsXVr7qpgRk/06lI7KY3lksAkSL9eLthDlbR/ShhSyPXELy
uXukL7trsuI71IvAcnsDAwVTID2a0QdG2ihEpEYVr4+9Pvk8QGV7ogbL5uwTx0RwEAEI9848sxdR
34CsRCZOyN84+M7UpXRyRLlFoLKGYjN2/7d+pY4ItuoGb9d6IHux+FkYLtHGQu+eSnVOx27detuB
I8p8g48B1tFcxm8svRWh9eeslTxJ7BAbZGO0WXgCQYwwW102PNSHIxuMfdDCakXn/kFAWaYoffhV
a9C29n1bejyVIRp1lDO95nTQHtKJTrjBEAzJRt7mIUVgWWDVK7p7UErWy6/CYVDrUtfeLiKF6jW3
DgdLh0kajRsmEfcxfx2ciKxSoPr5BFa/5BH2SmZrppEKv0skTwu15IaRMRaukm3HPRlzwvfxJ2AA
UrzcZNBr+nMItSgQV5dL7dKlKZr1sPXA0E23J/DeFDF75FMCcNcMjXQGH/JtKlGYuY9xa9HlrG2p
eoXsQU/5PX/gv9EU9VpOOZuJK9W31lFMJUrQhV3xO6ghVv95fVZfgxlbwj/EKKuCij3Cv9+Tr/K2
3mTnJZpE3y/uwjy3+QYJ7Pr55lwQiW4/ox+ym3uNdnIhQMwvelzLjxHjzu0cF6yGSCjvwlWYhPsx
qG75dsodSvpdX+vztlxqt+YjD9K4oQFVBFtK9xMoHzR2KD9S5kh3Sjxz7DtHtmtQOsZWCyeO1nwt
a297a9jlo2n8NLzPjXcMfZOSpvwVxPFR0laMybX/9tKGx5cao0t470d4BP17rOwa0ordTdY8Q5oO
qRGtinTJz963fGoeDzoX4nC5lo4TARWnoNE58bVkXqM02n6hg4rlRI+TtQ9Q4fkFPWNzLUGEGebm
EPKJKjR4UccsYEIZN2Nb8G3Zsn3l8bwrTc8Lo9k596OXenI52hqF0AAIr8a8Acie0nv+ASkPdbPn
9vOZZg8zBnlv8NFwbRr4zciW7dTjL7//MPIjf0L06midKUG4mOOyFk5jytnoCv+FpH3QbUFxo8gM
xSoGuGP+a5YAoUcUcOaMrGeSjXSx8U02kG3fv6+v1AuRZsi8ol/+1qXObvfzNVLRkHiJHu0hbtRw
M+JLXx3Y56IIVyzuE9e59Cm84MtsT2POwxf9XVhLipMiukhg2Pmflc26bilar8GOsSETYZFoAhk5
+bSKRJ4wmYE9NFvRbDCOVr+3N7i7m6LtQVIgT4KhSI/iqQaWh/LABsRFTKXk6ZPCeD+Hu62cutpP
2lIAwLOiqIWbzJdhpldvio41t3CfyJ8uJa20XVjoXpggP8C2qQvxygFhFIfeYi7Y7K1aUSD+0/C3
FSdKHHITpVL5zlVTFxrdDTChUzAbPQc8m16HS++q1DKbcYl2Qi+L7IQhF3AuSyAnQdnR6ndjgyiB
zi/oCVLCmRq/ImqDMh7712ENFRK1NSZvvw5Anlh+oLe35/MwatZ/LZ/Rd8V5PtSQiekkV450c/XB
RPJk/qzfa9ZYHDXyFRbWJPUy7SLKgB7mRXFeDHyyGODjvZZGKx905zhnV8xgvTthML3cYdGFEuRF
W1Tkvs83wq1AptJ10Y1LTEOz0+E9CJoj0VO14oWDuJwDsux/3FZ0LQF2mVDmi06rE3+Vud1Qy1Cq
hJuiyydE4FdgyBymvDUf34H7HDDf2uHkByrHScLVRMW5pBzYhRAATuMAjWPtpjVQQmVr66FHoo+2
u+HB8qaHxzUw/BGqO4LqNhjt8+8MhWsyzmkzP0Pi09mEeERoynOWMOHSB6k7FPHS85D/LGvu3mux
RFMO3kQFUWkryoQntyxazThZsKutr2qJXkWw78XGPgVm0zSkU2qoWAK32Ac9X2ggVURTxT2Crhih
kacJ4QWNSn9/gFuHsnjZOvrl388k5Xk1hjDlcUMyXcY5z3M5xxsOr8iTeDPL3/TavJIvh5MQkvEw
ikrCjnjROVTfPyO8ikw4V5o0pQrWto9srSWOWXwnQXgDNmiHv2+705OIaUQjblzAjqbki0XgNPc2
z/civol3xrt/iEhzz2oitBw2A1rM1DOIllwNC3m3VTEk5PFOkGH/EjoEUQwJ94gxRbsUUWe3UAzZ
2FbVkCX9sN4qmNTZUTxBWzobjhP6kDAxf8TaLq+g+cXgWyvJK/b9QRHuhuDDrohDGFP7W3AI4xK0
VV7NSpvReTAJClAacea1swSP4li7nP3jKKViwemNp1ssL3mFwmGDRsemYjIe8KcUMh1IJ2GhjXJB
HEQ3md8LJpBmAxHUdxuXoBg89ce7GCaVEnj4MbdnQ7BviAbpFhNs6TcrG9D1EYDaMbDM3te7ud0t
2j6xq9O3EtMgiF8V1WP+Jp5JsfPXQQhO1KmDzrQbWUoSSA2Gv2JcgUxPIrxbzY7yeUBPbm0wLb7b
CIQ3+m/xV45KV8Rivbsa28bZ0WMVfMokk3gsDNGzaCaa2spRP52uRKaYa84KGNg/nd0pU+dJkSK1
VxYPSH0ktqMY77vzn1oCcbQws4PIf7fBdrFvChxbqPpCUSI10m8FAwHy4O/XeIHUe8EwUmjEgobS
2Pw/lGBc2mKsrwWNQ2Q+akoBxC2vIVIJJ0ERVi2iLc1xjVl4SzLw+zyZD8GD/BShsCadkQGGIbTu
Q/FR5D6HV0HIX+sCmel65Sdm/3SsKdiAHi18QR4A8oR5uISW1ShMDLkC0Ik9hHQIh7AptNtZnsI/
ShTmDy+G8YVggCKbtBWEVTO1VngLgbWJaAlPxPYA+UbmVsd/MD0Kye7EUZCYC2Z+X0PW9q7TXqbK
5DvMg9hD/z4EdDOurmPnG/Xlv5k/Ek+nfHabfVPwR/avjhUFjsgzufiKA0FXGmQDOsZwdXkB302B
UpsM0lzIyLsLV5SMWIu+0UMTr8GzryR2qil5tbdDkTfTekVyBjFVEJ3qLWQhckr6f8jjpjm1VadC
MWQWFNWUsvYKNBJGj1ZpAtcS/byACUtwks6AqmaR0BwlbxNedDnM+QzjlonVt5eBjVz3WGl0PTGk
D0qxF/55UdDnWL66u5hbI4aINtBKoOdF+HBQduMQ2INHMGw507N3t6LwX7OxbC5Egi/0ZKXm1KQW
6dWJN3MQqHHByb2qm9QrWbPKn/uUEwy0rm6zwJRaVVOl3MrGkEvfbbN1UpQ6rifkDAHkahazJnfV
llaa5XtPWxsIQcijc/GmrazPrXBvVRCdNu7lHBzhvqEukOsdApWfDJXVcaU3O00+ukkep87Uxowo
gDAlBkqa/UN0lrfr7OMVLvZdCge4OPl1Ag9CPHlkz7K96rBK4C1KUag328XSjiyR8Rzfuj5Ny7Xv
ma3+glPialfO33TegQ0+a8P8MLimRhG7gFGZoUROWs1rl/qOxiM1kWeQVy8YtxSYVlrFUd13h+Ux
hO5QW9AjEIZgDRad6Wx1e82XV/Eer1SbwLdW5T55LoOz3EevW53a7JfNT6qKgiItwntXZlwTb/mm
FhBTnwMMr48T5B52q4L/7A+hExmjkSuLqBUf3PVZGjSrKk+w2XcI+sLef7zjj2KCk8eMktMU4Ze9
KwEhxyTP3ET0orHyx2fx0I0f4NstfOx2CQRq2GTT57zY3ZhzsJvWgUxe5tBZOkp1tJEfyeEj78pF
y3QARd+2RVoSgIo7SzubDFHmuVnJqsUyxoWtAJP0/rmPmqWU19yK0i+dgD9FHbTeMGkgGE5YTVFF
DFT/QDW58EPD8yc4dP95TSrm8JKj2pJvd4E2UtGtrQMzH5K8FSapJYDL1ZxC+rSy62myHUxux/sf
bextqa1rE76HyEu7lDM4s71fy9uQjwT1Ys6CZtOcCWf5YlxW8RQX9y7yPJVOH2N+wPfOOIQnLJTf
bH5mrTQOxShXAkxPBpzYDUA7L7bzQ2kbDv9434YgLQOFzrZ3O03o7j8YiWHJmFLWnLtJmU3AUyEs
6FfBgsLcuNUmRd/36zhQkpnbw13Wi9z+q+nM/aXIB/evw4YeVG+zKqYce08nDe38xOi6BE8gn1gJ
2x0/pr9rsEwjnQu3FXGYydGue0nXYpBfZFIrWWvwROFUUFzVAJpIZlVlkH7/EJQQyUadCDUtScJL
RrhXV1Rl+0KU/LHjJ5h1bHKZ/yMRihlRylnhvxS4g0LMP1oiv8HfkqLiTv8Z7IMTD7Dw12QjyTDw
bPh6Fr4tazsN723HnJSprBnnCkLn8rG58puuXRwDJCJkowvoJOUHYN0nPbvgWqXks83DMjpZ3GnS
qh/lPmYag+CuvOxgUWcJE/kODOncWr4ZLOMUVmGI9mH0GjB2Ahz1jCittV5pZukWLdvfsBmy1PYT
0jk3uDl5omaeQknKgLBwSiAYsrjkXBpPhGyTQeERmE5MDcSji1AasgMWjJ+ca+Sh7JEZWW1sLguh
XsZ0O7jcyMfncl2V6mUQOZj4twnwlt5c8jY2TxdRh57BUjhuoGwgi2suTaCPpRpKSMfDF53e4GCI
hvPs3khnm5dHc7LZH73Ai3NMCRFokLlGlwxO1RD5EVijPc9mEt+C521VLl99bZOW0Yp74REh0Ppt
I/3N2LOH8KZjwca1MFfioqnQHtLLCHQVsc42LwPT/vU9mZgrgBR0PdxBfKT+uLs73KAtGD2Vv4j9
966K6e6/V0GgMmYsnNopgCzTgH24MS3wsA/cDmLcbUx2aFSlJYwBp7yKaRz8C6oUijzivwCPqsET
wrb9kWKxbakEanMTCBJ/RnhRMk00PAm0mbIAuTN4cQcfLZuB8NyODAVFTLxR3ZD9/YUYMKbBNhPJ
e8S/7ke8avmbQhGfAw8siAF3PwFUDodZmJpXlL7Oz93m6h0omE2fuspebOOlgfYETMu3X0987Lu4
lPkTwxCfFQWXfGKu0IyI7pBRmJnZ19iQkcFQqyxuXxvETmTbanyJ/YDv5U/og+bbu3ERGcHN26K8
Bmb7MURR13gQPskEFNDeGg3WxryxZ5b2M6zoGWkEjFhfJf2yftERwqWWVcmNcyJhT9Ysm7vmlqR5
3YIQyz5BSWscwINztR3S+zw6ejue3+zkrFphtWqK3E8X74XESpwAU8RXnihtQHas1uWYHNGjCozv
JOM1IvIkNr8M0xMxx/5t6L0PM1LJJAfB7n8vJJHOaTNZUl39AhbC4MsC2/S6AzLQiVlij3VwdmKb
/Gc53pVzfc9/CxVn9ySihmySAZKrZKE0XxcDMbgRrOSPMe/nfn2wPpgIlN8jK/4p+3nKRRYoAqKa
1j/67XFDv+ysFFijj4KjwwIYqKWXAzZAzCrp6MSXeBY3CXjXVsDiRjCgyBkzxBYn6l9KImL7jq3c
UVI13C258j5uTQxxlmGuahoPZzqjUZpwWPRw5F0VWnfR8HY/ZUdgEUbQerTQ/zxYytcwxcDDsemk
AcnjHqhxP+1d7ccuGHfX+0IMzOIGe7GNLIYWetrwbS4Zl8veZIsZ7nsA1NGTNOHeHdE/vgCV/FWk
Hce7qnmFu07pZRq0crgKtbHXaVdSFFDwLOf4hmBWGGsaZF0NU5Q/89I0PTT/Hd6sqybqwMY+bSzb
n/5VAZk0g85ewcAHn3a0QXtAlg/r0CmGsDPtU5AYfruFvrcFhaYr2zCuBJCsLMChjlwtjzmOShn2
gViUkvno4v8oaESM+d2tvfI+3+HGAn5vunRRCI22aJjM7u/kn6Hj3rF5fEO8MOSu7V8utEmOH6b9
8kFshpvmlRmrKUhXtKc+XaHf7+fQUs5rWmFL9yZM3neL3hIMFHMF5tRf0UcHmNdQ31Hx+t128B6h
pub+qM/StWt6FAg61ze0zLo53em2i4Jn7L3bKgZzxb3R7y8rKyiAwDdocCp74nOOLQSKZhcrbGAi
LsecMhzouSjA7708R1/R3mdsRWFijvtJRXG644F7PRphayPHkCFqOIkuAGvGIItwc25oJytjL9tX
M7Di35LpQWNoiNlnlq2DyWV/rOIs4go+l8POhamiwZM1iohI//t0cRHq9GHU39LQbralp3cYip37
CcT0rgI2OQDKVR71s3sj4ZwYLTchbcYCxrlw5YnLqrBa9m8lnFosNl5GvrRwCxVvVrHf+riLDFai
HdlkpiZbD3YfOttvS76GWMDraNptsDd4tBsDud898aEh1XqzkYJ5EsP+Rr4qq5pjQ8Hy/XehqYgG
nblM+okcrUqzrKmQIYeJAyDYD3t5qxdbWECE7q3eDksjzJTjGFOywPSzqQPFbLp+gXVWs8fQB+G0
xU+1MgjkxB0K8+1J7bzWVOFn1FXkRWvVkP+o6mr9usZ43M8CH5K7QBoV2heDk44djcKwoZ4KD/lq
zWdKCR5fJjNbOmyl8qdjx1//QYBFMibBSOvN9QtG5UKmw+KZiSdkU9CqyEls2s1WDgKvCyldrdfZ
MvKHrMhoCnBf1gOdWo5JK9l9ju0RL4+FZbcqpg5j7abBWeLqb5Od5W5vtI0OYXlKOnhSMLiRRqaH
9XD8RbQ2/6rYszNZqc6h7CqpJeAraxQCWG3NPdCkK5xSHSSmKtGQeXSubaEFAC2fTwdxB6Px3NLz
ofHe6aXn57nPW0trlYW7gZE86ncggKg1dUy2FWlEUME9em5o2BIsUv8JA3G1FjszfKkhxvfjEJAf
uxlWr6R/h6t2HBQU1C0MJF/LMan2RbhpNY/qNn5aYBil0+jNeU7mqzjUPAeloUpf32URE2hZKXMi
jPSJft3BP7hoBrff0w06Pw+93SbNZYMYdFNe9ogN3TROW3KBmPy93J70RgmJJhldMs2UqzqkKuax
6fMfW/ro3sE8EvMyLny+CzP/7a6wKz+SuZ3VP/jJX7uqUyqmA4vxvfAEQv8p4q23u0D/6naGIxaV
0kdHGRMEBjPw+svTakplr/0jylKN1y+64jt3P6hFlEKWuUdnaGHTu2Vt2md9PJ3bR116c0yzYA+c
ADHH6AuNV5IQNm/Q8G+Hy+7WLLc5c6SZF8hEkRoVbEgSxlWJXhSBnBKL0W54zCDtEIC1rwWZ9jNo
WHMEnuavTRST3va44CYBGwU1u+UMilzVnWaC2RJZAxRJ6qwnck2ETt/9blAClnSMn7vHvz9f27EN
7CU4t6zEDuDHrruRrMi2Kf+L5ReH8mqkA+1NFD/RrN1d9DJcyJ0LME4B6LSpAzSlAw+b/KtWzhgf
uNI47xpegteLFS13LuwdX58r8XkLHHDyy83vL8bdrY74Z2WVBpz2H41yqLH8FjAHg3Pk8bCMaJUZ
f+lt4uoY5wZTi0s8qXacHUDnFOcfO5iLYal0j1mieTcgp14WYbzJscZDyaWpeDVLokeiEhBUoWpl
9blU2Guig+ifUExRcnDQIf3xfkMoDL03MF6XHAP3d85IJgaDRTXe4QvyTNTZk6CZPuSfxQJBol9V
3I1hWbFBCgR++SWEPTYRhA5hEKF8DIlZZno7nohsgaoAoV2rOvM0nHxzndthNhwo3Ivd0EMWB6kH
WWUCcW+piIolxy7yPAxwoTZG0Klb003tf4sjTPP4WdR2JvuNgEohCmZoyLxiinC392BDYlzq641P
aR5h2CirCJN88gcKTnrSbRSskS7tSav3FDM/KigCqj6gNHCmYQr/TBb0yk5T29PcVOwL4t2U7VnY
noBLBQ8Taa8nL5LWc8zNrEmlURhZ+XPCngw74/jgJD5KGJc1vTXolnh32jPnp8fV2dEOQPEEouyQ
Rxb6Tk3dPsoRq7IOfjWXv17IpywrPfEp8SckTcv+2/Hq6DmhPFpJAxmZqM+iIiIJuAIKfizilIdf
r1qeadmujMFlBzQuZe6zMDU+p18nEcQcwt3fpfJIq72WxUg6T2jVHPBrSljRnqOvv+6m1UNTHmCJ
IqMjBUMeYh+l5EAz6Dg0aTKjhwWBgi9RcBxR1YCifu9b2WKSDVSFiI9YMhNgq78J4dy7I6pKCW7O
mqY0x6z5YAxDRqZBw/WLAh8M4w1WDg4cA7X214mg2pZ7j50U5WajLaTDdJRAMlekhp5QeJU/3tNZ
eaiD9wVjSdxckepwGg8X7OnCTHQ5JRgg6OucgR8Jf/J7tPo3D2sPhTrKaMIG9ZxAGzkSEx+g+kpy
G6BgtwWZMgi1ZSKQTvh2bfqdz6vVal33npEXLgCt5BgQWlMYqh7+65ZRMswle/T1ib9/f/tKxVnx
oK4Hvz1OSTeAYRjI2MC9gNBMybluISw1PG3gf8Q1LPN+OmEGDlJqSB+WivLXB4TzlQx/1X7UB4jD
PGvD43tY23d43yyVcsO2FocLT1KNziQYYrjA498FXaZpVY40CVCE6Jx3+5PzgzWkNiOktIr5YyVa
TFApKxO8LXgKzHaMk+XcxtQVvmSSk4g2yzK49vSkCWHcJGJQHBzFiI644p9QWFWGqkBOMuxb/dvO
6sVdDnePcsdwB8rImCmEN/aLKm23jxvSXnz/zp7GLFt7npSepqhPm5XehZHNU3SUsFoDqnA0c8Nu
4jhe7X3zdSnoF/yZx0W0uNU2gwsiMQOEg29lrDAhlew40JEQYHN9u3it80aQ8HQh5fMiZUGy2ONH
mb+ikTo7fttGYaeV+LmRHOYGLNg4TYH7c09QuHQX1uMkNx6drVmmAXjj37y2kpJEwl1TgXlgSXsg
bd2L7ZGcpnDoTUQu78YLC0E6UyUlFz8HWgCRzLdfARtCkCJ52BGSk3DPWS2CGYqnNikLnatjd9EZ
WwTSOYWfSPVRbaslRYID/yXCvijIekYpsltc+3XmZ1VycXHIG4r7ftHWPK5hunpSNGBcxJWnTUJi
jj96xkfSaU5mU/1vznf1/alRS9G5yKlEco0QRQhmm4mJqwmNtTIk3nH6psOUuOLaLE1l+nVUZO+p
uGVDTuW3RySTqY0XsTfZZ86S9VVmg/c+PwdSe+WPDhJm96OdQ0MN5s+3wJkwYEIozNC6mob6hIqq
wpl1FoW8tfwUNu/tOSkV0fB0rOXw3AKswyE7uTTg1JuS1mdw/mZAiepI+fHu+AhtKa/MM/XypiZO
HvRx9XC/MrDSqpt76IT3ZQTXLyCucqQKqy58V8UMdB8Z6uUkfz8HEhCAZflemZ5Z/YI+VRimb1yD
ER1lqlTMutC2nOxHj0BJdNhmVaQzJmEZJD5uei9tr8Ae1Bis4MLurfHy0rBrn7tH2EjVKevfQd7m
y2nAzU0QSgTq71acOQPaMewoHWczj8b5c7Xpx87F43bLbniEmxrSElLeys4rgRwq0yofqjDF0qpV
qbw79BQZkzuGJyyAyhOBMWRiqTArFPoJ53AEGfoCFQgM1lK8titWfRN3Gj919GxM/GRHwcRuhk5K
Ckf9DvDzQxbeIdAimNOFOD3bMHq3rf0e6JkxhRDHHohtszn6BLGXnuDUmn7b3ttaAZc/1OGFtwKP
la4HgX0AgHM67ALjbZ6XUchGl4Pia3GMreSQL3y4ozg2iDU1lYizGV+EcbzxpwHIcczWAvNq3zGr
NBVmjIlcl32kbMO1dY8OMbjOLda69qFgE9KbQsejIMjq7h6RMNpTGO+15cR+injZgTXAGsCG+RZZ
DWQmkZ0fzkU7Ny+Gq6QD1gW2OZSkKNa+EOs2i65D4Ly06Vu0Y1Jn/ovxDf0a7f5WocbAWV9V8UiU
aeXobyd9OW2E7wfvS7aNDb45gJzLfsz2I4l9OPtIinXPh45OGbMjGPKbI3Hg+1sgXIZlwnUtAgYR
a74Dhih+jgtoCz/52YhBDFyAihommxnIaqQykL6bYFTUJOQyaff5f1Vt5AJO1vRRGtwUdvTR8cao
XqHh0CApDKkmwo4uHUEJ41Qbhlxf/2mAPtWwNhHFDcri2qHBNHYKM9tnM/IEb7kxQzO00ulpCOJa
a3WDvzcBPFKw84l4PpbCvOsN0/th9zKck2ACGGXjcZSdPoCTgDxI2Eu8DgXS2roENbCWfb7yYbr+
qEAVo7heOx4aQZTtIpYCo0dqzYL61p1QnAv2lhKF02dYvZrTcxjf0u/WkcG0xfj4tV0/PDf2F4Lw
GOODyS/RoaR+uH8vIc9w4JPTchGTsg6y812ybiFuXJAknl0hdmRcqlqJxX7Sk8tGOJ9pr3QUVa0N
qKZIKyTkOByRmRV/H30Na0uAS86Ohp6ZagSwSIrifwkNphXV/8w5DzT1dUBhrrs1Z5UNW1adEo1f
TVFGlSdg5V/xFfuFADh5cMEpH3QBKFR3bdvvRUkJ2iLwVfCGql1ctXN1OwZmft7e8xB6lPqZqkRU
3Ky0pz5AQ2/cgfApqfQfxazmXn4X3ijzab3OsI1NRDhvdgTOSHOAKB9b2YFdAv8CGsvQvtNDS3F8
nql/CjKRqrHx1hwibFcP08Njd5ySb74gjS44zQuG/lgrFsSsob993nvuD5rFdKeba7XeBO3uR4MH
4zCjGHMmeNpuQgFgV6get8unizKvT07Z6XUptJ32enY1gyIq+frLhEjsb6bhaST+SgRtcI0IABU6
cJyOr/As1wt0MWB9CThFHPm0TcoHGYFTE8xHrcWMmOnN3o5tLh4zkhS/mOxvi/jsNjMS2ugApxqR
yF33CgY56XqwZIyuXaVRtl7mcMIkRAWDrWPt6IK4W8UoNsMbMWi5NUmmMSWm/DwXUzU9+ypQScjF
wzOD59u97zdwu/czNab1MIYgEKRCZdVIyebF2h1uadgzvZlg2UlFOyZrncmRfjsa+J+m8DUNCRLB
8L/J02VYrW8CgMejp3vOriGCIY/PQCXXP4YuCzLJ/A5cpGH0GzMQnmwk6IAb8vG6hudGebGZXJER
/LDSvkkx/N7eO6CGXT7Z7PmYbAu51yrpzBpyMR+r99n2FE3nLVz0frFHuVLC2lJYp5rewtDYPyA1
uYmuywJlyWr5noTWvRicFa0T6gya0+CYSlz/w9cuQYUzB0x5MU/DR3ryU/HtHDkHthvt0X/uKHKP
l+SgNSqB8clsZkBzJFSnO9rgFmGuvfo1d9QnDQ3eEebwG8E/lThU1Y3CDUTYvC/BFGghDMrlx+JJ
k9pxZ3bI1UWxEqmssBwflH/S8plBglxrAYsHQxLSYCtSRLl4oowj+42RI2k4dLx13jX3+ptINtV8
n4n0Zt0XSj+84/WZaPGYRyLjt9juqQbXhuqu4OuFgFmO8Tj9MYXMs7mjkvpdk0p9kh8fYA6eAoq+
YipThJTHz0LelqXBHz3Atr2v8B4nOXcDpY9+YDrFcWz+MwFz0AsTxmvsyyYsMFMhXZ+WsmJBQaZE
jepHY39jzYbO+2Qa6XvEam434oB0Fxg+FDdkTsSi0rtvNABqs32v3OIl7VcXZRFopFj8vNP/kCAC
iWDcxG+b+oAjuURxYOoY3mluKJWqv+QPm0yFODElyh+UoDtWJFy2hDYvBuhfAKLNhKl0gqi7zHqw
GDt5bqn7emHkDvYmfCPYZd7i03S4jjL7VLPkLuJJKdW9iJdUOl21hZLCvO6zGD8kPNCexEpXHpuI
GCchSJfLxQctD6q2vJf4S7bu0NE7unly0B0wcGWmT4vDk6uj3fLTZ+1pavpBzwWi/vrAkcMQrEV6
cuWOFqx+uAHtZQOZv5zsiH5Z8pKcgtM5f1CMAqTsoNg5Gzdql0VPpesWxY0nlxqyzUFXJFqpkbjC
92uIfDhSUSjQX85bDUcww+OoUVM+i0Gjk7DHCE3vZvD8t/a58+/QzkOTTDUPzRcFy0PUvqOEmFop
wapDl7qAl7CRdUWZg/4egQJN0fS8MQmAPJIPefYt2lSs0Dm6cYy3j7wvdFU92mResTS/QJN2k5NU
eNVzu8oW965HrEnk1DRoQMDhh3sV6KP+lFyVneOirsoBiWTupfLEJA1sqOLEY/4KZwuUqbjSuop3
8OzKJIK/x2wN85gqLYP+1UfLkv6CQTgG7LZkG/BlCODnNVl/IRCMQ+IAcpeUzMXxY3qAEpaPig27
6ThuEP6LPRYEmIhekeUtqzvHTJhAQ02JOHqJIXb6XNdxmAj7Qzqf1ibAvmVvRdlzChaZaL+0XVY5
M/sK1nw1r5qisVuIZMwwz+tHx2lgFwVXTGuhk1lIK8W1NxQk7u+EWWSb0yRy2+HnsYgY0RCSqbWd
StJAdaFDkQD4mDv/kXUZGtWJndgO50X7Z9bRMfWcJWi2At1imI81Iwafi80xGMnne84A0T+Cj1Ie
7o6LM10QTVeZYUUcowsEEOa3eZAb2s9GYMQkEKYYLB/xBjxTTLASTltzVG/yS5cnC1nsc4mwkb3g
enLaiz5K0eLa8zlVGa5wZXO5L7L9nWya5jwzfGeMcvm88faTjH6E9k3mPVU4bBHHK9L3uVXaF7SI
16IA/3oUMc72rxAvXjTIYFIUXxDLM92PsvIYmDc8BX8sMB2N7dcTGer8fVrEAG9RWvyG7+7DtsCJ
GiqqxieJXZV/7qczVshzCilIww+DohXRS40ioZRAKvYywl0cUBeI/DroIy0MxqjAos29bOpRD65X
04Z9D4giGBbpQzINr9/YbWprOeplBgWTnHX3EO8zoUop58WT2c52hMKcZNFTl7oqWcVdZtf5cN1b
G8EZe+AJiCrLsSkV7PJhqS9czgZDeVngz7D4iDCz4EgSnbaW37iDoPWPEETgaTuQqCX3Qgv1/p7B
iz1NV40mo+Gr9eJDOjDfrr3jlx0ZiNEJAK68OsRB2y23AfCOB+IQNx2J0Njrkw0rqPnSeVbcL+GR
NK2pxxoU3o/YapLt5aAfTqyyVJGQ0ccdgIQKdwklOD5y6+o6uWTEmdq3ZI2YrHNzhvHsepJMpSjn
FgJTQiFSjPx5IYaU4MgIJU/ex1pmP3l+bqro5ZzJaxntYf5tO68GYQn6TJfH8Dj0hZYN7HrPksjp
wCIIrOBmivU/00QgsdPWpuPtUFQd8vOb1pHUzUrfU1pUy5TynsSn6zXFpNCOZz+/yAKhNrGRa7q/
9FqWktkZ8DmNqT3tveI6ACWzA1/xoI6pqU/sij40VAW2B5VhmY0xyP/Wg0isofCu0RlnuWQSdZNd
k2kLF1thbsi0yZYPOIMVhcAaJTC1L57thnjiNPK6TI/oHhIHfQv87P8WzlbFs1bn4lnivJqrxVVR
IfvRAEqMF+O0D9m/JMfptTKYx9fvUMbB613ntNBsxp7IxdVvjUNoyuFwM3Iqq9gbsbiENkf10bS4
F/a9J25gKkaSSYP+XgzuWZ/JlcrcgnjN255LBbDmOqORtd1y7onh2ipSO81nd5koypupaofEnFVA
/YoevQlmTPogjYh7SzZ2OcucMcOWa5ZNt5Ax14EXwJDt+aqXmhwhMnkbnBd4hg7leuhDFjkesW3Z
MD9fas8wu/LK4j9eoJ/962kCUK72ui/BBSX+/+kQClhCeEXWHnHSge5wBdijaruCaD2xC9ebpweD
SJqNYAkDKxapxa3wWc4S/NrsGfoyCwyUMsy7MCWSovwVdi52tsiozVtsC6IPJvzm/WQILT7vDsys
SPrx4VKUiYXW3AzW7wk8UvyhGs0OxkGc1VQ48AJC41j7/ZNdl+gnTvXKJEPTstlu3xh/lrz5bwTR
pBNXQprGpBDX2WiycJVBiD6E3BULeffmS5V1EyYaEdUS+EdRzDBKYs1GTNfrBUmhnNASv62Mf4ee
OY7FtEvnmtRJqe7pDaV4ce8YBBGndrl2gemTJ7MmpXZJwi+3L2Z4XSp440F6H6bUjUgeewsTTpYw
QlaCX0LsqMOKenBXHNvc4Tvf5Y6XYjLqfPy1tutxRo9dfoW6kRXSi7czixLxNFKLvdBkiq9jPbUU
tR5+wPMn+/VTIFFaqcTFiNWBopww3+XeIueOeFeVXq5T5T2Yhj2nQWviM/+sqzJjO0i70+p/NoEE
YnUyLt3PgTsLLusuXsKSBzZY+QMiBF807XOv3wg3rjb761A66B7HF+KkJ82B+UnByoPtq6mxVBBo
NqzBGIx1Brg1vz2E0krsEj8sMQACAHIohUR7xvJWQYymTGdbFG42o3qxVMApCDWKsvj/bhiZ/r8Y
g3TmP4FxnAcaDaBaJ85hWfUSvR6773nMDMhrWQgryxiEZg9cTaB7O65cs6DR68eLr1tpfiZ3L/NZ
sfBbO1kHKRGPD62BtWo4fWvB2ufW338Qj9UC5Oq6OQ==
`protect end_protected
