`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JBGcQy2j1G1MgfMojkzBno1qTN0v9S3M9iWkK7KGNBnnOk+bFsnU/xy7X+TZF7bYaewiAscUKC8p
Uy9THyao0g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RYXQ/3NBYzjw1mRA/nI/MDMgox15TgJVSKt5K0AwQjFaOJZ610sx3QhFiOGRC/S6jheItfU/7HwI
A8Laohq5PdLQeBm82lZZ41APVpmsW5DpYy+slPxXaGekBd0VK7DjdP4TzDP0shmDZDioXCXiGbX3
TLhPwo9VVbTlQnGoLYg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VsrzcQLVu3a5i+2YFwmbNR+9sr6j/26fl7FHVb27gQMQoyf7e681BU2Bdffqo+l6eKlBDITHznEQ
ZdxyFqvl9ZSMwDbLxQyN15/wbmVXh7FrltXpgHWn9hxLFFwF/aw1DCk3qAJAABMSIZPcB5YoEcyL
iOzVyXAA0To5PhAEj+f35mWI1G0AoLutLJ3uwR5UZqNRnDcwnpkbSmwrGPmlgVbUCaTlBpJtuK01
mA4FrBsub3wScHUyAGou8zAB/OPWwCZlrR20c9vdN8pKP3k56G/QhHUEgx4EhCjm75VgFAv4hBmh
dzTVS6RTI1Y0c9hY4MbMJtHZcd4AgefuMZVGiQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eU+kHENLD0InHp2zQEiVQesaxqCh8y1ZJ0mW5aBJb6vZedMNuKr0K1EcfH/tOmuHC208+bCgcEBo
XQrUEY8GRkuYdHjyXb/xjHRLsMuzfXmRln5a6rnpb3LXkpKBCYUSfGiQ+lirXbtT+096nyhuIJUa
suoxpDAZvYgnOwtdFvA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fJWfokGEuIX4wu2EJ//Pmg9MBw/SKlenwLPoaOzVxaMeT7zzClm1LjBuom6X3m8zZCKj/gsQFNzm
5dxj882RlB1pdfgaCwFItwXHM8TCcNNRUF/2nLm7jZtnlzZdEirVQbDaojNGzBlibsW75LUatPhT
i+U9hx+p7v+1H3pLclndFeO2VU+HWFpq8t7C0MHi15CvXyHr2ti0SBBNlHeoCgFYLxuiZMcJwZhk
bqR3V9HHQdhibWriC/1bta8M5IZ38SLE7ZOWRHF8XZ6woovx9Y49JpvslPykCiEDgrBut2UQ1w/G
1C3dr3dsq1PXpjUoibQJqGmKFF00CIMNwEPmHA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7392)
`protect data_block
JvYFg04dzOcdRr50ZC30bz2R3rkqaFdOlRN/miz4zlwwzxUTX/x6v3PQA09NGVP/L1Oi33laZ9u7
yxSNMU6UUhh1QqYZM26c3Hf6/iv9aivgFeAkA4aRgwO5ertRKz+R4/Oyb7Vgt5tPuaBWHpvcVz4z
uSScYG/vBPsJp7gXXoHaTfuGCf5p6p9UAYlFHbJFuilxJxu5Umvgod+XH9cYRyWBV7wC/P8vh4Ca
HBSZUoDxvLC/VpWhhtqMpbS5mJaF06WS0EkxL1nQUcw6qGAVt9Fe6/YDwFBW0ZmehdNhJ9ZrLJ0g
DjgLCXrBQ1QikhCBhRUtK4SI29oCVMdOf+VHlW2cclZVL304M650LW6f/fVF1ffX9/j98ZtuG3s6
Yy87r/VBVbaeOikuAJ2j2WzgMBnDB1zHsEeFgJ79+5/kEVpDL0bCvrmvlCGS+VvxhYzjTkdqeSFF
nlJP1Wszy3W1lafnrvbeTyPtCiDmpfBooPsAxgu3k+Kogm02scAXnGYz+dWo8AAfN8l5IHjS3Nwd
wwWqvSXQejowTsyg8QhXUJG1V7kY0bINj4owBabYVKqEm3xXkGIeJd6eXQSIT2WredRLf4NHeQvZ
1zwh/6MowoWj8ksZG1ardlOpt25dv3Oiy2bxGPRZiiLjLIxrvRBs/6yxzxKW0Gp4ZMbA26ittI9P
ZD3ZYptRNF3oDwtNYFo1Q0p7FVBv62VG4v+DEQhe3oGg7WsUc2FHNlX05V5F9rVR0Z74+aAgX71/
loYSPW3N64aDPQ73h8fC1IHlufgDR1hyXHN3DQKWdaIXwGed0BYT9aNDUA2U8uqFg6NioxC8/Gdd
JAUEjhXsVGGjXtA4urlDWaew5DTkMCtNcLCM32C4q4UIfcKh+Rgs2sERfeZlghlMcTRSkRgkifnA
mm1E0509erJ8xNEG90uYq+ASeYpWEZeKKQpgyE9UAhy0oEMY9yIDRhZSaoasw0IwByaXz1HM6n/c
/fOCK/x8NVlZnHuRQ9HejzO+VsBe82csnlUDmwYfhmsnA4+ElFVRe90K/cgn8CVmGNVBDv3YsHV2
miQKFMEZeG9yN9iN7+TFnr6X8vf7HlQ4Adzc/Htno6NzJtLkmjLwxQNAOJpZAbIyjxU7fqq9rfVR
c8+k6oY7nMItHJuIaLWNiHsp7lvWGHdTCl0ftKOy9IpDgF56i7zWui35p3pZFpseaxvTUl7n0aTJ
StjGhEeS8Kk2y6kIkHJaeQxmIAPgxzfxa9cyfoAPxao29PVnEwncFYYBIFjEUrFWLiIh9gq8lGGb
/zlc8pkyzZFxJMRkvg4e3+mYWwfWoXfGF0/0Tb0CacoLrD8F4T12CVvtsFjzDIC9AW9/G6xfE4A/
S09JBq0TTp0wdQyEq4qDnSEHBi0X251Fb7M7mJuKNHW3SDpbZcLtfi40PIzXWs18I9Id9tXbn9ts
5CwpAofEr7QgxFOjUc+2Yr6WsK16zQL6eSmIEiPVCP2Q3OrDSa5I2/25g8QX8vrraNayN7S93t9/
Q2aPKAo+ZHiPDUPlP/X8xIjszPR5X5C6fYtcPdYzVyw28BcZ5YkFuf6lTJFZTm5gKA9Owlm+tqsk
c8Htx+7ZYAnnjPy2lyC/V5GRFT23n9DA5SnDgl6o5pdz73xhIYY6sF+bipdNFWRWLPh9dPCZaNX3
zm8WRSR1OFRJ2mahfipxmDdXpECbGhahu68X0Zzad6KigmVbfa6pyCW8UGthllmjSMYAKAgBu0Ga
bz2Xz413SyILsmzwVocxdAM7n82ExXuS9CKOvRjS6ywXPc4wiIrF/qk6XSqAv6Q54pIqX4f3c8Rc
AeDErhE+vI9Y5C2HPhUIiW5QaO/DPe3U0+2t5HKTvCtzElRqBr6WtgpanA11QQ3Qm6bJ17+IqtSU
YmuTa/W3GsG7RZcZveF6vwp1IE8L4j+8mlHJpu5W7PEb4d3I1bcB3GtnySA50YJbL59Tmo8sbfRz
15fLjjU4x/8bprdnSiV3HPXeLmaYU+5+TgciVdWSgel8PrIkbzA/1QyMLTYugu+BQcAg3m5WSXf2
gB94u6PD414/npB5Y6TtLwdQMNftVZQCth+xlhoYCeDh2DK+YXxlxSYzKWH4sTmKhtqxMDjJgjZm
HclOSmBJs25pT+Y6I/QWm4Yz99iqGZKOccNlJknXBZX+GriCrWKTVDeJUTMHNmACFpt0WWHlh2Jj
rrIZklfNTS8uiezS7rL4EEiVGj6bpSixAomsPQ0e9jwu+ugHi2ZH4RjCehUul2w6bK2H86LP/E9A
kXEhCilUwAkwKXSLdiZdpA4uTez7hqGGs8kUX7eevfQrWUc/ZmeFzAspRbeTToxoow1Xc5TBYcXR
Iom1XhpLG3k7EcFgLIsASJQLiv/5eSPR8FKrLCgdGRLUYL4Dshs7zkUYnKcXfFftohMFDx7spqOz
PUBzvArSS2sNehMQyx2DAv+Dxz7axwrtjCsQu4OZpxmdwCqfxTd1zoKLvLB74vHekiZwDEJ07CBP
P0AOJjRsNvj/Wgq6gCUK9y9dj59t1U3UQa6jnXf540a34AFcOGww32+Dc4ek7EVgOwWC7coz/p80
JXlDj3YCw24qL/YADzF8lpEtrfsfQgCJYN1NYe9EW6gtBMIKPsy6ho7TwrL4R8y5g5qNXoDqJbBB
O717GX1RZ6/x62ZtF3amPaY/YkVi+cUPAJMBT6jxf2QhEv3P+V0MPsoW2NC0V3wIeK5aZLtnTHFS
2/SnhG+LH10dDr21henpciKYsNw35+YHYa8iNUUSN8uh9/9mdMhJYiFSyOGiJn/2DqjuMEXXCRG6
8SMauniy07alSUti+Z2ZsHZZGBR8KXDmJluIKRdp48nnFYw6RAo8dEwAYS+/S1+LTFJYnstv2o/P
VnPPWV7v/IG0UhcrNCElVz+iF8P4d+3J1BDr1abRp51N08eMuHMN6LwuKE4d0WCo0/LD4oaIVI0J
Z8BYPeMbI1nhgp5DfGnkbZLfF81jC0phF3Q1izsfDjVJ4UK8+GWKo5OOH2wN2WoLJ1x/oOesVtK6
UFuJkM86KNBngu921tYSVgXzAroP/kOrEO8XNtCTAhdD0JCAzy5tra/SIltYklDwfIJHf9+4dGWH
4szHBLOXx10JHMm4oFYaHd8rcLjmudWfTyBuaE/6grpRixZy1E/rqDkfhE4QcZcBtzajks/aOC9m
TA4M99ztzwbjIJUPttUjSIs5FIEeazwuAMReXzwVIQRJSyKY72P4ye74mMCaIGQ5cJBb5EBLfJ+Z
XcIWThEhc97iY+xkc3nhhsHyKt3MQFVF+C6WUO903hIkpKbxhV7ZXJWlsMOrWmViqmadVaN/ras2
lDn6h1sNwV99BqvZfqp6NgFBCL2gUODw3iC4rygY5VaU5QwZELXJ+dYZFl2WPGLIFdtW/wWFzG4K
u2D8Pre5yEWPVSDcxqiaaSrbfepA0HRiSjrS0N/8JCykhoZKrQc4hwuB/1Qogga7ZDsQVkgghmyh
yVUGAsJ2vgb0RmmgfsNYSIhsFWIDEKZBjlN2iGLFTuyfZeIC3BHoqYZU9PdE8NTzPfbbQ1OEOZFS
WsiK6BwceW4WMwKyXqZg7Nr1HB9/4KYJFqcO7izZDVVJ9FKfSpNBWL5v+SFcYrDMDwZ+GRHRbHzI
Hp6B1254KLp/EZUEptcFbt53K9TsqF5VuBiAoIqXgclkJjXR/m1hdGWLdlhXmDVtPq8WLP9Io3w7
bAqu4dyVwJHlyt81dMF3t5IgdWpyaNKhyA0eyG1nwpvt7EhngPPi4Q5vfKb8Bu7vNQbPNgvscZjw
GXbF2Wy+TV8i8vnPGu6MtLYNYsvtruljGZqQZ8WYaM0beD21J7WIfjmWwydH8TwBN+o00CPX1zbP
stBIsikq5HMXVwirAJmOWZSisMZKBooakrNWoZtFRmJT35OwGn2rrYRv4w+lctealwKRqdpcVbOd
ofbO7Qt5X9TKPQxithFjgFiN4l/M/M3S40E15udSHCHBw2i3rlJDETQx59kooLGh78WYcuWgUSWG
tWOWL0d2r3UrCJLbGKspNoFFKrBRkJInMtXkAkw9Q7YjaKyr6WRq9iAZaTX98LlDaOg6dgZiJHAd
pJzvxXk8aBxJDZNM/+6JO08VebsVa+jF7PUWa+ak1gMSYC/kkGHb2FUSG/NfJuw6+RcxbradPZgj
FwprHk5eW/+XFbnQx+SPCfH7mkh62N5niazLaHSY7jKZW9ecfCQKRwT4hHOKQIBBGFlTfrQ7ncA4
NR3z7in/7t5ZlLYo11kDNbD+jnay8k2IpkHpBJ4C0SVlw4h5eg11TguZ8Rsm3bDQFmHThLucHcIH
7b/wv33v583IT/ctcFgR+svvSvo91V0OCdsMLwVavTElcb7M3a63VVuHQJZERgw9l5Zwy5a/LK4C
OQIvLXP5yxFqZg//E+Azho1bZXWog1I86I8Obhcprqb6nabi8vMBzqbsNzsH1iEp908+86j/zSPV
Nzdz0EjgxIJl0nCyZJsyTsfcPw64ukBJhT6AZQ/TEfVhSsAN2kqZba3v67EJm8KDOI87CO62jfKH
/sToDVi6WyeOi2oa3f2WtdOpRFb/PF44m+dMN+CfqlPm5Rgfz5EJkeVcnsTcMaAVis2rUHm8fRMV
2PDYIzU2IyTGXjLXK4lqPBwFZqxApqGty1zJBMIs4OWrXdzfO+U0peJNR4vQwNRjZTzWY2HYc2g/
pKy3TIoh81EVJUunEG7cxBKQFpqG8mmWjK8fJJ+wozN05Ke/65YD4R09sDn7dluNhvfuMGUH6ryW
3QVwFkfYMaZ5awVD3Ci0oOEabzqhaICEgry9Q8RWHS3KabJ1mXAL71/6ldi++EVjf6Be8DFkJtoQ
xIe7QwrEPWCwmuyCXdw1OZhSeL6Ib/tZomThbhXwfDcG69qRHC4kGgwOciXHA3cL4ktSg5Dhptnm
0x3M1StuXlRVxip2QPkXaewxgOGP/g+Ff3csgztbTaMW/W0sBhKFJryvB4pmhWsJdEH9G1J0yzik
2KhMH/t53eiUPcIgKh6GHXcbQ8/tPhiE2nR2CVnfV9TY511wijYxmHJhKTMtFfzGPlQr1/JeHqmU
Upua6a1P6pz6o95QCgE2Rr4mTW6h3LXn0mavNwF8bXKUcz73bB6UGFHXPXwaPktRQwypJjHc6Gt0
0eXYiB7DaYb0Ah2PyydOqHW0iyolTcsTegmEyd0LuSj866+bO4+sZwOsK5pS8oNS/pItyc5xPKmV
17u1bm4Lz4SZibEyNmcOwj+7NWuLnhKl8+HN5bCtrxG3OAJ7x7v4XIJ32+2FtwPehM92JWjrXb5m
Qxbnfl8KuoUVZZbLOOm2SzsFoz8gtCWZoR+dbF0oFhQMlXYkyL+tH2v2jx7tNUpPqb5VzMITmXuH
Mm6nDTB8FkUOkDGezGne1Akg8TgewgxMfNvp636qcR7Ot3NmzCMLcNL4SyaRgCLel6KTdaoqTPBS
BuztvHBeYFt1A+NxeNT6bVJSs3OoFgVFXVdSptudKVWDp3mPh+9yaSvhhxv/jJ7Pv2StkXJwvmIy
3d/Yx5DLo518EOGQsg3ySFoXQvmpUB63Zp2uLnmEXZIn0kHW7H7jrJG871x1z56NirDct9TJg08b
abxGK2W2YV9VDb0XF/G0Iuwui9JrdaIpUb0Z//nbATWCWfA3PjIj4MHBtjPCms3jXJL2e3k+XOSU
HhD89KqYIxSdoUAxH8NhVF0Jc1JSmnbr/Bh23vp2Et4Q+xkss6mTMGj8N5ppt9z94gCPTLYfwPR3
8IcU/JIyRW/3Go4j9pCWW3S35AME4yPfnBdX4wDrDiMxtX/Ge9Yot+DJffSyV5+6b81B/AWQ2CDL
AMMOdv/WsO5jhBUue/iFRbxGIrTopftuPwqv8kRJLGGZkPl6SFJ/Wi/C2wzh3v4tVj+hU2rLtKsW
+7QjeYJiWz/VIZqaohLBg/7eQfUyDvBHGT8Q9a7ub1iGGZrK4sablviSopezRkcqBfF9/GIs+GCe
4a93TKqt3GoKsfV8hUTxxfYyZ8xN5DV92OKkgp9++J3t5sp7W9LTqejP4hbocsy+jrhBwb80+17q
GOkCpYgXG9k8+9xB6UYdlitMXrQCjPipkvcZ7g+TpkoN4WsE5vlN6a3YADZSuFDGH/ZnDySiYQdw
mAIR92fjmwuDT3fSx5poKC2XCFEv3gy9EprhtJ9WyDuUYOVN5IEmmJH0QYTs6cA3GjfDsFCBr3C2
Me+8+5h4M+7+9p2/zShSatMKRXgGzqxI8lcefQNm4K9S9ai8GokbnSp9dMR+T62FEXTanDTC5Rzs
+Lnhqy83S+WwbzBd7V+rvSDNUBO45fA+O/WBZ+F+nSWgGiHRAcBCuXRldwFM76GJwly6ueoWUSCh
P6iBcoum/dQ7YV8mKTrk4YOOSl6EbCZ9zfUMrDdcfp54fDkfso7mc4Ipwm/Wstd/MccCoUGIlmU0
lA6WBawgPJ4Hp4CsWS0mnYtHP9On9PTmAFRF/tK5JmLNQSegiuY0Dt2nU+CbRhAzvzodyvQI8z6w
8CsLWTOiYdNqIFAuF/QgFjBGiXPF2ABYrSJfZ5pV0kRCSvRoop3wPCfEWrSc5PVBkWR0j4Wl93kH
QsGcMDY6tKdJsn3Fbj3hnFbcHfvzEvv8H4ySRfcL//YLKI9lwI2hp1AQIKWO1y144KnWWlm2SOIW
w4j3wwfjr72pshDlxk83T1NWzJUKPcwEqsVb79WhNE/p98uuD7+N+ycvb6/7h+fE1Xs83VKgqAQG
0V1QFDFXv0HRHLyrQbu/jukgJiGSTEHIHDeNCvaEQKwudWhtALMXvsjWLj0xQlgTxVYZyyBNx+2x
uI2O6PBC2QMRtyierV93mjTMOmrjuaANmdZwevuoZ8t1LGjbpUkCq1V6KXyHWBVO2cSPbMPnfJOQ
MP2qOCdEejfJ/MsZCaineSaO5v0S71v8tBXCPn6wsuSAtAHGnXPQyN81X4Z5VAlfiCBoOGYptbdc
wgvxfBeOaJ7VkcbySmN0NlVp2iTWWEzMXQ1yDkuoKd87mmPr8NnyAOxPg0dEMnzX1hfQIEHrP51p
AIa20JZjXkZhumSlxWmbbdQCmS9oB1fHXF8s8VWoGDZXc/AC6ymSbrXIK0Enx+cLvcke1URNmy2R
CGgl3th5CAO1UZ7h7Y4+YCIHQLMXAO2khb7s52F2EVIrW1M3POaOVF/ursIOv4ggjzMmra9UUlId
tyVmUESA/lthix2IvjIMnlaGEQ/0goIVtFOCBjVLb7LD/mVrCnpDfJiftVvtET+7LPwK92HnT+JN
BLTCdBTZy39PTK7dTEsaQmTfD1EG/RB2AJQPrWMOUBolkEuBE5sx+6OJAeuL5a6UK3SbJqABHWKn
IT0HUv4mk/pT+1EyYznspc2Yj1H9EHNYAmt1eDXwCwwYzOc/u7y8iKWXpevykfx1/QB1geK0E/+S
bCnBVcJQbMcj+w8hta0Xzp9FwsX6bPOjQTVOzAex8nTo+rJcB1cqMiOv8qNZW2HEtGzgihl6Luhf
1wF/02VDCsIBOZ2Yl6Cz0sqi2k/F5dFEC5FB12yOFwSOjWUj8pSHLg20YmhxbsO/HVZ+dgSgblyf
1JfaNrVWhiG70tfSZwgAj6+aosyz5c5mIWt8xYNi/+lgwG8QMwQC+N1vPIRepM7WJSQIhjVc5S4O
VrMcnRHEfrpBjab5uHhrG2rH+buMZFlV9nWoqWSeNODvTG26gZHUNWQSXlV7LM1vtgNtyEB4So60
TRMer5AfsEsOZnUsDtBuL2Ae2kl6QAqnde366uGeTF5Pb3jRrvUjHuOCTN6Wv5LMmgwgzPK7XNHV
EaRwntMwxy2DpsTPSHoDuW9BxR7pZvp9E7SQbUg2JCCaWd/CflulOLT9FsRUZmxfKVl3YhsaGv1C
GeT/S/GxLeNFm/R23Lf9wTydj5vyeKkcyh60uWR5HLU1kb3h08IIDx6bYYCK5zmKufZVUVS+2TAE
07/vpsMpRDZgepKWa0K6B4duzvQI6Ft4eNtKpre+zzOkKaTH2xBuBrHSTNVY9tbbMymurpz8nheY
UPELybYJV23Ok7vK1f2+5liMe0bwHBAjU3qbUDwN2HoO8vMY8sIosyYmWtJjhk8FP0RUpS3w2Lx0
gFmXIbOIDfECN9I62nB6YYCTmYushOh5uACCkYAxRe8TLZ29SuyqYYs8YPG1rMdTIYRox0O5+r3L
iG9Qrl1I/H9cNqKrVTIu8jB1pCVjlwWPSlwvV2P3O4Q1vADN0nhEFzGXAklBKjYbdWiEp46NKfDZ
MUFpR7JRK5nqtLUjZyQsjIjrs9lmNypUo27tBG6a0H8j6jVUroLTtfLelQbwZ1QLWQwuzFmghN2h
1QsgX1G1nwGHYQn0CqNko1pM7H4XkTI8Jv3wj+hrlgWstRHm1+AhUMnR3RcwwU9qnYaynAY4BCF5
KzWNSxcv/tELsNf2iyHlcsXoajB48d7R+OdmpZlazribFg/24giBe2OWvB0GJ0dKaliZYvHdV4OA
S9Rv+DqUU4AakPbniPPdP+aSO6/SAF1jr7B++s/kjMv1czdMRDlR9egqKkWIbqJ3kbRel0HyEZ7q
I1deIEsDMLUJxJFoeWjIKT+0yjQWfzKMhuGDiRbo4wM2B8BLxW9Oa3ZgW6ol6+T+WHpdbUNnjYab
/ZDGyFCC6pH/Xe5ZCXwDBPSIToGW0l0TKHhUabuxfjPWtilPTkMhUXuteuFYCZD9q54NyuTs5z++
RMC4ZdE5/AKEFYExbXqYKQpFfCfgfMDzeaA9x/SttBgXtSl9iFGrRDjlvbAo0tD1H19lHdzg5kbm
iNnF3G5QAq6PoYbZZOPSgWpL5UQuQA2FxsoNizyZNIs5ex0qA7rSgHZNSTQ09ySi1ksqKHNMgPqu
rC+jlCP5lLFTC2j3uGTHvt7Rx8hqJBcuIHO8kM0lW5/j/gPZ4KE6LpjrAC9Fzi1RJgStXHo2NXZ5
b4GxTYStwtXzA1Ol9cxyfohGls36H0xkGiZhvXkzSKByuHwZdfcmV3W7B79ABx4a8l2llvVqxkFQ
dtGCros43TIUyPeiZVpQh7Zbdn7NsKnX741PZ6Flsc42jOqK9EIVhBG6aM4P4TbuSg9loEossk+k
AVdriAypnqzePdL4aoq/QhZ+jAEK0cnnCjLTHenTYlc9B98al/wQ+p6inG+CwrKTxhXzU2z+Suze
FJ2PNZubF4YFgRuV6exTbGSWHBxhRMX0RYnCchI49bokqjkZpNrWYSzZQT8PgemGwsNHGaXdJ7kB
C1exnvHBHgX0kgg6H8pccsPyld6bFa3Yn1JyqQq93ZYmqFus8v4p9eB3Srk3pWwCUn80E6E2k5lU
UyXD+SknU5LGNsKJ/+UAtSl8L84VjlrHxS+SJjAB4kvnGjAsY8yMtP646Wd4BJ1zKS2vuOD5wdc0
dbE41IkGz5UJpWVWJ6BRYplnoE/MV4ZzV+9GqbOUi7Rpt9cXQ4FEkPUcKwG8s0U+XA7ia/F9YAA2
PO6MsGDb02s6Xem1giSwtYHBgJVCS28WaXKluC/PcM04TDqJcfn8hbKjeLhcJUh799iQVlfYY3Sw
l/D96kdqL3fyOR9k7UC4j/7pjCm9AfhD+G1XEjQDu/0C1dC+gpzdYTHz1tnd4Dm595FdrP/rqR+c
3L0KC9kfYgF6nZuGQQ+gGKCjegK0oWGsc7R76LyyLMRj/+8W79k9pVbRl7Mg1HylC7uA2hNRfqQt
C/iMRignhGTRTOBg0AXBFFJxOwgRM+4cZy43fauZpGMMbucNLumLouL3WK/d0Aef4sLYiiH3FvXf
INlWJGTUXgX6OasTy4vHiXvxMQvUuBmPo8gsXCqviCzkVh0gPnzq
`protect end_protected
