`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U/TEXQjZUaRM/9cgwpEP/LBYfJ0jLWbWRkeNi7iB9W5NL2NH9QolQkR1qJ5lgrxH3yll4V1asg+6
sGUmIucWuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WHZACpkiDnlCGXQ9djDZpYQIIYvsuuU7UxGXkyZaXRN+rkiqPmodh7r0MHZcR2eglLvvpI0+obtA
UK6khoy2sIeo1BIy1jinW1H7bE6QLhgkxKojlZZURK+McLWjsACWq7ZGuV3o2KC5yNiB6q+1MvdU
dC7XhouA3JpZ45svpkg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DP8K4+95dnff/lZasMTEi1gqUuP6CfXWoLK3C0sXkPtHmvo6JCoPWeM29vbOZ7/oDa9WYFdwfFdB
cbF9GQKv2EN8q7LTB4WBdZU0ehkGcGnHhhiC+VtlMQpgHrUWZ8SJVsnaD7Jh7S5h078SZyz4TuOW
Ht7KQwRloOCVjcO6oPGONig0zSduxs9Pvk9v/fcInd9UgldZSSVqtngTl5nQ/fCtjHv+8xjHuXZN
wOy5RrZXNDS0v0tsH/ZRaOS0Qxcc6P0folnJTdx8XqMDptdRbTu0peQLxE+mdpPA8c0oxqNO99wD
n/e9fg0m1EQ2wFTxTOwsL6AS5rF+YEQK/0tofA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GuK4tPHwUfUSGV9ixlOfwFWcu7ftxSP/AKF9X/+3AQZ/jSBj8yr829fZz4TxW0ZwxxVMdjZdGp5C
krDjuBN0rDNF0NKt5HOno5nEEmAVejTa5KjGzQoWAi7kzCQMApJvZLd9vi4PkFcsfjQt2LC/R+jT
yP6wAqsO3EklkugH+Io=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GSWDLNoq+Dkh5zV5QPNn+l5h8EmLq4sVXdBWMKs2IfgibuWoAS3mSz42hgc6xfN5wPiZMs/9UPpQ
sHYQ4gVExqACJCXlxaHx5KZNmIYV7UACMlu637a8dMnF6DgTxEYYsIpXdzNRhSGNWBS3kP8Px4MB
XIbrHud0LYjetuQ5ziUaFwhw7n3FCl1Mvr5emmYF5km24A74Rq5lYdeIsSBtu9kGl7IDI/d5Ve6C
CMuiyO8dYzi+4btJbQVpMCv6bRm6QvuBNUUhYej/V2kdqcU9ke6Gwp5Tiw+pY6vdpoe/o9e9c9R8
p4bvBYoW7F0FoFNmI7yJsPcA1LtrVmHXzlsXkw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
3kPL7ncjniNY6UfiWYt7d1+Gx3b2BGX7njJviAL8exB6Qwd6WIrPUu3w+Whci0xyIvebtE2vTu9c
N6X3xtyKY0d6QHf5PKR2FwZu0clbHqiA/vbMiN4Mq9lWQMTG8N/jye1TYzUQwmzAsoK1Rwbp4LVf
SjTtcjDykRPdendwJET8uLa0ebAq6nJ0JpntJ7Amr3DFIIQqezVzSpm6KsIe4WAuPoEKBCZzGVsT
9X1gufY84SD+XPGmEnJGAPZhIAJgyBq7BJRGXyRbpMKT24dksQCqCuyn/kkC7l6dxRK0Br81kpP8
QzYFpn3lAclgFqHJm1xtjg9ifFG+yRz0XegkRPbsPoZsCCQR2gN7bpbwGdWCp/J/GiONnT0DVYk+
YnX/zoSncrwxaNiQmfDVZnfT5zQaPHPrg5w/NMsW1t3w+YiVNs073XlaFmd4nprZlXQCTEbZDtXi
8Zg6Em5c//guAuAiSl+bt+569h1k1KwBE5SHDpab5nt6WOp4GhPdEOrNkY3NvH7/BmbY72qDb9WL
FCxfmnMKabzJ9YH6ixXw2QQPjM9NWcdBhl5TS456BbAoFDBOXVFJNERVBl7LDv5BMqY4baYirzEq
N+NebQTZnmoFT28KDhlmV2iezXYXtxChzWtyS5S3HVR2BGi1aL4OWjOh5VDJekXyGZ6J8TfF5B3h
FTQmzfbSTCpQUqGiitsGEySh2aCGNkc3U9RzLY8GYLrR+lY42Pik7C2xaNSlrM5R8s/p5LyjQ9wL
W5JGZWaw68X2+HmqQ1Mb5+7YYFbxP/27sr5KPuiQ5A8Kl9JlesTd0tRLeiNiRWLhY4Zvtq5Kqg2F
ihSwOowHVnVzgOuizSSrTjsKLagt5GUyGctfTxNWcHM92OYNCmO6coTwJdxn432yiHkGukw9NR+y
dRIGArp+I2Z/xh1AewU2Yep2tTlOLnoyUbw7tW21fIkCa0pTGDc5WnEwn85yoCplgGlP/MrhAfE3
v5w7PKwYM01cGxs3OF1Rc9ZR/wiUU1pwq/BhKXOZzdm8V0uAN3EAJofxbVa2MeEDuHdZ3qypiNBj
WwpYW+F/zLY6SU00NJhzOh55OJM3/5/5ITyZSR+h9w0+rBkghN09yS3WuLrLkkNDx0yDgLJv7vMY
Oncnb5FmRPI9MbOp3iMGkP4YcbKZetRaDVtIq9VTlxOSqcZCwRM1e/VWEAJ8ERBHMVsWPEqa0yMx
B6TU4xiq7xTZiKXxe35VmX/wysrlofHQh2u9ilvudUfnJnuasAZzOtR2UkNq358DjPYvHKg0DMCz
QAPGOr3wkDLSVJxr31WsFHKfaOHKU/d4vDC3Fpcpd90K0lBA6dKqgX04CA3ZI1SWOlNkJXYKc/p8
Mi7kBzTqVl2PfYw6ohy3O9sQ2or0H6iiYoVHRo0qdRZliff6ipE/ZovQR2AqOx2zb8V70RnbF5tu
N2dozWot4bmGsynN54iVcLSgXtqWpYTrZPfZjmHIEh6bM/MjBW6lMNciLlzxT21UlhScgyP3fUFl
3Ymb5I/lNDfZxVpeNLpK+PbpI/JjJQTEqQSqCiqwuEWW57/NLKVvdMQGKeYixSxwD/1ZzIAayb8d
PO4UTKOYPRF7pM3NTmd3yngTZIG1W4UZ++iu/xcUknMV2izmXPP8wZwihJ9vd8LzeC1PxYSCbCEG
JTRNGbe4874YNZBh8Q4W4bo9+FmmQB0wQMT3B8BSN8xbqHBVVGvdxNhzfKtAh/br509qhB5xyEsx
gNz21Xn9xzpb2LtutbZ8sGk2hX/Ef9drx8KCJCE4mz6MkjxcotFaIXcpZjHeuLP4Y7cBXVgCr5Yw
aUF4vpFlA5zwmL3ybqOA6cDbcF8QGQTsH9dS0lz5dkscktjps4ak6tL1qlS4Eyu78OYx605aMrT6
ZwQ57f8USn66/p6zA8S5gXNa8ZOfDSsW7vF2YPNfnhEQxMIJfzOYzDwbJ5omcxFk7wHpAm1/b0hm
Cd7A3T7In/hPzlQvQMR5sRkDxCx36U6RxwSLawyEGS8Lj6SuEc5yc0KWz2cxUN139M6BX1cLrbMl
yDKDNDCKufFKthsOiziVjs3ir6NtYKPNMEcsUmSP6d7gxs0KVAHu7Kqxj1FR7Jbd/CqVOaqGH9tC
pX91p13UmD8LPAqGfjtmXnll1VM+VVFUSmqLFujlGBRKWz3rID7CatytQZRb95l5WpAgSYYH8Xml
dawByXtq7mcLRjMDv/g1ZtT6frM21ozY9Yw3545mNvF3BvhHXMjlLfx76R+aErnWoQss8bF9+NH4
4jurf35dV+OLTPV8SpzyI0EkZdeBXhRMKDON0HEZrjPq+FEotl9msiEVIKyKNKmU0D6nooGCzt3F
ucKXd8XSiZ/yNLdMbUXWj72QycShcV60zdgZ4Mq4h6ujPekQme/vxtz5mRWZ1lw1ET7yknA3lccP
uliUWnVM5w3hwqO0DHgzxOjYb2jujD5xorVgTcNk7Id77XEziJBf1XaPQXP+LnBT9fvEuaSERwkE
TwqQ4NE2BwHyF49mVfPjnUiRQIJYTd38IiWYqDTGzoKCgPCAYbVr2TrGO3X6+5L+MXqM1Xsshjkj
LcVaAxSe4tdg7zqW7fiY0QzgbVMEWUWzsnQKG6IgQMPKEbKPbF6gQzygbCtZNPixAx21aR4lJpib
jRlzvBbckYv7ZxuKrTY6Fox/Bbj9x+wdoY5nE+ykEnzgILLxXnS7c6Han0P4/YbBj9NQkd0EVy/y
O+XuCqC5Ve2tqY0wLj85ddhPiEtpHedg8vaUE01d6T5pDgqGkU7DsGsHKmAFU7kSEOtKb3sBDSro
uKyerGBCe1XWersbkExkbHhIt79/iJL6nP76InlhHdMPIAuy6sSeFWw5v2xgVtq4QHdGiNtVdEZb
533rYAph80QTXZeNHQ8/GPWkd9Pvh0KdqsOyvBKptsFhA9tkrf/Hom+IPYobgCT7Ih9lOY+fuugK
nNWQhrKT1XsN4dOmk7vyBhGjEwBLdWDAPArNmWjNynL+O/TkssPr+RUEL43ihjCp2YSCIKu6PwSk
D35kkc5AwL4aZ9lPVfO4FoBJJrq/XPrb9x6iLT/cPCKpUoR4T/QLePUwkNCqs2xHmPKAENJdnXwe
ZmvYQm7cuAEFvcU5WLL7W/uFJQvQhcHqtMWmGyfVXDsC8xhaG9nEjXI3lBaLftptnr1t/igs8Iee
UIbqjEJYSCaXxBwyna2vMdy6Nhgj1zGynw+GIO6DztXIRQgy+44HT23pumsQmO0O+yJntmlwWnRa
U2bSYXFrSTHMs9cbfXvgLLckYgoTHBtKs+YyBKryCsmtgl1qIL1EuW8f4rPTLZ86wLCVwLTC06EV
Jxfk/87UaUr/J64W8T/MW29GIiz7MPvBwQUJrlsgw48AbIWPC2oVNNEUUdH2DG4P01RvHPT1vQ/M
xtETOxVac8bQqRJJgeUHAYUQwOw+mKgnJ8SmCZ2uNXfkJEsa1VoCm5HNJ6VrxzDsM9kt6AjWORhL
VTjXfI62Z5KaFVbCT6nqO1gnse0M/VuCJJip5egnPl3HMoz/uEA56I1liiBqXyZImVpyHRL2rleY
uGQVwqJM2L+OsmTjGWJ4rbxPyIFcWRFEN6N/NM9FysFLnNAFJ9T6xPV5YaKYzZDNNSRSl2Lw8E7d
C2X6FOLmUUdDBA1ZBC4lfLuslIY1S9KZdiG0gYgnd8CSOxTQAU3oOrgJHTX+ajMSN3wBKtVEGoL5
ciLZKSit8WOFK8eqfJ1YrWILcCxRKMGehFjvYXfuYe1uzqiUn7caE2f5BdKf3yTbO760ipnpcxki
NXIQZL71dNUZ+wyJwnJwkt8vDE0C0Ze/NnHcHuVqNVfy5YTbzWChFhsAHreD7OYssMeWOWGKLbdL
lcSXVyiIRjE/ERqNItW+/ODD/7hfKGtxBQszoEX4WojUvnTZX7Rfsl1bbuO99EQOkBKHceVA2ctO
L0++PWec9QdB3ZAS6R2W2m1xiPMmP7SwmPTV2YMoEXvfoz0nLtN+OZx4ad8y/NgTU1MO9tdSa0uV
oV/p9sZkJXwmjmbSmwOMzi4hg4K6iTN8A2iaTNstXLjiVOB0Kc8JGxy/bRwW3+3Fg1kTfXOYfNL7
9CLf1S3Wy/PJiHz0jVNF3hIl6vVMTjWB2iCbUxI0P1Nd3oTgo1MmPlhNpG/F29+dQy8Jxe42xjgq
IJ/pjPJycc7+uiC/gJQtqVIrfnFCzP83qW2y79qmbAMILPq3ebKya2zqrMMoTl0w8wU0neVoh/L6
dx5rFgT0lfj4p1wKo57rq7YB9F+HfuQUV0aFRlYTGFCmb6SevcDAvSedIyja5vXWvHqX9avUNWVI
lwhsqlnSPsC6qVeuQDoGR525VniqZfXiVeBcZyPgb1vjlI68BC+WrJAHB9fpGV35ZQ4OWWmhyDx5
MybAJPPnDKWYRaGR9z8hZ7b+0RSsdGiQ1fbOwWsngv3xTok8JuEYqxQhrnkyWRtX2yR/9+6nvd4A
wXjLeQY6KBUwE+/Z407/++ohmjyppu406lydP1GQW0okuMFfxmNsYS8VJ5GDdo9L+DUx0Vt95nA+
4aMKgqHWey8v9sAcB3hTEWdQB5zXaEys4Ewrkj3Y+/XPTl/8YR93wLn/pMLKyWgrTBExRu6CMEbL
Ka0pkOET2P/IadcXXH6WIqhc003wlVFZVNa1eyKUBwZ+zi/+RT81UCsWA5GX47zXKtaKIuSVL8nm
iCM+knktKrovM0GhvNBmupVB/wa4jzdPjqc13BXTSsYcu/sfhLrtKm7iIk6YrBcvi28RRkifbUiY
DvmUPJWo09Y2XmCfUmxwSKwEI/qSCOhlhe1m9chdbmJMKZLWAbejNeevHuiSr+jxqr+b6tDEXMbJ
vv9iTSQvGsJAmvO2HJGhkD04i8+t8diF17gkpK1wyFi0sT59b242JyWCcOumf80ZBUOYkMpQIDlg
meg6MXL273N5bg/0OJF5Omd8mBJByqNk8R2PFfBCvG1k9BDO+8czTdNN7ZBWgJ08zqsRh/d5weg+
10GgvqBmYRuydVZ521l2LI4kMRanPrPXXcmxWKC38dNNIHu9RCj7y2bLEl58WU5XotvfjPSUxNc7
YcAMfLAkbun+EE7u/grAOP9LmFo4MuZDQB1ATLiMD73UmyMG37cySS8NUzpLWqCUSMiaeyEPh+ip
cZYraPQNK01kd8gv7lIIx/+eWSaZTn2M7bEf97DW0OmD2AvF6PcvYM6XSbUWX6ZxLExKTr1av4HF
XMGiySq79GS2wjlgQngzZTUScBXvNUwpxLQ94puO8zev+dne3BevpyM5dggaGxSMF4DtF7veFQQA
Bw6og66Z7pGiIQqA/CFT9b8TEZjXcRvPv/ohstsUqXMsbYYG4QAvAxqAil5Dfq5Fyu3PVIG+OFdz
4A6+H7fbjt5+2nUhbcaNXbMTaPldvk1duTGtqJDxod88Rrc94MhEG4WB9fUr1RsPqkVcH1Giim+2
FSj27C7ZuLH4oAy0pIymwvi1cuuUmX1csvNcRSGwD8Ve3YPso9ScH4qlND6bdf2KmPcSy/fNgCao
95UU5WsPAKWK7wMlVoGMB8YjpUqMZqkm6F+tKN4DGhynHigCABm7RhT4jCKvM4jv94uhGohzlqlO
5bZ6XZ9Tc2vs51Wrz0lwLQybAUvbnXb3KFq2QERzZAUnoMMKbcGF6kIrY3ZlhbxSGPojoPB/qbFK
Koaja78JdE2RnjklrFWfaOJJqERaWqNlCr8f4KrDZsCzAtQG6BsLAKikVSJ5EVhdhqUFcBaA91LN
jJX8rB0+3/WBUsjvpVJtiICqR6wfYMO2bo5i4Nr5XmTwxayfawqzifcqEDZbQGi2qU1JzRgR/7JG
2wrUCWvPo8bSZn0TwU9YUHJiyKNt3Dbc2zRbsNMZzavYeu644BCvvhX8+0lkZ6xKQRgdQRDdLKPu
UDPYSAypUB6/t98YpoC0jsVGxPLjwB68OrTDEBj+qlr5cm2upwtWPZ/0rzEIfOYlrDKcuho1biiA
Kyr0K33q6pyrUc0B2pubYnfc9o1wbeY4bhtilyku6OncAbSjGVKsikhuCnuqbFbxMP2JUXCbMdMV
r8hLjTbyALG5gMiZDPkvr1Jjp19ibEOLS9tuo+8FcZmKUxgmzUlhQ5JUwCSrWI/p9OtNxzdRWULu
kR9fBGcHwA==
`protect end_protected
