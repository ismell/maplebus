`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y/l51FFDy4EG5im87XNcmL8LAM+J6ck3LmPLutc61WOG0Wgp1Ryu7lTyRxlkRoBBbksz7nXNGPPP
HBwhB1SE0Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HEy63cTkByJaXFv0zDeVS2Z9R70KvKBdmycA2zZ1AaaOxZ6nGO40qyjsPOJAStaMRVY6G96B8/2I
J/EYi0o1w9JlwWcYpSWOjpbFO/CFlP6eBytwcDYmNqcN6G6ZWr0nMtscaIun7OdbgUeaiL8BHbSk
/AeracxMDAeZFhGAEcg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DoGiEX4NXkofGvMke3Q6Jk6Rvm9x07kvCJ/RC+a/IFqbl3PuvRjbuDQjPNAcP3CPWi2Nzu063wyv
k/vcgMh3Y7ByyqtW31HwCtJZo+yWLI92ztIYvIUE5aeozSk4F92Q/XJ/VU7p5pGFdUZOql7Lc7Lm
WaqYGTdaKcKDX9Ra0mPVjrBNrs8tnhO9DGjIIP4oOwbGruZKZY9s+Bk/8dg/6yKJ1vr8I/mGzfeg
T7j1uP4v+e2/DoKP2+WS4pIKMo6KQNiN8K785RnpCE/dAPV+66MlcJYsAvKkrntFxuIV0LC8UPtU
V96zQqcwmsCloud2CwSXVrdYgxNo7pd771aMgg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pqlvwfBRP807PGy4nOaVSMJT1vbp8CK2NdIJdGDxXDc5FQOHAGJRZxbcg29Dc8SeuEkcnoDgPT/E
pXh3CuVR4EIIsM3Ks5lW3tVzZu8dRB3eTwf2914ULHWZTE2zEvsuWEut+DTL7TtsT7bvB9G2kU3j
Nym13rNlu+leF8R95JQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PFWy+niDgehlrmQa6uqO1pfacyPTbI2/5mwN/NzeU5QZ9F/jMub3NL55cvAGcoZRXB8YTaj4ugSJ
BcCVa67HZHJ1CeSsJzcJT0oZOjYsXsiXNmG0FxylIzbekZdKLTwkN5HVnfs4NAULe9eeAoVpU3yi
jkJuGqSI1Z2eG+mUSvcPODh+gxXll4fRTQbA55REH2MlAJ86YukG9ph+a6qwLImsQZzFQQcvO7df
ErbGiHbkoFaV2MMHLrivQvnj6c3RmFug2dGd8/Mo6669AI6Vl/lAC6A4CiP0pPmrPIeGAu8kfXXn
o3Qta0iAcsmEw/q9hai7GGTP8BVzHiooKScs3A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13264)
`protect data_block
rYfpseLxZ2vNkNiBIv1y1fIqeVveLO3HRvQH8qcKoCLVBu7Y86oVpBm39nMiEj/CQosCdjDJXiRj
YhHThJYZ5I9fzE+AaIqMfBwsXgQ6KNbXglXpjRU+Je7jOh3Fx7fM5+bqHnxrGlMvJDagtNwPlVvj
W7NJjRyIzGHFW0ZbH6MzaVGMEdIXl2tHIdOOOzEEKgZn55SDtAdTW9dFgyBnhe2i/fAWxY+w2Xrc
vnyhSjCgkLgyPvP9VDBfGZ0nvLCHOG7X8mFjBp56ycqeAI1KwZKJJmUaiBNwfi0yNlTJfHBuqbkw
1kDjG9AqPf+bMJNJjdR//ON/WyQT61N5ItufPF0xnBQ5psPvv/mLg5KV9GKdAcxJgsT93hqJcB5v
26eHh53+yPDsub+EB1KpoPDnimWGeR28LpM4I5LPnLGvWF/9E+7xcliuyr2XVf0mVJXjSb/TnffJ
KVdAD1LJ4Ec6oOdaa0V2T37jvsbBlFvoy/soEujVbm8sITAbZy3djL23XZpayWscpWlyH6ZYSVi3
OSyeaUp1rhhEcmnpQcY+RpiP4eQ9dKTQpNIdUQKf0YN13tAgMPpybHfxDsCbEBQFgyNmK5zl8JWp
q6IkBQtV5vVu1ec2fm1e8B3cGJ4zqraOKG1ZLmXejUewCYB3ZXIFVgD425AeRRb0uMFNYK8WSUKU
izYWcSxY0KzZjItw4NDfFa7Uqw+hxbDT6ZMbaYgypIHSn5TTiN5a1jUTQsY4/3ZynpcYpKpuIjBS
z4FjN+1zQgkPGLV23tZOh7t7tN1ZTuDJo9925HtCwzLXk+99MxcMu1NLj+ZsabVkU1yNDijr/BaS
uwdVkNkjRYFi3o88+wuFUeL82c41orLd3QgY+9ie7YQoSlD0PXN0y5UrB5Dzs8T6mfaGByAIfCb5
x2JvxXp12b/1F/w7J39Dk6ygXb9WPLcg3FX2PDP9DlslVnEMYFX3tRh2g/dROBNPv+kl+PhGFf28
NPulqIIBBxyJgUfpfM5gvpYloGaURFcQIFcJhmz/Fd4YnfcdgC4F6ftlHj7W5m6yZdQ57nQ7PZbD
YxZcySxdzVvy1RpSoxsL7SqAt1Pq+mL3XgvQG5zrOVk/0Z0vQQ6BCUUDhglzJO+6adh7Z/H9aMT1
WaVcW1okXsFLfC+ch4kwjAAUJShoCPOK89Bb1dcZWi/r+7SdlXKaXux6zffhv2NQJ2z3B/OfyLON
tuHz/6x9S7V/EQc0WRTnuIaFuB81u+aCG+pvExvkv9wdpJpfjCiJGsRABd5dJkMtDhsaviX7EDhj
KZMtr3dYoN3FlBoS0PwJ4JCsf0MioT1BgH5+879S5QC7bmBR0V+n6E6aehqwClRxGaSaT2gUVyyF
xVWkwdI+wi+yWnFFZwUkHgylA0gyJpoVfnKTtghMq0+cY76wVXl7Aqvcg/K2xKZSd+sbRR9ZFBh0
18WZUwNS4uajxIwjbqLg31+einCVjr9xMVXnXt4p/nuveDZS5QkAh8z43MSl1HHrbpGA9y5cn636
LVuHvUqVaIBHbRRFX+iWrTvGz3N1KWxL2rG2bY8aojMWaWnUKo9fumXocTKKgg5YajnFZIhfiRIb
GBvkuCj45zCGldh4CzQQgPYE3Uqz6kz6jOVUX7ezAzeZu7cN1pUPkGXXoXkAgg/COu3kHoGe7YZd
a16j136+R0vgusZPpLj8V/KKeQEECjgP8gIda7UXQmFrHu4NI3Iqq2XhBzhPRz4z3OuWeExeVUGo
rj/yxBxUGVNFLJBAAMSFDI+7vdLLNzSs0Vmv33QgwZ/rQdMW7kizGNJtRTrZZDxPU1dNbn3zdmgH
X6NwA4IXD6LBZPSPfVeozFzfjOXdDHAyjZMwBkXkzZInk0woeoacfhgTg7/jzIVQstJS7RMmWXaH
TojfWREqhacEHRJjQ/50m01avFypYSAqfFv7c3tg3X3O8daS+FHc3FdmM6TSy3KivSZx2+Xd7Uar
2j8MeckPAd0IuwgmnugOlTtke8Wtw3V6MUi+rkXncBQWpt6ZRPRBg2rkpL6qbaPiFgNYdS/FCIUj
CZLq2KC7iOMd7njPuyXX8Ep4jy7TIEu4lPex036NIwXruKY4P3jIoBXwX7HKpG9tXPNEd1Fabqc8
lo/6aJ1u3Hn/2iksm1T3s+eeMvc1LX0KpuGbXAlGTuygWhvZHD3rOtlSexLCiS+u8JDsPuc6+NEI
keUe//+JWfMVZ7vq7mNc4O1T4AYGI4wooX2Hk64SiibE1J2rtvfpqtGtEwXAcq1TrePbZDCkM5es
Uq9Ks9gHpWGFXvA5POAo/m6xdn+xzrCvmKfACiUio61PEkQ390wbE+DJFX9P+9eGo8T75+1n2DwZ
d1GCx/qB+N+C6fZMqfT4ggdnBQiwHwwtgT5tQphLF+L3AAwsdxY4DfyJmM+kWDpNh8364w+2NPKz
iTdfOuySHWL7umHccnBY5DbGcawR2+WL5GHpHL/R4PraXO5U1zCAkCjIhjqCfvj+i/C2xakSPGBz
mzWoJpCAswNgaMtw2ws1xOTrhJ7RBseHSPHH82r73WIiR+vEFl/JmyBhbo4NcCvzMLok8VoLkyp2
s500ILt6gFISIF3h8gjneBOKMACXYQcsmXcObkiQkZZqNYs9O9VBJ/iH+IfxiTUSPsu5z4ro2E3Y
FkgXbMG3xfWk6xve0ejTpD7I0g05RLyN9QwBLN/NTd3Y3CCkMlOfb6FjBip2gpl7AGnjl55yP3It
WSgsXtUa2Mq3y7XV1wxp+mUHH4/ngjbSAzBuPOrPkFopeRXnb3QVPeKibFkW/XqhJwXXo5c+SZEA
Ont5BJcjOMhLMraQgdy2548hxgL01nIYjrEuWX7WS7beCtABW2oJCCNlW0BwacHbAnQONyJi3y1F
WoDDYKCPePIKSztzPJG82+g+pY2Ljr5XzLnEuwite4k9Z0rsSinFR1QE+WIMbt4E9kMARm/pRJRh
0GF8UzkaIT6WqQlXwEx+2B4OlXBbdAG/JEWtANfHMOztEwJ1Wecl0OsA1U2iijHQyoUzoQgAshsT
DrWzAuCNqrKRcCrNIYPThH9pbF2it9fJvQ/Oa6nXcG1TecuF2L1fMsxAcSKR5R5CXQavaoRdmSl1
HWfv3+TBV8GpFK6WQkNzFG0+OGKj3AGw2UmtkvjeJtiixDdOaOKM2whC2B3q0ZK9Wx8gGqhO6Xdv
edvvGQsm5RIcHTcU664tLulC8ka30mKe/0AQyoE9co4lhjNxEZGklouwb7X+RamqEgMoNNZeaTZD
hiD6UELV+9IRHkZ+d3G7yCFRNmDJyi3T2MYm/XZbPf3WcJbOgu1Olen4UF0TXY4wSeGnQ3knGGYe
csyGMnFo9hnnYe/2IXE+yppOFc19ZA58UyBe/sF3K6YK1UxTqQhPumKoepORK66kufzL4znbpW6/
I4US/twlsFZEXV9UQnAUOvP7BaDm5oNbBNJgCYJM4sZ9aXLsGUIKLUj4S5iY03BbW8npuorC2nfC
lKbPMvIw8PucekI6B2WrmY1KOU6RBcR10mGx24m2DJESVePgJhwI/nT8oLXWlbfljy51IXB2n/w/
RzDgw7BpJdvPdw5zWLBdjvuXRbsDloFDMKM0cAgYSMmou4QRP47RKGTNkTTiRpK3aAIhXl1ur25e
pIehELdIvlBGf3QruXeWcH7bdvmg72l3Y3KCuRrR4QxuC7FFWAsYYFWCR9X2Mj5pgRGxUde28PHb
hkbwb1nL0vyH/ainUQGRNLPcGw4jif8D2ytutVzjcqnHetZcjSfgN0HtIS9M/k77IX79mCNkdzax
fwTBGyZziHN2XwhEusV7gfWMNZakFfZy4uGLCJ95uJS1pIOzJMZtRJiiSEDvHHLR2KzNI5i50sTB
uk3wXU9xx8Vc8s0wi5OZzZ3LNcD67hA3Hv4Pn9Yq+cTGsjItWcBxCCmbVW2SDsz82FJZEYNmVkfR
Rnw/KlO/eoAONteq0Ro+hB9HbFax+cOKmssGc+bqfs3vAsRclvwQNfEEzvidV95WaozZ11IZH/ae
bJH72KclzzgGnJWnnSB+VdGoNEyV1rl0uJHf8YnAAH6DFITVyFO3AXwN3AcNCni12B+Y2n4x3cwV
/ScHqx4owOCBe0JIet8Xy9fymDQYcVpQCtjeU/0tKHS6u7zl9qLTW3qA3scjdsgn/hiI6Qem33zE
K8UKnMQ3mHcfXJV1n+x87bSrRwIRlouPPqdp+rPgMTxe7JuUH+JXdyApferLeyv88jvVmurQCNKI
Frty2dIegvNhjVKYT2h4xFRJSDFJ56GZLJpwEG1L/YX3+DeDJlFIn2WeJ80KF0yqVsxik4kQw7wP
ZR8RswZhLLmj0NYKnGtSHSnSYedqvHKhWmayPjal5S0ZU3ONx7h9LmjAU06vl9AQ1+9OiwfupzM8
Igl2mO0NIBlhwJ0eKi9Ztx0tpoCP5ZfZn9iffDmmT8YMVZKmKD1LcR4toPPxHiixOR7VQFf/krFK
kweoloYxSoKKvVKTDoVXKsuM0C89ys7QLIuFxhQBKYNQ6i4htHmiIUtTUSqD0FYdLmB2QxZSdhJg
DM4ssRQ/H0pxf2wtJTfOojDMuqjigd0zmdj4MxFzwPmnkYTtIwcBYpJxZwr1Ljkf56dj+k7YmhPw
PwxRcAwl6mfU9zWUuaZeKAI2aBhNA6hf5j6ygNsFSP3Wc+rZa8dCYh8bjiIb/TxC8nYIjrQghBkJ
0gdsJ+kGSOT5Sw0AZm/UHvnQYjJxAnP6f9cnPay+6glJuHGoauf8eQVR243apEpjaKNoK4d0vKC8
NzFWiAw0ilduS5ihc8qSYn0RMzIgR2NtZqT3M5BfsoDarrI30u1xo8rxp6CJBHKBBioja60i7IoQ
gqFEgxvD9C4XQXlVl7Qtvs30bRTRmw0FxUGNlmjMfSxwSBy0rbswfWZsopyuHEchYm8FMY8obofF
j2OwM/oBrSjByGUZwJDoetj8j5bJhRtyTLIiyxJ8a76qyVtZMnWIL6Q6LZjXAGy0QPQV8CG5nUuB
XX2f4eWUO0ZnZgWKk53o4Sjwmq25cmX3wBcBkK6roqpSySdcmDFCz58ts5raiboFUIGTz7uczyo6
ZsxKjvI+j+/7dHHbHGIs064jZrHYcFaEse+JsF2q2a4T0bi+xZWtOgQByOfYF1env1bR4G9Rz9u9
euL1IvusGuXeDHl3H008NQ2g89ahTC1akAgZGYc8yfGkgtQ1W2MbDEpSqDxXiMOKSanoZ4dFM6wY
E0t7eVCG8DtZcd2Yn7HXYp/ZjapGJASiFDz0yYgqM6VGQRWtx0Drzo2K1Ep/RQ6ftV9+oJm8VBct
wouGdA78cLEe5dXnLzmFSj9INEfPGif6khT2yiaz6m26sc2l4qV7VPQ8dY7MMROwDHbazaGEue/G
4kZ6/sMGm3MzQQCebRLVBxm95zPptO5rpBbOLbjTvj1eenMvUNOKlmNFFuVdtMW9GlEx5p5gBk+7
qFhXb+5L7TiQjbXszNyiOK9oiembaiRxPkM/btJiS/sWa89mGQthVYgKigwetjRMaH+Rfh4RHBhD
cIEHhq/1LlOqZ0hGPmbdFC7XrPw3tZJ/hgi3O9u535/ee4YbiSDzVvrEE9SUGyBk6U0GXkISz6m0
d+yhlFPkFVkSg0Gi2oznmhI6vKYlCl75M/OP6dfKpYxdWx/znxPxOs4f+36f9asHF+QqnQBhLhVs
4TcDssQgrRG/IekuOMsidP5F9yBu5nPAvnMYoaccVakDBxV9hyym+h6800qLMWyn2k8dyZCxRoI4
PGZ0dwMVE1SPRZpc97OqJ9M9TrDU390ATMZKUS4SI6ruz4TzjQZzCgnKidLmtG66vrQBwdJGFMxM
lO8QenG3ptbf8Y55v6n8qaJYLGPwf0tD+f4QUlzs6cb8yeMVpRKACuip3frXPFW71Uw0UgBBTo1S
kbxIg21xB1h0dAGQwVWQbe79ef9JShP8ftpXjlAlRKBPBPJUTFA/GRNc288VEdXZ5FVFSXklXMyr
fd+N6cFe4iDmAxZXB+idTclO+bXD0Vc5LEzS/5Q12qSd7jENcbGhr7Tq9BMQTkcNuoQREv7Wxv5q
KDzFmdxzIMOfmR3WsjqqBWGXiiE5dc/i0YQCI3ro6T3QNht1HnhO85qYehGkd8gLrJ0cVn2wTiG/
RlNzYZj25vvVQ6LrutnErZuEvkpt8uJvsvejacnRSbvhLWCmxlUGK7/S12YFM0ZJTnj/QRAXBZjk
owVe8I7OlaJQCSqCw6XOQKi7aFY031JdHe8Vhc9XWeKntLT94iIWmtQTVaK00ZdGZXOsoJztFFUQ
nGKifxzjown3YNa3DQmeLMlkErYs/DR/NNLdU9ZVSB/KeSJfBvTnGnrvTJ5geHvJy2mwJxZ5pfSj
B4efJYJwS/Qc7K/4Jfm5O4K8f2wvbuagl60ZkouzMtTkW/u5Ia5uFYcSwnZFgev7dzUPk9oTjxDK
mbR6ba9rKnkKT8oHMFhWEM0MosEdX1m7ieoWJIuI1h7Ggm2Ps+tR9wB+nAjHqsyDrez0AKkc5bnc
hjFxBmg2xKG3zleQiwqp6GdvofLhmu7jIZSF87LzF8in+/w2bMaoMBMThum9Lna/DrYQWjg/gCy1
z7KjiELOPNTlBm8M6a05OC0IvjjnaJF5XXGjLyrDWkM/Iw+yTWzbdHoNZrynWeChB07lf+6s8nkx
YCHtb6bHTnNXOS6YVx+5cT5qyekjZ6WEyQozFp6DcE9CMZbilT5UPmi6iTzeBpaRpJIzocFlh9Kb
vydfTAKe1ur7r7S2swYC+NmMzob4/xOQzSzz2Nu6KZxNJWUunzOOQx5cfssBZQsIRma5CuXdov21
xMC4CV0/A2pknXNcyRGr9D9Lm9h5Tj71uu4Dw0y+biQBSEfzrzVIiImnaJfSPCQKxjMcbfaCcMD5
riO2b+s4K/nEnqgcJvbrO7x4/cX6C5M482vZKCCuq0ortGxaKuWQpHJQIjJsml7WuhV9jo1+cxll
NeGtGDjRw4/5oqXhiwLSoZ8XOZhFhjYnsoidzWYqVC6oAHK4WeFX/8g1r3HFSwhh/zPxYSCXO91K
3eGPw0ezm8uvrG7DxPEZ2lRpEmEPnBhrZZdtIPVLS5O9yuUR84NxWwY2Y09307H30S+ML5T1Q8C5
vH995NB0xf7j1Y5bmiy7itpxPDSciaTGIVIv15AZtptttRmCwJkT/BJqHR832rFdQW/1GrtwnXyc
sTPdUy5Vc5koysKh81oSKRYzyBXG3xAZJ6KL7vOmQIko5+/upRIoTC36C9/Dx3JcI20tI/X3XFsp
wAKAx4Cnx7FQk87LPP9ijz+y4hp6IvETd3dgLcPdEN6/BHX+Mm8eSGB70LUdTGqJ9D2mfUTM0a2n
jZZ3QU7SCh+0RXPX841xUH8LxKW6RXQTa6LelG2OohLWTn2HwAnYX0qqfno5h3ZnOcnHe/sPb1UZ
hsB6cnckGKUSTy9WP/VHc82U3CwOlhwEel535rVWu1Wx6tazdOYFT7UF8tRCTPQ7zllzk8Js7DId
AVBrDd8GCWbB76n4a1i0g2gdJA3nywCHm7qEF07kOy4OISfIfO0qLAKBRAL8gAERzgqn0wywQKsd
R/x0AJBo1CDv1cAs2QvKQq0fO0BqxGwUfJVr4WFB8pmmh82M2sOPH7Kdne+rldT7zIiIIH2OZMuV
v0Tviasid0etL1xGhgCAHPiOxry7W+kI00+oInd9q5Ib1rsdlFtrFE/e71P93jdHHrfrMpOK5BUI
zgDqZDzeMsOUgdVijSLY9bgwggnsZvOXo5f9+557IhMsdnMcm8ULYEUyGI0M2owMbYAowjDaHGPe
69pDL0AiWnoUmn0mmiaj5kmqLbg8KAoyW3ps2UbQ0mZ4zo7GvK3WEZp/O3+o0jsqEsfuRmr4arxs
fzyUAALJfVCvKwFgpnUMr1Eox7jPHvKiO9+UlrQClODJMOFyLpcqzOxiYK7vA1pwAuTCCyyUEg3e
hg57zhRvkDAYlkIGdtWhkWhqVmipWl8GqTPm9ykTqIelCDjHTdXvT9tyLrKOT9UxX/M3QoPj5uyA
DRqnT8ylNpBUX4Hxr8TguzlUSerXzWXHh28E6zhuOEkiP9QCfybF3PPlmOpYAT4yCAYdd+4Rh5Ea
2GIND/OqtZeIPOb1YmcM7o8mMBMu7v4h3oN3Ulh5l3s0uq3SgiX0izZ6Ej1DMECxn4Te8t/FHgY6
Gpm+xRjEQTrhSAOqWnGxp4OK1kaH5gyEU5ynxVaMZ/EHES0kUXxsmZQVkYJ5LG9nnPnAEF56T4/J
lLKT+D5+XYCb1CU8JSiJ0euQeiBMVFX9VpFZHsl2UYGEoCxnkUHDQ8YRpwb28KzW+xuSPiR9MK3r
65t8qaMtLrls5NnABFBW24eJuhqIa3YOVZQjDJfsAFh4mMDhcGlfeh1egRXpYSS+neCphXLcMxR+
cQHgdMfZaO5ATqcPxp2/WmALmf9mX6wEeunsb4v5E1idYtRQnRV1kdaeEWJMmTBxJK27ZG+RIIb5
wKzbYRQjOXFz9nP5fxBwebV8DFLRAHfiELrR4W1+RCEAvouZ6nXWsjIA/1juyGFUPP8nmd191qFw
u4/zThaM2Qg6BEzMToH9cR3FBZkBox3qLvOLOEa0cY70wJh9gEPtMsmZUmDSTw5YRFu3Y6mqVziU
ZMQx7RrLg0mEjz91P7v1xKw6ZoXf7CLfV50HF6TnMkeOXHuBhBBTL4waeYGPJMzyk4Heb4broXYv
oMUwfUbAQltEwwaRLfSLbplfTGiOyiVJr+W88niDKyFbnxb4THwhMJebaVQBmgoaL+cVPnBUk54y
SZMW4RemsK/sVJnh03Q8bwg8bAjTRArnJ0+GDdRYEQJu62XD+S6PGgVSnltbcXwXdkgF+BSPM35N
CzorS9rT4rcdJ1bF7fvAgH6QnoHIYR2/pazqk4LGBIQZ48chSYLN++2EBBL3bNA00OIiEIEK/MNK
77w1rIRldr0e0RGY6K8q/BOR9hc+aNFPjDYk5quDtXTJqH7pznhtn69QSLhW+gt/OgHhijxKmdfZ
84KLv798cCByo4RttnBNiSBfApuHgAKPL2D3Qov1Lb0gtOES79mXWO+ZVYsAK64VSX+IiClZbU4E
r0kNjYdhgHWUhA2qTQ5hq9upCaMf2ECMNezBZ6fiCxKG885ZXSWcJW/h3HQDKetlr2OmdSwo1epH
pNQnmhWdvy0J0cOABi7W7tWiAXbDUBgQYi67Q/5rrr/yZK+WjHumlWOjCgOCkJsAaG5czkaMmK1a
mqBlxNZwAwNCDoqvngQ88qqH4I1a/VJZpBw4CygM++fiuKKv9BHI5GTOKsaUhmMQjWQJQyVb4bu+
sSK53E5z3MXjTdvArgsXsi5CqAjqX2v7yHmHp2jSQ7QiobmP+iZkRqZWXt6vm8u/FJEX64c04gr1
1IZblgdGTG218Qqz9KrFpm9zPfDqS2AUF1jdaCy6l5u99n4EBjAi0+9vMEaCqeXSp/DONj71gA3O
tvROTsscwqYigpKnIWLQgt0OWMf/PgLIL9q0OmBtbD0cbmS8VzBl2pUm4ME4OGdKyDeHW7DCR7v3
UQ6/gULZssKhurNV/5T6bd9u922jeZTJnDxS67wuZBZPImxg1Y3lm6BsU+Nbx99xey6Jj6TWATl0
bpCeHQ/mkbDyeBsHhENeAppcVtOSgAYcN8OyXLhZAr3ClNdHgzylHWZiFklUjF3gaGDUqfNk3Zl5
PBShuRKWu+gxukDdBolR8/nfxLMisVkbDyOstKjkzdIOfKusBZ98dghULC0Xp9/Dy26Z97PJW5p0
jhbo2S+8BZU3Jwesl/wTY3tztkjojfdRVC/8b+Dr1ui57uOVfYmPs/w47u3RluRTr7avg0POTPjv
61ZBYOry5xLtHaTeI8OXixqYBvsAovzBp3/O66ECyJP2V3F1s7fP3eNf+YJ6CmF6iVAhM3Lm/+2d
zHo6Mf6gU1nXPKsNPR8bBCjJqMs1AcAtVYiBSc990flYM2KDmqwgfx8z7rOybgat9sdy9YkH9qhB
VA8rbHHU4nrjjnus9nGMjoOqaQR1IUsZGOl1Q1ODLH1vjqgDIxRg9y6rNgrnUiwpvqOY0Vt0UfrD
0PaVc/gwDxnawIZY51KgS3UzCvqiJpueiH/7D51w0JNdRULDsBo1X2qxrHhUDcvWA+iJMieYBRXC
2M0UFacER8N6FOyxiWNTl30YRMpuY2t0iOls0e1KuNKvdlTlThmC7LyetEQctpj3ZaKl+eOoXAC/
cgr1cPyWKMyy7ywrbHJH1iBWO0PtKv10VdqRfRlK+3cdpgnjoKx712u8KcmkPhvGm/zKqsS5U/ks
HwapiuakpFzvf63NedlawArDgtql8R0bihZYqjRbqf4eveyQIL8cJhfW1Lfel5zcLx0L0dIQI7Gt
hZFfoJmQSA3RTK2IyE6NuDNjxtp9hu/CxREM5GO2Vz8Xm6fydMMwpdezZgWTrhkF+YOvpx1a4Zpy
GmwmdT6LRhle0bBBmPunN23EBM+M2DCFQ1oxqB6n6lh+36gNysPLz3TC8YHxv04Bta4FA/DFUV4G
fmDKa6v4488t91dXaPDRKJu3kRAmM9oZf0abPBMJ6GpqRPa8feRH9YD9penB2esmeotX2awoz/VZ
5nLq2QV14489fzhGecBYOQiqYkm0Ve3vQ3PXJ/TVhTe+T+9ii6+240sKgS3Wm8jD5cKbkObLiGqB
PINW0czgGJl+EYwAdGkeeAKhNJXIw5y9+GA03TP2M1fdrIq593fi5hkjQJpWadIV5k/4hOw1FQXd
I1Y96xl23R2kW6+XWQ4ElaZQi6oy3UeXEekCIX2Yrznxw7A3CThUMg+96LA1hLATJ6NUgoi6/jPi
S7cZp8oqDKM9C+mcOIMyVO7zauksHaCAUkALIniZ3UlShaVbVRgqQT8OBzn6LnH5YALsGOg/znWj
gAtSZC/6AEg1ZFyQXjGYZUCTvDWaHo2MS5bpKP5luR65FxJ5G9t3eCMCNCYE0hUPSTEnKgPsnyp4
9N4GW7ArKZIc9fv9gNPlcuOcbXs1xN3Zo2t9u0+P0GKyVqnMQgWUQWKWg4+t3kWBZJNOmi9y3diu
hJS2x4ZA15T8r97rbF4LkazJEIWchW0FggY6TKUqoTlUDRh22zff5Z3/FC3pL26TPLV06aTd6oAM
q1TkUmt7MC75RKv7M8z3kV08SxcKeeYc409VZGed1n41PQcMWQIGufaz58Vg7r6kPcm5hCN1aVmI
UskRw21HdEtvNvGgbIiv7ouz6mFwyQtiw4QnFx7U96BCLs2IkHza9aYj9JhrCarlhz2uL1PkdHcW
AAD43VqCYrSnuzCpw8zdg7K9fQuu714zuYxvaKQ0qpVzcFquVh6gKH2QqZfleQdfTshivWugB60i
yBoKdzIkkvoKJ/Z3tdOgo1ZVNANGVhZop8Atiea74JgVPAdA669caXhVaycfEMXjhKrwnXqp5mg9
/KLaF/d8iCmjXw/u4QpBAKrMnv5BDLMPao6KNR3t0KPNpy62PDUkl51wi5ch9g8ezuaxJmJIjEPy
K55Yd6sjsCt8gdThsHaaTGeKWXl1xGcwt7M5HCsNuHxwJ0OoxIoNQ5RM4SrkZRsb8lgZlEyfSVuT
TaulQFTZGIkVBITkSWogP8gSXCdLWCK1HxFDOa17HVZLkFAI7qUgzSkKLjGOMlMj1qzfzjjZLp0G
pInG9rdb4t0XPoOA1aNy/CLJaKdEcPI9BUvkpp7DWaxKIz0Dn2ExTO9ICTuScbXtEEkBAWvdUd1q
FQ0GveNXbwRP8g1aoQy1+fPMVO2dXWttrkv5edoamAxUqjEPaZ+9eI/Us1jfaGx8oAXukqDBhIif
LjBGXcMiQB75zyl9H0DMUpxsA7UqtKZe2alOxEV/DSlYsfkZhFXRl4IQpvAm1g7ExnTWlB+Eicyr
itcrrx7JVJ9uKvg7izaXQmp8YJuai7E22vQYXbF1FgKpGkXGnFrFrdil/nQjU2fvKzUaTm+nOA8W
g56WxTOv/Z8wsT66veJTiKOqS3+HuezcH1JE/CpJqofcOxrvhkIygi0CTX4NOnTGLg5RKBJ2V4J0
1G/C4Zxd1+5idH/sFVE2jhqKcyI2/yNmeb8EH5lJE8jcwCm3gXui0FZuqXZ2hcvHYSWYLAy83fVP
OZWCn/Q2qqnv8b04iymorp73ZBNIY14+nVx8y4RSzxwql9hrFCk5XhjVC9/s+3vGIVzULI8nZ4l6
ihruBE1Doan8pQ2+Qc6xzT1A6+Xq9AYByyJBM1zAkOVgPTLAojDNjvIrOd3+HW80hMVXaRWk349r
FQTpvcY+KD+NaoElFGKm0Rd/36yxL2NxE42OARLCucGG5BERjUUNABdyh99ta1hhAlImtF7FXIUy
Nwa/fNmhzseaUZ4Xuw3tQvuv6EJdyXyIhpu0dJZFm3trtXhgc3Q+xrht62Jm/IApIPnNYGjYS87o
1/ocXAoiNwZJAKryPhqLzqzqzjnaj1v+n4krsYkDl7k7Qqf8O012BuKv7IVzAfTPKFTiY71RpZeP
yZ/cwma/vDiROr8sj2upx7v1Rr4wwBhby2DEn2KcQ7/cf+7wPtY0KQ6XntWCQyPL+TJqYbHfGxux
NhlyRzY2I673Wv4vBQzrdx9bN38KEKseWPmgDMW8VMZZq4ofeyAUKW7KNavJlRVTkSdjIqArItMr
iMUw7P+ciI5SOuwvG/qyJ4Z392UZOCIrh38kQ9f3F6tLLbbv9gb3l1D2dbbf3wXghzc6268Hid0R
fs5ouqBqc3/850DtvfQdj6hku7VSoOISbUvH2WkuNPG5G7/ZiTEYlhL06XeyCt9CJZmXJ67KML4D
VYodhkwlDpXXI6cWL94WgapRWuqfDgl1NciSM6LVxh28bscKfb1fZv78oGEBfpC6PBHibnjHt/Dy
4FBfE0sfe5bJJkgngNR6+h9DCNWxFlmMgxFNx39hXEX+rqDL6yqsh4o3p4QpdTKMw+d5VAT4Sc24
WWKnSrMYCVhuxyFlU6VhjOplLZlmHbNsSCLPIvX5GYqtYr3DXxEkD0oxeu674olkFTqhAQzgEk0I
YS/YRG5Id3Y5NaxqQWyWvW81t5MABG73hOlY8HXzjtb6fhMpPW2w8Lpb/raAhbpQTsrY6qWcWsHc
8a/y6xgroVumh2mtwJoW844dvw5D+DN1KNiv6ICRh+eFqSaotcCtNiIAeoKc/AV80a+/LMZG+7Ff
nLh3RopFcI5YnL64kPEsZwkDpKOYAaPYBeq2ScMJQH+YNlzrQkV7W7eyKe75dHfFVVa+dCSSVlqE
cGFK0PhcUQ2vXRaX7CTQ1lMXjXsQElppB1GqtUTx/8fP0PMYP2ZT4rwLNctsiH07owbRWMXLyL5I
6g+FEwtOogCnpVAgWJgxMsoHBnGTFKL+dtKa/4YLReSgrjF1azxDV7b7wChBCanDJUcfkLqJQmK6
iA9hHK/rvmTCV4q3WT8sEXwLGX9CaX7w6R/XXtAmKPMdpSl39UugWEwKrnK8mCnftpa3jyzOMdHU
tp/LRqAQoa2LKCwo4CJY22liejhf56lj9SBGCo0PpjzREuRyLMyzg1Ezz9l21aeyISV2sZYsmGLw
efmo4Ph9gp3a8rtz2NOU80iLaxxreYHRwRFZa2cV0sKegCXGzA4JIUJ3vOexpHjsm6mfgIFvXoT9
3aNK4vE5IYAmpZmrsKDbgyFs2/re8PYo/4WdVBNgpv8g6v17Qr9G1Fk1u6HiuSV3+PS22eC9psMr
b7XAUg61dJYbe7brKswRYJB6ef3+4x0CpxwCnyLX027MptdKjlJilbceKb2qYEPbpnOa+6Ssx98I
NG5bUErV6XoMr3YnecCcbTj8P5HW3SyCDyXdRoEoBCdb0QbdPifXbnFPxC/5qV/aCSN0UsLPunST
Bc2/Oj2cU3T+4J8K1NTv8BpOI/ceo8RrKCr4CCjPJp6hSup8O9OTKmu9XdpnvaLvqNeOLHVmycbj
i6o7Lg5LSNFu65dlE61bOkSsUS3WFEo8ZspyNnnqvT1XB9u7e9M1MpkKVBXSDN6eapbG8OqRViqY
e3dG52pku4duMTBtf+7L0MqMFEeyBU/JbB84sk9UNNbcmmGpSk5ZW5aamI20vOlGVD7OeRCvXqBv
KLgd1VxKua6CaRirq5FZXfh7+vDvV0cO0ZX9pQSgH0VOSqbnkWd/9Oh0LwVagABfphpCkC3Dpbxg
mW2pX1XxNgrizJPqcr9G9SPAvm+MElnXRQcXFwtUldf4DPulpmSe8NBEnTjBw6jqhtjjeOgs+reT
xJxtChmQhLk0cjQ8rn8wV0CGPF5AyxRqddooKNBAf3R7ixqvqiYxMLcxawGDlQpTPFGb74VoC4a2
ukCoARAII9WAadjq/kb7zNVGYUqiJOIXC8qAExl3oZLOZG1SwClUh4NpAXiVWb8TdSokGedtfgHs
uUdwpd2u/xLK/xnYKLn4+iyis/n76+zQrBgxwYK0uGVPmIySAop4oYAPV40p7/ewrCi2sYm2O8uE
4O047dluVwNnaqlbZBSjt/yCEGdMs/l9DC4NAKU7pccCcS7GdFYljCxlGZTovSwQBKYqX9EBozt0
GbeI1v5lbZBBFTzdQY2dSH6h4PRrHVzAEeeAI88Qyc627Vz8gFpLZnBYR/iO2S5sH7cHu7KegJjy
aQX3o0RpevxbxLALcdYVXYvc02yW3MkB5LfgwkaqhWLFxMlSiqnheU8o5qru4GWzEXXzPzzXGPjy
Wa9eiktF6h0FCdXXSxeSjcAufQyt/VG9gYf9EjDb1+KmuQcZQ4fOeIJ+AlkgdPZG3yHZ6kM+Kf7x
DRbATlefNkndnC7RwgvnW5DAC+qb3pn4yVFnrDPOGT1+q0FPK2xkeoSWfBcnF/gDTQZYpy1Vwfr/
GmeJuLt5EBBuHdgO7UXE5rJPe7PiUJC+0xto4YrWv0eDG47J5O1hP70k5TLwAyuOPxWu+zJVX28i
8HTWxQeUfvJvY4vdb2uoKHh1WUozJTlubeZtPkcNNiSmwpGmIPEzd+sPyCeB05O2WacHv+eISCvj
iV94Nga3RYMOe2TAgfb13gRSFiOcYgpIa1lmzYOVkYHhyXi2gjTK34oIKv3dezrRJB9DBBTMcLM1
8OOLQGoc0FaI/YClzRHpGmtWEfogaBl+oblkQn5ujWgfGRZ64DC9QSAmQ8WS6X2bMCGJ0elvsGU+
XdKeyFUhtQmKC1B+4DwhCwBTPz/ES0RZtITnNTldOjr9GG1B65y5K86F0ocRtEQS5EL1FXPrvCzh
uIhRqzPv541msc3arFgmv9cHgTW1JG/73apatGoQ1Ihcbt0kKzdMXlnqXr5+MylfltjcN1yqubXc
FK1yo2Fh11BPnZGVaO1lR3yFcY8xIIlwljMRmIcJuNya+LziAA71KJ2HN3WpvV5NUr5eZ54b2HRm
9xAWiQsenr48g9EB196F4OYrMtmTcTTkodeXAe8flNqdslVEK1uQp07JSk6ImzWT97byXxigCXAR
q7ratHTbmB+f5N6SLz6T624Ub16Mcq668r1AqSI5D4C+wgL/2kQ3Qys5v6660JEtN8a/GqoK9glX
UDFAZCQJW0Z075UCH3NXpCqYeyhWcA4EcamZIdmh2UllTzn2rEmw3xrgIH8R46iGe/kPWKFbT6pX
jQl3NpJ0pExg51sFuUO9S+lADXnB51DSljqwT6uTmJoHbuadCfXVM9Ot7Oacrdt+XpSwEZmYjACK
kD3Vr160R49RmVyiOGtmU4Ejr3LY4A5SFfwGcflVRDA82NXKxbO7nxTiznaro769fr7zPpwrPzg/
iae8YNDeqdWc8jSEMF48P5tpNwNa1hD3yxZYLtw6ibuXQg/QLvd0frxzpsXmh9vzVYeThBo1Y209
Y8AXCw23iziE0RS/7EDX8TwQBc0Kr5cWEGYH0D6AL9bxety2Yha8A29J/JH8k8PXRtPzN3GxN01l
pzBooc5pjwkcBzERIyEm3VmA/RT1YQ9I5sCZ7qf1eERrfjWkVAgRSvhZU1jrWyvjnein3kbv02ef
L/zqzgQ6+nQKKmzg2DCXNhppZVSRyJY7hnw6aiKpzLPNSKp89EVuis5Mw0mgPXAsIFDxnlds7/Z0
AOTU25z3yAQVSvqN/bgIT9GG8XfoFqIp94sNVACnmqpffDRtcYeaP/MTmMxltN4qPvr4YIhHExH4
EA1GYMn6aFFllG5Xotk3EacW2Y6iGQ05eJB0w8Hc+C7xs5l3b3C7p4dWlcJR7hxFz0uJMQir64vC
61+zwgTBYXcf8pWTOKvPY6tGDkzKLGoLnqszLS7BUy5dq5Kg3RzimNh3tsQArzGpjhqsVE9QgaBR
5BtpO+O57xmw/OE/n2POaSDzLARPp4YTXkTXRcrWZIJ0g7oRqD6fXkL6gdyCoYOJE5tXXrdyobSY
EqasEzS1mY/Qc+mkNyvacK3wTHEjXCbjCO08N5P5dcWgnmnxHEsl9rK1wLUoP6kHxh1iI6USqi1n
oKGhBINzUJa+32O2+Xj1Hey0zp1gXQPzHJUOt+ap/8lU7NklTIimK+LGwEKcPv350/iqk3goDgZz
9U4k8HhAHba+bwd8KqsdNfAQBjVjdPoQVyJWfz/BpOWTgerl4AFrxNXkAgk5VKxZEC8fCRvStdJd
HdQmRcRGLgqSmIQ0orhIFolQBglCmYcfKG7Wp/okvN+KzZ8KsjovhBm/FTE6B7I2AtnFbh972NnE
/qj8sTOMl56ni4kd+oiWLjVdRkfwDOpa3fxBhw0Q8jmirnXYoNeZMyc0XMRos6iMO5yDH5U6UjJ3
bXXNLoYQlGCZepkiThiMsCUlx7Kv+B0lPzeRy6vGoYQwCOqXV/NVTEwCvCmw0ctPvlt72VDVkoOq
3ByzzGqV1/RUkDEA4C73eMevJ34s1CiUaRHjh5jgIpmLnirGChjK5iDlJyjuSQPtG2H+wwhjjWuN
lEcfpYg6vOaCeTlO+WKnfMm5aslc9KUlfkECexpv9s7QkUESVx2OoZaI7yDCJ9wS0ouqof8c3gXw
3kWAhxHPe5K4MGbxQTcvZQLQ/tquvLg88oDRuj5V1oEyHuZTFbDzb8rx5jB7GbBxAvETQ/tFRrYg
+WudM2Y/YAJQMRyil+xDzE9RnicMJmoGcL0fwaUX6OYuC4rVYpcSEHbtMVZISXnt1LxM8SzKo6fK
v2bIMvpbhBk224P71Xi1hPTrveHaqZFd5w374UOpmAPt+iLOmPSL4MlTepZDDxKsa6tgZbWhM8xy
zLlwkPWQuGDme9+Ka8qnGrGj+T0X4syMHJP/F7G8EOkjOayw5syaNyXKYs610SNj5m5gxEQiQ6IH
zBigadVlLOdw5dI/iA//niEztTpJxPYD00t0PK+VgsjuFtuLlaxDXHNdMSL+smy07eG3GIzgLbht
ke+c1nB69IAQ0WK8ZiSZnzyQ8htG08eZU171W7mTZqfJ7wd2D8mSTsKtBCt9DyIC8HjLJfHUNeqv
Royn/0FT00WaNysIbYJHLXoFUwzZUJ5KvS+0hUjRUH/xrZnWb2k4qpuXTdJHa1WFqe9WrmBN618b
Kdn3CREU59owSPjZtlrAhLHkne6z2udrNUtSSP2neKQhFSMRBjAFvKGShH5+0ojMF3li9JKQdnZF
Qlnm4PQaUwCH8UboRbWLrdkT1GmjCGYvXl3M5sZBvqTBfS28bdYVEg==
`protect end_protected
