`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T9SzZY8k9gM9533XtJLJJkA/o+75gJmaKuOMoep9nwkvSLy1Jo67di/zYro0J9GKF2MDoM+xdUm1
JbcqDZ75Hw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dui2pA/UhqLaXatx9Z70nDBW19H1lO7dKPhN140V07Jc0L2D0YrpN0+8y39D1dI4yG1WkpVSgMFC
4B3SffF3OHMOB5cVjgRcHnx54QL9GaSEGOH1LoxwctA8gmSzkvmO8iRzhOvDgcczXOkCt+YXoT4s
dI3nTAWBI2a3XCOvbgg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JQb4pHLv43VbvjLeiQJp3sIaVgayZH2jIbOLxS/lF33brBhGOwcZGs2QFJP/0nlReGUheF+Xc6pR
0dkN+UbWw6xe2SJa9THc+uqNRi/AH5TgC1c8QmhmmJH0AmEl/CEJfIVMvEiSRzCNiNuW1K3PDsAE
a8P4/pEjz8Fsb08sFGA8vD7Ef3K/JwqC+FBjvZAoW9GwTiUA0EKoFk/wJe0ynb+j+yO33vcxzMa6
/9MexNMW9TQ+cHK7/DRnGd0DNdfhevWedoIUnAonlSIlBkUYIOpQKkvomESvW9MMqDxOGYQ5pSN0
kObpxMZj7lAUgd8VISAObqCyIx7CrBKgM+zSaQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WaLpv7BCNtvA9OZ28TETtjkauYBgURrqhVIKwtw0ZVyfFTqKRC9mtBWPZGCDBhLuuADPOgHsX3jj
aS63izHd0dSr1OYNmyh3v9MtBhLsxdGt/epV6Qmtum9fYv3kTMd7bNQS3UmaA1I+CMj3qhjSDudm
Rw31tvJDbSg7Vj4Y9c4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
joapmiOHjgcOy6kSpCaLwZJOHjP2ocHYZH41A2gdy9376SmNad0bsibThe95jKeHRdlkisAJ6fCz
w/dznlFTjV5LgMORrJ/iMFs4Yt79Uie1qUVi074PrvHqPGKKfTSxn9lROaw3OUHGAyNj8FdyKgPD
YV75YwlpOqgPp8w3C0r1qyY8IJIE0mnTPypK0MDZNJmOvXqRon1HpWzduGOCuNJGX1tovGduaMU3
4NSkrflmvq4eTglUE1oNgna3N1wPuJNgcIDwEfYR390A/614GIoON5WAHBV3KLGiLOtPZ/uh7X2g
ZNxD8MDdyNduMSTNIq0EX+g2eoSUXElNgk+7Dw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
lJFbW3BScupe60htgIKGGeowbMK7NiFmyzKFVON7ExhcIEE4DbV/kwLrHoTJUbGZjU+Xaim4Q4X5
kMW1J0BOuWGw7UXDbZSI1UZPVoUdtK/QnOOeJ4ZmM4qrlVRhblZngRHEWks44USH0nebXoruCmKT
ieV7M0xh7ALkpyHfX15j6PJwMGcZXwMjqZ5YgFJJ5ukVR6LbsaKXvpQmR2cpwT/RxfkrIZR9JvC4
J4z9BQcXJ0WsXKq2YkUwLt1GO01L641mx0XP4LtCdpJLWgfyWgnMLlP4lDlwn/j35BmA7QcveIsP
5pVDOpiiVExTVL5dqYokH02WxBMe15YZBscoSSmA4WGOojV1e8IVCnLl8egSGMc4m/jm7oBLkoBY
qv8IZrKuRd1Olf744Xh6Cy1KdrHmM2cqRuTkmIEV5Xuby+etbuWM287a0Y/RAicS6o+PrwfD0edV
BwITEYl/QuGUeGH83e9Dd236R7m10fEgWZP6UBleFtj3auocaBOpNIBKCYGNt3JXo+gPVdHgI9+5
dv8dzKJZAvD7ukqjt19qZeq4DU0rSs62ORlSEKaT05SlTNUcoDACD7w1lB2+53w4a0hH0W/OcjXt
OV3MHa/iTJOjqdUOBVnGUyy9F/gK5L/mYIer5o8U7EXxurQ9C4sBNlI8VdegJo9lIUiP9gBbniuq
n3nnU+d5P2Ki5E7V06Du1wkjgxs7UTpgt16bNRIY+c/ju3E/hZCyq/IebQS/iu9/gS6GU1liYRW4
edPF0nvdiD8pcwR8hB35ly7cgqak6wgAV1hADT99X+QlIlPibmg0jCRXkqnvFx8aR+b844iXSyDU
7LAZE3Rw9ZstZQ7tbuwhMZyMbQoy7CIFCYcfMGTK7eOFPjz0kAKiv0h9xz94qYbrN7l1XUjFcrTp
DIPotEcE3cW7fiWhHcrysHfLzWI3baxUYagURK+PYA0TGTb1rEYp1ZpxiYzs79A/ZoRilQAETZv1
d4UjbMljwZ9WCSS1BJJo4u+EljZdwWRr7bKLH0VdQn0zQRmVbBBfccRvkQi+V01ta8j2hdd4fHPl
Ma4683IvUtlJx42uZeqnmo8DnSupxAQsVIeLSdXG8yynsRfs+T0uAaXrqmz3AWytzn5IKpK5Jfky
NbDF0OXhIcJzADc0hzhkNDDEODzh9ddA7ZE/7M9a3drAgpAKzRgZsxCHBii8tMQAYwGWt87SKER5
xZS0WZnsceouoCB0EB/iIAkuBbROyQhxVwPK66Wfp0xmF/a25yrHsgfSbVoCaJjw1dgqRPVjsbzM
Xoh5iu4KAGJgX5tqpE09HN4WG2a9q7jA1MVsDfmvoWtyKB+AgbGDi8z/cL6pgZo28q5T4WMfesSZ
6D+//ymSWKXsQH9cRpS3Rfbdwm+Ihj6xybwVVsWBVg+CDEn8PG2aRKEp5ig3AqRMn2oHrgdIVKp3
tL4AZ2lILj1t3sgQGEBdDSuFMa6pLq8C/uh/I6vH4iHUWKu0AvVipwa9YL86sPQiCYMXS76j5UhB
h7y2edkVFfmbz6I5n4oMkVIO+85+jiTAoWD7gi0/fD8dZL8DjKe+Ct+4Bibnd5bEy77lhn/5RY4+
GwSSD4CCCHXsoLTC9O5tNH0KViRD4Yb+GrJb9eOBjkh9caHi2+B/Tcl3AaOgdSUJqo2k2gV0WsDj
pMTkVWfxibnKHpQTCl49wm0aeW/66hkURa0YFh9YpC5+Lq0Gg6yQTI7gFnZYEUMilCtPkcOF80XP
e6FMhcroP7KLAQ+4YpEp/Z1Dr2JbbOLkMBMMoeZtPOZEjjr30GpAO71K5zcidI7kjy2Kk4835Sjr
4YlZzGNlo/tZv02/tFqRR4bBKwtPoY+ncOl+PCRybUS14CWWmEm59RMdwF2hsS0DprivtUvMPfZi
UU+OH4LhXR4UgMOVCNXciGDRr3OpYSFlGdypEH/Nk87v/3ypfNOLEXrUYIVOOjJhuVO/Fw858HQU
kPK6Vf7I+t37xVSW3aryH7B+TQP4W114lBqsRXDl7ZpSlfpopb+iVnMqj+ZYIkajRoUAp2JYtUVw
crlZQUOOkLAjnkuCQw6omwmCMOxZ2mfwfzkb8SSlA+ivxkDQDXVkEnh05ae54rYnMhQSQf9EVdK4
iJzdusac9XWjXR22FQpycUm6iRLjUXoh0laT/sMcBuRp6C8Q04ULMlfzS89QKGRPUmJVGkWLXuaa
hlFTHjd2maysXju4KutQkM/nZc+G/U+seVChCY2B4KP6/paLejmBkagHUmMtQdnyZUvNZBMTttm1
DjXboxnNv5BKkquRSwOQbC+3LFSOO7bzILhbwnYC09Unw/fg0uJNc5HXGDMmqKUqbIkxln9pPmTP
9GZCptIGQU14nxuI4B5bZ6vkdrO10tloA3D+XrgJZfbtKl5amkHU8uy4HaNGQgbBgWP2NkZnSe7N
CG9HKsBIkCMuJdMN2eZyORfWpEVgmP2Y2etTjx0L0XgKaMyRA7NxmfmLllagZKOIo2ae9nUVZiEq
JVfWexfcsKlEPe+IsfyAliRTK4dRpLsESi8xRQMnzZJqSU2aj1XWdOG2vcC9AhMjOJQBRsO3rKBP
PNCM50XcPu6hsJ494X+0UHuKwmXDLYtrAZp7Dsbd3KpNzoWxLalLHzS0MXNypfjiC6Y7wM+UHYB1
3ZJ2VZuFMcBuZaoehfZyCQ5UC9DsZuMVC948+oonrvIB3HoaUxC5Hw4LVq6F06ValUU5lbPlFS2b
xh9TivFBTxik380m4Awwnrubo9AI9vV43meJ6kgoPiTb7Fbaw+oNu+arvp1JkWxMo+jfwkv+AmV1
+gXSlfum2CNOLf8V/IenlDHlHAlAO3EcBz8yQi3WCJSat+CQ1roB0CcndtYEuq0EMZ7UnoLuDki3
7KHM9g6B+V2FHlau4X0HzX2/FnqE8uoaQY9tJx7DDdlFR/OP+X4WFDyXirXtdhVSaMK4EBD5QTlH
46/7fWJwLP6JIUQZZg7eMhI/SaKZqTWZNodMTRZYOjgJXmPm0L5cjDCpgeTDhuCizp2FPMuyvtrF
2QAYWBqcA5fwK8ilYnh9hos7FbcgY1i/yVFZvxAix91W6ZH6QNQ/Iet5E85JfnuqqCFc621lidnv
uD+vsDXiGbqnZJT2VycVsvtLrxIpZb3fdIdMWVhHnflI5Bx7ddp38uEo+Wd6xEx8MgQ7U2juRKPn
qlSndS8ili46r2tjCZwBSh4b+fkt1tTqgCCcURvSpSqQLi/56ZD26DeGZu4di329xBmJ9eQVJoft
erfotx06bVpU234iKwjrwJI8oE7D/Nyrwo2uE3eDHpiq9D7ykjEkoGjIkxjm2s/dVbpo/m4k6A3w
WRf0uqwhhAP+B4HfBGMXRVdJyig0loOu3EkKVV32RugnV4elxmKyyl4RjUvUVXtryYTu22zi7eFL
geo7lajlZ4K7AXvMjmK4p24m6hf570siho3ILQuFweGDkMm2yzsU1L/Y8DTa6oBOESABF7190AjE
cK+CF5JZjWtqCXyDGjPVEANEYCwf0AzFIYfN9uJkVYNxZEqXp4Vl6tGgk57l5YVdZoK/DV7DeZ3d
IolPFBQw/C1FjgghzAwTFYq+mQYBYb/rf0aOuRDKGLMjih6o72zO27lCH9I1StWgrZM4xSKkfUAn
ojXkuvxjZEP6+98U6hn9hG0DFrxekWJmEPaWGNKLJcS8axR+SyvMj/eBIAD8ef6y6kecDnaKWvPh
O0+JOH1L7xuOmqETss1ibyscpV6+UB4ElULxHuAMnRHfMIBJMJB4AaPs+hLcHNwDyEPgJtdyhDzi
yY0pP8DAkZm45lZ+hPe2aUXB+P7MqF1ksOUhsbqJ1RS6hOothXKKhb1YE0shj0aQavFuvjZW97KT
P3znRS+wcSDWcQMuLvyFiZiHc7KmUQcdJXAjM4Hjq6Xf88rP0ZYGDpxBHgwXYQJtVL0F/fU/ESwI
zviLR0e5L1XULqqXM+RPtdV/dMLqMkk8npcCMSsVwK6ZuG4ufYJH4a0vKurXXUaEslcBmjQ1zmXO
E56ezF/3RfGMBQmVtPiYqI8qqH+Rm+dAfoF2ZUO0cS68uY3KoXyQY6l5+zMMOBF0AOEZpX/0ArBz
YqHFhozbvX0airtIwfUg5SMqSickEB3A36H/u1mythHUO4lbIO1yGaQkSFeCSjkWT90ULs9pnHIY
SUzFOxqxneEyaBmWLTYoyLIg/X5g3i2iveuN3aBf3HciBOCIPVBvDebSDRzEt0/wVwVj8vFWEzrq
CyZuyzOUtL0T0i3VGzMe8aAS7RgCcpSC4+QGhqsHQ1GEmv4CAOEU6rHNnq/ybbzHd3jgPCcGxPzU
CZ6OoD8+WNLnXq97pmLTIAKtNYUZzQLNYoW2TO5BCaiHwedd/PORgqDDo8oBneN2FeUQh74wwSIj
NqGNAjwPDjURI7KyOzaD27SxHbtaNFaP9ObcpNI2ZQ0ZYrjZ75AQNwke8lD4kBcEjLYsMT+8819Z
BTqswvAk0NarytDXbC2ta6QwQallc7X6xVnQquCFJV+AJ6xkdHSrBrDBHDL0zNP2AUOQLjEB9FlL
MwkgJm3RJtlddk0xsV38u3qUOZ6SsGVNuaZv3BI3YS79ohiDru57ypYx1SfWDkZZRTJLL9yuuEyd
UvHmtiUtO/W4kNSp8sSHzuRuEZWWzSaR9RyNFmjiCHT0EffogdYUXefI2BFwy3202CZ3sXDH5iZC
yztFPbg3CF1SMG7j3e8gbobrucc1mgO182V2mnLwA0aYwSiaAAEIcm/u5oulZWeSadyPiAFg3F1M
EcjVdqxlc7w+/PmlT5hQb7ofwFwqkTiXpYF65ncx42XZgV0Ndxe0XFnmHuBAPblWkbthtWRCjXSG
t28+odyUcvKacfl9SFYkbsDTLF5gwKTjgwSkJVFeR0K37z4pmN6sBQdlo2n1euXcc6WfItQ0+64F
HlXRx23vWcaNZepNakUjcuEQDLw+iADnLDWvKkpwQMZUj0kX/pZg4p/2x30UdRJxMltvtYKv4gt3
0wGf0FpL0+m2biUE4gZiE8DainNHL8ovaHMVKheDPY1/dMa87JBixA5poYzYNhBTXwDgTYiiYhCB
ZbcQzbQFjnXKT1imwNqbSmnX8A/k90cNiDDcr8Exn9Wh5j/up9SmK1vCa9jBBA0dEFh8RHF5EJ5F
e4Znoo4pyzDtmk2vB3u066QZ7ase6J0bNUiP1MR26YOEQsO5dqFM9yIgo1DrpnoJArQ8wakTjUbd
6/xuHoDrphFyw8LdrWMlNyjf/AKfMTVjhNm7G2UgthmdTPa2f+r3Wz/X3v/TO4wh65OZJbmxyGiO
XmP6rcINevxJNP6EAvwmc1O1J4/5jRbIWBcnp4xes8KbsiS2AfaLRA656kiGg0ENiP2SeWEb3zuK
HsZKd5LH0Lo/DWZUBXhyO7xWZi6vN9hDpY5iarIW4LXFrZJqri8g1z41fLZkipNOdl/fWz3l1H9b
oKA5un3WVwHf/up0if8prxBSwuVfVmD6Qk8awZjn4mkPuNmOpH2f/FcXXdbCd8bPvXDpF4YLBWiF
1CqwgVOEL8pBwKmBb+4p6NgiuXTDseBEFIjaGaaRS5uPZAJK1OF4iXNiwT6crWYWlc6l4vA9/cv7
3QpU7pzudibGkt9I3nyTvxzD8ggYmVNuR1Z6WZrkiiMnYlKYeUkxko0rKResVes0VeLnQpgDNEYG
UN6IwNImrWsWxAUu2DHN1LSTa/z8efOo5p8Gxyj8bNjAXz964o1YX/8ISdEWIcV5XCWEurVuXNbH
EwZUWVYveGFuUWTridbT9Zyi+u/gwx+xNSIEeQuTs+wqF4atHfO/kb11lJGdQbvS58v5CUc0e+NC
yKbB53SkCzJR7vhFIGz+3IDyScbMuOAMNhp893tmtc7KJTbnUgRyeSx4eehneLOqGX5JwY0vDk4n
bffP1mJBDQ8ze6AmcXRwJio7VDAIEUDOqe5ZWzK7lHGyg/AWyiNk6Gx3s+VsQ2NbsdfWoH4TAD+q
NenKE4zPmhkgPj4Tc7JlGL67WJtU8xOeDYuKocx6ja7sFNGsd6ZomXdROipWScx03BNO3WJJWq5z
D8EskiTFOih6OZxohS/qi5ceFrayF3OU9PYgUW4WRUNZc2Q6zezpmhHyFMnb1Wn2sUnoiYW2fsGG
m7AP0ZnzEIfhXywQqLIt+W2KXEw76PkcY+NhyFYx+/q1AMTwg3gQFbbhgHQv/fkyfxTqE08ClVS5
unosOQ0+AkZb4mo1P+BZQ7I008kjPhvyysDn4vTQwPWfnuy27kBltcbLp8emjsjlaVV1GXm6rBm2
5dv8rQJ9/ovc/CN4hFhpY92QkE5ZUbXDRGXFjXrTivFbySH3DAHPZmE+lm+Cj/7y4rJ4aepn3Lbw
4ldZtsO/WgoVyb+ugbcGgwGGVmsDo2Q+irQwjWemfvNfACQSXi0cnXbIq7W5FRd7GgtyR3Ww0vZk
o/Hfu2jQH8q9TN9XR5pIgeePPWZOQrTckYBvLPksSiOpvho9ENyDqBoF+qhenE7z6ukp6w9VmaC4
IY8JQ+1dKcjkahuYwy7ELhToebN7W2SEC7qS+0Nk0PZGz2eLznOcz2rX4Femi+vmgsqCPu7sIhEr
nk9l4I0ck9V/qRMF12PXRTmBQzC9o+tD5nMH11j16aT0LeAnQLOppAFktyiGxHtuxxwnJQ6ub9vA
7+hVo1u32YR5XyzM1Ob/IDuUEu+WyepU5QXABJDCKCi31iRR0HYuN4bJY5Krij5pRwJdt3zhbBl0
sjQlW+QQn0uGlhT2IbNpxgXSRABwgDGjg5P6lIJ8zi7a148sCHSk1sTOeSh2IuzI8Xa+6WkflFA5
zLE9lgD/5HLPz/kBCt/6N8qDzzEjM5SiXL6QKUQhfAnlvEqHTQ0GRowAt3THI4vl9XgfXF8Z0C1q
kRbzqqOcis4pMQSsHPDFML7aCWCglPRrdUAMymz9GiB+F6w1Hqkhqpz4xq2l5aMI7ph7F5KdNDkN
3sQx0jHNsd535DBA/YoiuJJUMLyHFa4xM2mHDF4FwH8agw6vc8znFmXJFUOUm5ht0pSK/X/+bC+H
olTJme1CPF6hwODL+jsoKJ8YoqEnrYaUoLUthkbeR4W4tRg5Gr8tY9gqa8NYri5sKB1Suhbb2f56
E2kiGrnTk0A8ovuZO/+gWscbqJX1QDZ3dmMTp9ZMzJIC07NjkRKFkQZkh4+Ob1le6M+wBYjlvwcu
oPk+frRYYarP1mKjinATee9YB7S5BSC8a6b8azyKOE+7lxQ2fSmIurJBs2EoX4kFTAOOBjeJeLe5
oY2DPU1ctCxDOJnu2AC90oMa1adVHR2JThS0SOdJ1PY33dd7rVCzBMMpKdFtmJjds1R21ev5Skyg
HG8W7PSbh/x8wyb1OX2Ad9TatnYMAgELF6Utyf423EPCbf1cpAtkxD2zJx/4wzd/MLjHidTHJUX7
aBmPh1+uM2/q1uv1S8EmoSKo3sKYdgYRBA3LTtmks4HKO/FAI8zgdDSG1vhDqJFBPE5zdI9zNRdd
ylVqLwLMQByyPmD1SKnT7PChLK2pAigwqYRpbtLzWX8fhn54oYe6DySX1IbI8hpS21ZwgdbFvX7W
f88dhkbW2E/8SSNU9y5sHeevTSgnt50H+4x4Ps3M/Du1ZFqsVXpPYZ4i19kJzL36ndfqZAm62QU2
MT06Y5pPix1L+Gg6a8FMksPysuPzdV+KjbKAvN4CjdbFl+/i65MZbDyCGwTJA3lhQQIA
`protect end_protected
