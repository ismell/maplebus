`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Nph735vcwPEfJiMwGddBoodEOG0acsPojQBbpHCKS08PbAewG4oah31eUV1q2e0NnBpLI1FmJVyA
K+GCFHJEHw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l6bczCTB2+vO/FDn1u0WwxHss/Yg6pxGjIpr0z+F7Yr7f426L2t6kMQenD5BobhU7xvdr3NdtVYC
TX9B1vr2gxhpgS/orzuw7u5/CUJrjxIqggV6ry+S646KMho9tVJqlG8xcdZYCzUz39BvJdjsIeML
i9rH7jm3KyWk+23No/g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VtO19K1iZmHHH9bc8vtEdLEMt4DyHf0PfOgKz5k4h06KWbeMYQNt1qgBZbujNgqga6UA3EvDQ3r7
L7n56CL2WovskhVdBlwuo5yRMD/t5ffg4CXYOeu66A05FyKYOAfUsZjNMDs3p0npWC1U1Mxfv+Vx
h+bAIHknihMzrheAzvtv0sq40P7p8THogr14G6sPvCSrgWKbM/zSQT4lLAiDehXQSQKFCgT28l9j
uOGHO8R5T7LmwQ6x+y3mBPK3YnU6gFRbJTj/gynSf5qaXRdbxb78EO0/0IsZ2/n5OQYAVaILRuNm
fPyLxx1KTT+grUhvwK7JQi9ygtEXk2MnM9lBGg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jW58T5PH2727EQrzb8b0O1Qgfx64N0KKwJPbuNVZJd/BM7938bibGAyYVU3GnE+AB3CP3gyV7UZa
U8DIYajgzWaEWyfe53PoU/tAP36Pp52wtBnXM6VeOhV7J55azDiwaxQXL85u1/3keJlZvmWdB5YN
++Mr8E0ek50XHeUDfwk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XdsEecMreUbBhbVfOZXheTGdOYKeRS4Kgmu/2hmyaDn9lWZ3ejkG3ZpSKH6oGdzT9X8p0TDS24Am
Z7T6HdCNtF8ieYl6dQYg2snOIyGZqQ6NVTy2Utg/5WvaYUToAsh+K/Hmp77RE2UFc/D7p9aZcvmQ
Z7OT/OPHxv0vsW0I2ZYA2h2L/ZWsZk47Pu9/6zPLi6B81x3r1q6UYBXl6wPw47FEa+T4AAA1dopQ
60MnL9wUl//jr0L9TFhaCaHOw5LBTtHV695NYWE8Q5qi7OcBVCV3wpC8DaSXct3tpjuUo5D4xrYM
BHfq63o3GYYMDDiza5WcG/jdAqbyjvCV9rEVKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30640)
`protect data_block
+u+gFJeDm1jEnqyjOKhDlEkN++D8xF8t95kEtV48CvawuaogIUQUwqFMadsz5JXt+4RYj2+hN+J7
+zFFtQN/aHZQQhokj7ztHo2EN/70wRQS+1+JfAfeQz1HmSe5cSh86A/iMfpXt128YayF+hr6mJ7N
Hhl3sLQem8EL6IKyIGJiy9E6MPn5RRNU8Pp51Zu1q3IhLn/r/Zs3QxGIp8Y2OxYvoDNU+/vPxswU
OmZkzdz11oDcg8Sy1uVWWXTj+DltwXrETY7iAkAGn1Iem5dhbK+8Mj3yriepZ0xLOHzugflbzif/
Nb3OeX0xKPAhqnt1tlj8y9sUybrHirO/nsAxX9UR8/CRMYhZNFqKP72wGsiTbNGPZua6mST/l7Ng
eOiRQjKrGhavYcNrb6DkdTLOQX4esDCA0v4zRUfptX98xZcKIJ8MEIzpaoE/a8kJRSv6eH354IFY
djtKpJoH5Cb0jpleLGjuBDv5IVL6IKEVNFUNnSE8T0j9fNZtETrSZ6tjIzd6DM2WXK/ByaxQrr8i
WoX9m8BM2R6wrV4dOPvWJsmJEnYEpWK62rRqZbY+jENItspJxBGEORVKcF3THJZZU9S6ULXYzX0j
JalmPwramVASyqelfezP9Ajq3NSTBunidkwQHUQRSJ5G8YZrbIky5XeLMYtmLKvt6Nq401gJiTk2
3bfTpTYmzrA49BQy0uzJO5R+Xd9ymubM/52MOJOaCQEO10ZfG7XsMznOKvenHTZatQjiST5JoWkK
2wqSVNtx59dVjV0OyoczQBTreBxgTq/SnI28MeVA97uth4K2zAn4/XMeTEikO0lo6c2bMLtk4faB
tk8i7OtO+ZfYdNNqNjVY/Prz49+zrhg0k10ssqSIE6sUDngUpIbG3s7JBIMkY8s4qh45OSXECCQ3
GZBZo2R0JoRMhVIWqwbjtlJ/dInTKmhShXh+fiHgWIejNKU60wcn1Ku4EgXJvFZ+X100CB1hfX1A
GYm00ny3xyLRnAtAMKL7oy/0wqX6fY3DwwrVuaUi0yf+8vZ4VjEd7bDhrP88hrsA65u+vGN1nDbc
QarNwUQFfdgAN4qmJnZGKt6R/SH5dKe9l/nT5ptEttIfRhWRVl9ceNY5ncKDmwIyye8um2b3WTB9
WPCS3oZ7gcn/8R5MSHXQgV/cgU/4ISSly0nHGiRaMp6eWVtfZv9Dw5tN3VG3BCEizKDmGk8Yz2B3
Z06H/j0W2caLOa7iyy6M/gXNbOCVi2ZsZOcz0IGWbTa0SCkhTRvsinsmxq9wGMcujWhK3AWqVdrr
ftt7xqElCnzOibgJfzybZqoGm16DmCcxV4cLS1fcCbjNalUTL15l7xIErMl/A+c5w8gC5VOvnFz7
Lp1rhRnzHBG8DGrfqELMcsrNILN5A5+2Kk5I8UNk4VOgAu20a33iKKVVC4Rlb0RKsO7A9dJwjcqw
SBR3c/ABwhFCh0NJAcnsbITp+DDr1dP2Px+LvNtzPtHp80hqGoMexN8sv5BeiQq3+7WZU3XcxMc0
WcabhytkGONntZb9J00rov2LX8dtGWB1OkCctMoAG3qcCuaR1egIWL6SvPXoxdemKztWc9xi8fUm
BxY2vJibh/aKw2vmGqsw8XHLNHv/Fgq0hNvfZ7CitkpLPB90IZKtqZ6pIM/7jUC0HeAL05MESIX3
OIDjIkeVnGctTMAUBt9cJY+L2pDLMwKEKeHqHaB8sCUUmGkEs53U1ts8Lzruco2huf8I9MZIrRJn
z1w4wGBaJxp3WDa3Jl3g6k/UPWN+QP/qYewLpbhjJvWVm2w1Vr1TueZe2EjmCMHtjoBcnqqZ+AFU
dReUlzfWneqfoxQT1hi3EDauFn226nOPQxUFS7IAyR3g9anMwPg43j5Y2fxvXmR00dozAccxb6+V
1xVtJz1K0z/hilGD/WhpJPVHMhkWnkg6ujOBFo35eiVqDyI/2BORMPKN7HflgJNF8dP7n4twFvsF
xUYZ8fw91nJdnZr7TwMzzAX12wNHm0/vsM9It2X91w0+jQ5qjSMbQIJJYskNCLrEibfiRlhYXXr4
p3/qRDWCcwgW6KLT37D3IAmljGLfkrk4FNkrS9UaDzMK6Flh4AKfAmBSDIp1Ag0FFLgsJaBYxvv4
RkyUSh3Lh8cIk51IGSbEBHJ2dXTF97UYC9248SwYs0QPbpgisOMy5+bI4iF4U1O/9AZv2XesaPeQ
aReqsjiEzYPiAbLQLYXgH/2/Qa6kz1OIOu2dIshHmCP1SF8Fq3LqqZhBiLzWIVEbNb8nwACdNpgY
vsvqg9fiV/nPL7IyuIxJaUifjqKacnXl+zvUE9SKJ2ohfdKVjLy9Bd00FP+rh5vpSa1IYjnPs0m5
zf/++LuacVUeYdnu9Y3qAE1f611FselwaD1fRbztBmHG1d2PEV54lj6IODu3O9kIxyxjhff1t2dx
sNrv1WLEO/iDFkArt8SMa8fLphTUR8C3Qp1IbPZm11Tge3nfaQaU61dqQBGKLmhIOJo6zmb/Hdi7
nompBo4XNJcVKubXXW35E0spIXXyGnT5A2AK+tBkDoxHBQhBYglra/S9Zf8v1Dj58Nl0FCQeqZNr
qyoG/yRGvKO0TF6NXAszz54yISWtKNBW5FnbOM1zEeW4V3Ab+XXn0Dkw8XzgzuccZE4LA6uAYa6h
fL6MRDbc8/L3pErytbnyBCal8HumImCSVKlDTINhxVh3s8Vxf2TvGhgm264YwCbq9/j74bbIzfBe
X5lN3Ri744fIoexnEvUPU6SCoMNcPZ9TLW5qDPqO33rrNSGWzCWqL2AVwP1RqTUNg/qsRN6JGG6J
Y9j59n8QxZuKloQ8HKEQ1lUT9GyxvdNZe7LRfeRjw6paBi+NP0l9Qz46qK5hSJqA/l7GUKmNqdyO
/r3uxXQC7+43jQ2vxqAGL9VZjFGtqZlnltb0ys1ntOQV5sK0EijegXSTFsjzkXINIVlmi8c/RL4m
c/6TLiIZzpW4ZcoAUorIsaumNfTH34+5zlVfINk6sD5u84EgDzbL1mRU0/SUWOUu0MBuDap9ENid
Y7PfKMk1SsfB0Zjh5cW0l0t6j4SfsEQWllTa2dKlR2OBataXwru6VyjYrg8bqRb2ohcZSyamLcCJ
QClyEaue0yCzyE12Z7C+Z0BcuFFGZLcGjG30mhM087ZXC9avgq5gnHJv6TRzoggp8o/JlL/HYR1Y
LGdaTQTLK8N0kw2LpS9zDgswp1kIzEdcKlWX/q1Fw8H3dUNDwI5aj3Dunsq8HpZVjlbO1a2uYVZe
P7/kaICdLFQLYzlKeH5tz3NCw0CMMuJ/SiHdZugSYiHGy0aeFjoYUkZc17SbND7SuRgTNoi6V8EE
OV+eV1X8g66MdagkoVFqImqobWJmWktD2wIgEAyTUn1tmC3ei7/AS9mYscbcZjFRf8InElF1wBv6
DHL6U2Mj3CUIeSH1YgAxlhUELha4RB/7yYy5Tnjern+HSB4ebuAwzcMlhbI4ADPtqsAWtslp3tb9
VG8QtaTyT+49fW2il4idSfYCeWTgC5+hwJwPPKr9jEf+zX90KS/tts+mtNEGVHdyHMnJ3E0+wy2i
eOh0tP0R7dERNENx5f4nP/Q0AnWLxHjkw+dOzmXHXGtf5MQigFLExgkSfQICvO6brF7isqFJ56Zh
dyYrrG1DRjN7FsqmuKJCMYrEzxF89Axicru5du/TiLG7xAh+8wSetwEHzI05tIjUkdd/sF7Jyz99
Es8efaR1rey6DBbaauPgEA/EnUGaF84I0CdXPVO0eJAE8exN8363LO57rwAGqjWUXaaW1yB47HmW
AQ8jyU5c1uxQM8/o4ASXs8RnLlMN+q+SopOAUj0Rq8GpOM713kwf/f4SMFyuskUqPa6QWjkavqu4
zTe9ZIr1djP6UkPLrLnIZEEXokgTgPIcq9zdfSAfZ9A2tMQ3xCKSHh4SJT1Pd+dqyi/WSxRXf3hX
//GEwlGKpJAWZW22jd3OaHFGTW2UG4S3uit9JkS33mC0kwaWs2n4n28hVrJqRd2sOXf/MsYqjlnz
J+8ysB3HGHZcn5aw1g6sol3W/WWBTxKMjUk8lfkRMlnji2cW44fUj6QB336ePYfgd2Ih4+BNylJK
L5yK4gP5ZCshX+uYV0z28ATsmoMQkYbI1lA+eNho/kkicRz8pVvuk1Pq/NZclIoyFTFgjL1MYAE9
xPd6yeREy+g8ehjBwvLyESAotQd17LQ74iF36vHjO7ayuqxKi4GBAW2qLBeZMQmldKsuAOSqtyGv
MuaYoYZ/YQinhBRmFGUuTgB7Hn75o6AfF1AWfZlsUiDHv68CfLDfZ9gVCaxqlMk0yhh7MvZo/8Lf
p+NcrOYoX4IrzmNelFSm3wzw/KWzE9bF+PHtU7Al8oIJ6F5RMFYLBhjGxD3tSGKTAPs5obTOsyfl
RlrJ/Y4xVrerAalg3b6mklT2+R7VpA2A2NUXTzeqVn4iCQd148Srk8jdu/3xs+NLExRPUgIu0OBx
I3a6veWW/zPmli+suLJuKvrc8jiLuG8hlXdRxzG/yoPZtEH5w3kqQNb+NV5+bNqg/i/IyGShDG+M
H7c/9I2d8h9vuGrmk94KFrymGCm3KE9j2Ibhg8d0gOsRnw61z6Wsqt7asTSESCxOvNgT75jlId9n
KGqmQT+4SiIQ3X+lovmxBx9x6X1i2cGPuceZMWauAFjAUb1Unqond5Q9rBKK7Up7tBi5mVSmLuor
T/xA5b3Lz8eB3FOaWZ1sIYr9joW7Uhd8jvcCiELmFOoTYEB0goNsncdJVccnGpUrIPi2kGgrgJ/U
bmU4SbLzMesMDHMt113ZOYlCtTenNyr9TtPMHw8yVs2tP7xxMHVRwObzqu1jRIIiH+Al640THUGp
qP1iOLB7e/DH0zAPAb8KQRF7EEwxjz4j0YFr+2iFm/Z47ZfTOsRKd7ALnwpfnsprmlfh+XUj3njo
PW+UsxXuIWvDDFXbDIFCjthFAcNNUdHdE+hnmcljBm4ARzrW4G/a0PMfq3Wi5fmil1fFz5f7+TnS
UE8OFKRBq3wN+fYXIjz7WUaZANwaHMPtW6yTT4DLz6cvLhohA1/XoV7dXLd58rQ/HgQyO7lcDfb6
cgGZnyO1lKpY6zbH4PwVKtyb3d6HMQQSAOd+MCyQDN9vaG0JKBZCowKTMp8XK/ZwhF0VzUZlyseF
5ouX8OJV4c6i6QKFoIrk2/Bb0I4Psx6/s8dErwiOkwKT09cVw7UiQTpDlHUrFuo7nkEzSU0mNafx
XOXkYBtLrkHF2539LEMWHiR5zxkDipZfz/3vycwOYZydWFbdGI5R8vr09ULCStvLTaxOl89+euAX
bObAcBSlyVVe9gjK6MDvg/1+0hLsXcgeqZoJUdaSa6PjjXoMaSrAEZrRaQzeXQnC7R7zQYHJePMo
ltLc4ayHe2x0WNRZZy1po04ZFShFf0j1bKi0cGgEjeSSjJtVgsW2RK8+hhl2ZBW8W5fJFweKE1Zw
IrNiIiAF+ifbsyQWAXeXl7C3XJzXcoMw3ssFewQO7b5RpvAgWFfF+0qpTKg0ds3Oi3aieJvbkf60
IREQJRENPzAa3IleueCwk0Z6rzlexCSzZ+I7yNjlo79m7IoIGKGeXldZVoftZR1lLz9+o/PKwOSU
yD1EZXfzHQfDHeTz3CEe5/s4YWQ5GJGC8sEYtD/pNZv2RKnMkNKo51mIivkMh2Crv3T5G0H62qaO
rMm4CT6KejVxficFZqBFwr/wveMZgqo5GC19jEjo4J3UIHCYDmGirWxE2cEXj2EhZ+EfbFsB9ENL
cJ9AksGbWz53QfNbH71BihPjHnIWjpBFcfVGzQ1WTzvZdVpfxyt+1kScct/P1/VG5ameChLagbZd
qxfGuV7O2UQ6opasl7UjW4mUKYbJ3JK3+/xUXNNNmVcmaOCH7fv34a2BU1c7ZXExerjPaTkt9Lz1
ixjROYNKsVk7kCEeJx8NytkUJCsiWmcKJv2fOdOEOTZ3I5rjNz+wLCIW7E7x/H4SWQ3kLPey6S+S
9ZuCUzb1xJ6Ou61yhnUDeZzAI9vMQDt9RPYOcWOTfXDRr6N5L5nLRrwQiCU1AmyzlINGREPtqSLB
eFvvSiQpGzPOUo0ZsPwp4HtApdEagnPb6aPJsQ+Tsyn80bsYoEaVCC4YviNDsgSEViJGf4Yj5JAA
ewchw6gcY2s6tX6jTYkPUkSRg2N2Yr0aXcvRGHJMZ3amG/rhKKkiWQu+BspU99ScYM3Trghihch8
mowpsM+4JfCbrqJfby8bQ9JDPKKPXDLCwYxaCcrp1BpkuzJLXjQOGq1uiLx29jK3qD8cAsfMxgdp
4X6kUtnue8BQtirHpTHZhPbHjWPmAwLNAcKtjDZNmJODy52wvVaNQdSmJNccCgBJSFuuvR+L8rzD
D1QMw9acPM6mTkc72VLZVLpTIKaqmyMWLAxYHdiE8Zb7kpiItab0jszF7wMowfNO0HOxkUTJPCqM
s8cdVcZHSaBhvzl9T1Vm2nAqUNUBrADXpAsub2yXi7P2kRjVV31TlxD4in+wruZpoxnmbSwVQuHI
7w+cqSusAYkBvbuhz40+pZnOlB/o1YDmgTQAkckIBJml9iUytmlSjgaIqe5L5BF9blo4sEqbQkls
j400X1twnomXQkda26t9o30j37tPUy8q2qDBX+VIHI8Pd1CGxBmPHZ1FJdB/OWW6MRJXl/ud777k
9AJTD/mlbGk8INsNdM2mO9njAQ1IpJQ6LN2d+RANWwFT9TjmusxGac9PVO/+wy4hOum0CJlGSOKh
vxJ3CpvJK0BSDgGq2yRZywJnfH/W7ylegf4NkrTFfFwJmUNCsBSr15CXxtymggX9Ai6+IHArRF6p
5s5k7t6Z8IRT7i22ak+o1yd+HVbGPz89LshAIUK3PsazPBFF5jOB6n7zw4X9w+HSsjmtqvY30Ah2
5ZcElqP13OY1WAwVPTkuP+nLJakkZudwtWqd/cz+dQcl95oDQ0LZwtYbVd/QWpP5ZIeYTdy8zouJ
CiMq34NiXtGa4tMX0aWEQMaNiquVibRSopow2hzNOyBWDsOGaS+Q8rxmQcuqjUIsDHJb5R9vynPy
nxG7Q/shYjhq8s7FQmUsTrR5I1syCi2e0gWPAF2lV/B+xb/2Hh82H5MDDID9V5axzN1m+KTffefD
ivoWFAVkAxLTZOeenYnbnRd3Jpfk0o15lw0TtZ9uf4VztiMwA7TRHzXk4e+yyB52ZgQUCCnsk9fi
0MOeT8nCugfbNdWqzn8CYLVjcUxUfiNVNC+ychTcapKN02OCyqaaurCXgkFyxkTHPobQ4EJBGvBv
f6IyNWOFdqUVkRtB3DTnxOQUx4ElGzQNKFwCKROaKYwQXvbGhCp6ev3OYRme63+7hgpFWXpBlMzb
I0vfuLjIRYpUf64WFWNA+3Z6vULB2Z7NreG8MWehiV/aOiznkaHEHApZOxlLMB8P7UKC5XLbSMmV
nQLEW659pPcWLblBT9zFeH3PmBwJYZ9rgOdcQk5FW2G9uCgpaZmrPKWjRg5JoI9ftzukdQUm+iaG
WbkVDtNziXafIvKW90WXf/AoOgPYb3gXvspXx6IR7vhVCo4HwhyzM/k66yzijrZ2wn/vM2JBh0m2
4X+3CdjjJewNxrW2nNBzn7vc5YENUw18L9V+AvzgU3fLYf4wE251GYT6HjWX1s4pi4cXf0PeNkfC
N+GbBbG4XKZGffVYtHTg3KhWM0oEcXGHUKK7K4dCZmiz8pkWj7zSzwmAcb2Ut+6REG+qX5DyEZm4
BUsVzEyXuqV241W6LKkmJI5NNFq6xuUBlBP+rfVhMyiatNm6S2D/RQkWJE+VwtS25gQA5C0yYlXC
RYPJd4hE8p/Yl7EzAtH8lvBaKsnxKwKsHqja2BrOaIheab0iUtZyniI4GYctthfp04+He0a5P08X
eqjGVFsTg05spuqQu9nwaT3YA5nByTB/Hp4tNo6MOUPqzpvls49KEIBqo5av5feHVxBywfrxZl85
21AwYIjPJLPfImZnrOHjLdNz7z+A0j0t/AtFWmclQ+VGcTJNhI391SARbaMBzEGiaEW92F6GI298
Z6o+SHXA4yLCRbY+Wf5XqfHkf6Yn8sca9/s9rj9R0homWx1WHbHjTvbEba6BwNbZsCWdHAfz9rFL
fZCtk1YAKc7jGM0HqvyhaBnBEdq14p3a1c5OoQx5FS3F942pxO9EJPLqVpBtgL18U1LMxX2GMrs/
94WQ322gBH657fNfnN5niu3/VJpjJrjx3A5V2KxftUokfiHeVMvm8UGXhVDHh9+m0JakII7ONGZX
MwFJKkZq5WShm7gwcAtC20nd6zstuowTjYVZs45uWnq9jMUTLBuwPlum2Mgj+80wkhNEV5RO5D+F
MrDzPuctrihsFXXA4Jzs+h7ht9waVtQ14oQ967F6QQl5ynkxcq9XTyniUMeGqaCkovwj+d3i3INB
KjTAIE8MC/oJLfXnyEBmMCuepwiHPtej6ZO8I8BAs1vHnBTxWhe20jPOC8BSpIFJCXz42zky9hsB
U+KM0WYu0iFHjiToFE3n8WqGBy8lsO/RzbTP/uaBUn8b6Tyd4348PAGB87V+D7r7ulrhAYrfDvg+
iawjFfDn44JD8Q9eQVhwq3fK2hmesMUWzY7xLVmfKVjiumxfL4YBTSNWXI3+m0fm7hosPNFbu//f
nIIohov0hTxhx0j55bd1TRv5kfgAPDiLyJihwTQnYK9ufDcv0+5jaxJhVkRvy4epZIlfI7LM1v12
VpEp7/Lw9wt57ZYIJsyaE0L3OiA9ZI5VqY1gnOmIBN3DH2cYrw8HHFN92TV6+1yI7+DNlp3PKweu
+wqiRKTfKrgfRX7FQelMiJVAXwgom84tgB/1wWnIYCGQcBuPX6rnpr2lOEsZcqpkYPoTvQ9s9jW5
rdaIVjLHaOt/D1z28gnENpGWYMj9J5d1649wY+ayghWQzd9AUzIbqSX3UrbjTVtCUZ0yN64MZkK+
tBWl4Rv2uexr/kiOZf6vKBrzsvwp1XQ5CC1tCMyVuL1OPQ/H+Q+DBCPbQGr6iezG+ARYe4RaRS+e
KdUSwQm7uc0m3+tcu2WpchF7y/yApwSmmCFokDGAhuvvqVwPUdakbYmcmazRtGWOGBf4RMGGOVod
Gyci6tsJB+ONnV/MaJE2y7OkWDX4u98meT6K+PGxZKRV2sNuyWemlYyq/rFTyeMaVLVDzZ6gFPFW
Oq3VjdtvJ6vqAwcVv1fMEIyevjXY8b9zZ3JH5beFFIXAiYVW89B6nCX8TZApxNkXiE0TWkBxjmux
gvG4gvXgJ+iNdrWS+S18fBa3mWEaF4J/anqf7/ltbp8n9Zu1E3Z//S1khpglnbZpKtlNodNdzao4
BJVH/mOxY9oGvh+3w17QjO1MCo42ylWjM4e3Nb+SyGYVhf7tTRJEVB2QBrqh+3PyFvomu4SrnmfL
egIzQJZcXZGAwkbfznvkNUxmuZQMXZe0B/A4+PZZWoid2n3ksw0XT8jSMCkLoLACMj4dl1EWMwqk
hjCCF1fiSwTaq5vtnJlVPMUjDmFQI1QEHlhrJYLcGJkmGPO6P70ixapW1BUbmGZkgHDniwqw3WzC
quAghHhzpyBVOQlC4Y/r8AFOv/xk03HyTcAcYol204ft3u8L+OApLi2IhybYR9QsVJn23/RNMsV7
vJl6CbvOCi/XEaZcy+U9c4XkiJUe9n7CH5kpkMUxwA4Y66BUgaNAGz5KiwBFr8W9ADd8bZJDB/6g
NiGbjEb1VNuSF9o5MM9UTINKJo/ui/8RVHur2XFbCcovLWYxrd2S0TEecYQq+3zWUJyiuMXhmikf
adQ887Zqm9EJWJh2Wn3nSVNbIcLM+QJtKG9U7uKyZKheZj0gAP0hlqgS9mOkNRB7bh54BVly+cK1
JhVtbfvFTpPXrczunum7LT6ITj2nKmmELzHtDkLOgOhOcl/3X1tEkw5ntlT+f3yWw9dTlYQkOhly
ZhSoBozk7IFDviyN+b9ekaofumrGcUdw6fKqXJERFHQfNHxruJb/9zkdInZPsKgK4mkmbFmY9LbU
K6+gKcLXtztwv8UsJdtmFkWawUoKo5zFPWuzNyv71RxEwgKW1LnsaWEP580ncvCrurVtgw/3sPIP
UNzgoI9Gz9sqGo8XeDxaAnhL5ztIYfOXeH2LeXHrpUBs68p4d3Lhnpa/6lRKMaRUU6egrZWYY18V
U3KzVJawCM55lYVNOf46HpXVAHDOAntWq6cUW1VWFRBwD/Q5x+czb0WKhPa015FfQjiMzzZFjqoc
GqCjELRCsNsROh8RxA2SnFf90Sq9Ox37h3OeWfL8hjtiJjd/crUboGCENt21fwfyoowit1jnZjHy
F0ZQryZtLG9fM0cwghsxkv0yMPCJoVdwzYiMrL+Te1ET39d1aFMbh+plrV0zJ2inmFumW8xcE76W
H4gHYfbciffzPdP/xn4SZmGLif+S9iXZerHRhJsGmIx8MpqIs7bd1EQXdkjX/H/3F8g2lYvylFu4
znXS3UpR9MUwYq4FCaZcOee1a3RS6hrl+fPhHVfF54p1PzfS/vh/YWAKEzpihU7ad/UYt80lRBY2
O5rPp7gMK34ZknJ+cskQfu8mCgfw/XI9x4BnX/WR6M5ZAjpYJ4X7VviA1pCZ268CGOKN9NEa04wv
vyfIDcv3UJTKTuqykTO6I9L5wdlI8ET5hzvEsCZQfd2TuhFhuCpLiI7z7P15zGksAM7TZzpXKjbc
55vYTIMAFJDo/AOcemS8jcAIGrl3Nud1hlqZhRc9JrhX1r/qOPBmu+twkMRMBUHITP3KJxDjj9xJ
HhlNSt/T6immOTn4U/1apakvzk5fwujLSHLC9K65KApwyOdUyA7fKVCKA+ltK+XJS8DcpB8iOkT4
9q8KU1vjI+r2UAbfcrlaa5Y+B3Mn+5q91RIIPYdP2n2vdD+YuIe3Eg7wkpkLTIT7aRukxS07aA0l
Rf2EykbKm9mlRed6HGYbHZyyaG/K/1jQPCpiDoyTiEEDTc7dm28m1yNnKsjnnzAAfxodWSjUBlkB
9SsrBwNssrzJpkcOcpOigDESA8WgquX+dN4tWHVRRxq/a1HkSlfHR+1okRUaWPBdvJ07GUGIjqAG
x1RK3oqFhmJ8OmlBZ9nLTJRb935Ff4jno+HuUgPNlkwZPiGtO+CiBQ9WE4+fnMMxh/YTtsgIpkNc
ZnX+aE+3uxjgLwVkFAIbwGxH6nzFYvj41rt6c+YV84dYPrpVBcvL39WT0vNbB1p+OsGWjw2qpqb9
Stx922a5d5zDBOsX7rKbU4Kw8FmHXWNyy7h8OiglxWxA8PwwCOTqStrFmdS9+kg51LnQ0UdjBxi7
GGLZ/gFokgDkk6CggHs1z+wQPu9mm7c4PpSLLK9pKbYvh6U64K2jBisbDIuqTbHC/Pk9nJksy7qM
iJVqAheR6mx7T7oHM9BRAyGc0j6KwcFfPekAkqMjsukWqmj1MJb55G4aBOkl5xCIOOsIWtFNeNyt
+sNZ6jk2oktFhp99o3sT0wViea+CnGCicUvn4gt3CgbHQTZnqK5CP/3tHjs4BCgarqrxkH+z26l2
HPR+OffxWWddl69DJCpU3YuDB8Ts49KayvO9hvIOyVkwwR7hN2k03vMSbFZWe7OjA45huVhcucU2
Oze+85SYAZdwzq8SF0nv8ygJla/3AxtRxK7JErik/4N5fjRh6osrCCT8qjaWW0lIii+GJNzGz1oD
WkC+LEZGWu+LNIZLfYnbgI4NpeqKR/pI0X8Nd3xIktTU972KgslKnRGRmHWgXcC08ovBNzZooIe9
HFyKjnDAv+xQ7rR99hIkIbJYMBZNpMGRlkYtcVjC6sJwRQfzT9wueKmYyG32vEcKx78dI6rrvml0
2JeDRBWQuZSbFGmvrN6rtHIQbJS92PzQfQ6Zl3VVSCFoK/M5j9SsLShjA1TZBHGhfK0AwaM54b3s
+v7qfirnyiYTPs+FMuTcMfV/Q+ovOVyZ2DOolacOQvdb9FHdw0g6Fvd7khIIwql2x3yDJr6Rt2V0
SeUjVeCB3yUnihDkae6XDVbe9sv4GMrbKMWtF/XWnEY+Ezj5x3H01OtD9+8i8+b/7YO7I0ih2b2c
bLo7xdL4hPNjcvcquMsDXmZHNB1TSZsFO7p1GGVMzcc52S5VYFjEHagS1UL6lxg5QQ1t00eHs/Wz
m8Zqu5PuFVIeMCXEasNwqpV/96X01H5EdmMHMx21EJDXDiGB481wz5D1dkFdyHLfYQKI51hGV0rd
lLdXWoDDXv+YRAQNYCpiAensH5iZ3QwhSkFal41trMufSYYFSobnk/Gaot50emrti+TPkjbqhu8F
9W36r2QasEWcoNYYXQn7V0ZKycVfFNThJr8cPu0Mh4KOO/EE01uRay1kkIqbci/nd9l6l3us9M6e
W1WYwPL0uS3KEDLJkuJigoYI8oGZ4que7kj2QYmtRee/sObo9WDYsz1tq27WfZXrUA0YGnaCqbK1
7+KLQlASKGSlX7qgxYauFNceMMTM+SU1GrDk8xyFL+PLNMfhz4XSsdzNxCpOt+HMkMnmrpr8ruRu
tQEB13SyOxsXjCqpwwtaAe7+2X9Tuo1MWyGcyvBrfyRYMIv8ziy0q189FkMuQELg6NiZOcQ3sUGm
CYeF5qdRsG7eA+D7dg8KEEyvR3+O26lHukzgY1Eg1hVLK+prUPEig88FQtXC3RlNw4dfHMVYPBe+
0tNRm/TbuBe3PwFuftd7SHWscOhAbA78YgGnjRZiF5R/0sKcnz3nF02gmH2IIyxKonxAR++FnGPX
I5EjxRkxigSG6ijczfgkU8ryuxWfKJwNwFq0xJA7du8GVZe+Y9/nhEJDwuQF1N4JsTKDB8XzSM07
+k06G61juxyZFdqFDYJlYb3hd87rav2L0LgKLkQt77u3arHN0sPSPnSrObMOU9FcILFTHYyZp4Zs
A1BhyaXtR9CVkkOccRQM8qMN5VJiP6lr6IFLGRwsFcIWOCFWWUlM5hDHbkWeJpaoN1WhmK7BQV9h
8/sRBVnpp7Oez3oXx7SY5VLThqVl5k0Zbq2js6D6XFUApIjWo32hVlwJ5JWV3dEtVtGJK3PsyzUU
FzOV6EcZE4WPyNeebaAMGqGRMoLiOB/997OJFHuEpZ32ptjOTA7Dpd3IIrosJ10XfSpJiMMyxbX0
8K11P/IuH7somesNr7WELVodRrX0zXzkotLhkOJEgzFdwIskBUbzZJwHdhr1zZ+zNFwUYam7tNaN
KFACwS8Q5tm8+LgzptPY6UYHKglx4P3vys2/1lNohtwqi3gH0JWfobzjS3e0lhpQdSU8CCwVueFS
GLJQeqPeuHgWAil0YCDLytZe7hfH/EflM0lisfGA+MRc/Ihbk3CK8WPEF1J9EhHn7WJ0MQo6wTHo
X9t3BRIru5FKdpjDlQBMqjrC8/duS5abSmeZXKNCznwfVHHdBiUr2ylx+n1MdeJ4e7fh26C4g1p1
Drhwe9i5ABYay7NOjY8zItk4Z8FEPsCIgPdUO2EcS/zxTofEHtgSowjkfAWYaqZ1V2L8pvaOsXVD
yAFBTQGwoOPwe4Ydp63b6Cf/eoOJ46gcQYZOld4tGaf9+JzTpdg2BR9qm1LUYKWFoN6kvuG0WDtW
Rh6lBo7vnP884mn7JGpgpSO9QPABPbMz+nPibBIYnP/BjiatbNPm5aYx/lxSDzHFxHJzwCz1W5VL
yGAycw8JUH78hmySSvnDuy1WOBWoAVRdOirWEouvjZt+QigtW8OMafBgwSPcORUs/z5nrmb5mdgq
hgLN8eifvpSpgFhkKEICTcybaHsDpP6DQaGBb7lfIL9KcCTCjqY8c9YFwaKGCt0xPytcdKLCoVDk
HgvYoTdBldedeLqbRXvbrdxgwaRBs07/mkUONETOX20YTML2zMnseF0PFVMv/Nf8Ym82MCF3daBq
Si0IkYvxQjOnxR722kx3eEvAMeHG3myLxRKlM+PqlFfIP+cAIifTdmzNxa5KO6Xz/rELAgoCWueu
CSdgYZSmtLyaNY7tI+6LRZeBn6QyVhiOxcmQoZEFT5pFqFtkzhNV6P8it0Gu7FbuGYFYz0pVhvGV
1bx2w8ZRDZjdEU9xnxexLZUlblXQgnIfKEYCM3Um4Re5wEI/0BbJPjroMHYuw6K5kuSe4eFS2YjD
nEElr5kl2Dyua7ZIHXCmoHS/yD2EdUOsIooDuDLSvRoIWgVdFA23rtBJBXx7UZqeB1TApuPPrKfy
SZmFe6zuVw8EStiXvQ4wIvz9U1mbrpgBLHM35ILTyDWC2W5UnQrYyn5Vg9FqKPLkhei0jJq9p4ZU
NhUmRtgO4p72NKI0dfX73Vmf5qihlbAcHhlBbgtIrKw7fVD2qSJenp6QxHQaDtC8RuhT1vNy4Pdd
oyPnXNRc5pXrdr5ZXlL5WwnQpCO7u0baLahSZRElKb84b9VZyABOpX3CsiQ3guCjkY5THoJvgKWH
ruDHNPFdJQ4vEMQKEuHjbveL40s9uqMdb07myFit112UX7ZVmA9WPxqB5bS/qA3AD3yJgETYVsJB
vgqOdwCMoHVhEIwcpO0KZvyL9anyaY73HUlu4jrd7bZK4eQyQJK9Mo5qONtdzuOu3YYMPCYZzRC2
cPhTUt/gx8G/8Lj1zZgno0Nf5JglbtOQ8tuMznKOpXqbUbqsxKPxo0jINM9IRdnA/SLcAG7kJb5g
//sD406X2u9CgbRG2rT7Nb1iBUYyyaX1/0zu9r5nP6ORVK+PnoNm831JnA91Mjef/8GQAbLDEy8q
OyXEnD+x4MuMPT9494A6WuzZlU+hmV5iEK1T8XwQm7nakvHqtVQI7BxNIEc+J1E3nCkm3yQRuaof
QliRFLDVbEN03yNFmLjDVP9vz2IpWfZ8WKI5tlSjQPpOsl6Vr+msTvWz1Z2TGty9CG6U+4LA03fn
lzFAQNlwYXsByTREl6H0Au/zqCj0HJ0ONC5TO4SdvZEcQbi2bRyIPl4qpXbOW8WCCy2POsT9K3C6
TO5W/NzKaaRCePQJPv2hpC//kH/WScpBsp/Paq3KQk9hX+FmPvbL0Lzl1X8MrlhppUzvdy7USOf5
2qmV97AOBVMmxH96BlVz4PqXA01OhHJ30UsZb9pn512sg5NYgNObzL9OGkhWB5zJdtOlgyVEbrf1
RSTOkoU9NMk9RjAPBZURgZkerknirlpT0xbuYgod+lsO+2Y058GPhfMnJTengRnt+qwJOUS+YCDP
MPklFQtIBWS1tyNgFqeU0x2T4nLg9rpdRCZUL57xDgK7n3yvS+M8kUps97xCvjRxiB4o6aZNdQpy
CiEm0SJ3vtGvvR3ZYfz2pa5DwcpszBRRuSUQ5tSutPvzkxtkqB6EQrrNX4xGP/v+5Y6JihvorFAa
hyF0fEBDksHii44lx1cyJ2oeCCLURLUlyyhaRr+PvC6kTpnjcOW9WEn9++KdIZ/sFNP4uqelITx3
PGZHjapcfVWgSakz4AsFI0ovhR1FBjxqUqHowA9V6AK8kHQ+RZBUIOYmur6KTRVxYxeEUsxf/M6L
H1i0WthaOCMIyxh8s2F4fuHxeOaMtuIU18Xh/itxJnWNIk8DkAIuEuQPbzfAJUlO8VeDEjLD+ih6
MDA/n3+pFATTv7W0bvwoCSM7DIVyFkF1opI+uyK+isVcr0i6hV4y/eb68ZEntgXTrJ0AoYdeP19F
OT75cX86HyYa25ju0oOueD5x0Hcakg+edxlup3xOEqNXOHeh7hNZIwEgZQ7/IFi9r8VhkHX6fMX4
G5jD7QU+vSAIB1sRz5gLLcpSlDo6vP60Rqk75VWB2rnfTIYN9VL9QC+1+Lro0IdCE1jiewZdykyS
bLPcpGoxPqgaRB21jp7aNjuGNJKUgkH/kHaKLhGONn9qGVTtl3BWt0KBpMN/U0iYbiw0D08GNzH9
D43Z2Ufqmyh59ou+ph+oopWssZ9ebn09hNNOga7wvczBapvgZ2sF8ZMb0xiUpcsfuf9gPJV1izsc
rQEvpmGHGvKwBp9YT0To6PywRrViyGleLa5peuFCc3dba3t4rXGzB0sO+wtw/8dldGD0875r1iHJ
29ZG72GE/jEnYDYvYOh+xJ1qDOpNJTD//jP336BcYpeM3qSkXdieL0oztJBeSeopUwBaArAh4RfY
0KhXyb3sQ2l+P1p7qbIphlaY5dNlqk5RYd6dvFDVyrik56ZTeDb3RCzBYqduVjVtCcCjhTAgvmF/
pEK3VuZmtyGsdRw8KViDXdqyAXwGdD5jzhZQVTcpClWPnmc1KMMu6L43SQQFzXVFnungFhYJvTG6
vLBfHaw2iH89tbj7Iuvv+d01BYIw4VjYammqdMj1jXBwun0k8b67iyDIASvQGopBMvEFv15v+ZN+
t6fcDoWdaGVMadTMh6eYNw9zHiqbMbJkyd7mZNQCVzKfrf0IKiNjoUuEldxndEEQ3lv8h1AOQ7C7
ouM3jC0s+HPOPN0EDQemYlu0SeZHz82xGZuvn1iJmKi63jpTz2XY3U3Levs28TetBcPf2RXqAMkM
0SwMQpqm24ztYZ8/pBDzUWbr+73w2zZN/oyw8lmQbsMw5Ux3TpnsmDQTnFSVgEa3nKc59d9LX4Ks
pn7xGw5ef+YtW3U+cqr6Dcyp61+YDCY5lTPp73kFFF38LN881MgClJbk20xMaN2qWd9/L9vLFWVS
SNyZuPEPwmmHlJ5aU+2E545GPwMr6Z3xwu6myepG6f5ObX+BCue8GgV9Qr6mE/Lp0gS4ijZPQKLd
AyC+jux3RcZrCjbpaEYMjDKux5NBfs2uBoxaxNRrUfEULcaR+MqrjLMWRnLK65Ec8VPOad5xXwsw
J0/9Bx5B8WWtLgL4UxuSLt13qRb5pp9LB7ssrnb2j/wqVy0tsL0YGcM/K8qYrA96XptCaqQaqCW5
1jWSncCtH2pkUtEU03cD2LcjL+iX2YF/qWrQS4kLCwVdKCrgz8zpKhyLswmv6dFzkJ1tAjUQVNfH
e/WPtgQ6n5yXmBizHZebQudA8YCEM714HPYqd6vz5Hrob6ueWxKNvBEgsgwDk2TsG6ox0DMR0O1T
ODRN+w6vJxAdJqxP5Xa5KtU3j1mjvqkjvTsykBpxA4zXyfNozPyRyf+AYuGRgIAkgMeRV3v1/Aau
aoeC+o8vbVWuO+qXDkU2DYe5yvLhalX5fs2U3P6wjpv1dZT7ZwbT3kfppK9+mClVAZsdqBt1W2hZ
s9qHDzgHa2NNH2+eyMVNnQYw3TAZW+Vfuiwtdmujh0LlnFoeyi+BRGds4XIbCCAT7Vw3y9WB6hRq
JaBXM1uthP7xnsVrVn1efK/gCPcl/9rJ9zF2Cakyih1Veqi2XkdNWXF9SvWaXClfMujHnnWIRy0/
9R6gseqMfHxspFfE+Oe2IF2xKMn135GQhvRmuZsrtNSzCqwA+/Xf7vDcNtHZDG2oiLtE6FyTrVG5
kUj/yQhEoQSH7mfH6xxkChlRy+PqZM5NYlhF18Cxh+wsu/5hQAFH7U770DWMdKFr/f4o5uGvo+1S
kneRE8r6EjeDJIH3QJ6KlD+4CZuaqEvNxUMnuPQeqF0DhhI+RRarYxXNWga6uAmEHOqsnn5CbePe
dEsW0XOGEckVnVupd+j46LDaaCfREgQ2kNlBnAWzdH4D6QADTRYykj6tPLeeSUr4Klqf61SDlAyx
HcNym9riGYykArFxdJCJo01UDVuFVd/NmeVhwwGxtfVPdVZEaI+CsPMBZWVw2EL7mvhRS0iP69sh
R4h7bdhqbgjORB6yd70EJs7YTkTdAFO6XJ9rGu6R+CQJlOD0tItsL4rL8ABZOdLtbJda3t7Znw4V
4KLQxsAw0DR50pb1gw6SkX09/RbIQ3LhBH2xBgw0JIwm4Xn9UW7tRpukKgJtJCmYfV5QStt04p5f
WJLUbjHO8d7hY0gdfYMg5VkMtYY2ayWf6TNbUsAVr91gMl73CRrirg7qXxTKNujknCfp4hf2gNGo
56M13rZtOsRS8wxj3r5pVuMzlRwG/R4s5qHf+WDGY9Mr3l7DkPLIGSclvftgfsMpvv7FiiXKjLcZ
R10ewNw4Q/cKwLx6JElXhfwcGF7Ug1P7EVHSbfBrJp1gDvrgUTRg0orBkfDaIQj7gdBQ06ekJ9JK
tgNghSHl0ykU7KuF9xalRoDCRFBK1/okxWmFJimGva6LmJrgXPpGXMLMKibraCf9eG2e/t0Wbu1D
WftP18MJGg4QaVfQye6joJgIKeBbR18kx8CNa6qstm/5D9JHkcaQnovPzjd9IQZjVHgPo7UIEDvY
5ZgNFi5KpDxIwPmwyGGSDaWYZ/2tIQvpCze1jFnDsgqB3irsWZp6Sz2pO6k3oZoaKMPWg8sgULhh
tzol4SCy3EiFOuzwucc78NBVEKxr/Mo/JTi6upTPIkXqOtOhV3LRHErQ7lGBp+w52+n9DGrx2lUl
jctvNNNBpektszP+UZRdTKaODBoti6Ho0gI7MSuBUzusCUYP7aqVCFy9KNXBq/91TsWPL/iDkWeM
zta9Ex3IKc5naHGpNtvPT51jqxZlXn7Qauy5jiAVAjvhqvvlGdYSYB1V11fGRPitFAFOdem0ypRe
EiDQHgZOlO8/4jLspINbeV2KS8G2jck6c2pitL5DcHiqlG2+H+gZciS4kEXZeyHu04l37Jm8jHtH
fKEPKBDifaHWudIkieQ4pSCR83gsnfYlP0Jti+en4i89ru2gVGIt2gMakyrpAvAKMZpUc3OuoNLF
444o1vmrPbXsenhdgoSYkmTqg+FpAoGEKHx6bmDWPgcHfIiArIehvGBju+V5B1SJY8nYnMCZw1D1
lYHBJID2X9G59X7wIOqiHfoQhzJC+LmJfMBHwXH5ngzO0qpZt4yFhuewh6ot6ukAzM9zTrIolFeN
HCF1+TMEH1xZRwqDXIb0PdqOWdFtqOpm1dMBjJcUvgboF0V2aBuuotRNOdZ49vzqqkuIaZWp98k0
gLJXCD7OBzQjpSsfMZBgHynKv31S2uXl7VFWctCisTZEp8RG/+gdcvMwQTXADAdfZG1EikcwNv0U
X5m+2SG+78bNhb41WBMGGfYsOIYArDgFyF32XbxRBZ9S8VVSfcL+HXffbV9WT7hM9ZeVtkGPR74y
z/msBd++gkLyTOTwnOBBAL+Sbpow7pqUMA5PF9xDDgpmbLvHopYK/GiboydDRFzI4zEcgv4xvTya
Inh06VL/h7kAYpc1KpUPBTy28XeH7eXprowEVW5Jl31YQj0O9Wya9NV+e7uL6s1NukccOHpHsH1v
Dc6ooxS+P2ky3ydIRqfOlmItLjU3UCyfUYLn7vH99Rr9tXlw8kfNWcg4kaI5cWctVrbYbpkNsz7R
CbWu2zYUptQvwYDHIUQZ+QUcA5pLPWKLEHineqFu8vllMuxuW3sII1Ct5OlSxgBDfQDypKt/RZlr
VbT0ju3ndyVSm7NRW3yaUZAGu8XIkcaS4+ClkHAGa/mTcW7DVfQ2ce/wEVXwQtlg0VQpy9ymiXDz
VPGe0ESOGweYL+v4YmmHM8fzljbdiJRarkFVPrYrfuo6XWaGBSAsrPjS8x0NiSkFcjAou2Py89tU
jVPxz9axUpGzGqUnspCoU2VOE+rRYLdxhvAvwlVdQX46NL3aBLcwiYkcKgo3AgPDTj4ccBkahgpU
4H9QAx6A9qpigmojIBPWzRwm31E/KbBL8krCqlZXbkNixxQcSZEJEBayqPUkzz4ORD08yhpuuaL7
5MDqheF5SiycRR6ZCogr7omYBZzbaEj1ILYmiYNB6E3Oe5mZ7dMf8Z9yapWgnEX14hxjlJ3ekuUs
a0/P0+EZ9KUz9xxcsWLA1ZoKIGCB+XMm9kP/4N4nsVHaQ2o+IeWMFkpQi7Ga5zDaSG3inFHYlYZl
bTqmuuKPSnQ5pyiXrfeYLs+pofvc79jzcrWU7ypfssSu+d5lVmUGyO4MmH6EHwrJ8H4FADAGAQG6
6MV7F4zg9OTRDvkXAwiOx+Cmpxr7YsKSh/BsvstPFDKsuRtVSdzBBm683HVoWjGIpbr8sFBO0ON+
ESu3k/KVigw21sZ2FXUV3ltt/u6LnGuDSAl4kB8b7fW1esAxqBGZ9AB+CMjstMu3nX2oyNPGmpQ3
6VM6aXFxg/2D0PSLAo9F/4yBgtEpIClwxOxkiV2xbzeT2tfwuOz2Xp//SgZWF4QytWwrDoOTu1K+
POsHpl1Fm2kZ1YSr8UWHg/+a1Ztt2gXRKbiuJQ+mYhSfozrQflvKdYSwhZQ/vOBz6jRdQ2rm/GX4
f9YmZ3xAdbb7Xtz5urPn96ovANPljO8JheJWrZK2+hmd9JFLbAoPCaWxUgxt/nWl2thiKqEBJLH6
32aWHysVLO3kgjRwCT50yMV/mPvFqQGVVUHvlRytPk79N9PhWTVN4v5J6LXCISqxu8OHh2tjf48u
1lEKQC9WMm8FSgzxyfwUagm3c3FvYZ2lqx86im7IKjyyu6epitrjBPmu7d/IkU9EwUOtnhnRbo5m
y7OlV9sc4E9DNCWOUYltvO9LDlLxnMjpL4+euVDGwbbKptX7F19s4nvN+C/90nE1zIgW2oQNWISm
Oi4QJhhd2hgmRuqfd+W+vRxRy4cfruEUfPiRd4m/5vNOfMWpKc5MhpBHmI+DyMZ4ELco0Pm+yorF
3q7qEaGGqfdurrsfSx0ThYXCywvqnsvDAjDx8g8Dom6nPSFYJfgDEU6qV7fETMxZXcyl54OIB28c
sadFGgqMEnhXw53srDBpY8vG42XiHqdocl3jG/XW5ux+op/U92R+VbK/FZhTo2M1xdnB69OxCz3D
bbO5sRbXge8cFwjjPNhI3b1AB8Fe3h25tSiko2ktSxsHZvk0MpeW23EM0zXH27POp3asc+HdoLrj
vZyS14oHDhCXTNHekCMcX+cG23X6brvX1bb9pqX8fq0hBrKMmOJgPuhl3cMlrP+I89LAnJEJ2UPi
xjxRSU22J7QMxt9PEBOh4pbIpGjXJDxGZq8s9sHC50SXOIT16CyOyTQg5tjvJKOEY13A7QvD5Pch
ENC/hFjKzkELIrB2g1JoUtXJhGs2B7Cqjded+CmnddITYSUcUIa9NKcmDk4K6IIYDhzuj6O3teJH
IXvDv+V3uN7qAUzBxi45hy3NQHHEqrhvnVBkBtAT/gnKGDrMtvkYEms2Hj5o0AHEknQ6x5iZSpBk
xsTJ2mj5j3cnqU2si0EvZiEhIdtVkNppm0RmBVZIkI/NxRIyEfBD+Wd2LMCOS6Pv26EAoVNgZsdU
4544IT1Jq2VmTwIzsfIYJ0WMFmOxJLhlK2oL4Ayqwici8MKY3mGQk2bnmv0A1pM2rjDD+RLgWDRN
jXNIt6zNyOEjo9aXnnKSkKj2Wy5/IorxeJ/QAPU36ogrj7HnJHd+VfKxboIq0OUhUlFUKHVQFhXx
o2juSyd4mQXn+XgRoNLa4IoxcM++upuq9lXiYsz4RKIAYkwJ8YzRI02S6d9kOFEHbViRzAITMza1
Y6GuwrO3EWgNykDb0TyaBgY7UtYS0fZoqzarndSHLY4rUBVE3ueVRxd+gwgPyp2mtM7R0CrDfViT
vGrbMWEOpdjz8Sb+1NAq/WxNXASfh7yqghgd7pSkffcvWuN9riNpou59CxGdglqWk8M0ZH4nUzLp
nDi0guyBxCjGSnCT70wqYQS1O4BOgrGLaDF3fplDCHTtMC05u1HbG8EE6OicIKVFJz4VoOPv5K7m
huoNQKxzcrFUzaTJH+3VKUTwJbELjR19YXF+n6e0xHIgLDg2ycySlj8mGMvwjDfDwWLDST2v1yg7
0Mn63woh12BK2NaaowvqjdI38zuNP2ui9JPPC02WufzIW4d+2T3aD5yYVHuKaPMAZ3maCpX/L7hc
zkC2x36LGa6F8DYUpDl2skYQTaYLdiqx4UDtJsHpjE0SnbKvsi8SLB9yEVECvcb9+2fffKt+Z5UF
iUVtV8drT3K0B445/TZewPycKrOaaNozr73ZYI3l7NuHTF+b1m1mm2GH3K/+LbjtINQWBrIMcaZB
++B+Rw9Rh2R4hJuzzfle1UNHB5hIf0wnijjLnb5vFrFSVM6oxjgLdErWBQd/5Aq7GiN7H/LULSiL
IXweyfq0kM+MxFBOQIWousoXoZwkxfZp2o5zYKItL7jy9vhBPRQcMj80nWzSmZSQlAQjUGGW/Cle
YGpfVpXA473jQjaUyQMy3yyIv7mU0rgKxHmXHXJDvox7XMy+GCELZb2poG8XgC4sDd38d0EeDrm5
0kQngHrojzCYhnwNnI6suTx5LCMCmMJImcGcUn/MOgddhaFsse8OLq31qsnW7UNkugcLNZtMVN7F
j7l2RzezgmJ3264ZeP/g2dGNgxBc55c5WYVj8ycY71rwD+5ISWYfIGbSnforiA154ukgTTJPCQYO
1v/7eKtvOitILAJuF1Mh4gpR8ddh7njA44iMvh1axYQFRUenB8WH74QeCFP6qfF8N4AZZNrks4g2
J1Pke47XvFp1ineIQnV9p/W/uKjAtkaIPz9hIaI8iJQ4ax9UMdX4CBZN6knHiqm2mYNw8GyNqpEl
9SbFqCNBLWHQ4yUpGuPK2C0FAYyrbMPkNO+julT1B3mLxYDlcyvNG0nPgvp8e88OXQcsULJ3T5aU
dW+oHpeixdkrUTdWykSo/F+qedlBBM7SuaQ1YN+uahH47nbtelCdnf6e3QcKx12hAzEuJtbp9R5K
bfl6H46rKKLUs6lzfdRF2Y2pDrqIW7Qe2S65iOtwnLXmmZ6t2YpNoAbbVOUwfk6Chq6ilLFGh3Oj
AtC+fPLkSFCIfOMsJVRJcDMYpCerPA546fyt10HfGGE002fTvupG9kEEHKdBKGiM+VKZ61GaVPLe
9sLVdDVqw8RObAVcWZRfAe/GtAjXKRar7fT+yJCyyVnn0jU4j3YjdJUNMXqDQtiN04Cqg4A20Sc8
5KeA+T6Z4yp+RiQ7aJDE0b7ItTPdcWWg7EKEKhID5jkcNYpqNJ0ZwI1wZIpe7p0ze/9FaUv2WH/C
5jXKZ8aMfzIQqe+LutHScSLJX4vkL/1YAyvP3K35wLP3m+QWp33BvOaqIIExpWDOSWVo7ARk+FHo
QZa6DFGtYjTWEfu41m1vyFfUh7LpOmE5lgM6ZCiDoVcBoRpENv2zIlOzV2cUj7XqpVbB6ckvBKj6
02LIenhv1+JR3KXWArEMa8HAy0MoA4ne/tILdOOqJr/mjUWkTtYzvD0AytTIBDUCguleW0BUOBtR
mcpMX0YCTUgqK+O8qi7BVSJJMFREIKYTfSFZgwW3s1J5leLln320S0nNP8ozmxjQPtX9Xr8XiIFz
9O3QoY/DwAae1xPCDt5CQ/5/Hplp0FqN4qILdbJm2iCl/4PEGh/EyaHCyx4WqUyyFUKE6ex9wv47
v+1KqJya3z2/IIlNUzwK7en7RHfrnjeY6j7GdLqYmfshEbIceZQyWFWVA5EWZhMkmhbMeeKxoE6s
oaTohcQF260/u7rhCjZD2D9kApAOuWbd2/14LL4vk3wSEVHLhMWUaxhySERJbgRXEYRkmxOcE2y4
zmcbxPYstCwFWYR+iv4ECTG7BswcxQo4S9tHIfiOnkTszHcfW46sV6WHBQ1hObqXoYVAh7KS7BGi
78gaDgTRESZo4FbQOY7n9wHVfdmgDzrepf9JiT9aLAOvCY2M1aGSdi2CK6QRxGYDwW5j1GKhEksg
AdCYI3IbiYGVPSHEi9+hQSj8eVBiC9RIeU9yFWAZUXc8sm7u9Mo1QIa5O7LlqiDPBMFexpun7/jT
snKIGIb3jl2fCuqI0z2OaOvOIkIVj36+uD7jTYdeb6TJHrhcUVELbgG6+mL3cLDqGcuwP4Z/3H2N
F/k1drg7DXRd8Ewlv7N3Dg2Zo98E1gpmrhg1yqOtRqJifgCxKPMemXiX29RIXjqLpNxx45ynRFre
HX0ZiTBsQIdZOuF5bXv5oDqTOfT8mQ8YCj8F6icILbCnFxUlUlz4U+tNPa7vCwqbcJSpnq1S7SKp
RLxfbE//r3qW1cbfDchNwpA/rBC/KWgcnQYK+SBTu1pVOJMg5FE4cKCPjl1XwNJW/fPp2ZYm8ZGJ
YDoXqut/pfyWJBqxDIT+8rQQYXqD/lOVjmqeALeiLP9JVg312DbuJPBlqGTxntLVDK4Qhihhf5OJ
9GfSizFplS85tZNd5xLiYX5WNNNv4Rb9+Nf15EAFQV8d1VrT3yRST8f+OdFAQYBr++CoYT3lGW5j
2Wux4NV/bCnqKijc/cckM76EkOWyZ8ny1eiEzcoRr54Brf+H6YkIo4zeftNDeY95QHWHSy8l0lhH
026iAjbBnSE35yzMsMFkZ9fNBTjGFYjYJKwlCmqgqnLa3rQqpHE1jp1JKU2h9qhB+XFX1N7Cex53
3Px7hp2ft6+3fsEgNgfe+tvn5sXWxgAo5KTrYHyB56qFghFLE6LrrpLRfjKHS1b2N3DMscs6A2jy
RgqwhWhxE51kdQNvisXt0ivxp8YIwHE59of5JegClPCbIN+1IXzrKCBlFWw/iyxP1HSY21zBY5gz
R/ehS059lOarPzGNjmXlofuH29FGtSnLQC93+X4IA4Q9q1fyQ6gFAAZirLgc1cNLXWQJ9UMx+aWZ
lyfhU8K7RPGc/YdTgpNZfzLLsNDHt6+Oj0ysg8ir4UNBC8LG0cYPRPrXNi2ahRLBprB7/fxnza6a
FEpWpPPOkgb9uUFXLdSAm0uLQuXAoIcg55FvJ6A916heOWosAQgtkF3NkfL+gQhJUUezqxkuXAQf
vtq6Xn+WfkbSk433ewsCMtH9RPIfUa0BvC5mmLN5DGg8iiB5yjv5nRhWa3v1cvX/4LLdnf9l7i+Z
hWM0nmDRvW8NqvhWkqvsLxQkTanItE0B+/Ew2/29Wp17cdMDkU4/6RCZ+fuhSl5JiVGJ7ZxPthKR
d8UnchgpktaJ6FBMUuMiApQuXuVKAVvF/g+PyYRfsm9Vb93HH6yYJCEpdrdX1jwiaySz92tyDPEm
m0w81s/L/WqzjNHDf2MVPsdIfETEkrYAnXhUTMTjCj7UdAsyDsmUGWCX12zGZUPz4zVrJedxLsdR
DpnFLHnNbtPMXDJc//46s7vFOtWMjbYdpt3DbiQAMY0dY5bJWZyBCc+8rFxXo7edD/ZLUOwXkB/v
nNTvLhLMQtMzmrck6H6sgFUd4ACl9WPPpBtARbDGoJebR/swWhFzk/OnImabiAFq16Ovpm4EjFZs
HViP9pOCLj9Enjp2i79OzeGnlZXFE9E9J6uNdnBStWISjJ/ViIhqKyE27r2f3nat7OpgJQ7SHSLX
YEoVHDbxnht7ufyfndqFUI5NaiWG/z+NxMqfOsOBsBaae948XBG2Dg3cGOkV6EVigZAYvgpbOh8e
cW56+G+AbOMrQdy03AFbL3rTds6CT/mynCCb3xbqorD+qWLPqpUmqTMlkWMomzKPYzR82MHH2zCo
nu3rNjMSmecnGLC3+sOd0zidzEeyyMPCO6KZXlezsCr3LVn9zXUFc9d4cUVUbFlYL4FqkRtVDWEH
UjU5y6rLqA6pXzXjEuERLQkw52n8hAaERNx1bucbIyhCUAanuESfePhRRQtkfrZcd2NwZfvWrrcS
3zd/NX1B6bdurFe7MPFsxV0KkdAoXCC53ox7+l6ms7zLwzuf+MV4tT1tlmV+gOxbEltQXqvLUmyw
gGr6msDwmEvOU4HDBdt0KoNKGyPnuqgYl6Ls5N+4+o7fY9xdTv4KWbfoMkJtGBlqqSUpxt+XBpDU
39zbKbF/9K2/myLCzrUDKnWHkBDgDTcnLu8Zl+w9glGTpk/JnUk1AvvPUEdjUTugOsaydt0r6zRn
UQNpEXEICFoZK8E6Ph5p3mh+znuprYBtsi5iozgVzNK1Rr18CG2N2d7KsKeZSlJ2sbNR8dc0ozGn
4fDeW/Rc+fA1rNXme/M4/JNLEjZ6M9FCe51sbWWWvJaotriCPnkYF1XaJ82opgZoMnLtukLYa9Df
/Z6s+gWikkDGpZBNLpBp6cNeT1V2omAA4vY6oSU2NMa02xGBRvf3CDkcdpBrWs68Nf1ARoFfkSoc
3PWvQf+PY5A9Y+njgDq7SgXequy1kYYndxd/vvZGuWNZBY2p7Ur8kIOwDfmhYHGhkcZJBNMqejex
Le4MliGJa6Uo68HAcqrM8ovBTXmcFz7rLJKdXhJXNKAae0dBWVp54LMfq6a3WyhQ3/CdXPh5Vypi
+6FSdw6eC9gsK10Pi+oQTgOdU5bbTMDj++7nX7mfuVubB7Vq4Ut+nsWD4AJOwRcNg7Ylt2cDsMOq
3b9MqX5DBJ4cqM+MqUY2vAC/XbyzPPCwfKAYVdxYc2nZzY8LjcxJQXqnU89VFXERgfFPhh7E7g1w
/kFBToJ4CTtIeBMRI7tpf1wuiwyu90nuDv/SZQWCJowvPH/be7iIT3a2f0CuBP6iJQnzpeQ2Bgql
b/Q2y/WBDHngy7yICkyl80+1e5S/J1JyvzGRggl/PJKzJO1GvrfIsfxLGFCop5VhIFv00O7AIfro
/6UK633eyCaaWy4FTEFxU5XxuRPGB0l9fVK/1thmww55kPoxSglvpwPzARWLPt5AOBr4SB4IK918
AvNVOgN6I/xC/GOezQkqbPqHdp+GjaB29H1s+HZIQIlfW34r2MVVSe/9iul2e/zkPoqEkqV29KRK
vZhYNJvsK82H9YzIXk+PGm3D7oRE2agqlPiFTzoO6DGgz+lVJma3zf3Q1AIHDDq98PsnVfCWDl8C
kHjlFqz6n2h1BYbseldIoQ+xRVrunAof4NUxDxNng9N8BO4GYw7VKs3vpCjhOAtP5epbrt3tsbpE
jQ9ovIRGkq0nlVTPWO0iKrgQ+xVvxPEYcv5uI+6+d6/5y9CzGAmnEQDYr21c8T9ubjAvvGpephOs
hdHZnTuWjTRSJSS1wL/0f+zgZBnQjEfBbU05y64QGGTXt26FtUkjqsyIJN8dJMRBjoBwhQOcllgX
plTAk5hv3L7jy08c2gisGjeGyp3imK4yOs7HjazaNii52nF2nrvXKvmg7aXYzpoEuUcwv586+QuC
iFU8HO47LZ11chZiCYv19Ssn8nlUPYulVQBpaGk/c16Pg+X4IhbS1iP4cakZgoU7Pvn3I46LJKzb
KtG+L+L00OGXuns35719Pd9feLDj0wfM7NUlLj8D36ESqeRbRXTht0Hyl4tIYsB4Qy5Z351uec3G
xJLQede4Gevya083HcsBMVzuXMdnLThflJlVFFmR0aeEvdcE9THHjHW99IOZA0prcQyWA+ZupsrG
1uxchLGzWr+kXuqIZb6xvtM5hV3R3a1zIbvmmbODwL4pSrleHg2nLuF9KmzU/XFAATTecDqmErCR
NaDxIGDf1xc8c/W69kmRyLqC/FwnuZ52oH7SP12sj3Z/fJduazahQN79rxWYPEyHKI2c4jX0kcdq
lOqMhPMaeGY9fbkwRZ+C7LoGhHKSHJwiQud825RD0yimZNcZ9v5wa+VY30EmUhAPnOvah7mpQE9v
ZoG51dJb3+z4RhYNnI/mGSPjNi3mSIRec1987zAxqGDdVVqvvtWTXRoiH6I5/ZW906yxYcjIaIsC
5EK7KuLx+qDZpJYg09dHEWcU5xegTrZN7oeXusngWV3wpsgR/mSOGKnpl+L0ooJRyyrlHmvlSUtm
iyWV0yowyllF00M8iq277KOME2dKd3AdKePh4tAZVKNFCEi4LmSdDNitSWy/g5Ghelv8E0k3zOyx
+eNh7K7QyuEYTW0T3/yDocHdQLWwpCM4hj/g8DqBgOO1h4+pLEvnAPvn1fXqKmvKhnwFJQqmVVo3
5ez/ZzDESQ6/xbJDWhd0AmmJoYa+ZylDSXtYTJUmGN19L+LNfSlONsmGsQIoWy7135LSsWDVYf/e
vpoEjzRT7HIDhYToiXH01Di4JnyClPGbDdMNrNzcGJyz7/U8bT+movPuDoPhVXWMNXdIvJCLv/I6
Yir1+e/np/ewyJq6Xjz/sBUsyd9VSmV7aUDxZc6y8VJaN48zFPrZILZUHC/mjFXuoZVzrZQ32HvW
v3wKhPaoV8geFzS9y253zQV73mhp9uLgeqURS8kGBpNKFVDYTA+EZwuDKBU2rGkR9kxjfWJMGJdZ
xgDRYQYBkqxGN8hG5oJ/MQbuHpqblAWed4+zfl8fB0f6M109FAoevYpyhLF4ZClcizBIcERbzFyR
2MwhAOihr0E5vI7IC2LlfaVN3yR71eDVWiCq1yV8r6GNd7BPStUgMcz0pzpjIrM5BX2rkscr8qZg
BoPlFbvsBzySG8AaXBQCt1lZh7AXo/AVUGlHz6S73a4409sIgAEVQa03cKf8QCxm+apfgmskL29q
+hrijohH07G4gox8Qld6LkiWj1fbEiFpt6hrHPUDOhiWrk+aoYzC0WmmMPyZlztrRd48G2U5+LU6
5ZWy6mzxraHLPifogL/X8yoCj+kfEcySLpWW+p9YMxuLLG9GBujJZHCZJIvaxo6HgoflPmYmkES0
pwYSSoUu5fLxicbBOnDYSC6kjRzQLww6QjgMeUKn07OSMVmCs5t3m1kGGUoSFisoxvoA5XghzV3R
Lxz75MtAHREEXCPWzz1BcUqeAq4p/gVM+xk+O31+IJw0Bk2JJzH0NHeyRVL2UEGMIo1l27J7brpB
0UW0BVVqoGZZCfWqL9pLC39osJt2qEOJ5ifgpIbXf8qzTiPiLHsZ6ndSvf+uO0iamrUomtXvtBzy
+OUepbsdvGOe2oheeYn9C0u8dvtJQBxsOKFOfIReR6aMPIOq/gbLa2v45yDLKLNoWbCVxMc6ebIh
DZ+Fj8a91FBBPnSGeJfDFFLnAYK2B1Vwza+vfhYMHfJiSytZtTk+ixQwY/VHSB1A5UWCE9/hQEXF
aC95waSZM0Hj2D6PcQwdFPkMNXM9sVdgJZV3q1VbVh3iZQaiW/+xDkkOSIwkkyqMOPG357MRWHmU
jdvEHXnGgncB798Q4V3xFfyqdQFheHw8jwk4GZxFtzYeRRwdgYhcenS4LgSdB1fuovyWHSni7xEv
nklfXYObVrXpTxyzfmnFqQ8F0YDifjvmKzENjKrLIt3lylxhdgzemnY+cvyqOYkUGqTFz31xqm36
izMlFqPYY/BUx/baH/j+wVese5kOPZ4xmaIy8iOyF2fZkUafRWtP8gPT831L1DbbJwoz6vkT+Ijl
y4dKwqOo6QQeKi/lIMJMeZQ1O8rK9+9gNFg7A84OrlrwyzM+vD5+GarX1bFOVYQLm5PGR2cbK9vR
EfmJrsyU5EihJRf8CowgnV2L0ql5baX7wEGnmrA3g7UqLpt5qOf3mu3TxnyNzh7SCU3cBTTgTerN
byJM96wcjdR6JOqkLZt1kZ3V/iOmwkkEsRGJW8stScKWOq37w51VZWKFN/T6cjP6LCfIZS/M54LM
0OFAzuSKHIBpAK9FiijrYD+aja01p8ciKVquopjEf/pdf7491SGRCkgxr5yjMRujweFjP3HrsTrb
4nNZ5MrFLY4X2yTDkMQGJjexGP/FFZTwTdy/v2Qwt69/Y3lWCFsk+r5L0RjiploH5bHX8Vo0P9vR
d1ADo400QI3nLqhc5jonJ4jUxVC0sHVVnZH/rMC1i0kJJCUQ8Fw7CBWLqLTO7i5lepSVBriJ0Qbo
0djckulCxvVouKAdtV9Q+tlCVDLrgd0kJBzO0IY7oiaCOrqc7MjumwFw2pRTKCgn5+wmFeHykk/F
qgKTfheeMKcT24my8XnxOX852ff6IGs5fgDH1hX0Pxgyi5+KMDL2taiTuxaaNUSopYBkvQYEePaO
Mn0KKYQLN/zaVg6HgoMVvLcEvu4m1pkk81GnxVcBHu4AAR768+iAy4+G7Af3P06DaPl0SV4Qi/Ca
zAgWEwnwh/PicACZOeNCgEim42sw/RA3varyX3THl2jjHobfqt5A5WUSuRRpepVnCWRi0Ofpd65R
i26KIOBf9uK4cYwxSfRI36FcfuajideRvKhb88gWb0NA4AtFqIedFyT07upcudx9aZMrura66VU2
h2tYJdNZVC5+WYzU5OxD3pPiCdJV+uUsA6eUsQSL5wCHRE6KLaN6b4v2DmaMC+vA9KcB7ZzguiSu
d0GHieNfmc68V3GwHvasWRGVWy+4tkKlWaYQuzwHpUJ6hHw8aEgrB+HUoC0x9lZOIFhGcQLEq8rg
sqDEZLUh+Y0Dy4W3Iiq5lrAZW3drNZ/B4ipnXBu2IECTq8AS2Y7lQStHgLfADJpEByFPujPmQAlT
VlPNYPw2fR2gZXTVWPoaWiCR3X3jSfVvFW3hReqBmQPYcOyXrapLcrf5GDcenkE2XTpUsePqKGxJ
sOZSyRX4M8VF4d8hHyp2z9LlR+WMOV8gCYcqPLbxId7b0NLxE2T7TzsN6eytS8+Cw/GZfSTh7QrM
T+FhQuP/DUqWaCJU3jbEXpIGm4OsveTe5ZJkii4MLWdEZE1o6dmGqtl4QB2VowuXHg2T3Uy2ifZu
enak1lx7COBsrt39gR9k8hConkBG+zgORXyXsbUvmcEuRiB8p83VkUnzmXP4Jhx4zfF2i/sbE9ay
1GUVtHXMX3EZYjAh545BTSnhPfee8oajHS4hCpuBs0YfrYuGNaPZlzfBfP5OKM1hSOouiXwpxIot
Hnc6SwGzljW8N50kBFTULNn1Ewu5754x3liMaJ9BMYDH+2Bs6UoV+n6WUmWC9hPDZft0szmf/QcP
jIhQI6wkyMZTLAR7LA57oWYmN0G/qaRKvLttzVGkGO3Us1uZsa4Zxeq+6oZVIi74/TJUPxL8qXJS
Mk8hyGd8Fs2z/TgcGU+Jmln0i7EW2qXGHs70N2nObojzh8rdZSdhekrtVBeT739Sas5tUY4rcqro
Frh7DQi+Gy6kJG0QyxDilOnK71fgMc2sozCpwPFH11qPA7XsHTBegYvydJe4V/WelaUsYL7Fj9z9
a/Xtjx6LT73I4VmGSXQdQ1i1eeQ+0ANu18HxMBq9y3oPUio4RqYXjJb9rqhx5TYkxLyoocGYJtqA
/SBp6YJ19vDVyqbAvDZa47j05BkBYtlTZPIQ/ZRf6NOe2vjbV/6c7WuekPbAnBIh9oVWMx02+xCw
2VVG1tdBVqtG4gTqH4r0s829uw6vQML4d6LdPwtJEboC/CI43tVI9o1o4DTMfSFPDloiqJiE/CH1
dKNxWin4sBuRbp7RNDTnUGnLqBroVRjQRRLY794c7qu7alt3+1W1R1DUiZUdarFCyQ1t4tbNu6xc
ZMoGvfrMIG7DU3PbUg8FR2BPp/v38figD/LfX4m7sFVS+KsVsxiObpy1ivVuh0l13oKvMVuVy+ip
O4+xVIt7yLNi7+QLjObAFVKqXarHU838qdXlGZxvZTNKYYi/0XfRCxWbq6pXsPWqD5Puvbkm2jg/
bmyn5cSjNNKugUlnwADYXxFlQsA/fvn0KZGWK/nGoSmjBSMKvP2OsklX8S+Cd4IidWc/NlJoBho1
TW9j1R6qqpe9VwEebq3EQQKQ9zbUOTp7fH1C9u9QSkXf5lOAc326bnJ4oh94msMZta3vWIVYpxuW
ly3fO4B6F3b06uTHTwiYqaX/SnRvi/hxNpBd9iivFEo//XX9N7C9iTm8vW1ZBwkuWezSlwUTY4w/
Esiy+wGP2BADEDtDggsl785TlRMhCtP4SgMQZB9X7eERi1aQYf6eHnT+0u9gjRYb3OqAUHzlNE3Q
XSFosSF6VRw//EVv0ClZIgQKnJ1YrGsgh/z6fs8vKQb71rzRln4rUPgNHgC9Vn+Q0agvS+f5V0Gp
/c0YD7tosCYdd53QHfWuQj6AG/6CynDlWS2U1zQU822czMyj70uX52bEVZMRW0XEcAyjnH/JbBhg
/jbRZOACkcZYBkhSvZXzyrHfINiNon2X3KTaFBn0o2TVjwwZ9DCAntdyw1/bosEKH18NJioMNhJd
6AC1ll3fyOtwok2oyE7yy98J1bczJT4nNPN6k9gcWXErkB8053AW1S8jyKhwxM08qaieDV40e8Ia
8yw4Lg9xD4ZhoREp8rqRga6iIILjAR85g63oGmht3oWVgo3LhYpCl1vWEvMPynnlPRFygAhgTU73
vl6YMttdq8dj96/3eoixgz2fVzWKSmJEncd9a53KDiKduFcq4fRpeJmpC0T1+uZNc8ztEJglmP8m
E2jubltVVMQgecJtBd6LbCLzKndUe/v8LcytzIQ5GCS/0CcX9RxOvxmf702DYQC+ZVm5z52gT3C5
zz66dIjGR+kzUBIpLfHAcXxENI4afGyNUjwE/Ks3dKU6tvuH0gb5ob3OKZ7Nh2BOnOT1FWmDwyDT
CDBuPUOMc1Ee0gTrkObyN1y60h2CTsKs1gPfQlPUf1c2eacgYB2f3ZHv6wy4kqz/dgVnxUN7E6Jg
YQn2Ng+e0CqvADButl7BPGlkmHH5IpiPtYWwXjmRJLHRADQSMorLBtnRfko+mMK79ueZY0rRcSs5
ups3/4EG8/U4/06yDSFP712yGFppHSxlO+OZt56Yo2D2Xa2B48n1bJogOAnhJGfMVoVhZw3zGAia
CW6z0KiTPnRHo99zJitx/tBqC66eOWgaKsZY6TYPh1xUptQ0ErrQ68bgA55b3moitJlElIpKMDAa
vOnwRQLy5kKGAcNtj34PvSW3zIzbEfuFx4ZRhddvv2AjJcrCDVWfsfWt4PvblXt3zoNxJxeOhx3U
6lsquhp2HxSnYfp5VLOHb/xcHheRbcMEx3SjSIMvC3jgtvoHTU6R95boTvdUHVxpQAW23nfPpdSR
PxYXvQlJCX37RHfn+kHfRmw3CdzdvKffpM23vkwIBxURs5osG5TPFq9nsf174fC3d0rftAz1p2zM
vp8cZLqL2rr83O46lQQ0pbntmdef1eDNOI5x6AVYG+dQun1/aY16QwUKU+BenHWEI/FHYtwoqTtu
7hfbc38rnPXlqZdU6ckl7oBCuUlIaMobfV/7nQ2VVa9FgnG6mOjmh1Lp1jPH87AlGRgyPaussWva
PY6D6nUJhuUObjoNT/fflH4GC43F+dvWqU3chIKHEgUcdwBH6dns8NVHti7fk1NJvond/7MNDijO
iKI6A9lt8fMD24mF+wSTLTM1dMrepcv5JGuAfPkS2jkGK8e+lfu6J50MYCYRpVmt6cMGL45A/lfu
nvEf6Q3qpcgBYRLxpNpMolWB5YaMsQ2ePmjFSbKGeg50FVicQR4d+n30Z4KkUElcLzecFXT5NAoc
pYsedkt0WsFiHPVSSEM7drz8+tNYHugNf9cnjb5QKUv/Ks2wrBeQj0d1O1VndV0Zp4w133kLHPrj
k3g6YaO3ztoYN3nZ9yVadKJe6nm0KcifCno2r6wnFvnxXImVlOO8r2D5+PlQOH7971yOjSwSsoXj
JsFTjgmoEyGTWN1m2tGNamRmLemDHFRJ71HenQUHnkstrKXZ2QADsySRC7TVq4muS+WA4GkYicCZ
dJJ2tfAD41ijw80Qv7MEGHSjFCDIAqwmgjYwoNoeWu2u3nsE3V6RIClSjuVVDiqPuD4KfhuDFRcJ
Kvx8lUD70FBf1wvkA2BlPRhELV1WSXn4wswDVfa6V/am/AViSegEhwyPaUmxJDkYprDgXzEcz7eS
JDpuDRMaWrV7Zd0u3qKcNBAxwtXilDuH72oOfFDWS7vXHLb1cSSqAulHhHR0tn0CQrt2r1FveuGD
Ue8V4pEelfZzOFfmgxgw0malO+bGUg3a3Ol9XWECR+LBY5YGBMPk+dsQz41iCuBrcTvaZMmIhwil
jlWG5a6KCsybKl4KNVF7yMcRSKjWjIpC9c0bD9llDoaZIql3uBUJIRF42djgz3rmAlNWwdrW5RoV
RoXXZ/CZ0Fxo1XGrGTsT7V1TW0oqYxiHAl1NR7G+NCQz6btIuYF1DMsbpSh8BdfhIWjDgC1QrENT
WK9mGcb/EcyOvtr1ObKCA2spiO9WUjVYOYn54mttocOocxBNPe+CKwHCKKwL2Sy08RU11je5wt37
LkMI+y06/yl2v10O2pyC7vb92vUsijFP2oNtosWgoxw0TzPuB8d0YiM4iKPPzk+/8sdShOK92KRn
uukA63XR1ywP2CRC2E2kZqYrjh+nLtAdY6FzCdYzRo9xr+q1pry+yDFFKj80X4CGBbPeBbxKR0o/
Sk1GT0LRxRRKaiyrXokhjwA9kBwZkqRVS3lqxOafHNeBSb/RH8zEsoc+1fnIie4NevCQ2CcNIC/c
QyynHR9w0tzMyo4WOu/qh6bSYJt5Hf5x9vBS0u5HigJICpv/3h/GCBNiMwKBH73felUht0GfZJvZ
3DPzK7ThV5nlu2ZYpDyBgnGT2D+vHywcHlpySv8dqNfya4N/TzQCuebvICwUU9ij0owBbOzusIwe
vQ7t1JWZS09XUhEAotp0CbiqDldSgbAnsDz+FaX1egpkoDh7Y+f6+P7W/jQ2A25wGPFYsBMo5iMW
Qw9g/skBhH3SKnyH36UE6yTgS1d6TLpNEle3eldFw7SuOAQFt6Y18gKgc+TxKbXMn4Dg+hSggg/j
LTivKSEwBSzaxJQ6YetpRaakd7uAt69caIe4gUIiis9iqU/8i/98CIQIeRXqIz5xjYq72q/kor+W
n8Mty6rgLz68iEwQoV2FFtHO1+cEn7p3OvERDHeY9kOcsY6GqH3XVUj/uzRp+B/i/G/9jSzyudgo
I+TAkDi6PLTQH5Z0ZjRJnEho0PHoab+UWUrbB7hAsczi+UmZk9KJd07tzYnXV1OInLstW+F1GOiW
OUoelVzlKwTEE1VUQaB/nW9kiQCqi6/UyHWRmKF9HcOr98vw2dkR04gGHvkAQIGiIjdiprvy+qGR
N/TpCXVv65YQpqujoOobliblfwPxZvTwFf9ub6sRSy4vj3TpaQ17k2THpq3NAirEOVPYnyDjkMQV
cEE/AqdbvTiY7BhXvEuv9yqw0b73OpurGyUTXpS237wzLokVqy5IvbpjqAMpT4mq/Gd7FCm5X0Pe
ZWiaxA97BSpWxHxkW/Egox6lyxGdHDrpOV6AY4+ZKOTX2xxiLK6tUXg7hquUdsoeXDJ9r1U2RJSh
CtpRl4M7A1nO3bdfRSXPfhLyUUlJQcUolOcP0BSSv2OSRry1jnhaJ96WpJAYU1iyuddLDrZ6mTDM
JhFC8FL+1XUtmBW0uiWFYG34lPT1uSnigYsAvrYntLj26jQoAjy6TDVJYA7RNw0MVMUM72dHK8Vq
HzlV2XKqbwS+OqwMXNYuFM57DPwf+TFu7e3/USdXhwqD4gAWh3+ugkOLskBm1yYAFtL/1zeZBLnp
wE+BQHvR3QQKoCyd1cv5Uyr3BPu+Ac6tZkd3AiuYDakuBPEKovQJvjLGBpiMaKSPyHGEbMopgvhU
fbX/pNp1E0/OhbxDnx9jJiLwe5fRmR3fYW1EbY9bnPrWQPoeMd306Sk/ASE9S4eqI2JUgQ1hDVhj
SL5WJOdoQVVMdoOB/rDDn7pZEgzFbxwgTgMIzFlbrDY4UW66ldQzFO3pl1w72EkxTV3xlaFIDYit
0Q1OWtukjfaAd46eTKBdUa2TjiB/rX6g0kiVg+43P6zssF+hTKw2NbSKQV7jihjF2+MFAW8BLX/B
sMCxr4urzuDOGdHL/0yASSqF4XwAj9x3phIPPwUzhGxtQzzgVawxgaiUre4AyeyfvUCuxmhPdyRG
Krnk0fKI9B4g5HtLDVJONIoWs58+MMPLwlxCNgwqTO+Npbg4fyh7NWJ7AJ6QX7XE8ywxIJZIJjCi
maXJR8sW4kbtNiLvF8yOW+IUHetu2JZKTuai2wTSrQ/iEyFaJE5K8MktceE+Lt9o5QrkCgUJrZ13
foV0FfSP61c4trKFZqWh7IPO+CqLiZxObg2nDP8EHH5uUA+LvbooxPWFYlzkb1Zp7JdFcn6yhun3
8qn8JQrQ3/4zKdz3U66VDtLK8lq4it4aYLEKyz8QYOW0aMniHY6uM+QBYh7gwoD6D5I93hpCxTAI
FlDhn1mvZZZzZWlVIumPH5nKQtKPle2KO9+4pyZZo/zriy8bhEYXyPEGlt8sjJoq+/bfuiT+YK9o
PFZz077Ue2BfKNjdAIBAwsEHwroJJX7TIQDKhf4HyLH5xcXrxu60XYuUsHxg1xGED5g0SvFGAMuy
tAOKXcWrbpeIgiSNRMTvNjd6XbdK9fcCM3ERr9nzGQ7OQlrjG0AigqNyvclfUrkYmAvPa1wbvlNF
v6nXpm4sevZ8pMhKh3SP7U+sm9LJkwA9JyHithj2HfdruddUQxGlsiI7HCmvPZxTX72WaNzgLs4N
76jbZp7WtnyAodI/lkHoCK2dQrZDHi2bauzG5vXVLybJsYpmMomN3JYO44SMcaCaLOIPRwAskDOg
GhTe0yz7+q68kcvl0dmRGDpkYmz5gTO+lgN+TCy09q46jPgiht0DyhLHiGIhWpDJWc1Uz9BMX6hY
x8hWvhyZnGolffS9RhsprtMLrrEegODrd6FIAFIXn9CB2x2GzqpzTDB2/ysH2i8PatpKODBioBtb
0DjPkwUAeM9nkupFvw1qWnWRuC7OMxfWIA2XNUrkXsrfHqT7gXkxIPN7Q/3vhkJPNYzcTaD7A5JZ
aGt7YAUgtMu1t4RkwOYczn7D/uoof+UphSJDJiDi+0rGjHt/OT+cWZCJtERCEJsFSn2gv1aN+iQj
ihGBd1mhDyD8EPCmJYIGDerLd7g8oGXetBT88Krs7LjAQ+f2mntDdqUxuTuMRr7HCESbaZSXPdH3
+7JrZilxHZzGhOPXyPvs1eI2iqGr2V2YOhzJoUEhnVIqIN59WVOhJa1kqDmq5DcBoxsAr8/QQzgd
4xHEGPtt8JnI87lgazq4XAkaxnRGj1WdO/eNNgaccad+wyt2kI9PrsKY7CvBJrdWKG2TGwCPOCOl
0G+6f8Y9bzsTmH9+vMpvL258ihkqG9EZOOPXHjnbRW/5t9iC9iWUBiLPjOT14xTSbar6LHtXGVcf
FcHM6gTtd0kIU0phOKp2C4vc0pJ/1zQK5L5IY3SjhJcUxDV8Ahlz/EJHoEHtCa7cDbRllJV1lZ2G
gSVImfbyxrd4IGXWA79chH52e19eqHitfSEy8qTlUSEFWqsXwMYQPaOc3yjT8tv07gaGhoG+TpV8
BqWZocN3NZdpRX1AHquOoNpDwb87ss7LohRZ7mlnCwZ577IKMEAJPE09AYSJ8AT4+CtJhIb5IFXC
ilFbMAkX593Poipx1iXZJPSNASBBH7ohZWfDJV09i/ztBS9vZ4GZCrzjEkPzNTbtjt5w2N1QYU3e
Q4SQyKFS2oK647bTnsI8Je9lK9JOqdCJ7wXASoFqanQ+UzA/Afm0x0FrgvOHdnbrnoVANHttjk1V
QyKHwEFGmGBqfmYG+3iZR12t5erxMlgjewkFSUYRRQGwReFuQPGdHKxX8MAXAINL2FYI/VaJ6Kjk
agYF/DEBRV7DIftu/SwkjM7qG8cSWOXtE8j0rhh7IuY6KISy96ag89T9zHeHby3OAPEwonJVJ73k
fsccXLZAm75QpIBinKgvprxMkN2D2qPo8yvyV1VenkmIO/9wLcKsvkrvZAN5PfpyyXE9cLVHFx2E
hWC3qoddn05KkrAC1AwfccnC+AeEoGWGRcIPbeXOyU0fYBLj/u6UuLffoIEWEO17tyNOrfLNEGPa
b9WB5h0bnVrCi8JFveNAzWzIu3WP/zg59TCYSdQ77IlPHovWML3ZpBiqToyI3NIY0b4C81aAp/Pd
Tvp2Sw9RhUwUH+DXQT4f7Kpm28EZQPd7j9mI0NCB1TPYEmso0KEdPYU+k0mUTB8nxEooPjiUDUgK
aHd2bFIOZnuJDtgGcwfEd0PN44geGrffeqhc0gSZtjYEY+8bDnGNXH/T5EYI4I0R7WoxP/rjRVTH
+mBLRqD89OEWXAAGI4eJsn559TcDoybCzsRVccJjudPHOJi3sXiphinDsrbH4Qpvy68Z+ROZnrdr
mkmgcp7qbzoy67Mfmp4e2089cjx98bKGs0+zVktAL+8N54g7VejQqyoxt+NRmGm9wLV59fmgzv1V
YFQAYbzJBVP/jxifEOAtXYzrRPlZ/A6uZv8Pz7mBL9UiFFE+c3nj5bU/6+Ii0GJ9BFhsmZ4IRrZM
nHV2mWstW0TGMHWBmpFXgGDGszkSRSgD+IL1Ajp7tnTT0Pj9wB0FVGYjNlpYAxeHhlKywScbSTZ3
q+s912dvTPNVyKqGEOgOIESNP64bszROpxqVVo6gtrWrVxt1YOo5ILT+Uwk0tAC8Jy/YQN+uV8aq
rHCIC0GrR9hYAbL4Ry6N4Pt/BDKnWsz9JQvFVx10FuooyWdhTrNPVxQcoHbsU2RwRd7A/ypavXs1
/WfsxcmH+v4txgy87QbY37hKfcalVvnI0lZh/9anKRoRKg5NZrbl+pRhRoMqRQxBr2sY2+mTVbhW
NKF+HQhXA8+s8EpbgI8gNJkV0kF726Hxiz063pYsL4B2NwBv3oQ+1+FxKpjGXuXqsJed1HO/YA+n
GoWICS/E5b1lmV+GxmG8PS1hvf4yuHcE1pJ7T24PsyEHSjMARVTqrOTQbgZ+WMJkjEGPv/sPTJzr
rXLrxw3+og4fhezBzg3+zcaUaSlPFNpfuYDh4WMKFxtJgo9zXYaftEL3YhFiEoOtqtLVXhsBhBUg
HFCJrwnXGOLC8Ud1oCMmIPUYuWU2MBT/Ms+RLF0yWy0A7HAVseCKiAlcX/zlVw2mJa3u2jV9d64v
NxaqAb/Nwn9jiwI+QpblzkUAxK/YEhoTKGQ7bbD6U4+P/08N7X76ltBjeaTAHVGorAtnVytE35QH
3YkPMBHbjO5J+bM8/wmO+A+qGmCuNX4vYLb4g0wazDiZIePv3LU3FbTfXO8b7RRgZuiusHv6EOc0
aytCegTYWqB7YbtWN3O7rWlOmVddLQNqfTUG/Aidn8o2X53TbweaHd1I41ru/PiVDwse4D4352zj
tBejhC/cohnQLxa3Hptn4NFsrQktmcFpZM1+4D6yeFk/YntoBIu3uU9lmEIAajHUjDdihKifYUgX
dWc21OR1djxil97LCfyRt/QausP3S1E/McGMSuT5qzuB7UwUeE6PXlJGEG7uaso0dERcMNPQRAFw
DY6+vC4faUtirArl/XPWI07iuoE2T3UDYQRF/AevZSZ53PzYNYE+S4bKEMJu9A1PfUnEEIlr9Y4/
3nrs51MGj7B+cf91AVt2Z2dOmvThEMXsCwpr/1mWiivnha3yvUfZiCDeD7JWn8WTrUWVJGbVeFj9
r+scQTu3hNbpbRdWiGvSmJ5oJxKWhtNsMQev2hTDKIqJCjoybLH7MvG8jH80mBgrNypZZ4Qpy0jf
HEl2+/+u8bTPvamYH1SIMd3m2RHxq1MjgggxH12pPDXj3q8Eq9T5C39ykycft1p4WVmnw5bk8q9l
9+tHD5xu1CZxhAu3BqpqqsXmoDlrJ5b0wdiDmlTUtr5CUfximlgwWWr0IALjU5wHnFF6GwQTkZPs
cBkqqpowoSjp2is7NUUteTJBaEtd9SHiqqZsfpg6kCElsSFgvW3eeBZYlmEUhQFatCAYbH76Pn1u
jwviujyfKKmh8H11cXUabNecbfPRfcv3V520P2TVczpkQNGFCG8QVRLoIEwzNIaJYam8Qymn7BYA
PTmpnQoTvFUAnO4nbnmaw2IjQwmg5fhmxVAe9s4nfcOYbNjbLnW+dT1cSFZDHuNkJ2gOIdLDOZ+x
HBY3rfzZjqhNOcZzJ+8KBuwTAT4xDuhvYH3MuyRCQiM07moqCPcSAwP4UTfZjggH5/2PhZYllTC1
YRSApwVqBoBfnuPQdMUWaq0PBWs8wrFqDmqTiCO9k2S0vMx+1+H3KyTpjQi7E0xhyUzb9/a/+5m1
e1bSKtbI4GnbMZ+9JK6wHpaTKy6Haieu6INwrrPaG9AtykJSoSwrBtHjHw1SrabMvq/TMbZAn6GA
JUgfU37GCZ5Y7q/IL6fJvlTNQLTmjGMgrnndKoR5CZ3lybdSZsTqNlgTVoqIcX2NsNTxYWXksaOF
LOtkDQnUHB/9rOtXmXeiHPOzTDwsjGcgTGTLaqVjHXEw4TEw5GaAEXy8CVDNom5HAa4vqkM8x9za
e5/PwEsZeJGELXKWIKhzQtqyaodGZJccOS+r/j1dheVIIVnFbaIUlMLv+5sssZVTZAykRAk/03AC
KzUg10vvyS/XIZZNG6Tw5G7PoiBldGfO5oF3Ltn8UU6rFQInsFEm6V7c4OaXeAWLsY4whftnPWRr
bnA5+wcDSMeIikLorLcO2orZNV3zwywD9XfK9SGPibilpJKRzdeiUeQIbWsLZoyvJ1BUIIn5z/tS
hb4yodYRouzb8Yi3WE3RwPZn37FuYi6cxGCTW0YQ4DEaGKu3UKjgmasI00N6woLDCOjttfDNBB6h
qN+3kiii9ukoGRTwgtE16B/sIydR/2THNEh4FjFTsuTNmXOK0olZVgtXRaj3RpYAl1AqjxMKxSWY
TkT8oJ50PTE7iL25aE9bs2DlIX2bFHCx7DC5OHFL4jWskrhyamyRXbIqRZwRV4vbE4FnQKj10179
dHn9kAtIrLReHPuMIuNVstuBW4nc3JvR4ZUzhbEpiorpppyK3cdbsSsxdanhMiGFsL+Q8SUQNibQ
cv0yFaZ5n+AroIGDxzF4nApOiNK1+mDAInZr5p8yfDGWTK98md6a8mlLygfrq4Jy70MxRZZLhhJu
TaDRDP1qhZihyFuQNQouqrCbC6Cs6SmEczeUA3xnx1+ZR8ED3931o++ycJuPo/S/5wsvfmM92uPW
2KNQoZdgC4JH4VjHH2yu6VQ857THdsIrqOKR9sXRfyRT/Tn2Hyw7LC5exJMjKsioQSZH3bNmsMoS
aNanlohNqfW3ghSf2FtboaHP9b1uZ04nalsbladBv9aWfm+3a0IF8OYI17/mZE+NI3wMi0xKchSd
Mhu1XJLTS2Et5J73ohiq8m9THoYA4TXK9i63FyCCDg==
`protect end_protected
