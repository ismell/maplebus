// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Mon Jan 20 10:30:28 2014

// synthesis message_off 10175

`timescale 1ns/1ns

module simple_fifo (
    reset,clock,enable,
    pktend);

    input reset;
    input clock;
    input enable;
    tri0 reset;
    tri0 enable;
    output pktend;
    reg pktend;
    reg reg_pktend;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter Idle=0,enabled=1,packet_end=2;

    initial
    begin
        reg_pktend <= 1'b0;
    end

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or enable or reg_pktend)
    begin
        if (reset) begin
            reg_fstate <= Idle;
            reg_pktend <= 1'b0;
            pktend <= 1'b0;
        end
        else begin
            reg_pktend <= 1'b0;
            pktend <= 1'b0;
            case (fstate)
                Idle: begin
                    if (enable)
                        reg_fstate <= enabled;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Idle;

                    reg_pktend <= 1'b0;
                end
                enabled: begin
                    if (~(enable))
                        reg_fstate <= packet_end;
                    else if (enable)
                        reg_fstate <= enabled;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= enabled;

                    reg_pktend <= 1'b0;
                end
                packet_end: begin
                    reg_fstate <= Idle;

                    reg_pktend <= 1'b1;
                end
                default: begin
                    reg_pktend <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
            pktend <= reg_pktend;
        end
    end
endmodule // simple_fifo
