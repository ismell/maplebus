`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j568ylTKCX1ijKCu3zCEYX4KzYIJPurwijBGL11yx0O4LKHLMP8dlqw1rKJAJyrIFXxSA8VDlDyI
zGGu45lCWA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Zsr0AQ+BVB+qiaA/LMGWEJP/NrZG3InNL+c379B92bObAE0efeTZpmUE1xBqjehQpvWUAwUx+nu1
ovOY8kEzNgIq2y7PBozDXLUFYCGPeG8YSvcca9nazpYZq3J1pYo73+j7dFLANXGQbyuVYrJ2fYen
tlUyhv+6QbaysUJuVbI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q2+tD8NGxa+F0Kpjcc7LfAe6tSHp2t/mfv+sRfVCSbFXzphOA7xbOWMnCZ2v11rkLOTfvtsY9E5x
egpSXJPwZm/DAmzKgDWCXDHkuVgfrpxeZMNdJ1lJ9SpDF+JD/u4nORV5Q5/DeeXs2+CQ5PqkdYUD
eIjqeKg1UKhzovo4tymm7vrVQtfKqVoXYUxWEXB6QJLlvWA5gOpbJ72hUPw6a0NzFAS3PM9gJRWr
+V/WEj/+m/HldnM/s5CLDxqiKGoTJeipBMDXuSfUTg9agdUBzwGsFCMZJSLJ4cYWQUG6tMY3AaLS
MOniFSWAyMTYTif8NQsspDwq92mtLcETXdUz5A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SIoa1SLEDIJ50U+1JCg5zLLYmPSw4kw2HFkGIoi2lK+mwV4W3mmmZAX326KwZQjzb9VWnIVFdT1Y
UN2hFjGyLs8z+rzG4Oy9dq7L+kkKeWNXb0jGjejfJbh8K9cxmEEPP8/IjSoJaNkIJlUxmJUnjyHE
IKC2aqKScbgxjZHZt9w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gJv7V3tQbfvvgMOdcWebzitR5f3OA0wOotRLu972K8EfTJsXxH0DQMQ8HCrhd5UEee7Tvs6urOmX
4T1c3Y4NjnMrZItgHfB/3LHHU5Q6lGh2xEHpVDRliN5nKb7uvF+tFsRpVx/0WaKIcOh2TmdQivVq
t7Ji9bC9MkBUU/jWx+WFIR5jbfz1A1FGH0+eF/NDwDLQv0VYxbu6W1vfB6JwqRtBcN5eqo0dIzII
v5V9w+gKht8MzTOKz4lC6isojTNbPRTIZ0z3i4bXGr5CP+egRZFBb1Rbm/SC//k6cCxEnR69Yl/n
FEdtLDULJEcs2RJeCMPyEljAhW84R0RsF922+Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18992)
`protect data_block
/LNCLDd+E99C0N+ZFjqerZrTN+mszLOGsn/YrrBpQr6iRSq+1TLQvIQ8I4MZW1kgjHbadFbYMUF2
JCnrQPJiRYvo8p8NXXPT4Vp1LuYBIFW4RIix1BE8qyHOpM2WFmpllO+gPiKBR44j9JrKIQtHpxfw
fKyQgXME4A17iniX0DSV60of7y3KoBO9CpjKxQ/FskJ6889lnkqbFTZJJZ0byVKaCg3pHXwYGMXr
7ufZAektkunU/L4x6RxQe98FfLcrVyJ8aHJYGz0n9jA3WTwka3Qf0BrCmHG0XZlovnpFyRxcN/Nk
7/ZBcfM562p/YUVLMO9vShQKOqPFwtsMEHamLH0uAE9xdcDyn9WGkglFL1a1ZIxnH0gB+Zizn2p4
Y+AkijoA4Mdb2Hm9f7QNJ3BLoAbLeOBp+K8EANooolruIK6+guYufSdRa1hmPg25EGj0bt+SbO6T
IJMEDd1DIMTZHWOecG81JeHlXreXW5ZNJOaVln3zd+iV9qYtrazR/SIQK5hkDtTx3WnqQBChRgxf
IQKR8WtCBtRI0XxZmGfr9O3Ndh89SKf1JZ6S9iCjQpNJTYX/Wc1CYORLXghy18HBAFZWOfpukBVQ
xZa8aCwo0NFOyDnuYfvjOv80T8jtPGbAeh3B5trBx7+5lCsGAH7UJaUpUg9PAns4/cjwwl3l97eV
EnjtdfOaZmlEwx32+/DoDWePmva7cxjQfZfSgKayXyUgUdHVdg95QMTEYeTdX12+lm15V4felJdG
LiLIYeb5CB70gSKEMqdzivjhJ5QTUY3FxvYFfLeNcyoFEFzr/MkG1Tj9M+CLXIEO0oWXy5SXppaB
lhWFk9sG1Ov2h5ACwlq32ArorMOqggi89tPLpjWJ2CAmHe/pzcWlBLx64qa20PYLlob8b2yjA2R9
Q+wMD3T6E4Sp5x2FguHHMn+15r+CKzBe/3K+bFxV4jrWS1Cp2DCdhE7VmABhc89kHcLWOYzN+M+p
CLmffa5VcMVRnLrlKxC67vEsH4frCs54o9iLXIiJoE9nX0wHRqUebdr9OllumaRKAPogVHmKa/om
BJKHvqm3di/wLSSlVNPKXFYEQeZl6OB75KYVzgqDQb993MhtI3OETWXaliWirm6msTnir7AYKudR
kiNXeVfgZ8dTm8272M03pxlQN0FJloCfMyTY7PPcMYMbRv5u6CohBMiyJG6ftzErf17ec9N5uR8I
4YUgAAVIMk5fusub4DQvvEtnTMwOpWZMlVsz5cH9yWrl8vClw+1+wfh++TD5mW5XzzAkZ+Efa9IY
u+QGMB1uq4vakiCw40s9lvmBJ2zrgQUIZMit+2oVLRGVJbIDqOIwwgrZToSWeFe1w6ol6XN82Zcs
Z7mdncv2Tsa6fziP3q4eLV0y0IaOOFnhCOTvGhmBGA0NPDXiyyZJtfp1Rnl6wTq2Eeow4Y97NMU5
suzYN9wYUN/Kk6Z8tkYEHfhzuGT7my1184/xGbgPP2YPAcGcQtfy0wmbnLhzNBVBI+f9CK3j0/X1
0+PpWGEDQ9K3PSm6OSweTdtnPJ3+iJEIrQ14uGFgMpKOHFfd60gn8zDVXhh1Kl7I5RMLbM71tOEr
ZtTkkJVwv9lPGmqdCTDFtvgPn51N9MMjCWRN5ynm/gO327/Uy565n5UfyhAn2tPL7y86CKmlBhpu
FScvlkfloqsNWwjPRa1ivK+MomRfoCgpbD46wwgFWOQ08rSH9qwjXYCHcx6k91SHgCUNVeaPlmA8
GeAVOuXT2pJbOgrEgtozlv6CfwjaZKI/AByWc6FENzHwn8EY+KPGW1GEwLcRhQdeB6j6zTAiAtXn
6MaXHHB3+FmNQHTp2kGIaZeJNQkhdZiF8UOKYo/ncAUcYCAiUWW78HZXc+sM7ko95WIcx9NGVmvG
hnpe1Ou7H5Z26HOzB8GTHzz1L9NgWHv3AXeFWHq1plMuzFVfiBrM1ZfkbdfRXi5KZGWImSBCTF3x
xVgqV12sHtm4I1YxZEecdyY4yQ3BteY7F0f0JNkVB2mAC3NewL4GB2ds3IDiJfj3/xHKJ0ACTpkM
ybfnce/D0Sp+ZjranGJK3Tx3yqcsjOUnQUoRittSwlhC6KR6iAR0blwJyuOgHlfbpJrfFFLgboyA
o7OGoeOst1bydW7SkKsNO9izpzN6YPotwSQjdYxPTPTbJ87c9AyR4S5y7MuzhtBiPyfDJ77N0Xp0
5DmW/MckLr2W9Raey3W425U4K1CY8ivBPLkyJi0Tl+R/3a+/Di2/kov+R7tsZbFv2tf0utcsdJFF
Ku3jpWOJEMNCnEzkv01kjygnYUuC1nXk2VA+pb7pO4noR675CGgFnBkeBFPZli8qbDoioTgEBCSt
GreFWtvkFrjGjgeFi4eIXvCtZejL7Zkhj39viGU9kaQugKSfJKlg4EsD5+GXhBqBIOsDynQWI+Ay
uyle1SnU3VaCJce8ueai2QM5r5BYXPq1OEyR9wkIRVzrITfy868rXnTQd1fkjpsPD6q/XT1CSvI9
jAttxENK6UX27A4xzgr7bno7YomKHlRlcDBYxoBNvkcqZHSIofCg8o4P+8dbsHzK7oxI2BZVLeKH
TKotd5CI0qsfBjmFqWpqrS6wCUriMweaOofPy5YBD//IN/eT5mNl9+skHVwraSVcjX2fxccxLa8G
57OaGYVK321L6LsrM8tSm00FHLUJdH87e4qfkugSQBgim2XwliiXTFro8x3a+cj5evSHbxL0foEV
ogku8OXJRG7z4PfFu6RZf4NuNMs+b2puxEJUpur6AZ1AvCrdbS4WjBKlfcgaDEHpIHAeugIFGOuj
DulnzYpBg2nka2hquBLHd+NBVbTLZIkgDbNxJPPQPAL4Q4c8du3bofqJCcY/5UIrG6XwWJgrOzYa
XRQsQfaH10r++Zbhkq0kExPVm8YKHzQLirmJyFIq8mR2Mcp7ctckc6jnF1eMIA2u1ePNEUyOJ34U
G5KIrlpcj5it2T1cxrnPYKrF537eYGJcwgBoPZVR7pFX0qSni2u9W0kxjsErqUMpepK/SWjLikh/
NVjFb6eU8rlYnOqlSb6yOkZzg1xHlPL2JlGbaXOcWNmNpQFeAyyjzTThB6+fCsz5e3y+FKtvVDHT
ybODXplSOhIofGf1ZGdNhPPbgUM8iGum+2AbgxZ/TDj8RuPUOKAWp2O5L7cdozqOX0jXvxYpuWNr
utt+9C3SZyFNzbtrOl5bZTuO5J/yIFPYjeNkNfYVb1RadB0wKfRiRX6mqGSwXC4h2uNHOi4jStWf
FToq3381RtVpIoZ5Ex8YU4/u/6yVSKGrueoKCQBtMFBCsdQ0NxsZ+16aYjpKjkIkld+GgsRUtJRu
cDg2QI0jayFbMVYxzXFO47/sZrC/3dKQ63EJ3yPFDGnJF5CEF1041794U+1ioki2mqjHLBr7v+0c
iYjjoOC/XsaPX6v+6/x+A8kkN6gc9TQI4LLz2f9oP3B+82TrmfSwqMc4dT2EbUWBT1unUI9O32WN
RM5YjNuawt9z5d2l7MpJqEF6d6JUF7d3rw8Yol8YyN833MNaHVztCjq4fdBqA1VDJjZsLFWCCOmr
A+ST3fjn9djOVSBTNGMMAjRthKw1errBiAbyHalFkJXaLGb2SxkRiO4boM2AiYIgcaCxttmp+0fU
jxsXTn7NP6uNE8GwT786ikYAZbqYMzdnRnrr6oM8WZ62tQQ/lo7yrMtGw9rLHrkiRoRIR+/F8fFr
DBauCYPf8PCXGOZKuvR7dPHvEAdOEsYaPgz0wMB1ypEGgCq4sm3b9PTsGtO2yFTqWaNHSf+kdiGn
M6ApLg/xO4svgCwF+rFAD9JMLIugpkpY5dqvCfv7eHkky4k5LspCYq6FdwcQkM4SCx3ZJfejZAHc
8optjKeYyE467t8dX6MxCX30iOLe4BJRKEsAsbIgS0RLjTFEwowahLKHpsSOpANY3BNizKDDHFUH
otjnb8A7LjErX5ECBrDtYfwQ0CKYiHY1V62a5iP+brnNy7pH0LnIZ10kDbD1VthbE3LBZXYM25+E
ulYqZ7b1Ou/wnpyiyIxitWu8qNFEmfk+7HO5hSCStexNvv/65qFomybelCVis27hikfToy0zqSM+
BpIJGf1gVk/PIiPTvKedXpn6xZUc9ZqsJoORxX9r25DKG+addeXf7pm8RLxZApq7+dCeUT3dgRbK
Uz3/9eXgY2qOqlhOagRfsOQMkbF/etntpONeCVCLeVYJgFXMPZgCDxtle4OBU5SM/9AUc+dTQNys
3Wfjiqd7rSApiMVlYDjVqMRG3fdoVG4YwpOD5DvtW/pwQOVRESwUjIVwj4Lw6hpqh3dwnwCOfDbH
ezlLJVspXPA3X1E8F7zuBA6fpCizKwTXN8dlfPFTIvkhArG2GC5e284lUHVXvhQ7tLoGFCQKEA0Z
3ig+zX+6uYjMmtL/7j29PKUSSGQ5KU/lamyNpJzia2ShzkNpe05LoruCnePOlwYDsrF4nZYsly59
W7KP5YH/wmR2TVwuHQQqMZfml8nKJFbc4MHU0Yl8IYztFLRxvidPOdvvVA8F3hdHmuoBsxPJoTFj
inSAUuC50xGgPvW3CSOfv7leRoFEylIsHYlxawqNEcRxpz4QwJ2Kvdg+SWPmbkIHyrvlFEriha6i
/QaoNaUDsds/tHu9RZwM3KAAd/EoIr4o65QaV/0/gha0BL7ToIJjfgjZlh46BZPFZjJ7pKanrI7s
uUUmoMNQD7ZtajeW37C8qMBaswRRyflIdg6TrOvtNuwnQGFpLk49VkmeSR2zUr9jcCCFbaGqe02C
YT0pwWxFezXeHhPzIjDc9dZQmNQMWUEgsyw1aN+emnyRHiFOz4FHiRVBoekFoklvMh4492avhmm/
aY+gNA7nBBqDgiriI/wPUJeo5Xi13skqO9hVmPfp7eSipIxtefMbSicg7C1Ink6y8A37f21JEdxg
3lq+Kfx+tiNadQoIgfnDVRVhWilAo5FBtvlAkUP6l5WXs6LQVZbpBlNszgHmV+8vbAOlhgv40p0r
/NEKBMcoNHDachPWWC0syzLh3GzPCceNjsy1EHFd5bm7sVwUDjJOKNrIKD/NjF0skrUHfY1bTyoy
bWTCiZpTIQhzbAVrU2hNOuTKP/+toKtmoiOaHqHUIgJHZaFk3s4voW19LSUzbZeQQgFvchnTj81z
9WG2h8QTJlyDekl4eNiTD7DRTbuEataCOsVW73TtbK6lWbj/GtYSeb/Rv1d4aasK0GtwC+ImRNZt
j6HC5gZ3V9Dya4hvpunlS5y/m7N5RdWaEpb/a8PBWhHEvVlCSNYHOK/VEXl8+31DjO63syqVfJl9
mhse7+NDrgn+zG80cxAbziR+AXXjKEg/G1J5Fu6pheQH/NtBNVRdTqXwPLQqZmt87pBLFtn9zfQO
JiMybM10PisT5nf6OhTD91tuALR91m5JbWzXAzDH/B43lSR5Tl9CoLApp6WHuzZyUasyr7Ux/jDu
ykbeaYvXYW9OPlx0XRSiRj9vPsd/v2pBTEezb9IM4mn+JhQDc5xFDpjQwbuHWxS2RbG9qpsswYbE
Bn+YVbffZ8OiXIVEMtBRANfvLYDbBsEqGt3aETYARBcTLfAQRoi+YSoUYAxP0ZDTHUqd1YtUcZlX
/wBdn2E1Q8WsU7FiXfkyuYK/kb2nNniWT/7FPiqhEEM2GhwVy9GpvfU0JXtaSO/q98X2DgB0OH1B
PeqD76oj+o4LBvgzVDcOdSExYyzQydUPHxVPg6CXW4chrAxKgVozFilsdaH0TUDx9C9ZwFUApeox
tN9u+T2/O+WfCYQvf75WsQ9PbigFnEcFzSUG85Dvxu3inNh5uPDxQEpwbTbT+cFTpdBRfpXoU4g6
9/maMo5UAwV8PkRge6UP/8i92+fYaXMYaTX7e1xmmzaKE/qSLbXaKydrpUPXOvIxpbKax3X5kTo0
1YoAAxJgPK5950FCNn0hT4hzRK5ODe1lGmPAtwA7fwcI8DxNZ/qS+IHGcCrdNXtH6dD8nVRdKFEb
EXtNVBYmJRI4SN4RQ15ZEqUDdra3QtpSFqTNtvlXLNS0We6QP8ZIvnpJEABe5v5Zrk21D3sm39zU
zBDu1dQbKSWuTOkGJSDP0MExq3/Bk28LSd4eV2Zp5+I9MI1IVDXq3rVgN70HMyUS1oY31h6x8F4e
GZgELoyJzJCTHe9PFCye2v3x2XUXeBpC2odZ9BI1aLqiyOl4izR1+xZjcXt52dAYX+UH4M74ppYS
rFC0pEK2rSGoO6v3BSC+8C1oLONvMLJHqYI9zBjOLUJuK5Mcek1MHcVJMDB0pyyfmNJ1eGMNiFLD
JcLA3z3P85CsdOUSlcUfUrHConuc0OyNIytH/yXpJQYXip9aXSv1sxybXAK4GjoSEc+WeVIuwiFt
7pvzSOQNpFzfhHBOjHA6XhRNILAVFj/F1+hpibVPD/LhcRTUAEIxTF2JHPyf2A7MPZcTaxWDay57
JKL70xGmy6KSRki0pOq5nwrYRnT3uyig76s+nNU9AlV/1UZzY9eFYw10Md89WWaaYPB4GVM9ur0K
GyhYC6amYB52v18TNRPXGIseUCu4ipekMcrBJXcNbz+m+QhDyTns7yGPn8RBHOFpgQvoRzwTsl0w
oVMW1ADcNC/pE9NMwQW+i3mvaTgrKd2au5tZD9eAFKdcCoD+ATWOcMxKGDCHMkxfXlMV0EXvStY3
7JlACcYquax0vZTqBndyXMQ/ItrAmMpnUcH4v6xPt+giCbvx8VdMDtum8JtX9B+0TU6RvKwOxFwM
I7w43vFC0tmr66mfksoSEOS+YINatrRf5oUAxF7ikyNDFZIUSUt0U3+tzbgHVQF/De1o7S/kN5PN
HvKqrzCoTrVERbUUDO0ugCeW7QGgl6o15UNhpIaBbYtq6EREYShk+XiCTW6gvMbB0vX88p+4RwlB
IznTW4MTN9OAmGkTBeMaws/ngnwiqISm2ubfslMYDteWLYr6HEBilZJmamT7oPh4qcb4irxxjVEJ
pjIWjBcNVF0tRoc2/oYMIUMqOmhiMa9TgzLt1rCmB2KDD86xnbZPLikcq6uzlUH/1p47Hbog5KbV
Vd2HYCT3Y6keWvbGSwcDrDNk0s1rKSYS4L7Ikaq+r3d1zhaw36I8bhKnSawz6eqVakyYebQTTHu8
ptYplLfxRjyz6ao1bN0qUmRUWEDmElpVMTSzJft0V3+2y4gtXPwvGocB0616ol06fabUIvVHHaQj
cRy8f6vgPlidgncB4m3pSqHEH4ZMsAIrbBsxq6ndqgGtqxnxosekyJHQqpLx+pdrWKDUkKMj/VO3
ljj+l6f6DxqBwhLHXdnS/SESrIHyZZLI3d4b+Snmn3fwca0KM1/BLF532mYmHCOHo+sjG4cJVmS2
jhpIDHW70Rvx1HIGH17WNJB/iPX2l981vbTAoU+JJ0zXjngBu9x3sUlrCf/qD6YlYXMoouEuz9Od
rYAp2aFlIudAVwQnhfKPHZSs7mi4RBawuDdPNhFLv5kIl+bSoBvRRy614BHvcUxBHBDY/UZjjAJW
UrHP4of+WLIMknJ5L8wT/Ny53169SthQKVZ45cUA6BziPJUfDW+iyeeLDe2MCvHTK93X7t2MuWv7
5o+tAD02Rx0gwqzJMNGrHQtzXfVRNwzspbjPQdBX5OHcu/ugc2NGJFwC4fea4fqd8tGDFwH/6DBY
27KN7kOEASPi6+tWtx/ZkGD/ue/f9h7sX4zk3y/dkaESUmY2qLaSU34HpI7vsM0h8DRPpZLSCSTz
aocJ1YGzMRP+ArPbIgWknW06D/ZIJbOF8+N4JUY9OULIJz3SAxu6hqOJFH8YR1kgTTQ72PlfFJvl
cV3Mp/Xs2jotbtEdmwbPHgONYNJFX7I9dIqYASieBhRORdmTWkV5Kyvu8Qc7ViVAcRMGfostq5m7
eHZ9nI/JcAzL8Pcy1XSTBjqOVHaZNp8AnGOIBg0HumvriGO/HfSbL4qoEkSvIOy/xalrA17Wei4u
2QwwxTrMfa3OMyGfa28bX5wSxgTJT3wRau3tOah+bIFZ84WMD3863a29VfhltbCdk0zXSd02oM9n
1bqt++SIgqFIJRQ7IMoeQK8RG32b+AooPPq5396As3dcTrnLE3T7faUFdsETY7A0AXnK9SdeaSZQ
wGwj70xKUvLpfWG0DKVIDKE8LDB5oFQ9ZytZ8ANMfq+I4hMbeDr5cG4AotqiKsVIRlLsrpSCBlDO
RNLBjYiopZhQ8sC9HNUM3BiF61soa2vZPeYxv4qfLUORUUfQs5mYa6P09mfRXQzlS0uZ824/bYw4
pAgrhnVI/kmZtcsmOKPJ8bFArsfvTWDvgeks/1O/EqGWgxaHS/llh47YlI8hNTo0a5OG9li+WVZf
pUOvEOPRxrW2FdeG16+SIPfh5tBjcQFzA6ht0cuor7g9wOX/HqFiyJzx7TOotoGqTlaZn+9kQAvv
yvrHUrVUQ/suB/aCT1CsWaRJGMGNASA0oVY/vlc/240o9r7Wx9tRlJhiVyFsH03Fsc4uMOoq3ecc
Zzsio0iHH7iv2+F4luX9+rwO7G5sx8S9Q9wjaxBsRh0GEyUtMZhjG/Gj4CWzfzQDgdkg3sDMH6Ta
8ik7+pBwctIwSUWHpuw8MNRBRr0Jqv6ZgVGo3Xqs2orFXcmF7WPeo+XqlwwIjBlFEJhFgRlyUEQw
+wyYNCJAGx2CEsvEgSgZK3j+2zB4vm+TLxbtciHToQvjIgh/j7/YwdtzPUfBNCyzJLiI667SHzb6
Xu1FnJvUZkxh/UXc7GDa2ivLino/hdRl/DQewUQAo6awWVNS4eFICSZXHsGSBl4chpv6RRNMFORL
M+1/IrZHobg1XhvxgeD3Z02Z88QyTaLx1MtKu+JM0SwTvAgHZm0KLw3qxAvE0HcZdO72VzvhPP89
rjXZCjeg5BIe39d/BWuG6zL1rimaeyKLVS+7d0HqGwvwkS+1eV4DsSsZzjpmeiViV/FeJ2K0liuC
fcdCRQXwGdOFnkRvUUIG+Rtr+3/jtC1FdBVsZi5W7iIQYIHQO+bIzHcH53bvLGMykHLvsRckKjeZ
S4Yb+/kqydvqBy09VPa1N1IdjC7UjavR77feVfkbdzxfQm98xQajVuMvdIaxQOBxAzQl6RtH0jYr
IDqHgCXAUaMf9b/Pv/BSfhf51HdGhynASvwYbhLz2VTOywLac4bCDgzavoPwTrvxM/QanSwgEkP4
F6EL5mR7IrVMvgRKHgZTJUKHku8U/OvoXYIlc71RT9bTWJniZbK2vv9QciDIzGep806ueThvZWPF
h/BOt7ozjZrq50gK5b54Uj3BDbbqSFOs0/uNUh7CQahsAgQvoRQyQ70Ipip0xzne7Ws9oYXaEEBM
AYV2qU5yPzphTTjOkNKTWB+9Qcmrw64yKYW+BoLL7nvJs8ptYUf4y6WJK8ZTvcIMfjX55+OFhIuH
j+RTpU2rsKEFI4CruvtFkBN6PymLtEFb9zJhx8/w9fNGXfrzu6QVuAEaMEnG0Ilz87cojo/D9qnf
yd0szHqx5Q7Yl/f3k+0vd07Vpq924wiAkM5U0NP+UQ3Xcud1lEZI5mVht0zT8NmQIsJ1qYha/iBj
vrM9+HuL/P7bti5DhEQkYD/8zJ+7UwjbaaMBlkJXhtyy0lrTESvqOyyFw5x3NVrsFZRZoBvWNYSq
COsojsQKhMXeJxFQ0UQTwL1JxCiQQkDFzCvTUj6YRqho/AWHMxqWRZNSNwqj3/S3voRFvOgaR0o5
a4KD43g1K3299LT99Pq9kccrLr4uln3kcddzwsb0oscWQ7KaUlHFZFG7FLqge1F4bG5+na/mprPU
A6NaAu1ppOvChZ9duuu7fmO+0h9WduumFcB296iTAh+KmzH3cKW+0YiFfcGGGIvb+ic5wY7Psgrk
WxRYeqTGYjjorNDWhBVvwTkbe28XEsRW0qbImxTJuwQVfcHYbAOp5+dUf0juanDVaLlG2bZwluos
pZVl0M61M/NIHwwbyJv5fsUuV7GKkUplBMnwQ7OiVyA4UJOpc8ElxvjPe9rrG+Dq461mfoE33aDQ
iskmtRDhfTOcLqkd8KyV0rFWCap8aM2tEWeiJOymRKoS2D8EtdIcTrgLQYeqraXBQfc04ssYnem2
bWqBwtWGw6cP/dVON64isCncmYOagmHzGNFWfqTUJ8qlz0S+m0OneEYF/M2GlErVXaLXEWzDDY6i
gNB/lk5jfhVnxfMrUfuTTe+9pM/j+f6xJMNWgDdTIlMxSPaO0+oGxcj978PJYqyvS8IfBixRx6y0
mjZbxO3V1+wEZuq0rjW3QmmLSB/4iQeIfOK9eKHsBDsUD+vgfuMC+b9unQWRYZ4NxY1NRkH3h08+
H0ScNg+js5xPQTGz37SYQMnP5J4O8BKb/zxZGAjw1mZ53G3gNRjuUJw9wyspoGL6xKTJXIkFsLxw
dz6+AUlv6uI+W+eQiMD1jdQlYbZE0pdImsjON/qd6txCeAJtYzdvR2klVDNt3xbPYKvZ4oVhCiyf
3/n3Tjd9tNEZaY79ShhXsHfwAe+LGUSRvV7+45MMT+RusBrszGVY9wn+MdAHKQTT9vYZT2I9LKfe
nlO3wTMJ2baCUJQ5kn/XyTN+bE6DUjq8q7gkw3xz/fjU8g/V+u+7OmTj8byb0uly8WQbW+QUb0ph
8puO+RTt3He+FRFon7ZKsKyNWEXZGITUZ5MSXwIStFMuMl6M0FpzSDszKbwA3gVA+RMKm00RfF66
N6jKAlrUnkraJtqrqr71SZSe63Mqp1qrgo4SRFQi4HnXZBs98Uugcw54oWsdwBq7mwCrPmmmRjdP
lPJGgdO+1ArVvKMRXXVM1rKxSY1d7L8iOWtGZ6XTeuw3WTAQtlwuauRl4LfMABuzqGae4VBe6C1z
Bz+NblfNbXIXgQLdnuWTBa4u3DTBbD50LAgdTykvyXSvfz3GJa4zTUNgUQ6LHTKbRnnyjr17JpIn
z6OxVR5klOwiBeJ/xnnEYAhgrcJx8q26FrEsjpFMO6CctHary+OLCVhjlJ1B34z4SdnbBHNsHIoK
4v4FUWXhcKUxUpaRcpiF6EA1CVvL7cGCIVz2ZsAqKSjQtR+iPXOB+kTDGb9llOg6vNgC4uvuwrrk
ou5WkyjS4H2Cu4+llZocRrPjqP1inx0Ifw8riCSeMsrAU8/sETXN9/SBav74wblpdrQsHAacF8Wd
JrzPrpWPXrHDSwHzNKLvWmCQUAOqENI13nth6yWkHWlSLmBeAn4EA5z+aOu69YOoRXCq356yRYDj
reiIVDeKOcWlHgDUkV1qWrwMfR4575YgskQgPhbOrP1rGTxB+cLb5zYl2WvMlAyTNU91chOv7lfO
GE/FajfQyWjaQ5DiNEBeELIDzeevC1KRma+tgNWDRsJnOKEq3R5wkDJy3Cv8CMZ3dgxckVK18Z9o
uPmXHxVaDUDZv7xBnlpSs18fGvvPLrUY401DfV7wiMm/GdKXTa6matCDmOJw5NhhlpQqDVEaprMg
qH5kbYEX6qMGAUW4a8HgNBAeL5ZX9hEY9hi4g85vYy6qpg8kE/KCLirAyFPydAav8e0sFZWuNBkj
jm8Z3Ez1GWKnxGdl6do5t/uOzBIKO3lJgnvhjJr6If5JvMMl5H/mskFl8NPH007w+pvqxvUflQK+
P4pCKMjO/9EmmQ4hoXVaffGZkEjcyPipINY+glkrYtXasrddJ27KToBi/4BRP6KcF6G9lensi28q
RYhErcbFOJGIaK+bnr5VeT51Bm5Xy13X5rF222V+oL3BRp6r0aQU//sMLo//rWZj0ELYo3RKx3p/
OxPvBjuPYVTWwZWKxMBFtR8ELDBTXSRIE0wSz0IWSXe2LhTDl5MMjESV5zI0gA9MwkbCliC2lkzV
ff9bsEXVED1zJpcD2lPos2At9cgiLyrfrYsXhYBpZkcKDTjvjBHE61r1u8mxW2qoxu0SuaSR5dX5
1yzM4OvYj73+OAybdK/UoZGwXw0PPkofwJVrV/U4ds12ZdnIUMbJkKcm7HC4PCpOySNVVe931feF
CWQ38GHsXPWM28vSqA+brOPPzdXiwrCZWVS710Z00JNGbVJ+9xWXIw5XjIi5VY2efaAFa4RbpIQe
Zm/v4RsRC+pGYNYPGu/Hm4UruGuC4mEQW5qN8H0PwYiNhABKfATxgze6cJG3RqM2dtRR87yWpWWv
lZK1g524B5SIvBUvkWc5IrXJ3s+MM1FWx9uSwiFU7YPkgYyLFYK8b+hTDs2MWjrg59EsHzcahAGt
QQ+1ZtoU35GpFw0YuOfLYRE3D4pWZ1RfXxzYGiJwFh7+jf5kIqEedSMp/hjtS1xo9arFsC9BTSsW
UEHcXsj8s7ZI2wUE09wZYtulTcLkSPDvHB+55r9L+eElontAOj2FXI2AWUxTnyPh5LBVcsiajAx5
OW+Sp1xi2baCSBrmMG2C+3FubI/NNT1zZESAN9MPvXyGJAPhR4G2j+TSTq8mRFbHcWelEj6k8nzk
ywvXInmos2SEfPlje/5xSAMtYQuAGVkf3ZTfxsnnB6V2K1froYjS6ov4OPtEIBombxlM3PnCEFKj
mCugJYHU26fR3DQFnc2hRleB1KqH1UIkXlcseLWEu3uIf+kX3EhpOSk6PMzZX7tVF2/210BlbGJp
5I3J2vGMuiydxqOlvXSzSE9QN1rx79HMaWduuOXdQHOf9dPunCUoEezfbbf+nQyBU/T1wT6IaEwB
mu2tQcLvySNITtWt+modRcXPzT1NVCidYp3/sy7g2GT2FIiACuYW43MyBpxZMzYAoSyJTbJm2TDC
BXsfc9xR35nJZIIeGUkeV1APPi9lVDkAXJQGOAhqxRTJyw+IXy86F3xVwu4RtzRUeq3R65ewfoT4
izK+guOQd3bHUCf0Y4bGEEkie6lM22mKZpFijVpZ3YVzv0cWvqAH3YzZhGVxmFxlstkwLHyuewo+
AFEMs9ZuYId3Q5JGmH6I/7P4N+rjrEN7s4jQnUEVgDbCJTUO48BohaAkhOPRSgoSqIK6kK7EdHSX
wS8zyRU4QghX60Na3khkMcJDiQPcKbNAlKfP9z05OM7/+y97qUV4Krsbg2Y2MtyL/M9tX0QrbTLT
WDw4HO8j3KvCcMgjzPPmPd5h8aCkmXKjA9ORvJ+cUA6jlPsSn+HbfqRKFY5KCzaZDCCI6K+lGY/Y
8Hh3WiWt6WmILE8t6AM+wMZpgolN0ixh0OzJYV+fVtjXEtRk+7lRvQ8WdgYG123q20QDWlPkcSFg
+Tx2LuQVFaFd11CbPWkxEJQ1skVNB2JsnnHEpwJAxDEzc1hPGaFpATGEa0dak/hES1Z9pEqaLmtc
+kwJ1L9t7Fq3YtATAk5XpDuZ0puxdqTz/j3MNnvVEhynQBOpusYnWkOEddiBR1l9s/GyPblgW/mm
KzeNz1QjwM6VRdOgdw3s0Sl0zcP+Lby++vkNqJOc9e2Oe3MdPR1IMo2RCMiSjslCw/H5TH770RzT
6f1xgpOn9Cg7FymT4ZUwRMGf25wh7e1wvFMtol6j2lsqyumkfrBwQoiUf1HOpy6IulufXlngNOjw
aJV0brbZ4cww48cNlab4HF0YFJqiomzN+dWODryOhuqdDo7Mi9LFH1twxwONMr0ctEUZvWg/ef1C
fYX+PxCgLqaup3NULsbwQCNsVCUqfGPSSm2DuU8E9sQhDuIKeistU+dP7nxUI/s0aGr+2rnbY5lw
7iJ79ZLv4poUIz1CnOMBHKwNLzpyAIsNmUqLimWVFpeLzRO6f/2cM6MMq1jTuTzFSIpix0GFnOgw
coY8amAfSw1XgyRZISB9lSAwH+SJdXkq7YMi3tgrLRt8Ml+ExL67Yt84lwaBszQgRzZUGF+RGXFO
P3HO4bmZgli26GsLbvuc44UObEjHX3PtYwu6YR0yZ8cC5+Yb0rsEln4kOdZVNA/SfTMttjMosd4q
ZVkUlO8kRqi+bkMAHOHhm5NgDVZHGnHNpk/9iRx1wHRGM2R+dWUIpGKxTa2eyTTZ1riduNibYNUj
gTSktKpJFwjSboVSZKiiAajD1EU2F7tLWpcEWOYlsup2nyCnPtV2x286oVgjTmsewZ53xWooTXi/
69jW0fF+Es6KEZBKB4hN18Rzp14xb3FWjL0ZbZWVMHNG8Umpi9EdVNn6S9KiWLfpwgyoTHCnIDOE
ud+HQpQUVDwoG7nSipfu4+pekRpsnwo6LNtFR6TKnrH6ITla1tcmNGiyNCajWBXk/R4iEraTCiX1
NI4OhaFzt9YDWMRAoaimhmj9SKgkIa6lkVCS2ggxULCEvi02SQI/n6TmIKHYz3phdbP04qrd772c
eI6TP17ZJPV4rOGrzGy1lApfm63LKcOHwycatxnmQ1J+rd2U9TmvnA94jdNMC1cBNAJrcWsNm6n7
AuaeflZ0YP3pg2+8jRIlhHpTgBKNCccSPJIO949by9Do/qvuS/LJnXgRP/8i6b5wXl9UOZmHUbo7
uWWoIQbuvs6a05rN+LW9OFJoFwtI6JZzKU2D3nrjJh5GqAiWbLdvg/WDCmb9C9VaD60z1zHOLrLx
+B+zRnH6jouaaXwcMalS6WRTl1xmNFZ8Zy7/8t3cJ+MHU37LNFybHvb3QX+bbkBR12+ncVu4Hc8d
RBVXmL6ca/GN0gwWNgNDmMPkb4H3t800nDdRWscaDbPkQ8vVVYO8Nb6VhYPMUOz1ygc7xTA8zsXA
MVP3kQk4WCtK5FehbUWpljPaaA44Vpq8X6w73MgtMHVdwf7GcV7eSSK4ZzuhgvDRvvn0pJ/1cXII
fUcIXDkXJanTfP5S3MrqszQdh4R+xw0yAT87UX4+NFrBqqz6IgjXQezs9hQDyAdObH2Ol2ID1cUN
zo9PE1Lnvyq2nkQwxe/cN0zVHXxGtVcavzn8k/SVjleDN6XRI10Svh/HBQM+gWrdQZKrTwKem/zm
5UnMuxZ2HgLzIVfFMVb/LNNsyUn8S/UrysZwIS84WFQ1nHWT5HKyMpR16PpHAAwpG0mt6nHbwLvt
TcsqEHe2gO6hglr5W9WnZFcR94HBvRUVRDzEytHbBJ6VuvoHxRVrCs9qYHGlF1hyOoxMUYU1jm/X
E+ylC7jfzf6Ys4yP6eO5LTQbBAWUZakk2RiDkLS2hN8ud99tt27Q2YiW8CytxAMXVzK5Z+T3Rw1O
RtYhq2tobX0m6C93N4eO1I84VfuVfQy9+TtUbgUODJ3YGmtwzfIEoNuEABc19UJHoOCIyNnC+yys
olGuI9XiCcgShvvQGszjkMXn5Iwk+2CbB0cC7iWGRd29fgX8ENAIrp9A0YyM7qh8+DXt//CZytc0
IUHiTZYnq6BiA3V0Lny9IvrMLRKO76oeO9l0nM3Ab9Qj9CRjE4st2FgRL4FnAmDJ4uJjZ46t7d/D
0AktFt5MWmfFg0ee6zGfnLY/J4mfqjVWPpbQ7qpCAzyDloKai3A5utsv9Tuc7y7xkOzny6nLrk3F
4jDdclXHZn473IehHtV6q+1FA07SySwO80GfmdTcOGBZi5DB0jDQW/I166pVVlAr3oIRI9hXIhOg
mxozx/gAXmX7rLvtLNubFtWeWxTjrUXnCbD6E+GmdqFzCmiqbxXfo8qb+ikJrZDWiOz7ygiED/i6
dviGIRaODrPZIFHmS/kfH5d8sZApv7hX0nbC/taGk55+FCZncde1izTIPtnxc46uSsZb06F8NVRj
09/ma8BaLwvYMNBIMsnuqhJ75Pja/jPeHwyOkV85yVpnBjOHr8lBNy2RncH2xOIp+VB9ey7SYeFs
HPHRsgbxH5WpJ3ZeLc9p443Mme/K38iIu2hfubG7pAh2ljEVAvoS1k3JyyhwvvZfDXiO/Qxc4a/W
diyxQ5sI1DQt3wlGerbIyYHQijf/bRZYBl2RQQh8ABQNtVlvYQ3pdFtIYptWxtnAOGneIYCDXo9b
Jhk65NAZGIXP/UT+UVHVQs0FfeHmzrf+IkRH/06Wvc3BNDfy5OunFqoGh2BSCfHxjqCak78eOn5A
R7iMHs4vtLEC2esMA7XatYKBaWjcVbmpUk90Kab3pZFhYdFjzhznM6cr77BvwbT2THfKdHWTDWX7
XZjxuQNyZxZC5bmeHgJp1XZS05J0w8P0UD4D7x6KF9Yb+t10kLM2OxJOYm49ab0tHUNzu7GnGQMa
UXZkc3JAO9CrUyo0oX0mB3kdk2dJ2txF0zd6+XBgaooXKQR00BHamdNruucplQsL8PAsZUB2Ches
yTjg2/2BP92B3WSD/v/Qg9D4HWDV76LsCuqXJJ4rXR0x1Fp5KcFEBozUrpBl/ZAEhgVRVLLWHbBw
Q0kIeNh017k0+eoEDMM6fFKdMemutdRorN99i5uf5VggvRJZZOYIYhWApWTn9+qi2OrMY9X2YT4K
f5c7a8+y5j2jl9qA65qqUUT/XcAGmY7ajPDA9sRbYxZClWEXsvUamU7CslTe8iYuaCo+4y8DM19P
VUZeQxC8w6Csl/dq3Hwm0lWhPKqi+CR1uvl6GmB5lZO7HGdma44TRqyRj6PTHEHg85GUcU5A/gsj
+1CKi+TFXqItFp4RVuG4+i8o7pRXf/Twbsxho7kPpZTVNiFOVaR6FxNW7/NmMBZN3VwVZNpaiISk
jJoWkn7XjAj2l7fDKy1X2iUyigY4XdG6Nj/JOtIC/LRCZ8kTC9hjarPYXkAcPpCbiqkMn0pb5S6x
YjJxA62xdV8LD+/NwYP2xht1kcE70rL0tw//lg0IFKnHbTTWFTDHVzHDQnTUEvWS9lg6XC1YTDd4
/aLwXtVX4beiRkqwFAknd56aua8OfKw4fAEeqxsxwF6aW0XezzgNRBxKVAa4QSKvOc2bsZgX3gG4
OdKxTcGnXq3A2Z0iVphb6CNr7aK8PL73oaMxGumecpQO/+uqCdIGq3uTHsqywD3BSI6h/GLPl8P1
P+pBuydt24Mwl7WOA9ZJreL14WSKNraXDy2G2s8I+A1V2zh7cIq24RMMAJfCSh6YzZrj3mT0HJwL
4te08PwNXz5Oalluhq2uutsGNP9Q6N0qm+D9aH+W4ejGqx0c821RiLCvr9KxAoT/quguPa7Qi+PS
dQQPIfnoCY0oMxg06wG6sh95UQ8Xjm/viiVSGd7ihvieCtjiHVhK+oFYzWXBYGN8cZ/XAEXb+2b2
gtp6LorZ1aHJWIJYE55f+45BQMkokRmi75ldRukfUymCd9l9RuJbFd1Zl7Pp3dCYS533uKTOSRKO
31eUiPq7h2raAzzEikbb2ECOJirhEvLTW5RwifAbPrRc9GXIGWmvMV19gzhWYqDHSPTBky0hiWEn
dZtrg+6SNcrXThD5/c4BhVjZwyvLgahIt2aKDFaJdrGbipUw948Cvuy7mutZy2MUdmN/Cmh8MGTa
x9ekLKSeP3JwWpb5BOaSWjs2/nzdra2LnZhINQzO427+a4Mv0rvON/XYYxQWi7u4eyH3MM7s8IV6
974XVcPgDinpSORHBOCH06TpGQB6Zp76Lg308jmSe3lYP+uITwMkwU1jRIHsg9S3HXOe1N84mewC
JmrlFe006Bx5EFc3K9+g7AufQZAA5RubyI+WxhNtsQZYqCAOFneHrjbUhtoYNRXmSjw37RWVj1q9
VjNyiDSH7oFCVborHnUkYQ1cQZg8KmGo2KVCe3nznCf/VqimYxzP2ANZpk2KueUdV8MaqPlE8iOv
iAd2M4tsqvGN/+KU7Jni6joN8mbyp3wGtATJaDLPfFhBjZq0HsI6rWxsSCmcTMfeex4e8eNTVbx+
WA6QFUnotTcsvf2YogPjHUa1bibj7m3pex5D6EkIT75/fpyjdfiyHi3SvviwIXWe2AmPbCDoo5HP
aWpHZCxUNZDAAqsZ47X279KJHGR1Z6ekMf0mu8BVUVT0464fxgHHvEw652OlGsBqX8Zl+4cWWZmg
gVnrRXDG07sorezDtmOBi04CwHvVzE6KfeO0xVvhDBA4BkOkFJPDzZ++GJ8UY/JaMj0gGBkyeP2v
M7mREGJoWYuzySa/uSD00edME/7XrLPdFRI1ida1UqxfZXVK27Phe8UwdeKMDkNaXa+HD4FCSbgw
QumFU8EDhNivI5bLE2TtBsEAy/loR4T6dqOgV8eadDaoPjG/kf6AquwmNPrui3IYiUCIZkH+YKST
V33uyUAPyY9WeMNqEsgPr6OG8itrSFWmBI0mOCh/KZrfszjsOUEYawGKDyQiWbuj4JYYTw58cFj1
1qT8sNz4cJpxjuydmAmDjWs4Nt7pfIVTyGvzuvI1sv+9Hm4F8uD/4LJm4mUOA+DkQyhqaavHXL/f
tJTXXm0gVXVgdsF3UdxjtOc81/C2MfkK8hcom5K2A3M6yv+N6SJ7/U9/W36l8BUjXImEcqJPKpPn
kchf29PTy/a5DCQtlqqfaZ7vt2LQ5dYZFxBsTM8KiIeltTgWK9I0U82C0iTFrfD1/H+mLcM48WYD
hIEwS0wwQ6bFohfLeaICTQWAEpVEX6/ZALlGRYp4unz/jQWZwWaBoyzGSTlQtt8vV3BikVrCY0cX
QaDco8uN2pyn8tM+2q29/ize8+fZGfKlfniWuymyOXuaVV9vqCTtLluUaZfs2bO56uf3LO8RqUle
3LWs4tF4cakO6OqquAgJIW/YSekUr083Izof4te4JPVvhmZhfIsUf6g3CqZR8SuZoDub2NkxLNMS
R9db+wtEfcrPpiTuJ0vzitos6lk3Yj1I/psplhuYCL4b6D6G665rhuoj38UMR1ck7rx7LCzLTMz6
/AZ1TmMlfO2s6uSSUIsZ1s2cIhhcAu1KlYjA9Z60BdjIqCtNJQQzue/MboOu60rHtdSHvjFUP4pn
rfU0+zKXDybTyHg8jzFIz5Zro2MlfMnCGHR85+0j6+tD4udNGP+ATlQWYvh+GM8wf5uBEy98SpWZ
59PPyvy5aPFCHZU+8oW5u73PEwt5RGqhWcQg8aQb8TruAbWQV5+GE0G6GDOTvpfLbMeK55QkhBvb
x74ToK1XUXW5SVyBri1uJUZ8lxfJbF9UXP6Y8kTn0fem3rKRQFuXJN6c9SSIv7442dixW5OvjfKQ
twXRBFphRDJ17mM7ow3uMWK9L8XO4ygnZ8mWK3yEDbQ7BaG5LQQ7XzB11gZeK8KUO5+rzDYb6BUu
8QXqfjurZUOtta29lMcniWDc0EGMbHTGRcwldNrun78NRRy0U6+ZQ1Px1ZWQ6v+R/KsC1dui1Arq
IHwNw1SQRMcfp7zyNMIdWn9cKXYhwNba70O19YTWF2Moe9H15pbs5ZVV2XjXXF05z/tx5X6dHhhV
5Q9MsQvEZ/kfe1ZqnhSf7lOI1GG5rgRP4oi8kL68J4vaEzgtamjbPioVaWQ0SmZTpGZQHE6rV8w2
BuKPggU14ZhObdOYwWU063hqsnT+G83ikCjwxL98oFgi9/41VTGO/j9Seuj9uMoEYVsehXMm02i4
GIb19nFQJ3nGglcZp84P2dti8oqOSFH0YkHs2Q/tAWYHZGl48EqR9pJ9X1mP8wIxvyd7BW3VeMES
eQc42v7px1vgg+6ssBmmf071wAn+/U9Swd25bKB/hff/COjWmc6oQ9s9XK1XxEO3QjIXSQft5erZ
kYIxJ/GYAv4oiFPcxa4dT3N7dnKmjreHKhQ7WjYQ9NT8GDCBwnekRIF20hoPM6IT10wct16AO0o+
MK9OI4HxMYo7ARuMFkhL1bl4SbJw1Sj3fdUfFr0RxFm/faej9jxF/TdQzOOiGlLV/B4kY27t60oB
8DPjuNfif6Nstkvtu8/QYUyrtwQw6Procr6lpXJxwZOdFZYmtukp03qymjA8zfrj7wadYyZgnGK9
RSeyDdn0oZv1567nnNOVsVYgQ3wFmrrJ2YO6xggCpXdXP/y7OA2zl3FmJFth7+gjCV2FlSVOba0e
Jtvi+EiRwhxnxpxShWvHE36bfVFNuWRSf5XegUieRT4o6wIpdInJ/25vio9IQcSJqojnv96DmfFa
KngAsTufyT9SgD0wzOtMrAQmTA08XX/+vJApr1PuF+EQ0m7u5XWKHdBgoYts1L5yI16Cwh82HuF3
KATrjcAcC9AKxl/JtwSNdakiLAoGA1vV2SoXBwGVc5DWtpw9Adzvpn/wLjLU0fHq9Fttt+jgSwrr
/U7hZjFv19axybAi0EvcAknyATo9mmi1M8Y4X3X43QPJ5k/miTs3WTW8BUTY+k+5zjiQTz5eOh2t
RRKg+tnmEeU/ioHvJwkYU5ghUMafx6yxFIE0sSto/aHtU04IQs3kUITECKf2LuhIJRpazQtdHQLX
swMUaVE5ekJT2lNk2i1AsNkBGiDJiXMLWAGm3TRDhr1AMnVunOyDukP7EySkqOi1TW3zrNkGB2bK
UcaElEhCXoqXsWCJcht01m/IoZahKE/5GhBj9maXLERXT7vUUldSk0EWv9JZsQHH6jK+RgSDWs0b
7iD+RRAnUhftJQAum2Wj9uc/D0kGk2o0wVWh2m4Ro+89DzMeXygbnnppf3U/aPLWooJrsi7Jew2m
RiShEVIpnVTOfjTnxscbgO4QktcfTH7OruwzdP4vv1lZXc8D9Quntdky3uv2jilR52Crw30HFBHF
+O7QRbXETKIAm+ZQ31cDepYYHmsMyATaXdm2FI/MQlKmDGb6z5Lzl97elRX8NdSpBv7BJ9gwp4bV
dRvju9nC0UgFmyak6IJ97ENpWMRiZ1EHJluwB76alUGt88UKOMFdNmYFlyrL90xZYQAY5I2dj3Um
tkq4isQKQxCcROQdkHDUMZ3BQ5lAufxyVksRDEiNmM+SEvOTngBS9vMG+Tu+3qzrzDC8e75OY47j
kP3BFoxpz81HQsmNZuOHgwwfyoIGyDqX2esjHmD2sSZVkJZXm4RIfq/RV3ZwL6FP5TjFa7SAfl/b
TJakNLnPvPleFg3r0Z6PkxKL2xsqw/FO6bk14iBxLghZn4Pwe06O8sK5ed9t8YylGKzWUTABRLBZ
exMiKOehV/bilDicooRmewJaIg08x3KwKYAwsS7o+6ha3DjW73epuXjyRiZaGjFUVHs389pXfWWt
2UDYXROHWzHgLVTVaWxxGHyYcnjh7DLWwFn8HPn9TuwZUntEH0KKyE1hqdpL2GZZkVbKH+mYKB4U
g5dJzYmFdBB6dH1O/DPHeX7/yt1tqecN2oOuk9fYKcLoAZMV8VUtz3IseKfjaLvL9yD3swe2N7XI
ezhSbKZ+8Q2PXz9gGbdlvzzxfg+iS7reIgGilHuemPFtBaYx5Z2XmHlxHZ7qzMtVe1HeB8WxN3C4
+lo5ClFcEUb9KjBWbOEXVatFw6fJwqL2gmEDF0IGobN3KnH+1XJR7utK5Adh6JIEDTMzkTskBNOD
riCtIXFiF6lxfOiriPNpEQuL1+SOFUAi0/fA2yj3BeKju7KDQTbuq2RXSK+Vot+b4K5qThWoXOpw
Jid7zB/YMh5jmJbb5zQBrE1q9T5yV05IJ61OVQiekslHbQfvQTleMlbi9wLE9SlMug5WcXDbnpTS
QAqKyyGJF6fqcR09etZSuqoe/Mdhukmb/Ky7xIq6tXRI2Gb9Y2NK7QRZPwZjjr0TS9DuDM+11+re
TDYxhW/xBxAltIiEocRxBkEdPCrtuC8p9bNuUMlTSuGL5BeCWcuNbC58WzRvCf/APfd1s4iVJniY
2spU/4LctxMWks14K6Go22b387D3qiUwvNrw0oekyt+jaJXwe3auxBOCbXKSAc07syyzpqipvKYt
88IUL0CPuTPHBoEuD9dq2tWXaEA9V/zNLg7gwsSmk8QKZ184p5hHX+9EyJ8K864P3DwO4AeHQYsi
OjDXPeK49+FDC0HAZ6qZufsgzyE0bsSJ2PVRVdP/ULCIraWVAZoenWRD0OsD2HDA0Dal2Vz+wdht
/Ewy1ggJnpwHwNU13scqlhVNT5yJuDQ4N8YMP7wC/S/4KxjcWPpzKPArh+BPBDA7Fk5BRu2hREmi
Mq9d5m1n8A3hDZgWogDNkuvXNaVf5EW/jGj8oiC7I+d/ZFL+5TBZcCd4PB6sK7Ijd7fOfw8Bufu+
3oDrsul5+WtcvBxFDw6jDIYBEhdgts+PerEHlt1bx53o6+BxP1LVpGL0mwCwiPpnIoRcT9GRhPF5
rOf9K1WZKbZfjLWbntO4IbwkxTQzZOn7+AYpQjQltfjwjRNzJY4VEEW3ktk+JMpfShCu+QOq3R4X
nV5zQS0elTvDbzeRLPrme5ju0HJELdeVljV0VZl99LHcwZGJwaG8urpCrIn4i66bjgec8hqO/Ts8
zoqQJcl2VuWMHYw28CwoIgl4Wuk9aVBi5tgv+9A1HZRhD9nE4QDnNJw4VirwHbEdHgM3J6ULix35
n77XuDbPI5jqUIubDiMuj9ewSvIAI2MTxeUYjXjs4jMg/raNSMWkK+WcrhOorGY+2Z8KhbvoBxKY
dSuL8PKLhFmfBU6vPhp6szeqyr0wljeKSAAbuES0wevca2NjitgEqmCUBhBDw+JYecWybkK73cls
rscWO5WqXPLA50AEAN4USTi3g6CnIgLJuKyWXgZ9QlkXZ22ym8MiWg/C7Gix/qWuMxZ+RZpOJiHt
Ie6VKsihiWuGCF6CX+H/+6R5IvyXoaJzlLkX0vvYPMFifgo8DMQET+NQHGQfsw85cpFj1qW8M6cP
0bkW+cq2CCvpmpaJBBKU3JP5F8n5559dCDgN5/LA1kGuLhK5usiDVFVs+ou0YQJg5S86JoT2kqIw
BWHihiMgjAIo5S8KufXh0G/qLJrBuTr4pJOMXAiyyHSUG0s5kkeFBVTX8sHpTw/l12r6W+HIhjHR
kUwT7PZrHZkub3wooLk83urz6NpjpcqhbP5WyLl7CNhRA3m4dj7ffyDSsXk4HMPIwpHiGhIvrUVF
KiSG4zQWaUa84EaXnRkyAtaRhqrtVRdDFho9IhVAln73qiTU++BTVMzjvBMFbPAeVFEgUo/3T5D+
3jZybHHYjNqadFauIG4tJYl39QYrO3EpDCv8jZGpFqYIjxH5pBxAoXFiKQMQ/a8DayPt+wN34VD9
+jqt2Dy6qIF0Glgdp5CwlLkSmZL/y1xeNFnjCGbVyFs2PeYwH4hJ1hHOFBkYLfw0B3IuIImx3aVZ
UM06qWhVJoL6hdk2sHU+iduFgEUS/VpU2RoMRKLL1/kCsqFqiDKJlPouHKN9VrMVmM5pzTvkhlVA
6/isOq1HaI25+t/yEjXzulPeFrvjLJ7KctMDar7ZHMfRjzszpCcps5GW5mV5jpGyRDGOInEhVv9y
fMEYqyhZ13C913LaxHQhxnDSLKEZzYpyT5A0Hy69AL8UheYfAE6k5xmcIIB6VsqQ+Ad1CK9KPZEq
QJN0OlBuF2i6SJmb+eSll/VPPkOAoTjPxbIGt/yED6nEQnnjPac4ruGYTPXdxFFqo8C9uo9sLTjA
5Yitw6dKdBOPGzBRp+wS1zcA6A9lqAnpcUm3K4yXHMPRLrLsnTDTq8ZbtG9DUlJwYNSAwc3u04xX
5BnP6vXbkECOgWEb6UzuAEgVRUd5MPyEIvOlOSvVsLMgBt7g7cLxFexI2KPSNznf0jFLhrk9AfNx
f61LnIg19At5lWK+w/YRmSNc2SsIhq1mzXLSxb+MLeUUw6zZew5Dj0DiPjeoWB8NvZY1xA0+LoW1
0NWEe7s3ZiAtXmy2wVKYqUWtPfGhG4gAgY/jy/MZwyGvfmlbecAwkfKjGg9r99TGVcpyYgrPWFZd
2RODmvHmHBlzZd4Hu0y3FEtydcyOkfQu4fLDqzd/v/UEPgnP2p6ThaC8qypaj0QolqkSjPBYoWwK
Ucg7K+h/4qot1RzuzyGYWdWRv3oJhukckfLFBWacRQnqZxwMfg3SDP9GILa5UgeOWdjXWnaYMxc1
Qa7QwFQxSUm4q+2go971kcHQTi1R41NLCKnwk8SeqzTgLIZHSff1NecmQMK03Bm+mPvUXormH4Qx
CtYYfBBlvvkDdaKefGamOC9KrhdBUiLzE7TWGrs0NKEY3t2BHFU1bHsRq/e+gBrEw4ZK/GSDeY7B
zVGQhdhsw6N3DzZ7VfPl0mO2d43yQLyFYYAe4RpUjhcG0Ipd8EHfXyGkmiG+KYPcSh05IPXcM27j
GcI1Ek+WI2raUnj0N+PqywELoLr9L9NgJLFEYh6FSTAW1wIUTWKUD+/iP9kL69uBgHRFeYjI9nta
9WBQb6Ia5I3hg9KSMQJdEOJIuWpRK4Na4Zzy6H1rtBaRUnfCXA3WCOguoEmNE7SJKqXkj5Bt2Paw
jLQ2I2z8iGQmXCwCIkV1BlLHvfdvCoG5o/k04gNuhXAh97qr9kZEiOLMJP9J4lUUBvm4W1i5Skda
VhBaWW2xL7T8uz5gCmc1Z6X21Ri8WlF3or+bL7aofKmjPP9UBIThrPhgYEIp8JLsAecQEhDJ9WrI
xQEeOVHh4us9rdqqOqneVyaMtD1+klIMfXyZgfJpFxSjhv+AJ7FRNrjepkFbqlLU/wvoSzn2rqtZ
4xbPbYCvOoybdeMXPopfZJ4Eu0yJnku+op73Ra7hJbonov5jPRqRsYdhRxSiis6EYr7ZpKhZsl/n
2UROdsFXqNiEj9hnlHLWgjg8HHKP3UCOe2yiEHpVBG7QdqczaFRIeZND6GpB9oDSznRGT0peSju2
8YvVMcMzKSUlH6577WdBgFWxopcGTTQBNBwb/G1c3+Z6Nh/vMTAtW54mcCrU7BbmBQCsduC4886i
U8EZtabVpNHcfWsBQ/xX50uRbvBSsXSWDtzPHJ1TynJOBqS+Add4j6vj4pHOHZUYnRXTKN+zflB5
poA0VHDFTYJ5nPZFXZ1XNvKB8DivYOqpy2NqS4SStCo2VPkYIfx3rgbzwYzYnKVtBDdk+Is20qgh
Rn1/hEupNjiChnv/tn9oCYqyu41g0435BHNnQCqCx9VLGLSRN9SMMIUIJepGy7y8LWK8TppWa6/w
/PRU8/lhwuHXwdKKupQibJuQjsRTBOq4JknA93BwRfpR1NDh16qICrae8n4j+srSSco8ViPeiNiH
FRtf8K2nQocksiTbcqHWPqjFyRk0CtAJRUDT+YtXvR1DWvF5+bPA3j3UMl2vB8zA6PK4+Axh7lRP
oQGQ2VUpo6R1j+Nc66JSl56l1eBNKZ7xl0m6C0ZRiTnBHbBDQXc5KRt8OiCrf6+Txu5m718mA9yw
YC8UAKyiV+dLAY5znp4wfxH82Z50jy4QkEzaemzQZitYQz1A5uWzSm4/+xKKxga40Ned/bd65+pl
1idLeUW2V1srkIhC3n7Lq9gQvMb9gjdYQ7bHZZCSYM5yRgD2VFEERjsRetY8baxP13OXTAIWTWDq
uTy3qGs6fuPq1FefUbDfnpnCvIUYW5gwvm5CGS/VRM5MXJL/QxZKaAJt58WdEgho37WONYw3OLzv
0v35Mi63cw9iL4A=
`protect end_protected
