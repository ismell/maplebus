`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aoaiVYtNKEi2IphLWpIYjhvGKL56iz/1hZrHOqzlyh19Tnzq147vxUgLj/EcxcTLR51bcs5dOszO
wlKfbCa4VQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lejGYRNobHIkkh7AcLRdJgDyNmrlmFzcR6R55zgS3CXlES5RJ/8KwMnqbXzIWfuTKb2xwqA/Publ
ritBFmk1IUZfNdhlN5elCoQ6cAJiogE069ugAOLS3qmNg/lXlDeToZFO97UDDHA6Pt/4T1hGxQ3R
ViWNx06G+gIkLYtoiaM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fXY0SCBIfBmx3C+PAIngrpitGp84fUtrDM3GaoM07m/CqZ4bE1nhNZePa5i9ju3W56rRhWqZxF+K
w0TufAJlbcT7yC6lY4Xt3pnRw1vzdLBRwx1IOkHCc4/Fyeu/eZ6VhyeIhfOPGfVtzapshmhcH21Y
hJu37LINaUhWAWc4waocECWLC6YhUjtjmb5lfvi1PIK9xzCgIzebnl/OPFunVaEV4GvTJ2tEDPYa
yMKvOF2Z87c0ocAY/DVhXZCbpgoezPS+vCDL2PjtQe5QuElrABhwbYtHIL/kDtVi5S4sHHoa40g+
c7GQWmkJ19H+WhKrwgwn9j6/ej6j4oX6ALcLOA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qJ5QYH29KgWTd3pRXcHFFJQRAqPmxVl/Ikmgsj5cO1yp0WvvJ3LqgO024s/esNqGuGny3F0ThToe
EEugA1rC+gsVSSJ5TES4Qpa0MYXN/Tn28KZuXOhtqq+Kpw93uC1kgFQ79iBlwtg+Pt/d6Gs3qOuA
8IvGyiu6A39e9BuaHms=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qXXJ2SQBq5UdS8pqGKLP9O1fOlC1GJMDsLq01JcpbvAYvPpDIuFgpnWA2MW2y5sWKxl0eFFo7n0c
0D2sV2PYINxxnSmeiHhAl7rjUlo2/BicV6mRP0CB1vdkq0bGSEmI+3wY7PTq1IXFFqZqeY55Gp95
8Ns2SwigIHSSSUclFogfWpynLrhFkjBAkzA1XYOdHTX1UKikzl/w58cor6e3pXqYl075iIwAABz6
WZU59++1gEuEDc9YAzZW9GtgcsRblmm3CbJoZKZ4MyQcgVZm2uRSQTcgD4z3jD+ZlGIXu9EYy3wU
ma1EpkWO5L1EZWCgb433YoR/SdJALYQc20+dVw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
rDuxC8F163jNS0GGKhEMuiD2cBL33FtltVj3vzQSFMiPaRdGFoGMKkxN5vO6DRcdXs5oUrr+luPO
VIK6o2akDZUXRM+a5cS/+54xYx6P5C/muio/NBgZUf9/VMtRO6UG25B4uJ5yaroQ+ft8yFhjDgIi
PinhhJKkR7pPpgc4pm0jRndAG4MziPwAOEYgGht4A3GVCX8M6TS5Z0lrwnHKYYfo3obV1z/Sa1fo
wMrzyHxuHEjkRTXTKENS9EHgmhJEJX+JC68K/N/T3A7Bc4DADj6WZTGtkaOwWZ945Wr7K+4qNVXN
+TSGXlbB+dC0TC7xSsZue6tJN2Yv2o1rwNedyfw+kN6wwP+f7BFpbYMBnbovmbCdS3zjs593KCF+
Jia4LrmWyuZrSw6FLKBEPA6bhXYJ4FbenhX0oFH5rJii1k+I9BBnuypVFo3vFftFyaIk0Xo2izXb
ty1nIudtCTOg3AQEFpSzC/GQsjYSZXp2IfMWEt7sVbBHu5D0KHJQIzW1joJFqlzci7eFdhV+Uz1X
5v8fycIxd/trTPJxYwOEdllnXAeuqK1ef4lj/TN+alL3BroB6ESrk1j1mR1V4X1h9KEJncUINhpC
8M3iLzC0MpwxsfLjFljsiOeH0On6P0jnNU1TgfCM3pezHcXHJ5vtvIvKcxL79WF0t43FETw46N+Q
hXZDPzOLw9w2wuOFx1gNrEJSxy45C5Qz2f3erkKXSZr0zBOcK71ILebr5IuscSzAmqUl89yaQai6
m6IfKL19RQqW5l3JWR9ZX3u367JGFC8R8DOqAoPcFeEQ5K6k1Z7TZ1iSXmqetXyaMIlj1s/fDA/6
gbgP1sj8N0KClpL84omws1kQRYJhgECxMLJAsY7qhqDP0iAj0cwqVxvdzMaL+3rpBlF2VXr9FLfi
wsfwdqcknfK2hes15FfuV4wtnLG0JH36h6hd9oArMAbfxmQqOJD7uvxMf2a/XaouyOIjYaa6YyiS
ePDpGx9fsbNcW9HQZphjxyW1/Z3pTh/lJ5HtFeBSZAkKNWB1ClLRC3PQPa9sbAT/6H4ynSeKiCzf
FdzRUPDWX2/dHEEX5kx3qJw8oLP4Taw5p6vsxwo84SUImE4TgGokzP2eXhCp1cT9OZjZ1uL/lScw
LPFWhHL8yXJiLI+UPeqL5pD3Yk2/0KRZVbsetDYP/JgfXx7O+I9ITvMmiTIdXJUeP/54XUHQnv1/
9+X+uQTDemfjXKpFg2Pwc7oJQhNete5qObTDs2O94yUuBrqytLZuvCq1QhUE6xkA0Y2ohMq1cFbf
zW13KL3Uh+hQ5CoBTeUb4TEizN+U6Qa0UxqAJCBC7jqWZboPhrPciY4ecCxBfhta4tcoc0Ctu+/7
OJ8dPMCgWuO1gc7IzAAAVEpq6MVvqnZqoGhm2JfoZPr/Dw4dBeO0RkhHVRT0tzqg8Zg4LyD+Prwp
EAFiGMmTKa/TLh0kij9x/rQbyhiVFqru+GxNZzaGA0spNjzoPYdO8cWtScyOGXD/IeWhrpS6+6Af
0Hax/9nLdf1DvGwBbE0s8YaoF0mQIgcQQGOWO1wTrB+IPNvOZ5r5LnpDnoLaeD8SN4loD0tGjUmR
dR0+CP7OAyyUARR0nBSQhgD/ESzVauWeH2Ro+F3A7qb9EAx3FUIj+tC4kwkaKhRRZSIfWYixowNg
xzRksKDK9H/ripzPBcMUA5LaGZMeZqag/vRXUmC5j6Pg7Yfhq/OXvC2Oiv+vU9f1Rn0n/e+NMdWn
XxblTb81wk1d97PNeXSJ7zGkSv14XNikMZkkyf7mWmfKKsfXVLjlI23+03ljPu15JvwAQZxroF/2
qrE8sq0hmyQ82XoXtfiAv6gBZy0NaMxH2cqfF4DvkUperIVqXu0GSNILUspnKyO4RF49ISJ721w4
iFIV+UJdyV6WfQFEBXZ+M0ayFFloUhdWxBukHP6R8Y4w7aSCa0b4xuvH4AILnfD8Y+MdNbKoiKWt
K7r5bdQbIV7bfX7t1Fvrp5QUT3TT/oDXx2NXf1CTRYES8kHNGGz6C+YMRQfKlxSFieLCTx+BLVuL
4+0+Q9s7tsj0QPYUdp4wvZndeVKFjkiKB05P+7CqNtoVBhxAfLPWHQxU1qRISwIMZwq0yDpP349b
BVIlFwF4o4uqyxm+dEc7MAFlDk7ZHOxtBCIdI+ofzzzhfXmJDDQZUaHMyyyOp0RB5bxbETUW3Oru
vEeGLirhRXZqnaiT6MFlYI0iiEz5xmhho/2q+yVDvkGFxjIfQtNXh4b+UGx+6ygQ/z4eFLbpsHGN
z5WUcUX9SeaMj20tR6+kEbxskIcpczYS679Gdpxee0XIZ0hkC8WjqoLVz93GjqJWsGpKJyg5UzpG
fLIVZ4FiOHKEmgeewwMEI4bNMMkSEGxkgqyW/YX67ZCScwHugVzF9niPTGcau+QlyC/yPUy4txKY
NFVzXD5U1cYvGdX4ADrPEbpvfiAJ+E6FHEhwBzU8MsjonxKRNSf/hxM9E4nSGqWwtZJOkcgGoLIP
GZXLhWMHtxXyUVS1hL1Zv9xL8mOpdu/MkRDckgDqEVg2loNMpnRskEhLiOHPu6JkSOZnR2kV1FkU
7W6WfkL4RRx74NisFFSF9i0ljLyGsjHdoTWDhLlbHKhef8t2x26PgCaSpSPbquBC29cobgy4iGM5
kEMHhuDVBVP8rhbCj0GvnNTrao0M8Z3suTR7sh5prjnRCLBEzd+gBg+LHkdP6ennlKc3xIxYsLoT
8Z6dym5p4U2jYmLQK1rlhEMx3oa210nom6+Fx2vprtu4c82HkxMxcW4YAZWr8G0fppTcs7ZWDohs
84MfuXc7k7AvNX+cQ8mE7DTwQ927EJh6S5aj0xvwlXAm6W2boBuJO2H5e4ZlCeC66W/Ae8UJ5Iz2
AMDzt6YWKrjJQN2x3H2MXFCpxU+3+lnZ2xCXVuofVMDHTxdRgMJ7IqD7rn62QMaInDfVf2PnUql9
94VuZnOCsj33frTN27WogL7HzPO/e1yYr8gzYzQDSfguM7HTJ9lX/U0wc4D+dhpVap2dFX+QN6Gg
xbiWH1EmC9memvCPpi1wa9viw0MmOdd23nbjBp9FMqh3ij6o2AMMfc91QDw/1Aht25d2WeBfLmUi
IHbZYUAmkZ2lCNWpeD0z+STzV1IxIACv8x2VT8SduRvwgZ7bIOyIaVEOHfJrZiRo9JHx/n807lPg
/mgjTiXmh4/wuQ5xlWo7bq5K5Cm6YhvCKGWvuNHCDMv2Hq6sHYMdaD1IA1qfszd/HijUmEHVza98
1+KvKaXtIvD8InBM2/pqB27lss75l4Gfwm9UjxsF8MCVhlFdev9ryCXeXNxTVA+3bu9Bn8axXmUY
3ow3vODAjNTm97emAzywJi1q2RNcKrV2QgTUTHfLbpX+VafDcJs4oNsZEzrt0gyt9EK34WRqRIUZ
CEbGahu9xjGmRl3pBmVealEqcfVcbPnfW69vyI46Ewfak0M6nu+sPlAvmusV4yLd1G0hP/p3RZNd
O9HO61Yt36nMAnkRa3kvc8UsxjnkV+3/C0bhHeAkYocMCsTUkzcTNmEbPak0rerakkNJmGLcvy8Y
AjiuKe9ivcGeo3OKbgYQYvKmYUGAlQP13wq3OTp9sGXbKBeYoafXf3Yg6uqxCa+su/DxaFfOkcbT
MHH8MYrEl55Z6ckLRvqyKBtFclO/nARuI6Jr5iO3Jp1KouZVUcHOGmXmrcklWuSFn+IuYhRohBtH
UtwNd5ZM4LpKrHeQ+83fcuVKPnuHqScQJyToBFoT8SsGlWW9lznjzQIPZHR5c4OhLfiXwtP43fBZ
4DgXLk3vAS0aPVkfVcOumbSn/Xa3Rpyl3y87Zh9kqRyLMVO74hRK+1Z3dR/BiFccMCklHeW3Fqm9
IbGnp6lnws7SyJPCCfOXKDfAVhSAa29r5rOIOb4M9Y4FNi54G1Ff96KbGdCW3IqKU5ULuo2OxOuF
35NGXX5nWfVgtNSLYWZ1N4iAlb6R8Wuo00nF8cVEO+UHjmkUMPKcoq6NPpGb7byryMZUWwflJGAt
kPGn2zJTsAn6f6R0zLlYOCWdcpjeJKEgPpe5gFfVY+bPeGB6CXeXJ+86yJIoiMQLJ5lp3fP33U2r
OR5GAdkQWDGR4hzIvLgH9h6n5vsQX9fnKoTZLI65VJkk4IZpietYQmHGOIrjgmR1odV0wlSLNaUz
/nDSPra0r2iFJL0w/TdCU7FX5SjmUHmgn/43w8nN/O/3d3OL3tj3XeWwVww9yYHZSq2RzIGdB0K9
Yo5TdZJuKZWTD1n6bepoSbaAnQk+5QJUFsFwU0GRl7k8H1xGaA2CYh9FGp3FVJQIHUk5bPQ7h4k0
7PLIl8U41WFKmIJ5P9LahtJcayyeamqNjptlES6pWKp9KbvCT7Mh5exQIVpo1ZxVwrAOBps1H+Hs
06ysIKJSso0ijgjwB7LbRA9/+WtJa8AqAEmiTcxZAXxpe7wq3ToRUZm8Hj9GBOck+oPeIuyusmL/
bCMM6Xa/7dqljzVu0zIDn/qb2XQeEhNdDOEdMmOA4UPFlMm5CTfBya7XXRZe29E8MeiYCpml/MpC
dspy1CM1c76yToL1Zfw1UMChyynVOd6S7EvanYowCLexIfP3Lk+sRLu+dR65SkzSoxudDpgtTx1p
NJOrMrZhRX03/EgO6Pbspl/Ejl4Wh2oAlFfI8tqgaXjig6rQGp5dLaL9k932pLtuNfI7jBFDO6pc
O/91Q6i69npJuICYs+fuy0cVlX+bMuJU6PQJpPA9MfY4WODhp/vcAGSILKo8bnOXEf34/WCtbARr
mbht7QZl/zh+teLY21WQSqlMpyqsdi+LB8IautFg0Ck4XWeCu1eHAB3ItKMuwlA3JwU21xweqJsw
gr9I8oj35DdrmySCnI0uBvSJ28LhlHCZma/MxUW8lYpv+8hKZdGEYQd9BxxpUQBRfyyDqB6UGLfN
kRtfBPYthYVcR5Atz9xkDDEqnR7w7n5tfY+rqntBJBkrDJLDPIspaFLKMA0sM15LBQiatMcay9Er
Ge6OrX9yCSI8k1kQd2D3Vhnxw+AcW6PNDldG/XHCkMXIQUXSLArgcN/oSPjEhRoVe9v1r4uJSaOw
89MZVTVesQ0JkNXyFlM5PsK4Ztjt02LkPRLKQcq9mgMr7VkBCseGXKm1iLxA/9sxH4w5KJEiOYTy
FcupYL/H337mtzuHkrG0g76XUys5J/xnzW84eB2fWRUgElhulrX5ltiTqGn5AP8A1xZDSkSzbdAI
SKbIQ1ZmtyDJxnkpNn2eursdmQrr0pIMEkuZHJ3g5jehGH/OKy/lQ9vg3vskvtlI5XT6gb+nEk3F
27w30vro4iXLx4X834jJzjNwXPnf8LD6vMFZOm2jpwqZOgKcnqPymJULtrYFD7hZt+InxNcUaJ8Y
baYJxtKuOZBb91Ud/Uo21s8FgO5Yb+H8O4pEw4c3ZxkrGG7r8LpFVJ4P4jspPRaROB38NJv5WKoU
wvlcr8/FSYzgPnLkVg6K/3UvZUWRIeJyDFA8lsmFbO0AYnTXDEfmGpkvgLdMCVENVmr13S02yujA
VkR5F+RBuIY5g0adpN9slWq4V0P9d+P8eBm69r/f9wSbgHRgiTIrW5yKtbAT0VpH073kON/KBsuc
AEQ2KJr6MRXRIDu1kg1kDnZ2phdGu6AD0HwN9wMa1n03rDJ0eMhATjmkL+O881z7d8Ki2ygho1g5
4PAMUNhN32+es/DppWHSl1K/gYGbE+AS0DGeW/x41V9D/LKv6vUniJ+bmMXB7+K3y1tbfExqQeVe
VhqBP6u244dswWUhV4CdwcdiMqPG04v1/Z+ZJbd1/CWBm5O3yZqtsJAqeipFTcbVbwucc3eVbC8e
DsQp8XwZRF3PCxOXc8OC8nt6k6IBxDOr+iaiqkOEjIt7yqseqK8PzUh7gABI6tpfoMOf1+4Tiewb
/Z3UWIfEJutXiJJ9sZevDrfVQz7T2Q4G20B4hcXGmrgsA+WwosE7mmfKUWHN4XwuT0aAFJxvdLBG
srQCDXrVQsjWgeQ3toaE0uUas02AkZ30glNCaGz7ceScygeJtzcpNSyDsVCmtdYP5hsYtGTMAIuz
5u9TQnfTdDxVFgZQhgSYuRRxLmps2uaLlxOsGbmjsUXRsSVaF7OIQL0oi1/mS7/O6tm9EQyQ2/XG
BGpauKbQxwkVDf1QHnVqbGUgzO9vj6tMj1hyP2FKrDaEXT/9203NXkwc9UI5Cijj2UhZd1mjnqur
BqIzcbegRkJ1mtEnNE8maCV8tXHrt6jctRUxJyWL7cHCB4+u72gXI0OZT93zk+LWAGlY8GnZQ5uT
lkAzGlIkW/5cDIuwBsN68clAulIkx2ZoRZPjhAc0lga+lGGFtSOb7yc/Mbd/ld06qy1LyRuZqJt2
3gqFe2R74X5wWSwd0/ECiqE1EE+WhRwvHJ2Lv7czOaYq9KW/x2oato9yMTms7eppVB6cGvUdoo/s
13VbB6xUxuVzd6q8Rx2OTXK3eu8CdzyI95+nz/kp9AjFiow8xVeL1zXbBLrJw7QAH05EV5jUrKgt
R6AUet2T0ImXSr5AYiYp4HpwAFEON/QlSSPq26aWA8RZKGPH5aZxFwq0Go+NPZS3TO7WMoSS4Yzp
JA1TmnY/p73xEOablE2rzSVIZc8HrY4Irq9HBdOaLuVijshXjEWLwK9FTsmrRGVxOKQTk/+nEFMI
mKrQifCut1axzygPWFT1GxbBhpCILE/GTBcNr6bwQZC8fqiBnUYy/UbuPGnS/vbgS/RIZpVB+Yyx
EaC7YAq+BKehn94m/+wq+YAjHrsiiCa9pftqzKZrM5bdRSuvoSQLfwJLb4EI/B/AWM7sl8GR5lJe
ZG6+OPKbMIyYuiib52abPf4Xk2V/pyMVFS9j4I/Oks7+8be6ZWmgr49C/LTrwHah8wa8+uwjUQFv
3/HJ1/ua06MRTDLyeZz1DTG2JYq31TfBT/raR5VbsMfLIk3DM7MmYcJKbaB1gX75WDRu8muQmfV2
c8LGyv82iXsTD5NHSV4/JLzx7xL4x0epm8hiP1NA/JH6O5shd82ZBzOQ1jqvkQ+9Hg5bjdnHrkLg
BWlYGikxuXrnMInTD58p1fmXs61+m/xob7sA3XpODOf/9LCo19IEPkWqdDfTocmZwPNn9XK+igU/
Iprr9iT7EpVVqaX58qlB/QVdrxWWWP99nSuCmqYgsEIfxJumjj8dZGh/O9ZNmxUKHsPaNEeYMLAQ
SP9BOCrqmLeodGFZtZIvubbYiFid8NLtdf+lLFf2oRjNNB0mdoElMHCoRiKuELaE8DjNjldNt5UV
hAYHwjq/ogXCd4jQSl3lViWM9qtqORZ6odBUIA+glCp79VX9fVz+6vO2Ij3ZRxhRon6ksfGlQKTD
k6dNDkCDPDCgSmHF+9lAXNAV1jc0JsNlYvNbe3XVBxyxPPC8ECD0qhh8HEnYiGmaTmJMMkdZt8W+
23peclqwxiwZoLXMcyJUIuaNFvC7VRXEjLeJOZXlIZIUiic6IkAoh9/8VnfDM2eqSezSPpLz2SbV
UauPMOKKO0Doa8oZmXtCI7wgdoYnnTiSUEyd/XpIFnUrbtQPjkITHEaPSxfpnV7nPqKn0qELAP8P
INZqoxTSWaRyZRjnmZyZnxE1vWKA2ng3clDaNGXs8eVWjxWDRWrNzSo3jbzSahsV5pPTOEt/Vrst
7I1VBwMkxMxBiVMTjlimTKeziHtHoKlEp1kxn2WKwbURL93cyBq9i0uPSHps9+gcjExq43am8PMG
bSdg19vo6EG3kg==
`protect end_protected
