`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B/Lc6fP5S0dhf5AflLymK9Z5uUNdzgoWNSj7j0QZJSdwUJ66uHyX0CvmQB28Bk/wxl/yV49htveM
AhXEh1hsTg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UhYQuft42STOBGzVFu4+IE+VycjI4EkEDO1050jHbDa3xnOcVEsAaaZ2lXYfhGCM6btuVqQNR9jT
6sriNyq3mNZN3TGOSuB3Dqr0nB/VEK485Vdxnc+oizVSx0YWwpONw4Ls1W6paOZGjG7VzSy7ep05
xS/qqGGxidEoziUTcxg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VcHUlW7/EZ6CsY42ewqMQ9996BSW4zyr+O7iNaaxe0exWNqt7MXp219e7GHWE+qWTdPTLG9/f7mB
m0gf/WqoblBmOnOPREvPJ7WB/cnuAkrI7vY7yEd3RViPzZCIoKG3p+FDQ9dAnLmpGy+02szEH+If
qH9nslE2e7tCdPfqwiZhyoAYOXg4PPOsljb7IZfqlURIcVy+BUwqHCGZZFjy7bH51A3yrLdBahHK
B4Libm/QzYRiXsqjiQsrCnraXp1BBRkZbLgQ2aH4LAbshGeASNn8gue6OXsBiK70LYK4LMH16yFk
aM0V1SjmHi6SetaQjPutRmWYjA8Zt8e+XMrzsg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zEZ7lFfOyvU8lLVBVibq2pjoIFo5FwTfYRUqErnZqlUtRrqXUEvqRAkRBVxK61Pae00fJC9Jjb75
d12DX3lsAH9bhK4BXTHdJNLE6Qb17kxDxDh3VJR3Xrm7mnRZ7SrbotinEC8JAy/cb5+4Ja+kPGdn
nV6IndJ5s/+548Ner4g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Mnsnw5BfmhO6ikiDgpnJhnHBwBz521caVfGfE7vKZvpBERbJ58+Sd3rOfY75O5d9hNaBDFxjiLgm
VLLmbb0Q9+8ZeROguap7rFzQXK5Cpa0y3D4cw6QnFS+cNE9gGfFbQAl4AQzFiRIrxQYhpNeXEKkZ
NCBdIYktabOLkEiyJCE4dyagsXdV8q7M+LT5+Yg30Cqmp+Lf9XPH6xCZZ3JHUgxm7ZImn24nYGBK
XDjeGRYLH6IVFYDq6IiwG9BPE7szd5mQaqtJ92OWi3cWU1lDe5sHwy63RLMzw2pYmrvAGlBh9Hxv
QKDn2Je7tMVw3YQIT5x7SKReCz1qmWbRkP8l3g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
9pbnjh3iqELv/oQfOy3Y2Bhey1mAzTCnKERzc1u8es5a6AbahLEsZcFLBsZKffuvlmRAGN5uolIr
R8+ZhWC8LvkSgkVa6mztcDwwHx0PnZs8Rh8c84ZU0G+O1ras4A5r+8eobZpJORPbjzqzdcZUBuAL
bq+a/xUitgXChXDJcSZSDXIBKnKYPQxMlJBr6u6HfFC6jMR/AzV7tJXBEyguIU18TkWTjItf+V2G
cipIFYY5GURKqgfKyXb8mwFnfc2TAjR6hHKmTuC1+y0d6er6aRvvt8pA+LzzS4JQuSzUHhWZxgP3
9gIcABxoIqFG6AdwZP/uSKIrc0KbwIlz7WClkLIMUsuGmANacWMZkALTGAQoEa0QY09LogLFtbPS
7bSjmoOkeacOuR57rqUHOjGkjgT80pvme592FV3Z0po7Kxi86aRvoKyJOukAaWUAJSk1ZsFlyIGh
xbbMayHeDows/wV9+B6wxQbaMk7iWp0MpsSdhjiKAf3evP/3kaD8mQmGrlLm7n9eX6Oqdg02ToKJ
MVoRfY5RyGu2Vzq68bZNPfhdfqD4R56pmIZi49Gk4YXrDePgX29+KuWt9Tk4oaXtAvf+kVK8hdgr
NPkynnoWdhflU2HnqsX8qac539kLgTSXSXj1yzzQ9ylwTTCeTBj/aoWUfrl1ellxWQ64bWmcEmvv
10xMyQR9PYl66uWasjxRrpOL32TsQoSaGO6//6CE3LMKLIfTsob8dnGXhAIeLnZK6YqiMkBZofLr
4WRnSMMU1b1wVXvtNoTZ3cPZNr9k0/aOYKkcGP2Jtc16FmAvD3d3uECU8JjDgHK4lJ9+poJ99Ptx
jUUerUo9CBfxUqTxdHSIrB/kgHlC3SyZLPaWtFSfMDeNEeQM+xjFVt9LSC8aO1rvgAqNrJA65ob9
ipjoyBoPQJygRUdnPK/GIBt5kOYDFK2tGMtK7TzsoiLc/oIgv3VB397oB+uZ3BCZEpN8wMUvIM6p
LWNmI3Kucu1vKjAu5RhoxI5BM34QFIjyB/aBqGlzZy1e1ssTWn2UJpWQvcqWjU2M1ixb1sqD/dGe
EycBzu2zIVxY27Sji9T43X1/SQyr1tjj8W5apVHPDhRumgNSjy/xuzqmK2XhnBl9hEPdCehdwmKK
lkv1+PZrJ20cwCPpZa3F7a3ho3gA3GWBbiuWnAkxZkWBlESAE0+TPNpSHwdPumDNahM479lU0n9P
tqooPHhzhtERXjFauKhIxC+JWb30/S2TaPiFMhMGMHfD2LecA5H4jHDq3V4cZV08vqiOkyCJBh46
dOT3XfwUXaxdZrY9wAy6qui0fnm3bLl+UiMImWe1Zn0kp61bkcaiZ6QWEOnJ1PjNMw44xO0uGeHv
HP8BLikX6k3HATWDSgJ3cxZ0dpxY6jHSVuBZ4eO0+BtBbH84iH+qXIA9Wu+OTgAOYjShkp1PcyyH
XM94Ix6w+EAcdMgYcTMLsexjLkbWsbnaZ5pKJsPgVWCzqL8UYSMLwijMg15EnCyfOPDVCT5WEztE
6Gs6u3+bOLtDlBTN89CptcYpmhgT7xNRBhAOSsSIBNlp6igyOq6VKofsNPdAWDCW+bmny4mlNkNm
q/HNT1kCHTZ79kR6w4KBjIsbIr0tt+yPya+1nufpXzF9Q4lg4OiLD+NGxo9/ultZsF2W7KoScZLW
y70xrJYBGimMk5v3XxFSsaSzN2+M+hIbK3Vh7DB8FY5ZY0Iiy6CiuxXYnvQgeoDgeGDKYcTiT6eb
yVaXVhvlj46My9hdaTsf+GrbXyr1u7uuZSM/shjdXeS+WDIVm1B/LtlT+5lfc3zyAyfa8122PATh
aECEWxJxIKXL5NbOWQizWAx3wg001O3F2wvUc4qAmqRdLu0qeiXvYPQlZ9LLFUBbmxZpWxKkVjB9
vsyPTdpQkuWWBoSbQ0a0SaEDo6NVc6yEf2qAGI30rn1eY8mU1DjfEdlHYlflCLy9LJJaVPL32piv
WdLfwCWRusN/2YrRPfzdqWFlp8tWPDg0On4Z/tZysk1txtUFmoCuLE3WW8+lFWGWUDcpMwfZN/fG
MxwvVwax12xFWSqctbyoJ4sntXYkBrq4FT724PWsmEY3yv+PbMo82ymWaAvCBqohvmpM9VCGJ3O7
d8iRCthQVGu5+QVoTxevfdhhUKB5tsqhdA+GEzxY4IhN7pRoosGVB84JG+N2REkx3aww8vH459B4
6Gvjau9aqgq6QXsKuYs36MaId7qzhXWzUPjld5hMtenn0xX6KlmGYpHjZxY85qzHUWyz/L1j1CPq
9g8nPgrloIwMjkXdYV0I4SMua3YKsqb2WvbGZbyB07zy7ZoGYNeRaG2UfGFiMJdS/HYSVbgPFzTV
J6H9yLSesbzizqOivcTo69/cuvOnZUJ7XpaaXodR4DwUa4zTwIV08ON8yExo+p4GOySaInqQ93zN
99vOpToV8SFtlp1xElByBWB4jDk3rPLJUD0H0wDz0UOJacJ5t/B3Dwots9AebInSAq2Atr1wfKdT
4TihJ2H6kz8APmJsJHErYr0FfeHs+/A9mDkXHpcoYZSowfSe/6Lg32Bdkl2/1nWkqx7P+1lreZuw
P6fLt4J62DjzqJGT223Ukyn5osAVSDJ9K8ds0tMpwEbhH96F4xz/gmSsHyB7hsMrW3jSdka/AY77
uePipqILw9mhwtZZnuR3waHZBqtSeSLtL/b/8h2EsQV0b7IOcGAbSaMw6U/U+paiSThgmJPN7gtS
9ycb3sfULPnJQZYeFYwCC5QOkeHgRF8Us9/z65lSsAP5U7A7hh2D7ef5Mxl6c3qtlhO5MdfEBVLo
aW5yB4DtK1g5j/L3e2ATXFbrl+75XdK0dtGewXeapsA7RsVCA+fOrLX9HQUzLGM9Y7fAHi8zB2sZ
bkYoccFzhwNKgSTkZZYpJ2afgkLG6tEDtS/7HRHcyYdvcFnS9AePMuSdpMy5gJUxyFcyY/NvGuxS
F4aQeYFEBd3VmsOtlQJc/9T7XtvrIEnTUj4w+vg/VQFtpQxQHfn+BtAj6udyOMvOTBeYFJqyDh1s
77RubNu1FUUEkEr0QK7+vMY77yggOTC9tD0sODZzalvgWr1OnbEKUD/dSec/4xiU8irHKuv604mk
mUZaP4xQmwcauE8jtJ5HoICRmUA2EHAtUe73wZJTjd9TL3F0GiFpv9DEIlqQcaW7wAwXg19+aDBb
JJOoF3cBs/Y2I2PxWK9kBW8VgSi65LG7JaQJXAYdJ2GIoR5z1grKIKCOAu8fR94LAk2ecASV7JKN
MDUIk7kvbyXX7Mpx4gmLXAfc0pwa8tcursUEuA7Jw1iTPobHQSS9OPB7xftYiROylsaDz/ntsVGa
rX7S6i62m2c7toCO7ox/qgzo4CykIVqg8U8gMWx+GIIdFRP3d8uhp2ZVZGA707ZwtlQpARmhjh0p
4rxVksxh8wwt4i5evNYk8fGjl4LJxG0ym2NupN6F4U/r2YRpXQ7sfpNpY2S3a4WmaLcnjj6FYYf5
fn1Zk5MUNsjRM5KvFT8QYGlV721+j1hFOKDhxE7jN2mv3vp1l49nvIqHzE2ROEi7kN+boR2RDDZF
MGiAVRtFJ+swrdZdRjB62NZRBjCYs1a4SDlD/3CnKbQSncaROnoLybvM5tvZE6XlcTSDauvcBkGK
OO90ODl8y+uuwgiUeGasYg+QU1MrOBe0gpC4NcDaQ1+j0AdGl1AUc+s+XdESH8HW07geE35qgGI+
fqCmMbx2rg/Ba2AP2ezZ5IBAXvV0dBso1n4eO3PHk860Y2tV6WhAO+tMSU87+0Z2LNWcdyu9lqgb
Dj8jMuBbEk4SJKHaf9vhs1a+7nbGifetkhMYu+blFBZulbzJkVO31+XOgGM5JuZ0c6HLm7wMsewJ
VzJGKalxo/zKlUIRB0Yod8BSvS/LnMfFXKORHf2deIiR4XmyGxrhSv5+5yST4R2i08mSPB+Du8nI
XOA89kebWXeTvbFE26ldED4n6iWSvN6ZB7K4efEz5Y+OMFs9tESirNSRWfIRTGH+Yv+bCRsrW95Z
6h3kfzsw3TxbkFIPHRmeILiZ47njk1pIXQlN3uCp5EnZ8+yBX2Skgi8eLx2GIsEgclXfupCz+xJO
V/0Cag5zQ/VROIztSN7uX4exp8kT/MXyOXZbYnrp4GQR4KwQSZJr19ur4Bb2EN2PPFQA4su5N8Wm
anaUXGZmyBa3RxjQybA3taItfX+L+eX1S0/cwwPaiC74fq/1TFJhwkBtD6hE2F+tQ7ZCp5hSMUiS
u6qfHqesnY1v7Vgr3fmwKISWzd7XDZnFxdQsIjSYjZIZk6QRmzJdtpxGAZzQNENp8XN2n0ZwPVwu
0VYsUhcLxKRD0Nbmwzm545LC5bV2yJTdouUKp/II/8eWG9w7Zy843eLad0HYxctQb71p3zv/cBpG
NPswWYcXG9jilnHb8EnBDDLrn3giMpN9hZBdWqqa4e9XX6zfPibk98GQaXIWw53fMJUszhX0PSqQ
wrMF+lVAgrWjcu76aUCciyRch+eXo4urwR4Wt8B8M9C0jJFCula5Hpk21n2I0NcjE2yiSUoVvlJo
57k+r9HkAEAmi6bfkhb2Mn/2k4ISzyymIZYXgEYZ1UUKO87//Ekl0Wkg5Nx+SfJEegCDdGZZIWmj
5aF2ts60kh8Bw3TWuBd+AyMPb9ys8s5Myq2uf94KWoMnxLtbYHPmrndH0I+1iOS7Ao3CaQyQ4efw
rdJL0LTTSdcg2uWJipbKk8c1yCcCIyRTeSsaJQlQ11v8I3pilqE5ZWoB2RG5+bXV0Hi6qo6vIXXj
+hVakOFY0IJRUw5a/hQWM/CuiRixgzmOGmojduJCH9ESBbX+pmwxjSnPGvj/6yDCxsFLwKigHOyY
GS7VPqBvSTUi/J4uKFZWRYRtsdWTLP9LGX8QXEN+kFKy32Ntw/j4JgYQnipJ5AMse39+5nv/UfVV
aFcUk6VfJs3uwSwo75AZ4bBAR8WmUx3h+4LtRdU1pLRl0bfnzuYX7N/AegIxfBwwwrA4y3j53YO3
FqCLhGCesjZ06lJL72hLCIfyKBGPqJjI+8r0eug0nOLq6Ge8lceq3cALmnVaOUjC7GSzFCGAn2NB
ZYpIpzvh+YvZoopg0tje5Gh3EStD7vaLlU6LsECcwGNNCaAHYksLPQDArHfK/9USAHTCg1/YwVX6
2nsCLhfwx05bF1IRNv9shqBkkGdXzOsr8+xMP3MLR1qlyEe+6ebpQPY5cy7x+ztWiM4ADBO4qzSg
wqfl68sjqXniTotnk8AnmjP3Q7pFKbhSnQQWT2jD2OmHZELqCDMKY/ieM8bMLPB4W6A6vpHJE7O2
GZGejVuMwm7JMxk9NszOXw1gzMlzzr3UgNoxFpjIfpvSB0UTcYakRltDMEnY8D8qqbl7gBpCwC2R
3W83n+r9kQXp4vKrnPLgqbv5C4tS9sPEph4JzpxNDZs5HpTkkiyREoDR7ntW5eiavYF3YPNo74FH
12TsuricZKI=
`protect end_protected
