`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Q3ir87Ss8Csv8JXx0hZxoXIMCIySGSVYtnqo+6umuqjo25mlLUPa83phb7YO7LBkId30dRHV2tD/
st0L5r1Dnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gBvadK2EP+ZGrCQXYhLJmScnocQn12Olgvqv/MLgbNyeUJmmh3evDnMj2yfMiS8n3RYit0KbAVqc
1k/Kj+BwrTL5d50bOqRsomX4+iHo3BrcmQ/GXnMz5dnFfvhw+W8Bv+iFw1vadySK+O8CQ3w4+Q5E
mZl8BVczP7v7l4BbabI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AS3fZ22RGlt6g33O6el4P9fgu84QpFBRzKGZmSwVYBjwn7fBnzBpX9QMhchCsxr+kvMq93A5rATx
+v8E4AhcM7/c3fTxq1DlHNyahEpWELGz3gW37NnQCol6nr5yGRWBsy+lKKJZbgWdzkPJ3OcQ9r3L
LOv13DeoAl+ZFygMlKNr7OlIEJDN2GV8qdyNhfB0XN6yCFPIctCMOWnxF3DM0/M1VeQdYYaxp5P2
FEdqXNaDQsa/j3WtsxllSsFAT9wcxOOVlm4hJ5QJH/gNUSBwTxMb8msfmGTfDxjelVZsBOSQ6maS
r+zVppQxDzTpuo7+WWUZ5pdjD/wZON8xQF37bQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G1bm/+r0gxybSLHEAtR3fEp5p2DQ5zMaS10rTZImokNE+g4y3u+4tC/GB7RusMxByiNv0mJZJg56
7c91js1nn7ciPatJuIPw6a/eQ+yQcqfHvdrbRwpwMJa9sQ2QsMbEHaLjJQoDbXgbAZC8O8UbS7kl
L9G7roOYQwOWCRC4T/U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hGKB//Gtat3sXJIkCT+zuaGKTsIsV86j0iAlfn3rYgX77lQNaIKWY5P5Vzmuys4C4eA2xo8syB9J
Cdjm5J8UiTllKRIr4gYPpep+3MtUUI9/Y1L9/q6G9mWWcu7yG/KU7o9sZATBMNdzujHLmEiI3xmk
DJes/V18hFrq/EeolbrCfFnynSZ2LDjkRZh6j+fLeeAzljhTXgOxqW+Lb1gThZGUcxTp5GYLmFkZ
+EO2hSnrv4tC6bBQYCa8kFL5T4XYwmsbV1nxlpYbuBrRh34vCbOToDsV98v1pbX7dmJNgGb6pB3y
moQ4QO/YHtO4RbPD+NBeX3bvGiShE3RHVDehKw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
/uj8S5Iz6cIhq9qE99qxTiUZim7wjGr8VUYGR6SXh2ISWq0AhGpmDFYEMe+WmlMTX/w5Q9wmzSrL
qonRpEXhR3Bby6BO4uJBbd+6NS6U8xyp3YbLEzYY8i2iJm+fLq1OkQ/PkEJBdVBj77ByOsyL1jdm
Yl1w/EtpUGgKfinyNXiNm7o1E8KPkBNreJWpOO9t4sL7Jn7NdhHsyLoNVZb7MBNrThL7g/b5q3mD
7E26LfzxLR0NlbKV50OdErMXAvT6spuaprferK8vMYTOhuBcdliAVTHhbZCjVMar2rIBHjiO280Z
2XuaEtgDJkzwe7uzclA1burXBZ+cTTmiH+16Ql/Xi588WecxvJd6rxGIdsFqVhTLbnkxROFcdMmH
ftUSy45ym7s3+xl/xnY2h/J2IGwOZ6SUSHZZJ8uFUz3XGtNRGhlI1j3o3h+QO3SH/WmvmmY1f+Qu
V27WQ/PhyvrtdFDSChQhJSkkiw8MAx+6Yabg3lQcGNYFGthhFPmS8NUXDHLPUI4d9T00tqTCRUVF
qWoLsVX93SFmR4XOqcVPAPVBy3KdXqHs5VtEBjyvywGW6x9qiU9hoCZsm3TdOc4kBIl2PAXDRKr2
vHcNZgsoSrvOcSHDdCsyCCtgj0jTO6PKlSfwzbWReDr8Hdbze7Bg8A3xHEXG7DP+a7pRVRYDaKFU
6rc3etPDWxS9UGDFwh32Yj9ZLLOBl9PhqgAivnUCWPA0P3olXKsRrywNi2Ewk62sxizCzA44TXln
mZQd35MwNo1/30VIX+F93f7LVo7n9r4duo3QiktKbZquLRR1XMhFXrDrFHnAlnepZcSjQddpdQHH
R44D2+RL2GT8dBnX2g7cVFBaGl3MLq4mZ3ZJX7z2E91NvDJBLzRRr7MhpdxeftPPxOrsNwV8FU8L
xbcBJURwRBOQbePv4gEUTTKsiKDCwoldoErLD0HcRYKRRzeManzx24CiOt8BLh72gAhmHf2nfgGX
Zhy7IVbCpXcK2SJUzBcHLKG4SU97qOZqM6FVhECvsP8N401tPmwrWw8uAMgkyGRSmmYH4I4y17Gu
9TtgVg7LJajex0xuN34XrfSjjRx8wtCbVDQdMiE1vpFZ/LOGltGmjES9pSNju9ofl+ytuBs8Q3jF
BSQQTuAkhH3SjHLsWjttRSSAjIU4FEPBPLTuoK6wWUxPaVQA8h8d8Qh4ko2zSxVeVyRQ+MRcW+fL
vDtLWMHn8VqOuifFaAt6MbTDsOccrFDSmiiw8DfcPSE1M2nAGAMDdZYKkhmI0NGlQucz7cIoLCqH
VbWzaJ6BKZvP9XLtp7k4fCGiqYLvd5+Mrdw5/e/1X7dxJ59MrjqRtMJ7wcnFdW+SwESxycVGootp
tNNofqegLvddTRka1j/RInl5dOOBTSdHtqzac1smRdrf9mlhk7lf/tumTeWitEfZcfeMXm90IRs/
Idpr5iPsgXP6Z8V2V5lcngOQIkTYBFb9ErdUzOwyX75QQvhoTgXo3Cq3ibtwQhzTwfmNLxRLviba
7emleRwwgCX/kLFswzN2cxPuU1lnfr063AUbfnfio+TsrBt7afJrQv/93c8hQKOUyZ5BpNoUzlSh
aP6SIoJKpALrSWtBC6swAijUwy62WtAV2UfLT4d5MciuVsLrY3obqwJZT2St2NeiZBt+qRdM8y3p
o6Ii52tloKqs/WgpwAxQKDVsZBkNlmcu1CrHTmYxuH8pO7i+xF4pW8n0/0deEbtDTDKbh/tdkj2+
g7AMNbI3q+6/ODb+Bv13gvJACd6BU/2IH2BqZL7G/N3TdpZF/uX3V2NbQB9tMhiYoI1/tnQbQcXI
Q83ff8ENzxm169yop75oHTWV1jq9aOT4XTpZtjyZqESle/B7QBMP1NyfSZyjZNoHiDpGbyHLcSol
cWsh/uAlob4UBJKN92hLczElhK/hnXWQOKQHePcvF2ta8EX7SPA0xYCjNcnoANGA71NP1ftIrYOU
nltzVmyBggLLRDxIih52XsXtCggf1iOkP9Tzm2k9zQ05b6QNeJvSbEoIJRDGbocl5qj8mIBDtlf7
P6AB5vJFhQd3mM7WwBP0hHXFAppz77rYORiLJYEHTH+okr08qoPvLJze1UHaStgaSspRO7I9u1vO
MBnJkH/KjftbnP464fltD1Q976K4vT4KkepG6ZimAG62Y/gZ9vmqeoWbo0pPfNK+78zBKTnqR91W
HLXr2n/+V7DeaASmHCOOaUrcIAqxNPo0OT5fuLt4ZJF5N/Ig/GMxZr9yLh2VH5Tpx0Tih+8S+32e
qUyN5omJxi/yRjjh1c3WvRq3Mq+WB+a2eZ0pvVs2crT9s6MWmasQcd2yuyXDq9ZfJeiT7mubGBNA
zNKWly3xVmsDMDcbxXR8wPjnvdyxja+x1HKzR6sLyaqRluj+CXxBw48wNbkvutkgQ0SSV1w/85rd
SJrBlBph2mRhE/fhXQC3M6AQWay4qGeMRUsJXRz5tkKKvGWpyXbIVj8JkCNXs3TioN4zt1GODBZC
oY2Jm4SYNdIbHZkDKOCaNcMsyPVWzc8sB1N5ouHIj2BHP6JxTkHkzOiPhs5FE1rRrrfLRsd1lC6C
7T9+J6pKwCHkY2PSvqnyS1B5ebr4VzbGibO7ejCa3TvpXlN7IDJWE2vSa0jt44NhZxGT2FRklRRo
WfHpMQ8xz0EMpV7f/dti57NygGOBHEFHUJKpJ6FzrTm19c0VAW4uFNaTJ7MNuCb5vnJ2ytwwZTay
CsmUrAM0kbBOZQfdUVhWMQUHpOJIj25ZFvSgvPV3+t+5yliv2nphLLp+4MlcFyQfejRg0xvWN+bt
B0Q93ZhfyU7JV0h7mhwbI7OdbJKVMBH/tykEdsRDj0b7GcxW+wY/mYcPUB1Jis73ELj1oXjSy5JD
lRq6Mvy46dA39cqqitLKk9BOX9Uwf8SdQN6V2mNIkagWvBtAYtuMnVZC6zk/qqAt6zQrPxWZArOz
fa+la9Ly3RVVqzjK48rT3ZTj3p0oEzEJMTf4xDprPjYZiv/Yv4mDWTpE1pEZ63NsgHZZXHSj43+1
2l5QGgGVo9zqBOJnPcsyCybeh9fnGGvsSlrSk61c3RyCQW0OVVDQnrUjOZ8Ks94YbvVeJgs2tvmY
GJUszxTAb1NSPfTGseyQaiRMhiiB28v3JT4uNIv9wuOJp6VvzSHM2qbBMyN/uaPXjQyi870iyL49
QcSMlvc3CiS79DVEwNE8i4T5Ke+rpP8imat+Y17ARvdx4WjVvv6PF5g5MTrRhT2KkhpkTDADbyiu
FOqeBVKM+Vq3AQyv9v3xtgsjMzXtXDe94h0+jmxC90S5luGE41O8ymh/8y/yVRlK2NRoJcg4XDlB
tm63UtwWC477Os6BwpUZWhzI3mdP7LyjAkinaraURQqYQcDKrVbdpcdwBKTU/ZhhHxOdqx3fDSz3
cZeHtkHUwij7tc2B6BCB52eeJRxETwGAbU2a2f9PPwnufczGkWIfiTL8tbeSsKzuJ8B+K2bzeMEX
G2kQakN693X0vsCNBZrm3ARSzWZLYL7ElP3TeRd5nrJAeDeOsi/c0946SV9o9TzcjXoYPnwXaIQD
63+I0VIi+wCH6Znk9PzVFmRiSo0qslr7MWO8ENFFnQIBAu7gB+dqpzCm64iUtnpCb4RhdncS7hke
DnS4pDhp2fE5X3uKHdqRjizqKSaLZs0+CjAhz73OF4UEOb0NbL65/z8Sm45QYtmVCL0KjpB3C5sa
1Zoy9F9IoTn+cDBb8BrRQF2CGi7A8PCVsMvhA8sL2JZC0D67TTsYdH8+D8/VgQBqLKJVE4EYBswS
1SDZgOZSfPxoyYMSbN/epL2MXKedpqumLgoyzAJCFAaqIOxZg5GIiO3rgrvA0m1h2EMODjep8wrI
ESpmgW/XRbPZcUP8vcQFE57UwhupEpMmJw78syICfnEeSUYnaNY+Rt+m9QiDa5EzOaozf0zDX8af
tqchPuoVcXiW7NcxN8YoYyyD6WJmMr1aU6jANmS1mWEvd2uV6TvRepJftAhY7MGCo4I8aPN2KP0l
qqxFDAP8171QMQvpEX7DI0sYgpdm3fxBFMUurXjTkup98fUl77/u/x8nT0G7aZjwS6Ze/OkN4JxA
rQCTakOua7Jb0sT456XG1cN3coKUz0W7egesPHNb4APVQe5SDKjp/FwA+jDP8rzyVt/8cH7W7dAv
ALUZmDPrF4ihq8O5XmlNa3OO9Yb4tW/Hsat4o7du1WBGzYnZGIsF7j6eeVlACt+FOR9mf8LT3ZdK
YM7zP+SSe74PptPHYYfNmCpY1CeYLGlEgEpOLf7I6zr6KgBpG4BGPlBI5czJdBGLRfKesBi1tgOT
YEOvyL05PH4wO2Qn9nk5/nlayGi5plXcDMXNf+NU+rzCNZETC8evZx6X3ouA272QozFo0WZ2set5
neHYXOkgwBCd6eMiWH0d6RIPTg+1qG1sFGTziYcvOZnSqeMIARwl1eHpgpOPBTcefuTVxrp33wZL
4niqhDaZ9kQniH5ZnY55GNxlGJVQUBhV9p8G+Jd1yDOG1hejQXfA1HcB51Rx91y+acbC+F2V6mf2
31cn4rlYYRnlWzeo61H9U1NeiCF6L97uNTzRmkENkhhtV9aBYCOuPMBP5tFnfw2CXs2ttTvmlAzE
rUHmsNpj0PHwgir/EtcHvJOqSJfcUJyT+yup1QgqmfsMp5FzwPyxrv4cOPOeU8PpwWxMySJ28YNO
0R3lUl//tJrO8pOlOzGIGOwBY6f4LdgF2HEpFFL5Sf+5mT6fY04vL3XOM++QiQ5ePx1qM9EUZM0L
T9SG2xYpq+iR//kTWZ1LTHn1u1vKIdip61lqgjfDbdRJiAgq0UV4Dpc32n8+R8FeWYy9RMf6yGO4
P7ASjMm4zMVp/rBT065zOKYeICb2U+AJF/1JP9Vg4F5Loth5IQf6EhKJjLXPZlIJFdOwfjMEKNen
45Zc2bAkmToaLQ2o1ps0OfH00UbazeFjWk9mlrE5MQAElvpYHdIVKttX/OcQyZ1bK+uNc7f90f+3
xt3oKmsEb6/fPr4GGFa7041R/IA3f2xq8IeeZVQZh5KuBVHcvqJ1GB8Gen+kJs8mkm+fxF9hTue+
J6fjNU/Gm+QoPX1wt2kGDN1Atr4kArXpTSQOwtcNlpjb33aCElRVpEREoq6X8/Ix//OdE0+mikxp
heV9ZB/k7RYYg8bJtjJUKMyL29iSd2XGnKA2NOAo8Zia7pi+CQWDiVksrSVxY/eUnHtAcLujUx3M
ACsNH/hsf72EZGOdnLUcmhQJY4d9xz/7btX8OoDPEf/XpHKmKYFl+85VNVfEewrvk0zrd8/daXr0
jO/n9KtWjdzXyLhhMxA41/8PlLD19NJTY+UdA0wxHblvvrzsgc7zGsRVXFM/kVtiu3pF5dKpw1Im
QHvro+ivwT7sJuZ6pyMC7L1iX9q4p7aH1lXcZCsAnnAZxvkGQSpLKz6JrHph6I7R3HLyNGJm95c4
BWMWVFGDh7YDnZSxauyreu8OtNpVE+Uh33hPiwxs9I9UP5mY0BWYud7x7dhbBSGdpbNoMYzARC7V
W8QkZPQhwzgudChSuiEiZ44iR/7GSVdBw062eI7/jOqrGrBVluyut/6hy0Cee4FNrZ6ImOyTltgY
+s6xzwj4TFNN/1AJJs3fT0WwZGCDl5F2iJUTju4bRzHTcr6pGYc+qkGK4Ot5jYtGaPdbLWfhSilt
8blqosmq0eSS3w1TunyteS9RVeNhdOaVIS/PsChLlEnGah7HoBR5uT7XdvQYRG2vdB7Zglc62Ajd
uz+APApkUZjwEO2smZQDCsg4xjo9PFaSvDrlaUJh9W8xe82/kQtu/fmIlH1vn0qBxoWIOJts+O8g
bg25uIhsh/mln8zpl3AZo4Xq6OaZObIhTvpWroQf3TQx+Z9lJ6uA9J47zPigCeHbrZY6CSWEn1CG
KYvVpKys/22WtRS19tqE3cs59BgoBiUWpJBQ7GiXSsFPfMEhx1nnEKo1DThzwRDsxhjNoga/gkig
rg1sBHnLoe9uQvQDp/AYXqdrWfHcw7UTFAuXpxwM9f5yBRF/gE/swvnkwQTbfcwB0EtsJ6usfL9H
bcv91GgPrGHYPGhEW97NTf3A+MI9wjxj93MRQyPGq8BM4vIsZaZylkEugo4rJK+of9//75jtbVe9
Nrj3HtbhU7g47qDz0N1nnSrpPo2ALIx8ink1HzL2qAd8nE0qOKd3qJTn5Ccqt4q/YcsXTK7FNCKu
wC9w6JLjreixqNKW/zHxwfIydAHY29lTR6jYOmbfhTYpUi0K1W8RLdlAZ/q6NE1k1TQXoio4ba4u
8jv9YQ2z6gY3hdICho+P5omU6tTKj2jAEAKyrzUoqaPOo2E7ruADsUM5hFVMKyusVWgpBW52NI65
xRNDxyY/dFzzjHUFPk7O4XaFLKIJ+SZSwyD825icfPTazVNCE0LNAdDFI9AW/K7mMsK0YK25GXUh
NAkySBRgiQACg3VgR7fF4rnkP++oXcB3maV+ThakLXThLLrIPPjtI8xNbactgXmctfVscU+4Z2BR
AmDNMXmVO8xfbZMQ+DZJPO6GW6R3F4m0aNGmoWjf8HVVlGvdkbyqEwjDJbqapOulpC1BWXyLwn88
Y4P3UF8uU3jYGFrirprZYlpIbkZgGvct/3NiDhnxu2wxvrAUVkaYhvAnkbH7jbggqQLtb21r2756
OXOAy7UCeqsNBXlpjPvMrNeLvUZ0OViaEp3481H4JY1fwCMvNmXpc7PwFzU3CZXWdYb8KwfTZB/S
dqolF/2x6GgL+2BdFAz1qoFBWIzVuCF85LNTp25V/eXdv2jjpb/WNNt4BJEwjCLN2DVIv4z/2c0R
3vCN1pnblWEq0AjSLWIt93NMEstiWdgTgMdL8DBcgLqmvfiiGMjEUylWy0KV7vxGyN2xNi88zL2W
l9YdyR9Ekw92yR9uMQD+o00reDS/wOJYYhG5JiwN6WxVc1PXIVKSECkaxhP1xM6r9ER5qbzL3IC0
aCm4+DAvA3DKyarCrO82g1ZzOPjA2JXksuqxWFO4xc7ZDo+Pa1igIFILtbD1dPGgDd9jDRd8ncmG
gD+Kw2XRxPSecNHLjmBlzJ8LFCSiuTmD3Fm1KrUX/tUcm3O83bRIlT1ml6/F6H7g9RHcwoHas6Ja
mdtPhlIZR44Adezd4sL6lt37ugNn93mOeyr/hYJ7rlsE4X67BBcZxP4xvcJ86PCpn9rg63UD4gGI
ewGLixYd0wuQ++WPYeX9qdbphBXyyDz18fBrtgBcj7ZFZhhYYEFTGGGod5XHdoEAi2blDm/xGZow
xaPfYX0ivdOjhl/3R93/uUHpsw3ZFxFZdob7g0uAEYWg2zG1otWuubIeSlyiPBd+o8RQEsJwbRmh
zHhfVH4TSdIbmHiJcHiQhAXTjmTlyjXzCuslmeNAILUlKitvT0PZctanME7bzBkETJvvCl9DFOh7
GtCoiafc52tAroPQGXWoegSgakOw5lYZaIE8ot3TCsKLAXfFcK4DXX2FWUrvZ8XVrZuJt+LVSIEx
RGCfYC6qDRA1YwRLcJJ8tryIvDF9bM2GdSBxVMoyLW7Hq2fCAt67pV+U6BIe9LjpgMcL8uqYfwh2
s0h3zEpzkKl2QkpsEUvDdOyJ0vUwrf3aFhW4hN+FwcF9MzqD6o0UT3qLtELREntckqwIJ3DtzOp5
VpyU/dDi8G8KqsA5V0tjQlcCd3hfHQPoINuN/FZN/Fbk+mx/Vqkw9HHdwwF4LtcwDACoHN0bAH1p
+H6lnSEajcnC9jpu0/Kf1h7e2P9ByhlbF33xF1YTGvARC9sw3LlxLmTeX1fUBpz+SxJXMl1nf2Yb
thmoRVhIOnDdgx5KkOWetZMDYm05cnJUNlfcPfZvDnSSBhmuVMYYUcMqc2/joSzpqMZPyMPrJpa5
r3/Dv+Vb7SHxEh7Nyx54V3L/YonV5/i8D0cjGVxqv5GaTsWitde6czKQ1EOD2MSPrKpSqouvWFVU
8Lrl7SxzhjoWmE4m003FBX7byEN2j0tNe3pzvw5jWBmYdR9ICPFHhwABGpaVSrpRiAGQCQSWLz+d
/Re7wkUHauP+qDY522izzr4OUubHsu0YDyStTW/qtRcXoE+IS2GvLw7JVkEjJGCz5MWiPOFTXyy0
OlviHA8Z72Abh0qW5FH/FP+R28flffwkDk8xOyM1KetsZleVAlAg+YnMP0xwnyxPwIU/J0V7b+OF
pfL1DByykbYJVCxFSd1JyzNkrQQKyPLXxqo57Y10RG0w+NL29x6M5UkTsrBK0BYIAZ50KZn5KF1O
GdbpyOCCO1WYsEK+9o0kAhlWya8h/g/M2H34ef6Xrs8Ve5usy01ICz8gXGYzAQ2O1Kur8LU5mSwp
IWtADoVq7VtlRL0lVVjZnnMHzlIicsH5OCKBWHGSO72hg4WPUfz885cArQPoaWa8Hml+1Sbad/3G
Nn7NdwdGEmosx2yTpLsX07UQsjowCe0CP6C70UFFsphz7egDBKKfPNaaE/Ryx5uRZhpU3japGecT
HYUniYzrzZxx08Fxu2pwjitvgRSCNrFMJhvqksOTK9rtDgL3CY2MwVZv+eKTUuvzpXmR5tEu6J1N
aQiEhAb06vnu9J8bYrdI5S2lFOcoavPXMPVPBHEJCz+iWwJt4DqZY46bZr62p0cPk7R2N57O5MsB
3G0oBRTVCimZtszuW3val2JFe98Ylen/lj02c/uAE8O4Vykd9jdOvHqCaVam+/cBHuML7HKmb2F6
0nY0IA6FXXU3Ms+vxruWGX7F4ifhvOL8eZl5uUoX0D9R6X1vNG8gd+odtrDQyaV3bmT5EhsQUYJR
36F3bctqgpYquQlX7nygnW1pmfQxBTXxfnFrRS28nYxcmAnOwAJG/uEeHWAGIvwg37Qm83AMgmT2
xZA0FQdw1dohjtCg3oO8RYM1Wz3qw/Ju7TBdlXQmeHOjKoR5DscdDRb14adB/HChFt59ofUb7wrN
F+C3lT6sSNl+7pzfkFOHy62PJX4PiVPGZcgSooUum5uBrHJfTmHxNcz+ZitJChm31ALzMD3UUYic
Zpd9w9T9I3t8KtG7wvUYrA3lTHB1VvJzDZZ3D0caUt3v6CW9Mpaj69zGGt6jCU9TO/5mspRU4+4W
c7W7BG0O4p6YbmaAOEU6cgyQDqGfaMVF+VwWmpRHMkkiuDWEC89gbqZXw15vz9Ese9ze1pAE+Dvg
6qhjNd1rLxYY7BgMfgBl+FTX+KV2BfM7sS8waIrDNUz7DbCqpPBf3btzldtOmueCm9CID+A2I9SU
LfFEGLsODODSy+rRBQNCYck2yzoVd8jntXH94Vcael4+dywcPEiBr76DyorLxSqb0ePBw6wTUEzo
qLq7qPW2h57Sf/QETXjXp3XRecXpnz/LGXwOpQT3/L+opa6aVD1ph0uauL4V4m8e4O7rmoJP4eQD
BKOJRhaAWN0NC8frcLZq+QaQEQ9wMtmzaKhRxD0ttP20iivd+KBmcjk8iNOKbtC+uMwAEHHcsGQW
NBcI7TZBU0vxMy6YXsDOY8HXHd6WskJ4+OQbP1h8pMPbdPNGmKcQD9HL6cP694aQ473U7+KlWBO+
7bp9egTaMrcQ9+8gC9jVS/52CKMniejuRASUyLcvItaxxf2XfW1Dh2Dhfp1kYua2+6VGww746mhK
yHOQZ7GlNKxrRVijdGQ6EY2WTntM+bdFZCeX0YhRxfZRkrkJ2OZ2w6tyVndlkZb3eG7XacRxje9b
26m3Qpu1oPLTOT/lNrebUDG9IZlCEmHY4eN1UAw+DayM3h3NARIznRlYIsC2XLCjOUZBDWdRbmw1
+XnjQdvj+IILKekdyP/BBcarCHiHqUR5xEka7GqXKULY0pvfiKgzqLnUZ71DAOUdOB7XaFNFzjyM
2k7pruc/kYUUAWKM375WGr+AYCUJBqXw6smH+ZYj+GuKmVZMZ+tPaQ85fnlN+r1rLQdhHy6onLxr
wXH1VxYeS/5++iqa/7jkTKRF9UOaF2JMqhYKrMjjkDAXZT95beI5HiWQMdAA+tdwgpaGo6a6ZLbZ
44qMtj6MGw/QJm7XO6Hy9HsZLHdLqZ7vKQ/+ldylDpjTAuWKt066rORyCPkAoFMvHYWqWUdSPZwx
lYi98VyxWLIOL+HWqO27XxMX91Zm8zHvX34xJu61sfoG7CR1XzegxFQERJIc7cMR/TkGj/WzHqua
PqluyaO5lD1xFKpjBvCjVh36oOFRypvKgwK/Rqa7Zraes3k2JcBJlnwUzqVZSU2uk9zFeMF4ZEWD
DebjQaF3aqARm/aHmvcj29BwD37KQdW5H2ng5n8DNPSZp8zDZ+Dzj0bHpGkiAsjzFihFMp+B78/h
/0jeNnxpU5upuovvLfcH6UfgBS/CK7lMcHY4lwq8O2X/Aa4zxcdiH+XxzBEgOjVOJ3ox8AuJHfyP
2hroRGjYU3EbfqzEGrSXsI3d3MbVrSvxE7R/otUO6rbJ+nzt4ZRyHuKkPWiPZvL6ryeerpSxm1Bp
ltAXNYtvMl8RI2tvaSUkWmYsNvgQQo5ZMw++AdF9os10O11RdLJyv3IDGwo+22sXJNuU/4U8SCRt
EutAla3PAFrE6aMoRlmJ+hfq7rjVtoxUu2BrP1VoU6W6weqICXU2dA7F6YRMG1QliUWaF2h4F2s2
T4T2TTYiX6VaqAoF9v4iiDv4YmmIquNDvzkrwz7vO3u4yg8tR/VVNT2b2uVarZQgjf7lyu6S2MYe
m2W/3LpWzfITwOJX+DHm1XuqKAhFbEfb5euYIaGX5eADqiTfSCHEUSJcOm5Uejs2u7vWdl7irlAK
LBumHGHg181oV1AwXFXCQVU1bDFBxO0mirF1gnMCo2VVY+LbnFUlzVb8pC7ofrz69xctaABohnsU
3RYh5BoO0+iL7cMcjO87DgPc5a9XbXa80HS+ICZZWLC6HZWhjHea0N86+j8udwxLs9CX4Y7ALhrg
uXqR+iCBlM5LW2Ihf/tm2nv417BnINo2tc8NdYDq7GSoAQM0muxrJ09S7SMxSGNJT/1yXPBlFR6X
AaOPs7e90AY53HrtFroWcgUSWk7SZEvmYgaC8Q+t/22OGbCkH9jMtq3/XWL1+Jvn5L9mxawxcKkX
EQxIHNqHpprQG8GTzuxzGSfrtbXIvo40tj36pZeI9RDTqDmZwSe3zyLTgpE0YhkZcy+ed17vnYlI
dJSodDmDLw7t2pAg1aYf8wZHdRNtAp5xhjJ77sMAJf0L92ejnVV5fqPrP7gIsIEHq+l5Hsk8fFkU
Yg40WNIno4V5sdccgxCDPZ0YSL/0ESd+4SvK9BtlZxR01bCgMnh5+zkAZmD/A1SvUTrkzX4R4L+q
RYiXnmJ4+dlqd2voCThmfluIrEFrxBlYQWbcuCmygqzKKcF1Y5yyCZwX37GXbzZyGEuF4bTg3T0U
3JBMqSRUXsQ1WSisDv2e3lnb6C2UbgDhc0ejEENxs853mN/XrHOvdWkDNckdxRTNPJxgr5fRc3ba
Qb4HedeWSlTS89NDIiMXxqY8DVVprlg24HVA7/DR1NiKwaz7fCdZtZUmDEmPn/jhfxccf/H9lbjS
MgcCFuk9WVqgeAsdztRrETqt4noAFesUfxMvDR8hdCb4IZX0wKLr+BL+h9K3tsnivuQaf2vwQxkp
n/c4jtteC/5hpeVEQp//UahQ+hotvl2ZhbqAsHcnc08aNBDAG3sZlgV38wYruWd38oGtiFA5tFpR
I0Cha/q3u+uvyybReZWiKvnx1PbWJTLRJUK5CcrZLejp0NWnHHOpcWfpsJJocNEIaFPXvghFqm79
6CVjCqDsElAGDISu+ID/Af7Pdyogr0gvdGTlLgIT3p81x69xFlrmURjlutf106xyHaELlFMC+RKM
Aha2be/AsYJutMDaIJOTOCMeFdJFySuJKwVLYKylv14yOqNGSFBP1gM+Hw5c8bxvHvIRynRVwVp2
UFFzGgqtDA91ClYaFHIQZ18v6x7PoBeiUptX2kLqqplzVp1Io80HPqt6c3gMa4AHxqTfhy4p9tsf
1CMDIzess55gjlWWD15oRblEo0DiVe7WeAJRmq6u06o8281OIfegXUxTIXWYD07rhRYPpF5WKF9O
R+xoCUZTkxb6VppIlVWpkm94Rh7YsszYqU8LdjDRZkzJb5Ez1gB3u81MLqVNWQNhCkvPmXGH7nMc
XHF1eXE26uhV/9/pnde+wGjID8aTaLW0Fy3UZ9u4KS1jJakwEwLcZsbWXi6NpsjNe1p2avR4Hm9x
Nyqxr2TRzgJbdtCJ8p9R5kcCHjSvwIbGP7jrejIHvts0bEjmP9J53eF8iTiqHU9C7J+TuWOlqH0z
9E0XsyO9rTEIvI3lIrz02C+prcTkEDNKD+GAlOwd1dLPP1nbPLSQTUN2IxFmNfV7Vo2wQVV6iPF9
Vc/Tt6Xvu4fHB5WFddtAlAfd3Id7EIk0mDHgVZV0RsleQbs7pLB7UJQ9KxaWv96S0jB4mbbjR6u6
7zjGKzd5XXCF2RPydKZ3hwPSU+8fe7U8+vf25DR/xmOae01XCKmNP/9SBc2T67BRRfiWSxNCTIow
mThxQSy+/xH7f+SksoYwAY5Z6t54EqAKAqmpNX3jyQZMeE29D0Kl2ap1K+4hkHRs62pCrmGminrK
eOHOm11CrPvoOplj6Tly51h8/sv+sFKi43OzQp/+pkoMzXYtuuHTRrhAWCHf/j5bYD62v1P5aFR9
7tCJUwOvh/Wjk+ycCoj3IjZ0QqGXaFvvS2947uOBSKkfHiih4P409adDQYg27osYKK2XOVHll4Fu
oWd6ASjyx8xqx1Wfxv+KTXTSKb6r9CzRDcg5AO0pkzzckMxOf5PMsWEddETmzqmqHrtKAp5d/FaP
sum8riujwLx5mXgGsnH6Ch1IeAlW9A9M+WBqtn85C6MAnCdOP1lY2ZHgHVUwu3LX40leuzA6DmmM
1AyNyyiUKk7lSWKxMKa0AT+wd+n9p7tn41khqC7+KzAEgqLScbZVE4+ieIbjdK56xtxeoEoVZfRM
zwKyInxeczWKBee80jPCYFOT+nd4B6GIL1STu+Poy52NvvjU4wdy8Ok7aT4F+EMCBVn6+RZdExxv
+9sWB06m29mwzK5gu6+7ZEzCgOrbRUU19Or3qdAXfSrk+mFTamcwznh/QnwaHOyq8o/a3JI3Oz3l
LOj74zHKfZxa2Qzxv5AovrN9d74OTb9lHQaEGcDhzJ9UhgzZHr0oCeXbX0ik6jcE/8CCVQvN0Off
Pl9Lgfe/2qyggCRp6KiT7fOMm9OoV8eUJQ0UQTOrO3JlBByHy9TNV7RcxbzHPG8Di9ciQLJe5dQX
pzD3AKtL6dIaIF9LUrdaQTr3LLkJl/CyZ90f1LOAAq9brcm+Vy9O8iggQAnJ8lLNmrxbyDUlyFC7
SlUzIEXtswx+UhrJYzh55137Yd14BXp+UIdmZy4HCVU+4TXIlPiNySEaRHICnuz4vN9hozXL6b8U
gtCFzwjDMkv7WoMwmw543u0tTn5BdLRWSsqNYK2f6gv+uk3UQIz16lgP5bKpnQy7yyLUpPJh8nCo
I6hWnMr5xFTwKHfYneA8KbacIcz5ly4YzygdV7dJDs8dyftes4pqa4406qFPCgHWSMgkPJYJvZzp
/f9yj031lUmn1YP8CFXG9H95qhazlF6oviiXadQzu1I4sx9d3BEkA8zoDjNrfdm9sQ8GFaUozEyC
4hXF6OLLs9jSuIwMM7OKrj62pSoH7SGyHdkFqKXAPh7y6JLNgattpR0zUPCNuzEAaXI9TenW9TBO
0tGnx5QF/6wwq57ZAb2/MkmZaWXZ37MePaRQYqe8A5DLR3a18YA/5GfHdZiJ3CLLe49UBshckAOm
dKNoLdsgRq1uID6h9mowyEX9tGItxVIDqfyKWPqld1aCb9EuxQr2+qCPL29/QsUwx78kZxS7Lyns
b0V0d2RVXz/6gmI0//UCejxHwGOWVDnug4a8/UhDyR6iHIQeUbJfN4qIKaZzZ1S5IgpkJYU7jKSh
2ipUozhlZRsyyWaQqAk8X2ZvmYIcgpEebljMP0FKaU1uicTOd+Q95v/2kRdTnn+R4jhtepJs+Mif
RPngkJjM4gkGy16szdy2IsjyhwLXNC8wE8nUDnUTHcb/RwL7bV2tdjS5URoUfhGNpxeDwijXM2Lf
JeKdxF2siMXwboq4vC/b0mqaTYzsA2BdDYNKjZL/FsVkWfxOryrS22/O95nS185y8hmNqcu1F34R
fqvhELAviKqpwUmYLOQEUe9Ca3uNcV1W+215cLVLal3ErZM9gnrltTmoy4YLit0+ZLj6TP10XFkj
ojKCMgxjayg1DHZ2EZXhPLfCwSyA2MkVomSSqeOygvOfpCJXZizYUNRkt3D4i1kp2QNtru8F8acD
0+R6Yv/W57JnED4nWnQzD1yojNjeehIclY9ar4mZM7S0ZQKdgI3sv5CVdzxWxjnGlOOTknQurype
5Qe81BNcMWhykVs7wAQkbuVq6LHHYgEukTf/fU78oFc0bLbnF9F6vQYxl5i5k1iYQd62Gf4OTvpJ
TBN4l79e+MNlg7PIQUGOKmIu0QKmtucuBA8Ir9WHzN7/rttaFQAjOD4X2mp227uBxthsH/H88ra9
entSXBDGcsPgWwG1imdd3B4dYc067jq+7QHT33kREnkDvHjGDflAzICRm+o7a18BG0SV/9z3AcrI
+t52JiDk063BNTKmhrsZXUfoHymsqTFtLxL0l6aMG6czSoM5gGkzrFxyyI0gQ2wRucOs4GItDYlt
UpyGmeWAJPWVVX5zh2gXygn9y0h+rsVYwwgjWn5Sqtem265Uu/yyXGpDJv/zxyjsZOHGwBvk/z9K
0UBht1CoelfDEnY7CIvigSwLUZVgvwZeStTC1ouFK6ZGwx3TTmLIRVs7ggzZ06qYOoXbFMhYpWuE
HP52S4r7xtx5wzzMjqBm1SCxpnACsz6oMPaoX+XUy3D+S0Z1IgCgXgfpB2jNGn0TJtTsHrxg1lLI
+6UPoZn6ycDZYM7y9Xu/Rr2yH4ATu+wKCBtztEsXQq5RNwO//qN/9D/gPZeMzjKVbwS35ukqBjTr
L4ViE0H74FLZtyV5s5GHSyStU08WQ3LtAzOSePfYTIbnDOyz/9NqXaFuViTJvLGW2F6+8qqBFCcu
cJk+Gk8XLUr0lwbj7Ntk99/N5LJZN3+bxTuCTuFuV2yPHPDe9nfYHu+pM4sDForBGh1iCmMKwjCf
dAJfKfLKClvjmPkBdnmpLaW6af1HaikhWgGHErWuy0Q/RHLXx/jIpEE2EPj4BDMsBF9Ibqy/PBkk
3APMRnvBTgTSLSYrz1qVH3MuB6p+TuX1OPIMOuf5Hju7LohJrIYfL1nAlxlJxbhUwElUD8S5NIVy
Sd7JLlTiCsJSymD3fjm9CXWPlGdLcBWqRuf4f3JP/S7vSjQHvfsujrUl0vGhB8sz4T4mtpf+I+bJ
VIPMdMlACfphYTakCvwCRNyKka5BIkiJUwpfhqqD3Tw48DT9NtpRL/jwBMB0/Wh0YBq2fUC4pvZI
jiEIEOtsMQBGQppzlqdadAVafOoQ02Yr8qSFYXxmM6/jfqBeGfN3pAgP9n7l5UIHmk5ljL9TArr1
HhKI/o2Iup1JSvkYyEx9EzFosrtqwMIjsZiGvqCEYHAm5FaTFQlvCEZZvY5FMEemTdc+HfOt4Ub3
MzCngwkSMGW7H7mjut1WHb+laKG9d3PfWi6pKyafsVSt1lZu9nOCOHCNjIgQcN5Lh2SCkId9ekKH
TVZD7piGHDzb8X9x27tmqoaI98CPispH8gTp5Y2BrsBw3scEfci23/ApPYmYFxzSdX1e+AYpNJMz
6ayUxiwFBENT6k2hRfzA6M0YoXfLwpGvENIu+BDJGkA0A9URdbUN7sxiQSZr9uaObAUkuCc0OIXg
pF2rdxfS1ErLAFSIw8zVWidQSqcK36H9y9p8aehRyVi6Pp0hqWXXpOMHe759qsAtd96r2anS44pu
PPA3mnDTvPXn3iDlhECrnQtb8KI6U8GTk0GCrX8MprTV4e0bsloT6WbCpRV52I4vBAoX+Km3R/Au
a96NJP1bm2kfVt0v4xy4WWXhv9l8WM8/bPjFmRYaNiIHtKoLiwf8EofCBwN5AWat2lIom2vjiMmu
s4bHYAHEq/0sznMbFrhPBk/ipviAsOufBNBJBK2KC2n4YzFBiWC+xki/xqyX6ExZR/Yr17bAcBU5
3SX6twwsvz+s064JC/Phglgw6dlmextnfCf8Ij1K3DjAEb+JuCMGz9AeBLF0zLuqcY1BRhptS2Xc
NHASOi6Y/MRfzi5sBGSmjI7eqmmrZY/TUkl4Fmd6P9Y/09aVbW3L3UneSFD9c4Q0ojFEnNI9pvSY
HyCo/CzpKaKpTGIWlGO4RiE7L/U+JNWG+bCKUIXXsxLwU7Bmq5pHso6aIMPjfQtCMfcycubSdkiy
8/KZm1avb0uYQxOtEdqUcJG3MTFzG5iTOtfmX2dSJiCSbTBn9ApedXe7W1s4qWxZf+vYm6AqZLrA
NX30LpiUIAmI0KTUGC2MiXvZ+IDzq+UwN/WaWWoyfYC/lYEfnKDYaKk9ipfozVVjP5aIMPa8Kd6s
kfeFIR5/lFP6K6XqyRnTumipHsWgSJgGLNuOCrwkL4D0H/xvhkDfnFn/VhhaRlLZlc4kjLD11WMr
AVhXcUuD5N4c36O66eAI1ArngdOU4gGh/KkB+CyP9kwq1q1QMVg2t/vfTH7rIu6vxh/ql7sJXqEh
ByegyKpQGFXTBHK3nYMwuZyl0DC4GA3gVXK6Nw4xxeM4aTkfqGK8ojBLIsDr/B0gnA59/n3PSIBT
gR1O52KO9xtaYj+1v59OnsNhsL0aAOAn3tOxtr0IcC3uIpP+VXVS/bxN3ko8j9usvaReabbmSDba
z6Rho9wB8eOMpV2DJxnTfE+YyxogPieD2MofGAA8uKu1wrTJCfm8/Ti8wwciF/354kbSbNfDJinU
5vClWcrvPXdLnMU0jJwIisVdqCsi47p/6o5XyIdbxNGtE94rzc9JdLFuEgwfIRvrxdclHkQVx18h
tzs0osIJdIiycmKx0KY8Zroi9rNM5JWD0MPL0UdZbKajkoGC1VqYht8ML0B5e6pPom80ZyydFzdK
vHrwaQY1C3RBlgi9Avx8y/MMEANM98E5M3bIohS1onSGD8fl5bR2yugY1RO1MwolSVZtB+Ij9XIN
dn8IKJ5q78QuUeTTp4ImOUaPOtVIkRvYVHXsaKxlCQCX3/ogDuls8vCxPxJtThNVocfq6DPTAFrt
3hXKFQ7xAhXsfLBBcnjqzbeRiDdJWSDLKlyly1etY6PjlOt5Adv5sPuqiLpDez4+tDXpAFb3o8Ag
Y9FOztD22eyOqAPtz5Sb8Oeko1HxxzTGsUmwl7k6e+Tn0TEsxUEUxXaEnCQGIPSZzIrDDdmt+Scp
RawPKlmwd7NZauFmSbT4vOE1v/zSFW5EBe7VWQA4yU/ImhHw5ebJkKwFI2TuOLQ9mSpN4JWWmLMm
GRVg6UZyzURQINMygm1eDgDUlzaQ23X7ruAQF3945O4cDaa0sJ2/QmwoPRPjTVofexdP/had2OlI
+AGJZXM5/fessWMzfuRgWBA5XJrPRaH3ATDIq4xXg/vk2lRNDrcr1xV7TN6st8tBxRJgaAz/1j8S
FfRbWuWYgqqfYgPWcgnFOLRx477eTBtSjtSCbmeijsOFZxx9zdkZE2xA7d8F1T2NO/KuvSN2qKQY
K7MDXVRdfyX+KwcQu3oLpqItwGCXNZmaed8rHri1uaruzMnRDO4WIYqYV0NCZrDwVvM9bCLcM+tr
KX7dIbpez/INlvnqLuVtrcJJXmO7jLmCSWLGcImp2j234VPj/PcqObG0UJGbr52+xTM6VrWPp/xb
1XCON/uUt+RyDVH4HtVMqiSRlRirLvgn/D+tQwjiihWlTFe12vTVbBMan6rUwWcMLz+FkMvrJKCZ
Jj2hVQmL70hhUFwBrbPz4ywJTwsu8lD81BdLlYMRtiF6oVACOJ733yrPOGv0qJjJjqTNl3JCsap3
ekpEukLBHxMw9KShMNiGUewNtR3GKBQxjAsM7XKDoptxOnt+FCGY0Ii5wQZ8Rr5sPSrM+FzIzw9k
7ffjGyDVwHGhfFyWkaB9iqZvzr2N1Wg3bsVzpLiaORj5VVGhP/1UNtssSvfD3I9RQs/JzfSPiTad
0SC9yV6M2GsZJ09p/VR6nOS98ONrI3BdiIbHIi6U9NUV9HgD1RQmFEVR5U7wiVCFmTC/fSqpS5Jf
06AiPaQ6Oe8SGcP2rlRquTRo6CcZGLePMH8Cwnx72W9SeBuZBF8HXPy4etR2hvkikfokisDN5FkQ
12VT3bAWjYW+E5ZQ/S83kiOxRoraVXp/fYZ6473Ga3YkN1yIlop1QCIU6QXA4AY2+Jx/44KKOEuQ
g1JhuO4DFuAplZ20pfGusb/Thj4V3iwx3WUFtYq4pHMeCZGYXlTTNY1LlmQ/9+7ljrWG2DJUYKd7
BvBvMT0LRG06PpZuIVBA3EKNLP6yzKGEVw7J7z/HS5/nHknI/Mf4ZqQIm8B/xMhMfUhvBzFWIaaQ
bq3PQcNut16Sh160ioyomvxS2OYlJ0bWL18V28W0L5M2NahFSWCFBPh1opDZSPuuZwV1zb5b/9F9
ulGvJ8+BHt20hz9H6nTNCEGt1QEXi3fNrg1/OBSy2BYcSUM=
`protect end_protected
