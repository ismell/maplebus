`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Rg/jCkZDq9XQVwyvSkbqPwqMFiozVkiZkieuMtMKuUzk8VmX/hw0+TpO174TPuSM0PxlEAAU7uyO
M2w5Tvmo5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XJgaiZ2JCHgJBg+XEwt/F33XmnOujqpHsbUskmUyOGVJSI7mYo/c9fT0/lg9NVGxq9LVciIe8Qz4
FRbupGTwjfLhn5123C/LzAsSzOpojovOstGV3na+Q2CfMhy5dYGSLTD7DTNtzPOqavyAb4jg8PK7
DuWc5q8uJvyWlEy8zSc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OoNZPRZB+O4fgbakUis4WpylVoMHusJKW2Vo3VUF26dKiAA3KHLlWw0kPMUjPy3iY7ATZcLQc9O7
gDpj1ypq3PMp59Czp/vVO2KlAdsWxqoaguAtN5bxvlvIIaqYnUL8ObkK465CzCggFirukELOIGeM
N16ICCtV3G4/jRufHQUaB32JKIyL+vFJXeHDZOYo2tMWJd1UH2UMTj29lbZeUICN9ct0tvZNZwPt
nmGzyPfL2+YrLJWMyDLMPZ88nFIwCIGFmqQN+kBm+tj8AxN828wRSNMcxTrN2L4RAbblay6P/Igo
40vIxQj/AJ5BkG6IujbEKjOhmlsg37SpKhOCUw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ygfSZz89nx2cZ08Cn11X2l6ZPEPFoy7mnJvs5QPsfp5PuTE3eDifbnCnbYLfh4oeIGmZjBVuu/vL
KHWuDWOO18gq2IhC4izWCNGY9NDQlkD65ZjmB8olwT1MH5OKk9M7Ekjxvzu73c9+bMfXTcFqkRda
VUQbfvr+/yHIq3tZwAc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LtACBladVC/Rz+Sg3p6gvjJNipI4Irx3zczEaw1fYWqO/7wU0AWfK8D2fJgtmC7E5nLcbfly82Hn
yziSEM/t1IM6+ln1nEUQqg5S4Fdn8pzmmHXGbznzZ653thyBFn91GwDF2Ov/SFgobjytYWi24y2t
wYomaip+HABXxxtB6PWwxbI4IpaysmbI3+6j9qMU6JpJ1p5fNjoULvfnSIkws6KhVX/1+gl9hlpC
NVOBjx9vtF7I5P0l1erRivj5MWX8UWtY8RmaihKxAfRQuKwp5lKc4IqDT0Zp1cdQcLIKYipl4K60
oIIQxMNI3b2eTiYvlgcbNmv7gq0AaFSXUIdi5g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24176)
`protect data_block
4AsPia0gGzAB1RPpwqbgVWC1RQLAkT1Dj6aee9dQNzVuohevjiGGptQWNg81RavZDoSYk3bbCnd/
75A/b48ggiXFc7Mp3Ivmm0qjUX9BAYDZJHdh2bIpWo1AFwML2B9fbu5lxDGrHA73SNDTPK3lKBwN
V0KyOIQQvZRVjAEuDxelUnIxwqGHgLR6Z5Rv0LKWma+Rwa5EP99fSl7si02v3vv2HeUwvtSjFhg5
BJn9Q3ZdY7BVWM41obyuVVlgT3/xkhxEeqWr7UZHtwLaqogYSLlZRYHgteCMuuP3YAVSW4gJaOHX
v7kfSdIFyXktYJQ6IMrzpuw11iu4mqPvhg3FYo8AmZagnN3aD1oqcS1Ck5dhjQet3+OYBv0YbArt
pIZ8RFXEzljZr0R8hgMj+R1eMKIQAuYcw9Scncfj83ApIaQKyyeb5ucqhaRnsy0n1aPK60rr9tJl
LKhNheZVOi1VYDDXf5Mk7TtxL4vzg1a7or97rD2effihz863iPs8/kCSMu8baORjT9wfDS8Trk9N
txlFxEschgzO7CdFH8C3Cdz8Sa1qxyZee9nF0YU0dHTNC+kWLeEYshLH11oHNMiYMqn/VvMf6/8g
C9O8srBEVX0YCmIZaF68yfW3q5//BMKmE+Jbyv/ag8w+jvHE9+5c9RPZR6z92BanrzdhXyTiYsdw
ppzvPt+OgWRndmgQc2leG2vNXDrUh5nB4hJmjo4FLRoVUXrPAqpKP8734Sdi9kYMAycIPrO2UAhR
1DtACdY/vmfzF8hmxRoNDFeuutavFpJTJFWX/TcaJ/wCpRE6ZvoWM85dcgoQJJa1Ujiwk42rK7gH
4hCgP9dl6Z0V70GaWFNUNdA5QE7kyB3KE6OS26ABChjdFnAuUwvnTPJpvphVZPLxsCNeeLdU7FHV
plPG9+sNmjVJPWCFrrQsEUI0nWVxR/CvuNFoFgTQIO2xn9HdOhQ2ls/P3BOjmJkbcjJ9jfzOsbEv
bz9zEHNbyLvWPjSM6P/wX2tm1QVlVcF7GVwls9npm0DzsC6wg2dmgk+mXtwplbYdKhkmp0P/UloI
otUzEmxQx77zA64yZRdD6YRgv/7of2wo6dek9yElBbWxIxbFwgCN+4KGINwZlwjSGlFzTJ4tMDRk
UdbKm4Cm3bZ9wevJmGLhas2zO4IRYxG7LYigYxj/zmJUpT41+uzl5A0OlXHm5B+/DHCW3cg0Fr4e
AaAMIjlcqsRG1ObW9Pk79JevU3RNnEqQFNb7w2yEIF3WvJgIqUhMob0ugUb0zLqKKXGpSD0GfXst
9A/zpwVbbWjc2DTXXljJwhEFpmSSLlEDi0G2nGBX1cc313mDSN1iIFSc4wBbeVfr+lcsxrSiu6UX
2USwL6D5B2/O8KLzxZiVLolnhPj2Njrh65c63XjRXyFK+abDlJLZ15lOcA4N25AoK0CT4kOqzYQK
Od5BNfKCn/v2LC2z5518RWSqVn2IiKfp5qmFvRnZYfynERJoztTv1yg/+yqXklD8AUdrwoHo5mdk
9CFaAWJOkAJNll5VFkJg+FE59aiO1x5YbHnI6SQRsXfw9jtKQ3z2GrRwMX14v3BC+LRPuSEUXCd5
/r/Xm62O1F8+vGPZqqZW+tF/S4KJyHhmqsPv+HL1LTLu87H0MnX6QPod+qquDUJFsFz/LKaaZrip
qf/NrGtEyh00BO8pvKbMh8EarmIS9NMFrYuJpd+4HGcl8hTYcxKKAGeL1D0PX8oUeezoXOzl4RZk
4NTld0ediNXjyPW82Il8pCKodrKJpZk3Ot+i6s5zD8dIq6PoMOAQG38AEGLJM8s8mROOlxFSppVq
IoUQ1ZUek+lVz2HRp4QrMwawPnr5Cv13dmzHSdEqLOy6LFFUtOmrnbUgZ/uKYeOF4lc7IYoU+o1+
sbM5Jm7NF9gpZvIvMZfmMRQ/zqRoCRrNGntYEuhIm0RmqBNg+g9S4JII6vg7iQywVDRPW2br2BID
+Ziz6BSIkYAaBB0cBq5fBVHH9bCSvqW61WCIjtXy4jpwzeSBTsfng19jh5Pro3WVx88nTw5QFt4T
JESt5Apj5WenwZTclBQjumy6eoqmfdtsMLRJeUmlmlVodcdY4SOspmG22gS6M7s2b4IeU6VPc5az
z4yMEbmD3rdgqSwOMNAbORiGtG0lujfzIKUaiZ2loLGr+l/03HuzEg7nhckG0K7lyUffZVljdD6V
0FSeREx/RxLlEUGszM/TGKDCLmMIPtWopn9+HoQTuuIc8dKHgV4X1AOzSuZvS5aObrdfz3YcCH6C
XQubZORQ9OcWbgaUeXz3P00K7nOZ6vQiDVRCo+GWIfaP5+e49CQzH9qSaww/ogv/krLCZ8mWtcfg
SF27PROoGoouNF+OyJkdZO7W+SXg+mFDFsG/0lEwf+RGZIJRibwz1Hf+AYBY3p/u4xLvpbf7F0HI
dBy8TurTmH47CFaVIe7IrpiFDobrCQb+Xu5hOVbVb1TKTQS4CEUDHK0DIpSakx6m2b22RDdZPxr6
PdeI4UveNDl2e5y2OJjj91h8bZYx3xUmYxCpzGyc9GBw3642zZdTK72WRu8s4vvOnn4ecuuXeiYi
ts24qUV3oN0i2id/Nu70aTd1Si2r6gu8+PnmlxtdW8r6MCKGmPHltLljiu/q2x4kxktqbj2U/4oP
56cEMFXWu+4+AUkA8LbYvRAXBmOdy2NBPuEeKyx9MBX4nPBMbWOeUpsc4FZi1bQsnKZ/QjoofoLx
1f5O1vMlUceajAuMdjA8MVjGYP0Rg71v7zO0SXQ22g1+StKWW4fk22z878LMDxifNZAWC97OQ3C7
vvOZzkMlfjFT+HYAM91V6FPNFlygfKbTz47KCeYRcLo4rKBwmvFnwOHi6s9kMZNRFJKxaBed1lc9
HLXpoC1PG6HyGHTF/P1uAH5J3AhGQpzfw5rJKBmotl14+RPFkhCjK2SKDbfcIqp8QHCQEHfX8Wzs
o8C9mrLiE5mcXKY1z3KSMyWLN1Mp9uAcKA1QHBBwgSFGTAQoxNVaB8JqKTgky23Tc3ef42iLqE1J
sbkmBftXDdFKyOpNBGtuWYMzE8K2WjxRtV9hmVnLeQpHOHUJ1r4TYiDrRlnDM9jg52Imd7d512h2
xrDR3sBwYsI6ZuwIhES+XYut7T7R2Qn0IcPnzNto9O3REghTx6g42byEkvMqhxm0RLnZV2ADIX0I
6ySz9AMFEDbKV2g/ENSrSdAxldxmQqZyIQliciBCgZFjbuRjOBjw0gsYGI4RCj1SHysqTtum/MeV
8OCB2REn8gJS/bn3sKQuSqvbpuHsYX1qObkeyxq3y9updRZPfQlIXe4+88XsJzLetBw0qZiUSl15
E9sRSUGhOCTfdA8ES8dr/HnYOvKiK/ex4CaV6h7su/6B9rrWy9AEe/l08pBsKgdf082XBp6exo3u
enK+0zKe19sTxj3WCJ1Gf061rBtmhgdR4z1ys/cme2j++91ROE4Rnez3nTZGUk4CDpPoEqA7kWRY
KIbXWTScaBAzJkd9fqaojqC56JYNirfvE3ijuVZhnOhLpYO79omeSKLpMI313bIALdH0yKyzmmd9
x7JmEi9SE5cpw4ztS6O+dTrDICOZgftpx4wNLGm4Lj2oEHDKh9dqcQQc32gVtxBm9ssrclo65A0N
7FLzHEXo25PW4M4HSYzkao0XN34z8ITr/sKG61d0VBidEBW3M+sSVHHZgHQvYCR9XYW0KRVb3971
qXomjAjmsPAGORRo5R1FxONBnP0JqM+g4LyeZ2Q224hv8QIhq9WqAfevsgA8HIxdBxdA9vISq8ng
56pPAi+vVhQZyIZtQuEAZSYnZQ8gwlShBxbj6kiVB8W7G2BygbxYKz4YQpAS8aZRgTnnq46TP8bZ
9iOguwpVWfJH+j4jZpnkFXDSXW/Ccgjcv2H0inOIEo/uJnmG3Yg2wYgZ1qRAV2Uof/RCNgojtyq5
l7BTw7x7uUOtfUC8Rco2hSgEhNeIjGmb8yRv+3PrJ8ZnyTUyai/qV5nJRZ2q/cBeqTGlFGnHK2N5
pGFRIv8pIt4Ja5OfeZxK2UyC3TMphki/KbCfqs2SzWDDth+mf4QtXN5LyhF85TJhgfcFs+mDL/4W
0VHSfwS2btaYDklNFJbfHySiU8FU+fYc4h5ED2dSFH3alrIWvON0a4dXBXRVnOBDc/Z134HHV+UR
3/8z39VagULi2fv7CwM/YF0qKKk1/CerSze+kteuXuJDE5s21m6P3wlUGz73z5RNFcCF2yYCa7zm
QAiPKQdtD8pocA+xNUSX54qO1vLqu8RDzHYj4mnGelgqrkdmsbXFu6tluZVj8vP1bF0/wiM3jx2E
4FZue2IDJTTzBilWcgpANItrrYHuM5LfB7LAxF77RKiWXK7tYRVKt9je/ugvx3XuoUTes6uCedNy
KHZfha16d2QAcxJP1Khy55viyIDvQtuYSl6FITNPw1hBeX5CLbRstVpY5gnyBttN1+nAAx9v+aiZ
VQ1uGP3+A1Q9Ww4GTbrE8Oiprb43plYZz2gEJSWeoSi9ffOQYsvqNk2Z9rBAapncUVRuI0YMCh3x
Juo7a2fpflU7X2iw9eIu1jdKqEMAQ6bMSmHqL3e86bPgox8Xrea19fxBjbL8HMzVCsSeXvUIv5Cx
1ppJfxCaTpcSQpdid5etDMBI0qAJRzuLGeHzAQLHZzPrSm7+dC4YxH9FCfBT2bbOMe2RGwOR0+Ab
yo784k2nNqU3FEt2R0fCWsa1YHMrDqLUVMiZA/TblZQ1WxfEmOC5TBE2X4aOKpgPsQutq2+IA2KW
WK+cWozP8pnL2RUgV+E6eBbpn/SbMGQ4NDtJ+ifzCUQwzocWFuiRqdBhS1ym6eDx51gTvsO573mm
/p1gyTg7SFURin5N/0Mr7343A/4fLGmVwbLRZSCkWN4l7PX1LPBDRmW5F0XdxOXPdxfZif2q820V
qr0IOZSGK3I6F2N8AGRZ6QdQ8MEey9S51XwmRbt77Qk3qsqjy6tLNHC3zbMDXMsnfX9djwEkemXT
ne+focHcyBnGkqTX1aRm1fl9U3GdIj0hoakUiArjBriEMsS2pxqWWQZxq0Yd8i9WrpQWrS45SMBP
3xVqL7gIS8kWlTrYjNBOHuQDqDKI7Xv0MGdWWV8GM62ApfxHMuBT+Pz9HyqLl908kBgcqgKnxbRA
l58P60F4Sk2Z9lzBuqEFsSxtVJjeTmngz7gdQhWMT1WHSSVQ/FKZAm8fuzj7Va4AokDoD15quK0B
m6SLCMnb6NBuB6rd+Wuo4i7P4HqD2LpCzRF5J5V/f/zhxq7iEdhScYg3fVR+5JZCGCiYXa2G7VDb
YKwlZWPtqyMaL897k+k9bOzUyzY3Gp0IkHIHpll/y6hjHmkbZnXKA2ChCQlfzzAkFdxD7XC5GF57
PCosl7FPQv6vjt/NW291KNxPtA9jcCl4Hu2pKpNUjClTLY0HQy3W+W+rI4YEg3NCQ10Vk0hXJJ0T
//IapjV/GLuypW8R/rbBFtLaFWXn5+/4yuv5FIiQH64Ny82r/qVNI0RrE9rFhRhNHHErm/rsBT80
V6GBwtqGKFoD0DcYTUPRiyp7A1Itd9bwu5qRdYh/5YyrSXHeqbkRFJU7jn+JQtd2sQjl5CMkOJmc
ngojRNwmoK5b8sgHJssYa00ZoxGVdK5RKMPeO6x8TdGcUY54gY7S4od44G3dVlTEH1f8aqy3DxMz
SSrfc2eVV4GAn2SXWCquJnXLCLrgCSR1ks4upmQh5ZnneI4kIckI/n2A+5EGRt8PRpF2zvib+eEM
PBUjoltf1Jk8BxvfM9efHFtWlEY3NmJ2g1jF9/5A98z7wRsJNy7G3k7Q4eI3Rjv/5miXE36HGEBd
sKBPglg8IZ4lfrPKkwSbfCCsRuP4Kl4X5lG5EfHk8XDRXar13O9RPVlkgeM6vqb1zoKg/xy6V2E5
dQnU7NqEihLVefvuJaTqcLBymCfoGqARW9Wml57mwR/T2QXpTFELafQBQGjgSG4iCrM9HvQ1HSOX
6HufQFY6WkQrdWqi09DOmkaxqX7GAN0UUuYFw+N5I4YSS+vuqy2snPa69w2EuRGPe2KMF+820QZG
ckaG/PnHBSHOvf1wxi2pdl8J3ZGNTqwun3mY+/dIAl4hU+2Kk5JezJJ55TH2vo8ZvXmo8xfzupy5
Qy4jQIYCbUkpzuHDTFr0dmIejTDSwELGlcAfX24dW0m1x1rl33XlrVZdc0HNzgqXxjL5oXpik2wd
8y5IcWcoU+G6TKWRW1WZPaH9gXbIw7QipquzvMQEhXf68vM42ZsMFnHRtHDqYETfcQswj8aNfRvr
LB3VZlUwiZva/R05XegkYat7hh3VC/DY94baIZjESPy9DKnzI5zA8luafacX8djSJ2Q4s0nsbMJI
6y36C/2m2n6p4RM7oUOaRB26qwYQOeH4gdOyDvPqa++ja2wguA2+KGLiIa4FiIkAPc/yDuIgg8Lw
lVrPdjOPuzPOXNyjStJCtv6/vsa5DsCyfDnq9C49wbRlcL82tuDogcMSnyVYB7ZCzxNSfxhkA7iS
cKRic1ZpaLsUjHLIoW7ILPsZr2b2F7yJrdkalk+/8WR0iekbR5GCviRh3Fe5ERwGvRNi1VdJkBvK
iPYvNTnZRs7om922OnIkWBDqLKCmszm9fRyMfaA4bvET1LRByTyjH95NUfe853ZooWqoNFHXzrKb
sB11bpWyhh5rnUU9dhR6wwcqPcywpnAIeuInaE5Mphfpdu9mxz7wywBoJFpeE/CVxnkts/UI2uSU
7ULtcnLEvG6pETu1VkpPPsJYFTQS1B6CTF5EnSwh/+RqljxxfOM2rx6u0wb2wu38IaiA2nYS3Dyx
lHxR8dZuMU8LT0tluvwqk1H3QS2dI9g2fjMdvs/ZJZukHsRZ+i8shkQ/7Tw0p5f1+MTDb7h0Pmmb
rtTFGBsed/OCmdA1WJweq5xc241s6RqQFT4Uahyh4GqhcqVFVZv2wQ105Vw9n1RDkPqD64BhnLpf
rWPxquBzCoWdTApqn/3S96NyrZ6Zw/rEfbTXp8+4H7s6bzGfqGayRDEX7DeKMi6WEtZBCtH0TfqN
GZsEAeW+YQLn2VHVKbB/9gmREoM/RhOuvfPwFNkhumKzXqtEONXBLQw8R3LE5tnJxSUEW7voZ7vq
Ov7Ex+uILs6DzqzXqaNHsW2pLn2F84WRq7B/Ecc4A9g5XPWHFesNTQpFGs92T4YSrsgfqeCMQglj
VlaxUxjSAov9Ty9gsJiAWQTzkvTguTKpAkVhDrxTNFiLYnbCUk9N9xc1TOl0wtpXxX3bRqhMqNcA
aDpkMf0udY/TPRpXvCM1H6HGXHA3H4splIUeY7t342C3v6MFCc4YoOUyuTHmxVeU28/Hz+GWqyaZ
XC3Iky7a5zpTVG33n58PzMKWX4pz5kPF32e2kfWOTd9u+SinbVQknWz6g0o3wTNKGPDAfh/xxN8V
x2e/2FhXN0WLIMtCJap9xqJ4LEpLjN2usYIFiU21OxcqRYCwlZhDHnNYpmsRQSJSZqmYV/6+Rqx1
T15cH1cYy3gXxhFD5nFLNZdIq0Gdz2Oy9G/5qjKCPdRGsXa4jwgsV1Kwiv8Cet+1jKM7U8b01QXa
XGqoIkDK0G+tU6c3ChXIy1GH+uClP7eoEnTwyX/rSSi8afyZvG6NIRYeJtOLXfZJdYdl3TvoazVr
+XwafXGg3y9yVmld7vy6ZwHJq9dC49VGFnu1Gmayh/H7a3J7Se8aePIN2MFn+E5DG087pNbG+zEI
NhCd6s60sITAsHdAwus9oJhc65gyYgHZftc2VpGVKDGwIPd+zB2lt4XgDmZNX7oTOxdmA2/izqXt
xef8zO9W0V08QPcQ3CYMkB1aOs3mO9aUUd+gnMywT/WwkUMuX7KenIwlyx7fsuFgGD00ufcfDeKR
Hb9S7kJmtDeGWbj5zYU2+MMmq+VX/Ch0d4dGUF6IQ2QiECR6VQblHxLadnr9QS7zhmNJ0HniaD5w
bSCbuMGTEDnmiwJCHpG5nFvrP8ci6Ev6VhtW9kxgLYOw7CKXO4HP8qb3htxS67WbosF3gBs1D176
Wtxxm7JxtTbW3Q/POJ/g+sWkYvQFhsD8pAjX7UgnDuyJ50ukTWh1LvA537li/JkZeZpFfzFfSwqs
9qPEooBuGHC0m4JRZrv9tw25/iRO+u0+cbekBIRAbMyyFRYEv1BwBgBWOGJX2IYrUvHroZh2+6pH
bcVnAzac1JUt4v9PnXVw+yhR3soXPKpeS/mrUuanAtaKc+GNzNyNQPYFDnI5cuVZpf1veTB6wpIG
MT2MQvaYQNVdRws+x9nV/fmGaNHpR9JAZcbDyGayCktztI+0gAPV7JE47ot1QsiMQ5Mrb29/3Wm9
PjZfSNdR2h9zq9Kcw4wpfePSEU8q/B9h0HT7FEDTXo3DozzRxvrFNRf1H+nvcnLdf+MKoDhdeP75
3Spbo0emHD5Yf+pDLULtHTwBtXXZCIHrbQq4wlRqGpczmi7smApPBnuf+Z5PqrIvTRVbOvXMrz8n
k0Et3mqFr8EJ3z6xFptMZMlOtiyp0xLOKtrnTBEKb/c1+QO+9qBlNSAgCj5ByDxzoVCphekdABDD
R7UeivLHgCwd6atqN16H55869XPiL5F5O+6kKtBO0sQGH2nUpAnghA6/11zuQLu7HEParsEjnPX7
SflzcpTyVKeMC8gTAMWdaV6m+LfUKRvo6nruPfy+QxcJVlneewTYNxKSVe6eBhlHYNu1oCKsRFfw
u+LhA2M+rsfXVRYZpBPK44JypYNzuQCM0F3bCoQUlhlMDBAHl5fKtmeTn9D82b4Q+rrdm/b4tUQo
3yMDBh/3vLtknZcQH5y5CT6B7FHonF7cnPKAleYjm+B8AuAPGrcYQy5d4597tENFt+wtEJyG4egf
mwm3UrBu8UVFflsXwWnkGCROHZAcB9lmlgK8ofg1pvYj5DpnX5Uqpp352TR4OABHL1OOIewVe3lS
ivD7IGfS26XMVQTOlPLwDwtC+nYEzlOXIjfk0BXJaqMRAYR4IxshgfV36Bi8YS+dPkDaWNLL53vp
9szhsI+D2018BdlYI+11ig7YJ8MxtvubLOVCj4/PS34ZPHO0XlPBFm7bAO83MxTkQ3NwM0hsViWv
9GZ1WZs+lzUBUACOmzv2Pz0oKm3FvensHtaoRLx4KRaShIepJpklxvxElNKOctK1SBb47gqq5q0R
7kIr61oox9ovixg8nKWIjDbBYQrRg5s51W5kizyjjjXHkYo6KeZp6U21rpZWUlVsC4acVbtfIczi
m/r9sKeB15OeL1roEWk00+Hk00l0O2Kly9ufIChhap24gAgIriZHMcKh+MdENk1IGpSSfCrUbR4m
IPF1n181LqA8dFoYDN55ocSaZQFGzlP/ZRov7tgDB6p0nlr8g9XrozSV6Hd6r0pMgZ70Ew6qdOgH
M1PvQ+aj0rhNyWH5+CDKliLEFaXv4VflUDG9ra48k45UKigxQrSJ5RrbtNlo3h43QmQ1nphbu9Ef
0DB8ZuFaq0AEraTHe+g618Zg9t+gkvOXzYo1XuG1lm1IWTwoXA1iu1cKVwboVq19JpLTxvby2GIY
aA9K31y8kBwf/lRCrD5klZ+8H102Di6jEila+fjL0CgXvJCVPyn+MD1s/Z9vQIbvUe3tkB3FxDuN
E1RBE47UV8ZJEFV306s0ocOijEj/R0UaTuj5LspuYn7pI7Ujh3dqX9QBI4OcA/nyD06ZNFpNgC5u
QQL6Ev4XSapEbHf1IngkWI8yjqdQEWjcYIZ4eusT31FcJBRKqQvb7op3C8lMS8WsCx0mCk0r4J1W
snzpxvee3isFBxyqMaLnecAFHLJJcADtc8WTWkuZNdXI1Pxkx1FY6fFo50HAWGq2UtgNhS/79MjB
1cSE3zN9KQKkR5kdxoTSiLg7yQB12zCedPuBw08gHmUOwNpdyR98Z2Y+dRm06sEixv9FrTLLQnLB
e9HY8DVsQAm2FYEGjUEZqQiB+PZAMPALVUtaPM+PZZELSYcuEVAtBipCJ457P3PJg/RsNupxli1n
qd1lf4wQdbU0y3kVCdNSHAiL2JOyb2EIi81nPpsQWIGDbe48AhojEttZ0YsDz3Mc9NNtSXHUknfT
gW25rAOtWtQDY+p9LCUvjvbi1GNA1hzmnD/LaI/j/5t919Nwigy5/aS6U/n8xFI5fgR9R9fLivLE
0AzCrcJVyr2kK0fNUInZERMnWK2voB027Pmt1ek9mtmhN3uClQFJiQsHt47dJRbEyv7JY5FQLwmW
w7pS1fvhzxjVfyVPWdkekpP5g99G14xC0T6F5NeKYnzu9vU5w3REspAJYPYGEtaKMBUAUz9Y2puW
ptzl7J4TNJL/JpHbLp5UuZgu7m9fr2qyI3CslbsOwv5uZAwmYQTrOpNWgtb26XsZIqdSRIuIV0f5
ffAAUjHaz7/nfIg75WZFEHe/KlVmAN0dPSC6AdQJLBhz/Yn4wlfBiJt5xWbXKV0olrIK5lf0pXtO
IHuRLFirA9dTS7L/5QXOP+YuKQegu5iFCN9QlpcmP6CWhYb+/NdKLG6w1Huz5Lgjs5mGBsbYgbS3
Ma0OLGYmeTKSpeDorD+8eHlkqCwMLKmNVCtOZxK1FMgPuayX7MzNru9XaOrMOPGtR+ZhmDEZDx67
U+iRDCkVgNQ4ZcdXglu9bqte2TaN1FVGpBOApQ7C46F/Zzx9+I8CXKg2Y0AAnJMtIEkH2UuI+r8F
DRjjrjuAhJmRYJtdxurcLAxJwbDGeVvNgQmTt4UxfueoYYz6s40yh0GD+D5iUiJkTVzwrcTj5mos
vbphSmXbE2aIaLPi4ddV/ql5zDjlQE9+2ypzowdXK80bvf0i4naT1fZQENL1Li+AYbE0V20UoaFA
f1Ldo740DT0Rhxyy8NjuTwSQ0JDnfKC1k5He82Dd+ea2WSm/zZeOzpfivFf0CkbhaBv9U916VvuD
55ymrVr5gjEUszQ1mEWbfKtMVob1FsBaWIaMq6YrZIGUB3G6ewUGnbeompAWvCweIEZfRwRgU+XW
OEQ0wff4bOypejL4JW7YpCO9WUkFxFCASGPe3WHrWMZAxc4KgT0ivApgamNmLLUy4OElYHdyvhdU
LRlpnDv+yLrYZfa4S+kaN8HtxFr/Y6rXGDrzPL1w+5MSj06SUy3LuMl8s8CaeiM9ZZl6ZyHjzK0d
BrbYe5SSIlIk7z/V1/F0A8uQvix/5RMqOU9euOVAaLLpJfrvbzGc2gTVKBJuzrm2tyjnZBPMFmS/
7CHXw90gYeuS4Ana9goyDQD75FBCH1mj0x5dspImkLMRqxui3R37CYrk0z4GGHlS/+ZFxrzk48S+
IMmwBpX9thyeMVOsC1JFPcKLsfCnN3E4ayFiIV2bBqVlxPfcQXUKFeNZtkDKGg/jYu9k02VPPSMq
6HuKPQFtk8657UzBV4wfiTwH5mL8rdiog9NIUz5vjrb9BJsC4u5uK5sOUyp31SeL7g4ZRC4hRcrs
clHcIaicOgmjB96zzGcWhJ8B2YcQpiDuXZ0WM+diriWiGkq/MIlCOjDqXbs5FedyyrQVEczucNwy
X0J9ZdWqMPtuNDUXkXrNJrCXYkqclFw/rvN5f/+1R3oJbN7nC5kjqZPwf/QeYnCpAdblo1iDbXFo
PR2T3+q3V2Qif8kfQBvR0DSr1LkEZN5fjyYt6P3EDiiHbQBCtNm3PXM1/38vcLhnIvQJMoOAVY7b
BbjrmcUPVTExLMYTxn0lFSQ8F44IXPm4Q7UUfrbzfbBLr3JrVYiBieKWSU0b7anz/ed/9asQU4EH
H4sClCJ0A0OiddsUm//gvVWTHkQgqXXbq8tJo1XFY+iim3uIWgxMROIo9V+0rY/bB8agr+lslVMT
zcUYVbXPXduv377e98EhKUM3NcKany08PGS/Z2GANl4iE2MIUgiH2KR0bNLShXM9qcEuY59XEJX9
7cAin40S2fsG1MCElJOCvwz8cA4ueGvvhPEVDyDNVP/h3x3bYOyIQrAbEvqNKBmyUD62+EpqSlIE
046fhFm0dLZVRI/D7e8xfv7wteWGVcTJ94vXlOFtMmyfIuaubpT/twsetDsFwbH6GI7Y78vv/9+v
4V7JBnxhCZ1dgu/DC1qGicECE8m6+na4ECZvsxZtDHOTJLG/czeYsE4xpj9tyXURRM/FrqOFOBxq
TW6DgB1e6UkUk5JcrecdlZB15PxTFEd6UU2VSx5gSo5Yc9fzYrr5sVLRfO/wtHSLyD23mNYwV9ed
bGumt9oZsUTCPAaVwG1y6Z7qCUP1h1th/gh7QulIGRVk+V+81QA0jMe0dF6QPRr0tXrX4qRt0v82
HhSqasaWxUfZcSDNr3bMCQBxkVv+eggNCecD0yCQ1RwBFkGg6WQTK7J5YQn3XFHPfMH7BcERoUD2
Y7KtjmRfawJz8pzIW+4YPE8qXbtow4/Y6rkOgdVDEvyz5VapjDepHX6jLQlB9hEeKMMQcAWKoerP
obkrGQPUEWc/asC4k4jDtmRW4ji7vykhlBWzne64CPEItXW/HnQCYkgJ9f0k3P8M65ep9foUI8kA
Le4qgX6xhqkyioEYcy6xOkwP78GyqUR7bL48ff4fCwHIEW/QLlej7+n61nuZuuUzCcwXRWkIV/Gh
XPUg54qWJcPCPye1oACPlmEsqFY6RX+aeN+k/8bAzihGp+nAWbXx/mhLcCr9d+wdRK5/NHX0hKSH
rxlh9DSwtyoVZANpBOgJF/3bUuELO1h0Zwikz+VmPtDyR0C5mMOUcKkSkwVrumSQQUjzSWINZX5+
VIFzLimMoLVq2T74D6bLJ7U/FF2vHDjYTERyykapNMP20maDzd6KslL3oVyH/AEHwZaXZjLe2x8L
13V1IewzYy3dUCazT7X+KTMtNB3Ph/UYupevb9dcAjfQc3jLTz8aUaHMSt2/zOZBHCtRKa6uUEtR
zI6lRzhvQ6NsGH707UA33wUngO8tWMxEhxTLzesdRHjIiTwfsWSBusecmQECOEUWo00DEtnRJYHq
SFSdEf44Gapx2I42aPSM9OKofqNRYOFUhUh/yDMQJOZHes3wEcSCBpxpu4pgqp3r3LhVuQqJ+2R6
PekQTxaqaa/TEtMY/04iCdEYCS5Z4ujxMK1VXZo0HUtu7t6pAdYI6FtiOBUfXokygegAJ7Tt1sL1
OrfXeBQAzTI1ViUFfeEmUbe1JhZG0+nfkzOb5U580HYY5VhY0N4QznNgncvB9tJM+b2b17TcO9Io
gOCalvZEcO3Xos+HCyaT5tyy6VYRd2tYAdA2ibNP1TE8MwhVFFlg4xPEXJQHe9UbA1cPxSVmX04B
rSmY8bOzGs4OAvcFCY1rWFfVT68j+zDR0rGgq9M50gsFgjgD3Q6Eu++KmLTHs2UlEh+hL9JmWJBQ
DV5bnoRVr92c1d4bdPSfs2fN3vTu7t7miE5ikX/c883OIKEzZc4s/F2/nYKnkCh04YL8XynK3eSa
+JPH8wML3WHk9BgjjJRRlmc80WwGo/uA4909n587ibiVA823M5ZcSVZQ6+oBMH/T40GnmIIRwbKQ
fJU7jE3rUwHdJ2VSK683WP3dJtiMpPafAJboz21B4Zo8XGLx4qY+PYdt0zWaVn1Ev7Z7ukEQgK+s
Obu86jfkbkvtYdjJ1PDZvmHFdtpUhusox5tvZUHCGbTxGQx+uOJHddbMKpM1Regl9IZmxZQ5O4Tt
/C+SJPCGIiXTPQU6OtipS7eNMHCPLCRwVyX/rgAKxBPx2JrmFcedLyOqV67l09oeux0i7vMGxinz
pzQaozUm6OVoZutc4Tp4LWHhbmKePPn9Dd1seCVcBWBvkuS+ktiDrIdWBYiXEpa9pr4AvrDpV92V
48vw7gVbUI4cOJv0dQ0LT/0f0BfoMGEM7CJ+lvA32pLHoHHbWcna73GbVZVJPCK3eNd+2FL1acgD
0DJfkAYVb6sqLblkpTxkOu0FalGTaZ+1r8EBar79kOOan524P4ZzR9TONXAfR8v4uXE3QpgQYRMW
cioPgsV6Co6AM0OQFZeQWIZzE4RE4SiuV5gKj7GI1eu/6mPAx4SEbhnhTfLvIn05a48f9p88XMQv
LsdtkFcIuQ74G8K4rcBTezR012vDMzJ8gw4EF9yJfScBIDbK+vRWos/GsDGEmQXSGnnX8qe19KCr
+TGjeoW+JTipB/QJfDM68Na3NuSExfGsU7OUtFCSyKLdlXp2FwAFSuOMphdHHthGqyHyWOnBFeuI
hqmNTTS4uyqGoAoYINYXt5MT/C52H4ZE0Zvzc7UzUpI9PsMt8JVPcx8tJ9Rjs6kN29/Sl97JLsFP
91bKm+a4C+UX73APXD6DqSQYiZNsYNg3YgB2uuhZTrMOgfRQn/7RLGBxBXVG98HKZT3WMYalsEqM
odQCo1BLvk2TFDn4fFWWMm1knz8ZHYXsZIh13/8yaj3lmcjY/RKlHHshE3ScoI4rQTMR4xVz6nlh
zBjI3MI0pFFgOTKC3d0OgR/2bdMnkvoFKjczF0U3FDB5tH1138OPOzkHR8barxOHqXB9I/VitLkQ
KggRxCxdT9y1LpR/UiFzsXDh65xRnYROBsd1juy0PWtG8OHpGFzXr7Ix1bL1tsU16Orc69sf9i9+
DjpVkLHEV8PuWM49PhhFq5Y9+aMJNPm6vqEXL1eoE90lVphd+UXfcVEF1rh2aUmzp09IbntNxyQb
N2HWu6QvHLpluoS1DqhVLaBaeEh7psf/0QKeL8+v2JttQOW9sNWlaBr7paA/pdWblyXWcYIWI3DL
4SuAi2jywO07fJWLDL8eKEosja1q8iOIlZAfS5jHkoTy7XjbISK80kH4zbrPNKDEO+0xqRFk9P1W
Gpnhq1wK5u509ivluU9pkL+S/ma9uubYKiCeWxuse2Fs+CMk4HD+B7Sh+QFhx5R8yuiXa+KNPwQR
upn9XmQ95jMHeugaFpNzJttQSEnWpHq6j7y9wJ9lQzsspHo0Oo4FxA92UVMMrBrG7iH9F6wl6sge
K1DPNM5Nhu45/j+y8I26HL75AfSDoJkyHkOzl+R9syS39Y8xoeWNb0ILUR8/wGTujRa+GesuxICT
bA0e6j8pxX+QCqoqVPl9Uls2DdzfxDt11gWe+Dp3zmf96UOFD3u3j2GgSXWkYHJIz3q7xiphOqKZ
tX6PK1z5P+Do1YN+cB26Vx0xr7LEF45EZajN0b7eg9Z+M6+sMd5DVEIMDU+wFnW69lmKKaeJyZaq
kfKB3OtBOEA+K+nPVCvoIq/Qkp8vf/z1oMs97m3zp8eXX7qgISBxv1PfPnvllMHCIyl4wZSFHb//
S+4bNyxkPDj/fVEO7ljQrjWGXbzu9qxynNll5NQuU+icBfPxvWajbDjaXCBjYq9ILD/l+SC/XUFj
mtOB5elYzIdXiPsl0FhA8/8yrtTTkTuJJYCQP5PGnsBBw7rAFzd5zWBr/k2FJh+p8Lwt6b+0Alox
80xtERBxr9HtZaLObUyba2r0cvLgmqtfuLsn5TzF6B8T9nGZenXKgR0e7z8nPkNfQgFOlosF6bGU
zS5RZTooAPexQ64bUsoMV0jCq/KHQSOsMYIktITnB1QbiY6ti35CT8tfoDHaismsXzhmNlEryp1D
+/iyguozuvrV2FDed//NWeZ0zGZRDa72Vr6YRWW/3QOG52YzBSj6khL8H9rhbHdtfuSFh+VDExUk
bv8q/ZucK1YptCgjrRLUqu19Ru1XHJ5qKrbguIwWWkV/1ee5Zg+XNjiWZTqJZatUQTLIZXh8+Tle
2lrGBiI5mHzxphXWcADBlz7ZlRsmJjaUGn+++JcvkX0CM+6ErkMLqj5WqkmYv4I2ssNLAdpD+GRp
nmFBdW4OAw7pzp3alNaQlIaMWoEJr0hH+3q3TTt3stYglW++RwLXHQoNgzIniZRs/y2t/5wlRDZ6
gUtzBPVye+O5+3enittijYbCLJOyOx+R46Gh5Gz/5lCRu0ZEiOneArUNxnvJOTxPR6roAA2vSRUt
QH1gm/13Y0BgD6NZcAxjoFdTwqt7TX+K+lRbFLH2ZisEJ16Jvg13APXFjb4EI9hgo1q6vhkojsNG
rYg6j6zhLf+TTLtPlEDU9D6pgNXIzpb1mAldyZJO6QPLbPnA+urZGFWeTE49KSbThYirGWCqfxzo
9AcHV2y2EOHqhcqVDcr3+aJq1PNEX4BE1sYimsP2lpRZcXXEg9092DpRIh29TlRA+nK/w8zlBOYe
OevqK6vndQGYdziYBYRsLu38kbEMDJr+obFLI/GkNGGp+clJQpkJhqCb8u3qJ7SqtkhLaYC3smTF
fnp+MOjmvyzNyzv1DoiKPeRacEaWIIhCu5I+yofy+keFMPun0u0+t2DTygnvfh1mbt5w9j3GPcqK
tpHfU9Z7/W3KN+9qyNG6L5rNeW4sNZnD2y+GkVx0jIu2J04rGjxE4hjszNtxnLgqvdcZhSImtmmL
DcmBKoA2kMUJexhi82EZMG97BRm2zGT8uopVl8pK1Hc33M5WBAubU3Xc3UsSFDAEQdtjVQedrYm4
X05jnp3Ol0kDyN3w659hwcLD16doW+KdJuPSOrIvXPOLqveqCfEuJxWTahGIQJmjaDBpSj8HLPhu
eoBEvXeNR92fk68iyGjwu0yKoadVXNtSlKLBdG5GW6eQxJtaZzjBstSLMXHV5zcD4Z5fMgCNhJDD
8vkCB78tdW9xBkDUQl4jn4qb6uSuNFFlnY21FTmrc1rx4NhJILhd02Uu+ony0JyVRKju57bmvB4n
pK+PmlCq9CpjaarAqJdYn7+ICaRfrm9i2WTGqcld3q+xNAqqCaHrBapXiQcAv5bIWjxeOUcJYJmu
FdZG6LzJIdUJlqVcLdN9tfVyBI3uInCYHQtLH9aYccNYFnh8kGfrArSKvBTw29vA1aMv0x89tQw1
bbYRYpLS26Ak2+K9U4x3AELjEsTX26f0FWORNAOInQBnhJkKx9BNtL4Qbf3pI7hJins0lv/egDjT
/FzjANmxtV1BfxNPUuESkHyzZsNeeedZFBTh2fclNhveZE8QmXsNeI19EDZL9UST1g4lMh5YbjJ7
BTpV2VffYC33GeAQOqdlffrpuiOxXGYFJYSS5LTK1He2FfjblIcFyKQ74iAwUTyNpt34Sl12/Jah
2VLh9doSVrYP5ZEHpIo6K/67wSh1YtNlAFXUmy0LNFRg4PU/rb9GDGXbTrnE1Rt4/ERE+ff1tgeK
W5xfAwf1MqVZgQCK8yp3MfriCWDioD5yR8mEKPo+zEYMq79mm/6bHILzCYyu8nQdAYyzfoSlWT9J
ErwhcfP7wX7IabA8RtuC1OCN1I1E5Yv7TSgzwnkYXAqE7ePLAOdpGzrk033SsEA4RK48bH43B5zy
SmYGmlfBYjYw5ef3JGVaK/DlD5+8G9+NkZoCptxYe42T5gBaKk9seplLafmxcmxIUr1/BWS65Tf/
CTD/WmSxjzR8qLMFs/5jq9nlbegw/jHW7OMlyoHR9i5csagU6bvJU5tSMs4+Se3oYkPPqDwhSPQC
YMUylnYccB/h1k+jJVCA6fYT2rnlBLG7PvTJZYZ4MeRkTfyA5H8m+VZK5tKhognKfzOSAau5sAAK
Em1/8WKjH5hwz/U6CwxcNAE43gvF5yNLbctqm7LPPC19/3qPeC+LSG0WR+Gl//GIuLFIvNCQhDZM
WvkehKhNdv+zSeKdGRlzafo7fDy7wJWDfwuZUrfF63eApAEmAGaysgFArwlvVj10TrwJpFwg0r+F
kEHUvlWzcd535qXXsc9J0cNsZt/UTRgZUcOuCGwYT8W8ZWamTWHw07fLi3qXrEdFqgS4VAIq+yBx
2hfG9bbbnxNpZF4+3hHnSMUoB/o1dg4cMFJx16NbHE+TQ8tch82oXMO8sN3+VSxLIcNt3VYQq2dC
ytmDOWkERGVs6uKJ8luAyCcIRKft/KWHG9eczfN4G6K+Lq61TV3EWoZu4Re8sPJURrtcZb4l6FLJ
Rvdws/5mxOJxPY3ecqndHvLKdsRRkCKTi0f3WRh3VrqUn2hozu6W4h++5tMAhA2WwAkxUPaBaT8B
murK5jRX6gyuhBNoi1rFZstBek15oNR4K7Y7WCXAnOpl2LjdiONYPBB+NNGVntwOOho7HAMxdOc2
1dymLSRj02bOwRwc5KHsrWu95x5pvAAbQLfa+jHbvNfacj94R5F2RgCOHiwEKPteYKxvvddJbAyu
/x3cdJxHsUANLOh4arIhP+1sf7syU+rnhIZ3o5eUk3IMN4PoNz/wr8V/gQEidGph0m2N5aHvAQkh
Vxja8SgHGL/ZHw77T8HAvp+PEy0tyMLh4Gf45D+IkE0XQT7cOCtaqV5kM8s+i7sskYkGoh0YDGtC
SpsHxi5MMxO3OWHgiqI5L6jN3zag9Quc4gL6/59L9aitqiXDFcxudHlDBc2/rNdZHqGqAzxyNGVM
4eTaY5Nr6N6+uAgWaNoa+MDN2HdzF/Yyj806FJaYGCB5n3MW1PN2SnNa53S9S3N9BTB0U9m6de/O
Y0knxMI1vISaqoGUryoCLY+AX9nG5QMRsdqmVvo46yQVmitDc4wBVPNkeaNsvTKtnCeyfnm9Nor9
zl+L7ztaC+iWg4rIJGGtPVGOZdNlwcp+v6lZI6m2a7cInk1acbhOcup5AOggTWAvOXFNUerKUoRO
4v5YMVJFfk1menzU3T8NWJ3tQkz4IKvLs24LJkKvqQLnUlw1zVGVB6MpQHHo0tIFjth8F7KRuNS1
ZNtu4+QKh/4Z5owyZPXbb8LG8ofAcF/0UOPaqGY0BEIq35yheqZ1ah53pIjrdzc05aMz8d8kGWXz
e8LWzRHZU/wXLy4E8hgrwca2XE1/lvtgvDYSkmh49WHTDBt7l0QigKZ+58WokF3pb0c0j2SPIA5p
NO9V5UPyR0WWNP+6EP5WE6jwSz9eIvNvRjf3pq8Ymq8N9iyPbBQVUiTWxYfMJ5LeLZ3Hf4yZLm1R
QGW/VINpEnLDFpLYzMhfyoyZCvpAw5Z2ZGe59FxPZaMHtasxkJ5Qg79pYGNIv1lemEJX4w6PF49t
FF5nW1q/l5wFWH+gMHiAsXNzrt2tLUcEPXYlb6nXhDVy83jVwoppv4m+vEooWtAnIgLLAelEDFfh
LsyOs/o1wICNshrYGQ8yTsXmmK3MNcnNnVbbqK4fy2IQ2ifOAWfZWJkNhIPQ/xq2aidTE/1TjEXq
R+vAXFQctRXHzIMacNbD/iacOBdrpE4xDqemmux4LCUlzYrhl9fDNeUlC9LxTu1+dZB7tZqXPiAT
hsSi1BovxsWzDZh1oWz/ovW1p+Lq5jnMuD23M8xwIcKp4feCjN724HkYWz1eU7F+24m/LqxQ3cxH
G4EI4gLM66J8KUzn4dM2YaD11g2VniocZNtyCa9hrJhdnJ7wPN5A0XJjrpLOA2SK6H+tNc59RVZO
wAzfCojEMnDrsIq7SQ5wCu+7QCZ6ISWIzAVBtRrNbY3t/myKl3IfnNEZ3CgwnAgQZySYkFjG0FRN
+xa1Z36xa/YXl+IXnXRyelvI9OgWjqC4LHfICJnLF8H2v1WCvILo4QFESVJV/uy9jgVkNvFMo1vh
/LNwd9rZS8olCaTz2X93JFGk7x5ds2EAUoJTipMSAWy2JcSRMuSOFgyocgTh4Hcfu3CbKnzEKhlb
+sYdbmlQBPv6ATHptAkTFwPOzpHLqEHVfnWfPoWEEtBz/IkwB+RncOQOn+eFY+diaCPsfDym7AOc
s4Nm6bSxZHuT03VbioZXUo2wY4ylQrhxExck6uRmapmxrnHnBVi0ZGjmFTUFlJCp1o7nWparlqYy
EWUAQk80a7LwcaX1TJOYzDwWh1wHeyJsAYG/ypfDdghAahKdwwf9/lGVjQwqXeLplKsNiUCvtfHd
rhLzn0Exx0XxahAdsgk8xqBeZDA8kpYTN9/A4140zpJxcGL0gBzPYCjOmQ4cLzYPuDi0Z6yzmlCa
bfcivKI1J/CIWGFugFw+snAYmV2ipB3T5ZO0QIq0liD04WWBzYW0n5S+o26enACcpn66Tmmmtx1b
EfwYgZcFZv2Iz/Y8fwEWQrzYVNKX7R5ThbGt6Q6kRlQ3+hacl8gQmdVD/KB0VMomDWncEKwcPxQg
MkIoF7VslE1C+Xq31FbjPpnK5JlMDPntSNk9eonE3D5n9n19H7spZzEsGHgr0uz9n817IkhB9TED
eAzrsCNW+x7ghRW7EuMlKvDZc5tarwxQw+9kI8NueglgslmQ5wqiy1zI+3OlP+Tb3g2hRWqanno6
ERJZfgMQf75FutnS9tQGDcWw+9rJTjWWLbddQEsPb5McuIOv7i7GycbwTkwzwcayQNFMVUHhEUXT
aHKTVJ0R/GE8CObrmkFIRGVgzytq339BhWRt0mJkEgj0jf+SGmd6y9d7lL9LzIx/lcovjd6RCRM5
2dX3UF8TFJOZRpRG+Fku0rSVNLvhTxXE3mWF1OrC3iXpquyYbDtT+71OLFimlzEsZcdXJnonQ7+R
iAf97aA3fLu6g6XYSCyob/0J0s77hlypH7W5xy1w8mguYn5GAMn7ShkZmvMFVd2Cj5DqGdMJwuR+
elijdtktIJgeXIM64+OxNCRjFuSeUXWSQPjBn3RRrRVj/ybFMCcZeCl5H43EJrvdaFgN7+NgYtCF
3bPCGEVAHGwX5yXehqM2e2kl04BpEo2Z6hebnCAxxRCxVOTiDpKbMX114Xu+WRXPmnlGyse7BC9e
92Qv1unS5LYDF6syNeDrlRMN9s0WIlyOCkWdw+NBouGhbDQRVdX/5oceLmxAcm/h7SNAdZvHwguU
9UoaAEvl4DkipcioyvEgC6QbL58PEWO9QkyXFXSV/zMbeYqT3yGW73Au2GvWJQ30JnpBb5c1XlaP
GADofjVRXGkmZL4dvU5QWpuiwP4Z73vrRb+p9WJnGprnUtx6HkTeqYQNqI6ufYsrEEhHKDb2Rbmu
UQWajRpbROqT7nJ/B5t3ILR2gBFWhFFXNTa6l/JAtcaxMRDdxwEHovxtIqTZYz+QQUlNDruI233C
NXNaAh4RQspkEvqG/uR/Q2k0lgA7jXatBb+fvRISERQO3RYXLJ8nUNWJvMzBOWL/3PHd+s9phHxt
hQ7h/DYvUspjNzvgcvVN2hWxQKm1GjBWAPMr1SzucKhZFJ/8eUTkiZXfLH7+wnCfVqGWkwUjj7Gm
S95KC6Q56/mN0Zpg5Bzy8zkWYolTAcoUfU4nUozrvpo3D+u6OF00tBvLEeVLIsX1zqw5WW3jLouh
yurkzGH3QSSSNtlqtSGBM79LAtVb8Kg2BJ7N4GUpuoIVczQGIbQa48J2rPeZGVB3Kr+BQ/xZLHfr
C431eeUBOWqimoRJzERSXY9dsrgcmgVJfW6wgzOt2nebVHSfhjyJQXgrDYMZXDFUDjfZvv7HTgkF
bceRtcUxzSNmcVacTai97vJRUE48D1Bsgis8M5FudwQSl5oGH3yR1Q+n4wpEpP/23FOppIqDE51P
bpDfdxoz5FR/S8ISAtAcns2kaUYPfWT67QiXX3dlfXXHdpNd0FAnHPHfZCNmjIg7hErvpR9raHaR
IXmiMVeItPs07d0u2iXQNxzo6su0cJAWR9lhev1WE0fzKRcoCcKdA9cEiJrmdq/Wg3XQoS1Pvsw/
gNuKUtxTo5efaBaG47O3lWjCsO3GI5agb8HQl7ZPe5k/RipDdr4tWKLK/unIsSLDpQu2wiW8r9JI
7T1bfaHJoXVBBRuitMonbr0oV8659Wns0lThLCi75S9Y7Ec7T8+atgOBSBt9cXYLZtwC9GZw6tfm
8xsQkAFVCDy8ykH6uikCOeewDJ26Pr8+WOTa0CHtP0LUTo7Tyw4G+LWnqjWctygZmYX1OBvQyqO/
8x38YD0o0wyZAly74jPeWQQv/oLxeo7QZdfV1Uz6NE9q1ZxOAOO2gy8w+psfxz349eP4tHc974o8
Qc6JbYVGrYY83p0rlZNK2SnddelNBuuwge5OASCwcmuwC5HYVsEX0Ctz2/Y3P2OpNXDX70xubJnN
xs9ZnB94S7aheKajzT4vBRj8L2RuNSy2FFTqgCYHQeIWfXYzXqx2r/p8vLsv3i9v3Cv2/+gByU70
s3Wjtpngoqu+U8rW/frrR0bgdUtR5CQ2GM7cLTEms3NpnuorzPB8jW4SBHB2CuIyWrC0W2dkZp46
Er3YdpFGMOu90TtOhW7a8x0Al3ru3tGnxptnLmhGpBdYzyMVVdRcGQyqb1KYvXidnfM6a39Od7OO
RVrSlIiwSJb4bV29Xi6rRwXTMmvgemVSdyLA89+SRUIz9rBd6mnnmzOq6LP0nEaaOZESMMiTlScm
QxC4pFsefW9uq1k7afnFHP0E0p/RJdf3BPSQUtqB7It4gwkGhE82AgysWTn8CUKi338u3LbJPaNh
G7KC462cFrRN6ko7GRjPShc3YPOwHGXFjpO76E0j3xub8mLv0rt6cPb9LkFsUWOw3j6D60Ii9AAJ
HbcaHUUCMxOYXiJTsqrzrX+qoSrb2dAMfwjqpU5izitLbY/XFXe2ZGawEUzlM17GGfBAeIoSk0GD
snIpIot6y3eI8iiGSMammW4Dp+oZHHGiGNuF2ViTHQs/JduwbBcQfwLg3a5CO5ePsD3Gd1qh3NRZ
V/wiFOwOKGFDUC20ajUH+mm6l3LPQVj4WnE5jUWneazmNv6A3iWhiOTkWbIu2qYJmknorsj8jat0
lwex/rb5azBWUlAgTQJWYAZftgyxmLBXA6E5gT2efx2VySM8fiKuqkcd7ofyINraoJbSrI4Qxnsl
yDtS22DtOXC6E5pFBZ8R7vEPuY5s7krNQ5orhbUNYHVgoenCUJoKTr+3hsZeukdx9bflQMCNWz+a
7KTB3UeanASIJLTyGd+8s+HLoI7BtLMRGbLeB4iFq+iXaIvlCaVygmIafZu6k7iTryPcEo1UZSsm
AI4i1FMBZVdWPv6SRBBh8zXieYYh1nzsUNdb+xgjZis/9TvAd9EWipJieZXMB9QD3AY4mFA5/nYC
joC0VihcOz2jEi0dEtOy6Dcy6cnHxurHzm40ngi/fq1TUodTIjmSuPHWAFeZldUz6i8CXGGlt8oH
IoJsQUDy6l49I0dxn0ACgKszMNH84oh5xPnn1oBHQCfSL6yYZLJw+lx+18asluQVEaoVD1LDqTly
pSkjtvtFDkUVe3h7/UvNGolZ66p9jOyU4GHHUdtJSIkqL2BHDiFrRL9PeDZqVfBz1mBtiF5U+a6X
QMUhFPfz/12uBYbSHm0vS/0qctOkkIagAPP9DD59nHj2B9iS9BZsqHhD3PCnKldSfwT/K8//LoLN
62EzPNA++2zcHPW2gZRKGaNJ+ekXtN1nFMaKLIu8Z51pl+rooNsLWm8j9CKONDKfqMrw3S8Cp+2d
I8L0LYcb9TIjEk28IsFtrslmKL0nJLvJRDKLaAQtEQ5B6ZMH+CVqccRROPmpi5TmRGEImBcBew1Y
vnETX1xTAhbQasAbi0W15NsLa3IQoAaHAyDj+gbHkg1ju3bvwuD9HqMI2lyvSYj/lL6YGoQs/2+b
G+1un/azd3jBL+yxzwXzl1U2FAEeQFYb1axApPsR5hFcv560KWVkUMGVtcxZ+GpebsKrliyvHSDv
NvVby8T3KKWu9KUAJSOs3FLnPUW0IV1/DJF3xDF5ZYJjgH7VvzmuwtlRDksy+oMpaDZL0KOb37pl
aq9Llx5mA4UJZ7uRd0XGYJPXg1HfnF7LgF/+RHtWzpHE1g3E3QCddGqctE3clGouT24O63W+tbIz
zWg2gu4R7B6PQ5haZatcFto1nKQkwKXPnPHPrufqQDAiRJcuXh1EGo4UX0sDe2oNHBNqPhcF1DA0
cBcKQYa6nIoDMek6t7NODFXo5cog5gVHRz6mtYK+AJOnsfTki19NUitZgVcK31uChBwSmb59zd9C
IPooMq1dMHunP/deCw9iQeAPiOvaQ1RYLvEDXR3MU4fSYn5O+eFy3karITZAGvtOC9dDW983pn5e
noxf1V26lAHees5f1njDQ3by6pQTeFp1ScVZuK598OP2i8VX+xnBmOTnyidjW31IRy+zEKuFwC/W
Fpn4R2JsgLSxCHtC9jK3cE0SuF/yKgWVl8YD3iSLImsoiRn5Sh0Q94zX5A+GYa+p276RPYJCswwA
qx4PWVCl6ZvgCygEZHR6SToVIjAcxPOh96F7TI79L5Z5xE7cAUCpoCd1wEkZA+KDZPZ90xUxYGsU
CdHbilAab9dCZtLH5893MW9k/M1Kcey/+3CTOAeYnJFTKnqMzeEDdH1+cJdbNuNz1cDZUiXEXYod
GoAG9QUcQhIltVr6vXzFGYDN3ihWdp051RzzKLkK1+y3g1wahGcy4b9hMfiEfV1FsGCi06nbit7d
ECnxYW3aR1UGRWw/zF5yPzgXHO1gWpqnOqZehoYiBB9f/EOgijz1xi0OkecBw/UIrQufvrU/a4UU
SXeUH1qVHYtUkMp2n6ZVsPWTd6/t7wQys5iHXFHrcsrLTtqHjdziy54FltlDXXErpLJwb/tznNuJ
ae3bsxvzeI2AZSO+LKfMz3BRs+/7AnUI1I1UPzl4wHGAGOndDLheritRHJ4PTbJcC5vGZdi2Cp/s
mbevrOZzBiIc8J8xQL6uYiyGPD0w3r4XfLyJNubGwMP3BbC38nARU08jx0vxA+ULmS58nOdpiso4
KJNMAp8B31AtdrrPzvKJY2MuPJXHg1LIeUtJXXwXhneC8mS8lfct6EeEAvbAl+yeFp7z/NIpXETX
R1XrL7hrCZ7SCj7z9HO4znRIPe8sIli9E7dt2m4xi4mBxKWksG8iZYBC+YBNvljqKN4mOmXKH+q6
MwwPmKELKvx44jlJoQFa5kLT2x8bIEUUmtZpj8Dq4O9yc0sN1aiKjgUoVRxUKClV1Bhj4kjRqyU3
y5plGPXQQlyof9N2PaeGki1s+ebhEhbByZs91R72Zl6aYYIOuG1jjkEW65sXPLJwBZgU37L8RSYc
/blnsVlHV0p6WMlp82H+lkYs0FGRwmp0EdNPupTh5nGlb9W9GSM6AHxL5PeYaanng5zxrRrBt2Lc
rwmUmvCZ/LBW8xSXbrWWefTGn40RfHndyaVpvbA7bTTRi/OmY/BU12RRK+WuKroelacjPoeK0oeR
2zmSlzzezYILOskfPgeg2quFS0U99psU444Y4RbIEX0MiJoaKj7XXLZQ4xnUe/LoGmiTBP1v+3mM
qwF1oBPRSimY7AZ+IVeMe1g5v3OGwJodmsc+p69p35WyFyTnbICtKUJx/Cyq/t2heq8JqDBLAE0z
JR9aEgiFRt/TL4GPzXntIB5IAaVNy+8WUNMXqyqzMh3KerhEYXvtIl1r6dH/mYpoyZDqzgh6tfW1
aPntqMF8m/NCHojzHpWe8wafKArLkQfXjvPlFJUfs0z1ZYfu/idntfKIyhr8s1SXk7pvEDRCkM6L
61QL+/0yAAzaSbARA4WDQYr/PmjhljhYiUyRroyquq9DgPlUgMokUMZdsXNc07d+1jLw5r9JLPNx
qzGi0dSMODRWVZDG54eOX+1CxI08ukutP1lz5msnqy44yK+mwTSoATykx1B0VeSRjAgL73dgW/ry
JZQD7dEQC3J6rCgnmmn+qSqv6xcrdejsfUcKHF5s2EotVCIekSCdxSGX0gnENgcRh2HBzTcjc6UN
Oj4co4lW2x7cWf6+yIwBVRuBzttcmpQ+o5Flh+2KJNgbjPuY1nqC2ghcK+XUiqXwd/5sfjdt1Jrr
LVl1LeeR5PgsD7T1KkW1GtARStYKsWrKLcYeAcRLQ8+epbrlRV8R7/yomYZYcykO8U61z5++msrv
GCLUgo4G2CgaNnyoxFrsHZtWaAAazlALrB+w7KP9Ant9wLIIel6ZU9k9iFIhfEJPpHCKKklwO6PB
Et21732UlPci7nFijwXtrECX5eWVbPkT8qRffhg1XoEQXn1j9puCMxAfYSd3ulGFmUD46jl82zdG
EVxTN0Yr2MfQs8XahfgKLzwqS6ZeJARlpDT+3/CCRl1uAE1z2dRPFrRFA7MFxGzitAKofwPuWHCG
P6zJ5VuvjVchrjFZh+e5LFog834NZjiVGQj6fEFxucdkPYvWPiun1kYhzD9slKFzQkk0AAbK0FOr
GCLRkCiMalT8W9aOKx/HGkmc1AEv+w6AWtZed/N+A7WUtivwh0QRW6DifZcXfTwYJHsF7H/4tjW7
wjga3j8WJyyudCG60kTAu65OIoF6SBrxBfoHSFgjrBNLEMIk2Q+nAJVkBopBnb//98Xj4Dr4EwwZ
kSURDnJy5zHo1NAyC13lx6bLDnqR1rkCx+kTQ6nm9silHkp2/XCRLB6y0Tx3HAKB+se45trUVehS
xNPwGnpoRB9isn4Ntz6x30ywfpm2vbPA8v0GLvbxRmQQ4CbjIMd1u42Gg9zVf73h+KbpF9W5ldT/
l4pYkDA31IbMk2n9SRQXSMors/fEtgqbcr3CPYhG+uViJIgV8+I6VkUYFySPGyncwlgYwqE+1g/E
jaYe9lhB4btHBW9Xvn4pIUlUK3f39H43d8el7mkaWgn+E5HhUGw/k0eBP9tieIBP516CGL/wVRzP
vh7JUxNRuWI984qSDaIFRFaxewz+kuRe4X5evEDEH9WHKMBmdQX4pAewwv8GHreVf3MsDBKS9ZI8
uXp2oPbmEOVkzgUefBq02sAIJ/nIq4HSrw/hmcG+QlHhC5brquQodt/gkOR4F9eOu0SCTwREX0+q
159NP6olundpA1N4xyXYvw7VqDCDTtQvcrU+OjtYtNLcKh6hMWi6djhnduX6uVKysDQ9c1Ydrt1w
aFxC1l31/LE41bUEzqc7VMvmTlRI74wPsMe2lFyHG8VG4kHdHfCO2f0+ICuxlREL2mkKhtGYvcxW
3EalIrCCT27Rg/RngAsFMxKD5xsZdfW7AIbRiVTiMXIzy9BEDY7P27PnrBJyWG2iifZSSzBllYE0
nUTnwybLp0vndPgI5BwSzuxKeYMZXls5HER0VKl+LdLRPloGn/Q9dAaOpQucnLXMRh/PT9l/Fx7g
XKhnGrECd4FlyOWLG57Q53iJqaLigy6Sa9JQzflmLZnrewMBGrtFFYcKvVOLJOfCwsfG7SKlAp1P
io9cZEKoL6xTE2MUr8naWELG8QXvEkAmwdEFFkrh9DLU15BP79ojweeFVr0EfVnK+1CzLz8iLraW
Z/W4Or7e4IDPfBijDz4DNbXSAOjdD3TZ+KmjNdX3xFieMQ3ZSvXCNLuufYEP9avRUGcfsiIpcrBG
CkT06vNZEgY+DJ10MbMrwczuPqTbMeqJDOZCr5cGkvVEB5unJvEEMqTpee847l8ABXqloWP3gK9i
iTz4oDxfSFjqs546uwGoDxIDD4HDZDUoG3e7awcJgEN+Yj31NaGYd9QUB1yXujxvP0Tj2+96gOmB
hGD0JeSNTmvp9zq+GxXL+zmH6J5nFMY8azd/l8/HoGos24kqSCQeHhUGRQ0fweiT1abzDwzL9C4F
JhaAP6TQvjfSkZ3NoRRoPgZ4BP0200pgubzkbDWRV6TIm/qlfMgLgU05DmsIOp7kIWYg8ampqrw0
VFk9NiscInOy3dPG97nv20ezyp7Ch5Wct2ITQGCD43iS+QSthH7asydE4v18u0SOXYvPwc88xyYZ
QMvZdKhae04qCuQOHiZjKL1m515Jyc3nExj9/J2VH8YLkF2TrKQhpJ92SgI/z9ECpy8s6IZVfSoF
GqYMLQa737ImTQn1JQus3bljK5EyG4KsON1fGn/2Pz1D8FwqgC0IeDpDai+TtrWAfsZcZJZ2C8ri
guGgPbbw7d2PvpsomfmOQWxdg1kDCLLtRHI0ChcLYzu9Tf6luosXwMTHMWqc++djS60vhRdqShIu
LuKxwieuJOXYT4/cD4EsB6npZiNh7PudEZU90XDCEgxOehXyuQqk7FU8ZIbz3RqFhkMBRdr7eMjV
yYrmGLbJ8MoTKZUQLnhjHhF4QRskHV4/pS5NHf6Ks96Lp4/Wla0IbF3edMCVKiaiX9A7iWz/VwVC
leTQJ50lqxHvPRLrU/gqEp2qLiUKg9xLwema7QLdVrfEDiCyvbpOWCq51OS9IZs63fwLR71qtRFx
ieABHDEt7YkdBi+zgkDSWOIe3hFbSbzVFlVBNQOifsWxTB+I2zTsGIDV5y/kqqWn71bIJ2dGFNdI
FEBYqzs49zFbR9hxPXaRZfd4XmRySSSREWWjRDRPrF25rq2y9J1W95I6vM+HmHIlP4bb1C38Aj4U
fIYumfrRFjiyRGprtsIIKUzajdz0lpdSmc6gptqn7UyM6VXKyuS2YSrGvDeSzpkrxDyF87HPgW0N
5ptW4m/YbXVNwieQpYvZMqfOo/8H5Fn9MU8QBkqPu+Dm2aOY4SduP5dLNOZvGJStZn5qLRdWud8F
QyXuSJ+SGuSuH064CrspW0He/5OhFsRSbWpPDa6WOjq5a6Q7v3gJgxaD7aikKXEcbVq5+Sd03mCE
yKuMvMbVPbseuTnwBBUVeViSjeEDtK21CgdFZrhwxCg+c/f+030+hYfKu1ezIKvBRCpiia3Q501l
El9qp6fsczCIbj2ZyjnIZVcwrzmcceREEPio7ME87B0a/f56PXtj/DVx3y748R08ELUXRhcIlZGR
TBCTZPmEHUJoDNhx328Fbx0tAo+WCiD0G3vF/t87Ug7EGJ7VAnwwpyvGbk5ifsj5ltL+z0Nu4qy/
hrVtyRggdxqEMRkol8Awws3NpZHZUZBiynlW+lDJ7DucOr+xLqksv9jOMQp9vCrai9z6JgysRG15
NdWemAacYpMejLlewhUTwUyG6VvlT+3eq3qjYOZc7bbtgSnuV0CYnzXBUamPWJWS4Jk+6jUzlg8F
fF+BvJL6dvfIxiwrK1HxQv0zDzblG3wN3yLnz8q/4F9qT+WwiZEWoCycDnEGajNlXVozUq6z2RZY
eOu3clWaPrv08KcvSjil5skl1JOZWOq7aRVmW41MPf8BtQu/o7YXd07WGcd21HFKQJZO/RzO9vJB
CQGVm39gt/Wmh1GukdwxYFoX1/W/4tTxMmT/TabhrfGvimBAFQwKJHVjHyzBjtCTsHxGtuNU7z2p
HhxmVaDPGp9uYRxCfU3M+mE9RfRBrqAk5f9tVcAe25iQSPmyZSyX/aa2cNLrsKfaQ8L0kWQ5Z5s6
UKeAbSgzQFPznLAkUor9ZmYvrwCHOs5M1jUlsyyRgk0J/qOCxnKWgEYne7IZAbjDtRFZTZC6ySZP
rjZdlRuNs1r1FODiaum8z2Q2Igy5hknYdDz69ZIDEvMncu6WMM/9ZpP1E38gYWItAIkZxSrZKN27
IfPMfCpAWFaWODNw/BzthfahGv9B5CN+osQFfhnaxt0HudF1X7/2ItXzmYw7vNmCVOiKp5wV1w4s
lYDF0cJDy9fVTxt9SvULYp8wGRxMe8+reA6IlRyXsZ2cG5MozEE4Nmb4CbdLcK2ggNQYoaZDLdD7
rUMzdXJe6Xx4DzTB5n6Dyxt9dybaf1dzaDdho2S5yolzpNC/vIK6FMbjx471qVHrXF7S6cat2ypp
JlDzpDEJcXfO3gLh5n3j4IjeTeHQ0HtWdEhK3ctSDYLjCLLg5zZlDg5pB690s00H0WGYUak+0kVB
LZhHWrWAxBai4/C7yePlvOVsHvOhm5k584lKSTp8XSLlrsMWGw51/6IbHnKexYDsfys6gEZvvMkt
FoEwoJ/asd4Oyn+/I84IxcMMGTXg/zz6MhARssVdEhDrfJst3kh/gVS6N6scDlsLqPtA+0Y/gxFs
gogw8dLeY9agyMmpQvf/PWqzr969ePpmb7BygtwNjfDa5Tytf5k7dd8lNw0g1kzJs3a5K2BSkUpA
qzqZv9Uxw93owOanR3+htK8MMG4lA24qSTSpIQXXyJjFGVGVtcRkAxitvLHYYsgKV7OlfQ06N+Dq
lQpuud5ajNTg+2lPn+8CBHMIwmz8jogbNgKJKoBCMZKcqDmO+NPHfzkPYy8GxYUlCeuNv2tz/vE+
Lpj2eMtJf0bvxhoVKP1wpPlGREgAvaki3pwwMyIHGjSzJsJo04xRckuuJRcpGzgkX5c6A5OKCp77
s6wo3yZ13C9B5cWi3lCnll6hXOytIrueQIBY5nld13qpJkpAsD8ud8meBWn/I/LXK6lXwf7GrFeA
jGXjjLFO+soyrcCPUHaT3jP6khgNyEpHgbsRR/5xzWXwXzxaLKII3nnLg3mB6K4EjD9TSZkLHALQ
L6EpQqKWfXqgAB0PHNNbPTgm4o3DSd2NL4dZExdu6xgZXl/Csp36/6op48SdM0+u/L8HmyCsxPRN
TmDAg0cKN65jV05cyGp9piHCpx7vyFYO/CFakO/8ZwiVsaynNAdhULdE23hkuQOmcexLQw5FvjDa
HFhYVOfu3VY8kNkDQDhJryy3yGBe1TqwF6Q8hmue82rDfdw1u/1/08MXY2MK4uefuirl3M1dz2Sx
6ayUw/pnhJHp2KniTwNmg+/0JJOV4CZ4fqu9kp2LNrw6oRyPhrFE2+q1nOw2bFRAErqjUEqDCA2m
+MSjew+EcfOBhG8NHCXXEj/2X7mHUU8DL+y7EcMpM/uqo6GjLAGHZlTLhyWwMiJLLh0N999SCenY
yZS6IFb+KJUu6q8spI3UTFYucLTwuC0L33lhdC3iIE9ppl93qGDviO8LQbDQyDPYE7fwP/kdhR92
nBKI+gqK4GUgLixHhm7K1NLkIlj1RV49WY6BcC1SG2dmqh6g8kql4hYFsfTDHKa7xBLMDrmPxQ6n
D/+11Io9Dc6900Ene8PM/at+zIOadba+tOVsklIv4Gkg4DnO/NeNtGZ8Gz1R2uE3KdCOG5Ujunbo
lOqh8AkmiO5QehPpKI50GmKf2NPvS6ofn5w3Lco6fkkq4H24tMXRSyBjXGYd2W3UGU5kwEml6BRI
e46vIeicMDcKhcch5oCSkgksMuVVMl+gUqPEU1T1EJ6KVmvnjDcAktbzZLaefU1Oce23sMZ1rWZT
v+z/eBIDIOpBlHOleCZZ9uDoM55wJs5KTpIXsLkQcFsRRu3jHHf+x1QHLcIvUxWN7teSteFD21H9
WcPp7x/xZbP5y+PDKRuHs1ONkeE8jN2nEqZMDyjv1ssvpQ1upsOQrRqgQN4p9CImkh22s1bWJ+Dt
rt0QbKFpHpen0KcQFPQrbuy1NHjRNZnKgQWZTv7xD8uRolElPIpmXP53kdOv1wzyxRCaPXuT0fja
d+gKItxW0W3++U9Q4lf3Pj5oVVno5t5oHMYdS53iOjj8EJ7w+5Z0N3WBTPQC1/kw+rwm4Ck6bxx0
MhE1rww5qQEBAh85JCwVnDQRnVrmQjBduWszBpv7NlI6GQSC4dFhk3n2ft8GS8QzDap6TRnvYru0
KUIeXJiKfKeMXkazXN1C7S9heb678xQyR7oiZrPCkMMLSokjpayXyUus6UefKsdm7zhwpeqt0GjH
lJPX30dCApuUZYAzFEjVGVx6wNHmnPjkjY7kB0UJM6ydSV99yr96Oe+ZIDnPcbLhXbSS9/hKX42M
1YezYVYDph4XJi//dMsZwE70ciPGadSDYtXBvg73h5Z4hOSvuBnfgffYWXJFNDmTLK+2xm22bcJ+
Jd8+5Ovl8OsvtjVkTn2AUeP6bpzk4S5oozelA0YzVAETGghSbo8GAWu8ZfaiJJe4OUqwf05EFkIq
TugrosjO2elVGMwpk5lIUSJY7TMEShz74rLgbOeYSDYuacbDlC/loGdnG+0wCveMaZW9hjHN4c3f
jKnDCCLeIi2soKpqlzrSb9TVK3/2cSTyYn+xD+zW1HpH/xPhsvX/WSBCgT0N/qccpLeijq4yrUDS
V9S0EsxXzVv5Osvrpcjz2gA6/DE/UcOGpB7hrqqsX7lVjGL1/CUXwkLTFM+XQx55qwDzCZyY6vQy
JyoZwccr+9Zry2MDGIkXC/+Edr6XHOt36GOqySjHQWEkirODfbufN/si/4NJ06Rh2qFhF8Av1h4i
rKrLKgN4z+xXAjsUiwZLkSaUkwhSaZyOgUSvNXQeon7U7JFqtPemuLyjWuWoAZYGMH1K/8LKRoae
sX25TciND1rW1osEgQaPDWd1PBW7db6Zd3cSoVNXf8FkGTX2jfB3BimzUM8JfdbQiPST+MHgtSi9
o2EbMPhJ/LyfReP6L+L1g4TYyR/QdYSU14bE7zg06um80XhU75gVKYDBohUBqaESxVwufX7YQJfJ
u5xuFBG1IpDpjQavcJWoUHqdhT1l+pQNQ9zpqe/hKcdzrS9kVbm2443fOxYQE7RXDQPnEZUcXgsy
Yc+UePo0Eog=
`protect end_protected
