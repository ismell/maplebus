`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WWtJI+hY51PBIHEJuMmabMx/exsWif4/+eIlqg1wHwt0LXqCBCF/9KMUuh0c0q1Aim1AelneHBQ1
OAUIypxCcw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LHWPiFER+ylhKASKVb/M+rPTiZEUFsSoYr0JzoMMS3GVOGL2OLFeqOogSRZKIElrPvU6koRPo+Es
YaV4XvTWQrPYaKRuwsx4NBG8Kxda4juxxP/rp9bkfo/lyl5vcqup7qHmHWRkyViNZaKDThZeE3RS
GK4cirCmiwfxEo4Mq3g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYgjStfBUMWeU3jKprSUnciTIMZZPy5txygzDux4UChegSEbbUtF3rfC3SvidfLEgr0Xx5YrKuqi
8UeNbGyLgV2Fztb5G016ybd926sP72A+bpKraAlbcvGRolK2h36OEHIbd1QCQ1CK2LHFu4yijIpu
ZCVGSRMDfbCIVdoIEwi/d3uG3uxZJ/MwcPNEV+U67K5AP1cQj/MZSgAHfDEJN3ny/eyKwQLT0b8X
VrJgv+gHNlk5pWmHGp1jOFZV21FW31bI2ureAimxycfLq41ciw7AJu7ntE0aA5znCk0zlIOF29Wv
FVMB4Roq/qxMuTuLdNHOyDamSc7+1ymlG9PNwg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IqXkpA7tC+yxdagm2gZbfE8KY/sLSwkzWYcxkLkeovhP6k5hwXB7qgBFgwiDFM/bCJ5ScHqOq+cZ
9SW3fwNmkWjldStW5jyx3Kj7D4V+TZG/OyzKcMcs0tleStvsDR1qcGkMdGgwTBnHkIPkC3uG5oo6
ZM4eXtEq4AXscq0m4s0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QQXOFVhuXbc80+zZ2htCYHYcCp3E9O59+Yl7ypoRWeIoCrrKiW+q/IshosljPYv9Rnj61yuPSL68
usz2Y0hE3ZS3oeK3PPxnd7ql38jWr1G6pJ7M5hierEefIrxu37p0e1dp9jw5djTq//qZTj1uTQCY
59J/r5hUUP+AP25sKdsRw6TJVm9uga7G9srmPkRIdoLPPfYk0yF5ajnsD7NGAlmU80CKSwU00Ofo
u97sna6z0bNS18cL5p3mUTSRYh3EhR8yWYQDBDVfjOUeffgGq5Pb9Fz1RotN+JuUStC+3C8AW9BL
pf/Y9/KyYenDu5RF8gCAras14scTUMduPi8Rvw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
oK7CZuHusBl4p80xpwcKpymTrw5o1kRNzmjX+ZhFa1GtBqHltzfjdIMu7doI6T8t4c0tLg4nBy10
0J1w+YaOK0eaIld1vBoTsq3bRC2TL/FGTG+oJU21MsXdgGGo++aHGllNx0wI8SgNpSMvxNd1ZjCg
JMUPr88kMoirDuIbAqvxRo37BYgEPQfMmLxeSRNhPDfISFMED8rq6MDWmAwMsqikye0c+dw264I1
fQwVR2hnoPglDUwOiiFmM2FHurlKNoN1b8g9gflsQNYKMZGQbREN37ojBOcMZBSmE7y92M/qXXVi
yj17Vbm0h4rU34ck7WjS2/eo7ngiAOj7ptA1Q2VhSkntfbtTz3fcUJ+nk5EMX0c0UshPOQ3kq+cE
bl4X4Im4xJbCWiRYbfbO6WRXcE71+bwMaxvD9S7oS/oI3TpuDzcUjM0fiiH7iU100Em6qOc+Qvi8
yjQL68D6n0ytumZPcsEphe8hyc/l8EtMat1Fb13wwx37NDhKBD5VjIBFM3D3GEmu+aNF4/+K/cSf
N0RUQJ2AOqB1b/aUGUAwxbGxAx2sLM6yzYC3mZqwtU2lwKryGVNxplP9QgziGaQxYffra7J3xq1B
rf6rgJbkpE4OAX08o0zPvLtOoIF7DsBWnZv6NcsPm/HYCj+H5rgKaM8vf5Bfq8dEC33UjHUfR63G
kxotSoTuTicsyWBtXDptqUMr1X8AZaZNBw3qHxt9D/9+yu8nYv0HyXRBO7MpaTo1uC0HYMmqII5k
AnTduMRrbJ5GdhIGDwNTDmCNRZXPiARr2fdl7UxwOnX3sl7EWcZO6L2MctGrwuWJjrP4tyC1L814
KNFnw82CLs+v0dj9vQ9xc7Ep8BaRpTry3A2zdDY8Bedfuwb085qqDzA5DA7rfYvebH5x1tB1q+c+
KNcoiXOOvapH5fTDxg1h8oKA0gkC4lgkWXro9wwRXQf6/dGQdttbfQgILGzuDf1C2H+rjgsfr+0j
Mz1YgMd968IZmBsJ/fgmyO8Bzh1km67LgXuDRSSOI3IOhoDeuitGCbOhT112pgy4f18NwECUf4I8
pFPgQLQ9EmKApBDhRD53aeQeaUXZCC8EyhaT6TUqADlgoJIShlslwcysLYfSOzH/W/DHKqIXBOou
3W3s7HpdMvN8UJiVTmeIRLrs81vlI+75PlaYZrJjbZs0wtcLqYRdXb+qMVWmqwANfiJqn3zPcCE/
a1l4lK76Dhk2VHVjCTPsPILwzGsBysPoZlwLxKUm6hVuPMLi/zIl8QvZyH/DAwsNbffqv3CbifAF
28xnpGwBuoxxOW8C07rJ3Pk+MBvCIyXRGTs9ZMm+XIRGqp8J+ecb1qvaG5EatauiDazvw/QQsdsR
jXsb1w3vQH/R7MnfZJSB/gi69O5th1OHFcpO004VoA16GHIImZgXAF/26bshmcdlcizQXH9sfSke
oIj+yP+UR9Ix4EKd67P0x8uFag3v03E+Lp+kyCpqxh3dz95kAXrMSYaczX30s+TjGHriTNF/Fzlc
SpVcE1OUdN4D062mqj+HT7kb3VE4mNtK6kVksbTKDv86Olf2gDS4yyk9wAdmzSW4wpc6ONpUZcyH
/IZTJPn3/GLA1n42/Eqd27PPZWnR2HNWhBpT36TS6WfGBykInNtOfIECai2WeKkeukD3zTnBJEt2
7p1Bfyervii/AyitcwibBBxS+i5VTyYXxr23oTv8HPdptL2VYTTJjkiB8dBho7Amb1wq8rh33mKg
r9C/jN/ticH9S4GP72y3NlnXINA1inAOcGP9YArsGIkci71MINlIAple856esMWt+vdhdaO5WXXQ
H0LQ/DrAOI5fY22LFveIcDMClhD1Qkol8KuZlRttzGpj+aXtRKorYjTsG8x0h6aCfT5jzIBaZG3C
fJhRK8fbg5vqY+NPebj0j+sGdNCqaoR2wcTADecn2d5bKUWHLEj5JYnoeks+SKVIVIsNrYX/YRGG
cy0Yr59KeQZc2hWsJ89YajDTi93WD78tAMI/RRAwsldj0FWupgmvzk655NI247uW0hLzjSbjAEcV
fXQdB438cDS8hpMSmfj1P7dGP9eYOERhQQlo3ncAvDoxXZQcqzp5B5dn4C9n4q7m1IWhbe6ODM0Y
L37Yc462nVgTcBT+4eVS+VLqAYlWTqEAllzoVFWT1MXW1in7GBjVgtR4091CmTwNcZ5zvMNfUvMI
xOCcyoqX5iiVD0TMca0YFJatS8ssamEUwhRJw9OAy7I2c8RQy5v0rXgY7dYb9F799S/RvZOHQenz
Hi82DX9anD83gVUGFQMNy/wWVcVJcoFcrFwgOtGNkWVdbjDRaAMwRg8LKeMcSASJSZGsDUbUygZ+
tcnGmePJTdJFwCjHO/zhNhXnYmq/rvbaOq7m12vrsUqroKY/FIK8Vo1OPF7TvMl/0kswm62pTCw9
57ZeGvd7njFmj6ClUb2rsa2mTmHW81FpxDsIl2Rc7LVKk9judawpHyioeoJbPpnfK9fSMDoi++DG
6NNKikN3PFXMfpj58mH9AhAym3CPYkbHAb9cE29Hf1gJ1X2etCJNK7i9CRU8dnNknFd7zrC2QrEf
l7BV0ttsAprnQkkeHxpZCubazUjjzR/M/arv6pMo/VUzC6swpuJw6QIsysUJ/58qzDx0EbsxLBpu
uam/1wm4JDGp2DpwA/vtyV+40iIiE26HIRIk3saQBKQcpQ8oJb0oRu3WPRc02alKjdsD+OvXfdCu
cfKcenhqCuUBcO1m3fgXhKVLzIGAMbINm5NNSK2jtho2z1prW0Do05u2k9eeifJUQ2WdMVYv9+Gx
IKTs6W1t/G3mUysnPA1RXCHQ347olalRlQWOxetq8aqSJTLQIw64RbmOoOw/LD8uTBF2VytbnZXy
74Cbf5W8ne3HCybAC0ZZMUqRlw4kJh58D50z3hdU/MWmxY6dSRGgrW/cDWy/KY/S4+zNYONOhb6Z
+MFvm18oD51gdObBk2MpcU7XO5YZLdwlSef0ZQHdH++AGqBnI5Zm6ibXT65R9CXkQ8Ss2wjz6bba
IB6gA3AGh36vy+xbZ+SiEoZc1rCt54mVSkktC5i4fJz9cuX9uUwdzjT5tn90mK22CIQVxtJjDCMj
pMtDBNFG/U3hr21JxeliIPVEmtCTQhFh86fZwr90WBCdA9JBaYWhaf9kRZyApa+c4MbIHbQdx6pa
OuGGxHz5pdCPki8xF7ZkLpfxyKK6l6N01XHVuEbXD0kJy7yALXfLAYvNoActQ9+6oCV91FFssFt8
s+Rz5Ng/17MyO1aBow/DzwFch2UhCoU1z3QzbNdb2oEKZNX1GMhE9+wOovaCMB+E1sSWZp/0w+K7
t6atjBUTvWNzzrfaDJ8CkCertEdKjRTK6+9OD/cxq0LqNH+I+lzDDRUXACzkODGf3nDep0wYEUSk
irdDxTge25tOGANzIQDxCPy7yT38E3EzohLUOksYGjx51SyHkmitQCWomNy3jhibulMoR3vrd4aY
O6nDC7VEc2M6LDLx7r6ROT9dlhTPIRFnr8iC1wc16VS0neEgmTxWgXDLSBAvw0G98XJ4glhh6V9K
hJOzBK4uCNDkmAFNmrG4+mCwxKfasLyPSki2/7CI29VQ48BMeUhEqEE//YyXXRYGXq5be+1JrUjV
WfJ8rumN3CHo4Owah/Boo3NeQhqi6tOiRq02htjd0GF9Iccg1wPW4V9OSZRXSV7a3LQbzducZR9N
AnJ56+ATTF7byKXvMP3ufg5VvteRPnsRlGOfWpg3zU9088L1CNEu481tvMt6s9+COnQMLycaANxQ
H06tKoemk5hbb+rRoQCJqD2uUGIGK0S34As3FGNx6oIVduweSNdDtsD0Ksn8dUjBfrewABFfJQB6
/zMeLzC3wSV8j184KKh1C9wsX3AjMM5sos+a8C2tflfSZLim15o0lLhgbU2nu6uLccselSarh0MS
P+STtwmqn36MavzbU6NbVuGCOmY7P27YC0YfPF+2nPlnEKaTDnPgO00k09ptK41dywtjDLGVHW7j
DnOAXU55B8WbiHx2U067zLRBgfulm7U4MpDyFjfAYoUwr/8c63CtTGRiLyhdri7N7HIaHz+eRCJ0
8eDpCcGtg8+YFkMtTxXAkEtC/L/NXkjfXTT3PBK3/VgbyZwQZCm6pzhOfZKj3i+3XTGU3jL8UO76
VQrECPbLhc67JIOGutCPl4o1o76xdGao1PECdnLvLvMrJRFVwjXJYJBx/o1NjdBCTaLC7jqFTwRm
xR9I00PCiX7P5iVVFC9WVodNARTnyfyuNJUkpRzEMU7nmJ9/OzxpHP7ZKuIuPZjD/8IP8YxDGnXB
9ZbYNInJazz9PD18jKwCQ/kU9P3qwHnXElGxLN2qzC3Y5pK1n6ZTCXxjfBdOPw83vxktKwSde4wM
zjXOYIBe8+6W+v3WmTQflH7T+DJ3C7TiHpaR1rhRUaYcZum9iKD8ElV96sfPYQededXy8zXrX98w
b3+ctK2oF4kkrSchUqa7lcECg0325EIv2+4qwMfUu6X6kf3p5PvkCCnwwf2TNcJhZyd95qpPnKj0
2j0tO4SfKa7zxrmcpXqhbVlp1CdN+Y3q5a5FBRI7LDCOadYSiuKV4rFnuPZR0upK4OXnhZdBfdq/
Znfx65EvbdCfTe7kM4Y81ayN5zk2J/Glt2mVeRhs3XXn2wxgKnRIIkPiLgCI4H7qXiIKkWJ3A5OY
08YaJUSM6L8LMxwZd4l9lCDw2308oNpDThVn7DVWizerHh4KZuwJtI9JRhhQXF0OhbUK6SxZ73vd
o54raXky8Cyl1yAcySZyzN9aP99X5w6uiogx4YIY78QllP2d2xP9JvlTdJid2xtivt4bGRv6G8dy
iL+ONyry/6+f8T8KNDg3JGCvyo6WB+120iI1lZMpgi6ur6lOiOOA/bC2zMvEuxiPxe9L/zhVbuxV
IrWztXsfHotqYBpqn7PQJXTxz2z4CeLdyTf3LVWMb5KdZ4nobZIS3GNGgTjPdpDk9RBIzc0DCSbL
xsslowZ3lqPf8A1jU2IAxPq7CjI20kDVvY9DByfiyo21UuGQyHudYPCEwdzjhXufgvODNraPi/5C
EIRIYD0laX88L6D9dh8xxlpjcl3bD8b1cuVYsUOIyrkkDffTQ8bTFD6NvV7dqgU+JKfdtNJqO5KT
g1NBDpG6a8oGhz7IK5FZP5yg312/hcOXsNUJKenubHsW8y0RNQJoVdqCE8nHv7O0rQqir8sRdBVi
vBL+dKbzMcY3ind/4R6wTJXMavWQ0X7ATQdVqZLyHcTxLyaqe9JwH9mBWbL9Cwx69OT3puq9Qd6v
FwtRFrfxHzPkmfmofaN/0kuMCfGvtHTFO01+O303QzhzHBpRfSiDn1upjVYv5yK7gQ22QpsHI+X5
QsS0aFPLsDEajeXI/S8U4rp7Ob4Bvxo/jlGRyk20UONQ+9t6N2Iq0gZBNOFiV1F3VP1XX25oyYRE
Xph6o+26Ry3TQJnsdVb8vUomkawUxvhoKj+gmzf1g+1hlUkO38uKfp+3d4uBIvtOjrDDF+09vstQ
MqxKN3kMHNrSgJBBf2VsnNhMuFCTsSHDV39txhUzxflLL7G5SilF/MAHFplIEgsY7v7mIOpjJcH0
OJVwa4Fl5RemEhd/gwLVnng8tIHKvKwjr+DCoM/Q1FlmqLl+K9/Pv79fmFPXvHTFNBzKH7x1Yhqk
gsDsDY3GK3eosjAwLW0jGQfbzgANbrJZaOCQs+YLjBy+bSSpLj7UgC3KeaBaYxwIyrTuXDhyHxAH
h//hf911PdFgJWdJxu4sOAWM6TI3tVZKoYGSBbHeIBv4+8oh+njrJh9bu8eJxtThme6Ss9M3Y6P4
YqrK2lEs75vgykqtMBxVtLIPCZTilyLhQx2NMWxqenfwnt3CZjoOB28/pIzVXe7IhqPu+f9NKMM8
cLizf/QolJr6GVfBhrSc+yZ/rG8CcuaZ9xYYa/i50Q/Um8kFRzob2cK4k3hYgz43hyLXOP7uLkyp
73/7UXVQDuf1OZp2shm/RT/X/yT+EYxYDiYtJwQy8X/A8gfhWxrWWGi6hiIAVse4DULMSAIyqlAm
2vCBfix+ZGz/0AUMm7AWZukPp9kkpJRfoA72xs2CjpHennA09Ie9OQ7EXdldv3CgB3z999RYfrrv
ZnBsu9ttKRfob/FVeWO0qPoqskwNHWGNApaMhjJcODcMMvFSqFfjKOFif/XnTudX0F6v3JizmIHz
W8oFLWg1bR9lAAxKIWOuqUo8pgWFUBXz2avopXLv4DjNUhNH8iAUrOWUg8ajBWW0QcWetn7OTRkM
4HcmUJ7euvyJ5OOrkeib20DGr8h1RyVLVeCMuuXSKHm2eqpFw07JzFkSiIo/C2Yk8bLCCFlY81fR
as4wz0wbwV3yghSW76gxdWPNQsdU0xjjcWJ8H/LlE/B6VriveVs4x4QqKyNMBFs9STMp6RyZUPeG
UIzm3B0XjrwZdcHf7A1Lwp5WYpltp8GHYYMC0eRi9O+h2JyOlKxJJGDbZ3EU84rVxkr2XrZqLED8
dSpAL+QL5g+ITFicZRts1sTG/rMT9T0K7L2x0vPH6i9g9zZMtWT1mF0vFsUUdirTv1hw95A6UIXZ
fVYeAbx3h+lcZg8w+z3lEhAOz1k+ckXKBVdDMOhlAWGTIzavnKGfz3MGRxtAXXDoJgVUBVMymR8g
hu3qBPXi1D5G/1zeQelLgXNomx059bhVsYzwZzbi8FsrowZKBHvVW8YrfkjPSeI9FyeL3/Yma7i2
6Dni/D1mLe3rmFGD+fUsLkDqolWrQesg95qWi3CU08OaDl7A/CB7DDFNzpTC4d1jNuf8IKyR9BBa
Y1PqpcpcP6LhvmnWGmvHMEvhu31eowpT6LvVJfx31oLfPjf98uvZ2bS2InG99k+QB1RHc3OMiLB7
q/W1LUwnAkrtykaEqbfHWacnPOEXeis/6HEdOUM3EwFOT4AVQKgOCP1Eebs/CEPX4gSnJhGTIsLY
1ypT5OQeIwwjQn1Ap1C7RWVRjtGrcpERJ/k5aOE1iPbA7MbU1iqk33cnhGTYscNeJZnjQ2eNg7qA
DUDBbkI8J7ggjoN2s1G0a5P5tJWwAyxq4xZ+OhqpGwSX8RXDQLnr8Ylg2PMURNgjHRHgW8P6qrqs
6lHijPOeIc5j88TR/C7xVu8Pgr8BbOafuucZpofDTEXM0ESRTaaHjWsefqXNCQk91T0r3XhZMVQ9
LvZOf+wpY/TPa9n7mExyGHy1ECLVs05Ig3ajpFbXktORzw3rKWLc8gPGhZDpecOMAZ4b4vaEy/NT
qX8u/8EOSD0Owj/5KkVcBQcJXjcAFSekL4RfU5anArWol6s0qKVn1ceAL7BpK8OGOxcZ7HRxf9n3
5VqsjWqV9R9d7gmaS930Q79ZnWLWbqP4yE3MBziIOAFGBKmnzdi27GSckDlqq025L0NY9ehEv11O
XPURF+jaCAN5aanfVKy+bL9WDAVdOb/wIm6hZyMcjenDj1V7VOpfDZc8q5VMGIkaL7iRpx8czQUw
PqlqA1AHBXShOc5Ql3561oJn4wghmkrLiFQeLvuZgR6A0RXQmYdvNzpZdgrImEkkWnJipuWFJoMP
NAD4hbxoSa7W8Voxs0u+4uCJ24v7ccQRtmfl8C71CuKEzS8gcJMuXfUMWVJwBPedTapItRSKy4ML
7BFQl/Bq8LLLhTCANtMgCMCMV4hTSOGRRS0FCCW5h3jAPtOVC0rulU04Do8BM9sfanaVuGO3Ojd9
EQRhOEM7ISOLu59GEAxV88aaHLz8rPDg9oZf0cbjKE5KLNeAfbMiC76idyfcRjqYIgzmngehFroW
dDTm82KAYsMSNYGLT7F1cCOO1LRSKbFJrlJalV+V3Qjj+CB1HycRk2oYJEV6/aNBAY2n5TAlimrm
IAjzDaPgMAsjQs0/953zXoXlURX/5xlzoYD7osldr+wH9D+B3/6LA1Ub+KssNhLPkUXzJTjXpa8g
lW/CssuzVbDPP7M7DfgO+snEJVeHa8lYVDXYge21yxdkvM8MFPt2D+WHLDKAE+QbEkoFVKgc22Ii
eYiZUMpepe/4aPGx1QaEZ5gLkUxl9qD5du3tIUofttXcspJfgzZdmZNp7RUpjFCCvODK+IxjSg8f
vfilSuCl/Kqla586AvsNc+/YJJ5gfK59L3CC9FZWRwcOeoM6Rstlx2FbEmg6UjpEzCDRoo2QUwwg
YtXIpLZgJFRThYHgUGU1QM7cymSInieENdkHXn6OpIktQ01TDIKQ4WPwXCOCDAW3DOhyTazXDTZx
mG9vRD2rqt4DJVVXumqj1cWeMOxzOYraxj8pF5/Kg/O5BtowM3HqLoXpE4vXisqBGGtMBPhdG5s3
VdYg2fmCrBAKSF76ctsBJCF2gIQd1u7rkmq07FEKJIX9Jy19mr4joTk9R06GOFaOq4RLHAkis707
QpbVK250XOXHyF9NRiDDcqGyzmzfZbNLjUwYCaJQhtBGyI4vWr3e32/6WajMsoP+VIJYbv78neHX
W1CI5ruG3Tnd217ydc27k6CfB2r0dHlMxKqLiNoNc6vOpeqHXAAffLkVKR082M/g0L6RkBF9krbr
VG26nCzeUE3Td+S0Dsbey5vT5vjvYFU55CRddxEQUj6ABy0uc9ihE8mYONjsysifrBH4ChDb/+iR
pyILhj1WDaWEtL3UggCgSzl1nL8AePemY4VvXuqikllsYEH5yC0V5yoqykql3IxwbUSkFTV8t6Wi
fkkjstyEc66mV25npLSNefF6KJYNunWTo1AmaBKbnuclW13jvXSi9/GeP7MPbB2sei9NrdEZkj58
dRSdIuBXLSQi4NYWgOMbUIcA7uQ7/0kwl19FkVfmfo8mfPq4unua7B7FEqQRTf4G3rJlGabjC5sf
Cdymaaqy1vopdm8D0p5owXI+9TU9AZwC1DQTTx6k300LfUPk3rFNiaxDtskpZqNxPaHTYQgoiNIc
Q1OCicNEF/ecz1k7/q6gxZinErr/49I0RnLt0VtyNpSAWQDAPuxNmANs0FIR/fVUMvtEQuvjDzf/
bYbSkJnjmUj58LXqegBqXc3xLb/LDpeRPUlv4f/jjuMaSrrrS0YX8mB/i/HJ44qhrbnFLP727Pd8
eOn8nHpyAqNXjuZWKe+jNnCmIVtuLqPXoB2dvcUOq6OuSP1Jp5v3fPcXohiQXBbWNQM8tNu1yrvZ
3mDPlUtYJLBwv8+wSKP9FaTLXMZ49l6JX3SEpP1mWcej5VbeJYaA7/0JyfLHr/NHAXFsCm0Ezy6Q
xo4U4YWq3/sg8u7yOYcPuNCmTI0cynbPL6KHSetOA0lRgKx7b5gOsVO3jPMw/Vjknzo/5NBvi78y
PLPoFK8Mi6Qxo1vwztjFP4KEZU9gFjMB0iLbbPLL3PAA/nvFNEXsLzvhX6joDxhFpXkJxLq04+Jd
Sy866Rn/C/z7/jLo1fR7G3GpBQeDsYgKErl5peZrePnfZEsYdBcjWdkHYxYsPA5twq/ojPQ2shhR
/Tc7MoxgUPWv5RhPVbJ4dV2VylktX+XG7i3Q38cXN0t9Usmcg+2cS9B6hEOYCXY2DlyVQXO5pn/D
WKa81TEiJYq/MXhcq7nweRcNLaUEOPU3W48m6Y9uE8KXXPEjBe+L3YGGVrYHosbxU4h6VycQNxXE
dAJR4tnrsGZa44Eq1rJDoUDzF0PPH3+izfyEbmIFfIb957NhUJPVS9EdoZsOqIp+jmumiBRfxjMo
FAIJa6h6TdmAw58bOfAhNm8/5LQ3cTpnWhALNLvHyNpspMl/c/X9F2MUTh4zJ4gizHDL4hWtX2UX
wyES6s71r63Y7dKd58uwkImkZfU5RuFxSK7PNuWxgqtVUpDUJt0zy68TvDhclRIfE11rRcmdaVSh
g6Rg0cQMa1GRXANxmCKRbDnrmK4CPlKAcwG1c6N/pmfFrhstmkzxT3bte/+MLDDXmP6G1/695x4H
zeJm4voyxOzK/AOB1+JNDfK9i4/EPLP8wDR0JDpVE0y4wJbwLFegifNz9TzWOyLc/BKBUOTdLrCV
0Tlqxk4f+XF2z+9fu10jrh0eCqq5z3FYtD12mYN0+K/0Vb5LN7Kwxzb00Mjz+SxcLRplhv6qoCAV
Z/2qPioy6rLLVXOo0A3t1k9D8vnistEUYaIqgImCOLHS7wZABYbQ84T9csjB/a7pVhA68B+R9kY2
s8J9CEvWfDkgh6x2738OeTI2V1wLUa7W6fK6CbnK/OKkP24MRcKFiW//FuZCMM0UpmJq8gp/H/+0
GlIiWMeKb/nUj6n2Ah0SH4inYRYh06eAPfQ5Nx1DGeKMnkNGRUw8ObwUxbaYmzfLab98eQm4qpeA
UWySEUAw/gRhugu0klCWYR6rl+pBdcWTAl2/FrPi+EvXVx3Yb/g1OP9gGVgzqTN5ovimh73Hiel+
63UJ0RhzwT19X/1zKzlu8Z0KxX1XXTHduEetCKrQ2PsNvGoG54rkWMZlQxUKM5FDLvHLQjmpziV6
mih+RM+3aiU1ELTXpVNUGEknS6lcp9l5qtrhlT+Agiawb5+PZSAPhgD4QKU77+0MFv2QkIvMvvPg
VHaRGrYXryWjmUAzAU4XZzLpKGpwpBvnZUxhq3KvSFwnvCD6hMgA/MkwALlrn5tQcOGwLFLz7EFP
Yyi17FKwCf4RTwScQ7fj1OjRMUkYvicfCBJq6llHkHVewcArKKi8fz5/fn+rtTA4HRr3J5kyHywe
2V/sJDhGHEnl+Fflwki+PPfFYVcrPkLyX1D9YE08BDD/P6nSn5e7gigH/Y0JHcxBEkkETtvSunoJ
HAT2MFq9TWAo+SW5UDKn3NKGe4hpNjPMwFUuAtiBp7zjZ2e0i3+HGyUE0WJZImBWGdaL8IWxV716
N8FWquCjJ9M7DrGakzJgpgTehvifaWhpZ8D609TIzOOSdD5RbAjjwN/Ch0tUorKBdCwEvhj1jcIC
BoSF4eH5RkyZ2PUN5DHDrmdBVD5c13m7cXhVznVTBsFIPbgqYyoivhDxpvp3LkHJOPl5BSPiCeg8
ksqfftrVsoCfZiqHDogHPiYIpvzcbfmfISy9KOxKjCCqbSbUrCsfiaowBrNsGQxchj37yLsD8D4j
rh2KxvAGCA/eo84+seQeEoLyl199/hXv/Epk2H5EdvQjYWI7VGNfoafHjPWKQaZGThiD/LCSERt/
NNKa2s9CHGv4XGXWPDS8oF9kF+ZJ3nJ2rE1ZYSIwbklBH6P3WJw7OBFX0XVHX8nWDMmxsg4U9e3G
jc8RiqaAGBfbOx5fTbpAyFywtt7iQ295O0ib/bGCElqtKtRaxjp/ZlExme9SYOJTF4OPK2z9wDFB
7U+ADN6zsGl4M5U2vHL8FDwCkZ5YQuPaEXJOLG83dMpSd00h6bibBtE+4+4Jpb7FP7/5N2OqCUd8
WIrE2KSf8y5/yRTUpUyKeReSmzNI+cc7ewQ3FtntVSJmAItQAflwETXFtmPvmOIMs0N3pGCD5XSU
bMhnIvA9wYI+agQYgPDsLGLEu3S1ejqTj5eupzlGOPo6RIiOvCEtoot+/7meFAN7PVLJvlo/zPTI
Ytd4DxHrtDHAFhdICfatvnfZYV83fZ1s1UmoDujoPneK9hXZL0jcpRxEfL+c+0sDBcJ8OEIrLKYs
k1ZZNc6EV7DZnkCXbDodVmxyWj09jSQDfJfBGhKQ7AfLOsL/E/VpSjwrtuQQZevWw1Vc0xX6I1X6
2sR+wEQ60d3aJQNdi5uafpjCLdymVQN2nvH6aySZCl2o4Bka0dT2ZE5IOONHzPjzav/4JabJHvSp
8vlS4Hscgl15tzj7XPRxRkGDFmU1tvzU42XPeCvPYxrkH2f4XFQfxg6XeZAd2pzeDYHCen28RBVO
2yCMIhCTOGHzbnLiQovm3tXbLnxStoE33SFlywYsFabaE/uvRJ32GtMcJ0bmEMLy0S+P7GLU+flV
PgXed9p+KFBawrfJDAa9YHipoCq+zkloTLDJ+0ySkwvuaedxNnyYm4aI3yny9Ge4ZKImwvBsiETY
F47s+yceGnbkW1k1ZYb7sox2TzLTFXdKCQBCPUnrqoFMsg+S/TJkXbSqk/J5zsclBh/DkGvZJo/G
PI6nh4iBwQeG2qqSQh5HoR3hyPm2o2MoAQ92xTAYpg4tQ9MViAB920WZeu8miETlKqQ1Vaa7fmsD
ao9n2D1fSErYrCGGcuIkTUQijjluuj1HbCj47c2ODkbgh7kHI8/VKceu31Sc6EgXZZyDCvzMtvUj
VDEt1QiO/5+Sk9vdIZy2URsJO/SIWzlE2T9/2l/rkuxK/XuoZ7qgipvfnuvFd3Vj4Gyv2LVq3gid
P/vRu+Tl8C3KptS3IQd55SnmNmLwgxUdk2v45tkZSfMwb5SqaEVPJvH0/ZpqyDoNu9TpZlnXAUDe
QOsIxMSWq+k7o/YQu0dtR3Rt3v94xHIFXvnYUCQ/7hvgm9lCa33N5Q/AjYX3T6ynDow+kJvuWLbR
CJZ7vqCZeDUORoESmkYSRsL00vj6at68dTRJu6C4uTdkCJ2XlALh/KtAX49OD9VCHwie3yktPl7Z
gluCOsNhFTXZgWYpdxY9B6KGgAsXBlKQXP7EGt0JE5xOqz25BiGjHepsHP7lWG1BR81xSkV49KE8
Rz7kfltegH8A33S/eizOplRi+MjC5iEgZmLbiyZeqNaKPc3BrqEY3+rlEULuGUDcAOVTC8Tg8oet
xeYLQpJON59WnM+jys8YzSaEKWSaIcW3aVVRgCVUIIRU1V8BXZlCjAZzePH56QDbcQaT54yAZWiV
ENJ+CNOmiiRB5RgaYdRfeJZvWciNnNccsGeZqFjymMKdcyYSCLISNx54vaHDk14p/qOa4gHV3U8u
RYkGkmCvGahIv30Ax4gIg/JlLG4tEfEf9w9Yzg9maqUJStUi0d9ahGlP1xOZEYB8EikxpN94ASG0
SWiQgtZ9HC/nRLZkC8IEBKEoRPQodyhU1n7wbu8y/GkG2TcB/a5/Jqz/NKwlJe6fIgIoytdmvkzZ
0+Lq3OGcS/Clp7EZ7iYpqSLI2/0tWrcY1wB7uwyHGHzdvdrMPNRfbjAEDga7LAHeOrEQ1SlfiCAZ
NcOcCvgcn7ebV/C5ugjnfZqaeJaPzrwKls2ctLipDjiqKKgWWq/dG8ces99bk9J239Vo4IFfnefE
BnHvathp0bAGGEA/rVIatd1xJqbVtFYID/M0B7DF2MhwhCj2cqRTDbsZY+SZy+ekmCQFlg9bd0q/
y3ZfWBJ4wBd5bboRmiy6K7GJUoBXtxMVazWPUu6qsScZAte7hsdMx4pXhhlNBsIQbQOkgf3M7yxV
BrNRFE86rMu4QfAK6EU4D3K59cfjJBxxk3P5dtiz+EKvwB418p4YlDqddeLARMHqsEGrYDrGX2Gj
92g/i+7DMIjQh53qleCA3anLXk/qHyomLzwKUMdxBduNnmySe6XXBj9YrvTbwvBvPldTFn0AEjZW
cpXfdaY8A3yZDzlmhoKIUadytOhgAnmyVNkAjYS4UWHjjO5ysYv0/nj6EL2ykEseIPUVm5hg6k65
d6N3wEFta6LVlggB+gHN7et/l4xSBJqRqPeWKIY9M/uSJZICR4gUnYG2Uw9o2YVbC+1J8dK3mjXX
mIm5L9BioiF42/5HEpXjB4zi/Ga93Krcz//hBL6TM8s57wobJRj8jEZvkb+ZLZclgUHXT2TEMe4S
0mmmmxX+tJtNjqC+olEx0Y3ucvujd5YEQ5Neff3S7dPj3/5jdMWPGndUHQ1zTInhcqukTta5/w12
pyeab2Whl1aRSC08eE+OUgAByaPlUZirQ1pm7ut3jqOc2HQcr/lqjo2HuYUJY5MIC6173cd0BB8y
P4qkQj41UTuugZgU1dGHYxpKXB16cXirSqGwShliR0gGRH9EVrc/ftEhIFS71jy3uPlDqs7JILV6
148M4Cp3KTsVsAOHBStlik8LIOWkkwIcsKLMHZI72XXWLMUNza+4AUiZqcBo6gsw/qSM8GHlXRHx
epJjBF0L3hl84XoFKIztTdKgr6qKLoSORPGuhCLVTrU2ifa1iFtXi1Xg0WlacbHEmpf6XZ7ML3jK
R0OpoD2AgtTeMXXd9TyJFvBz0gT8iYqcNKrC7Vy4/P3p+xqD1RPDvKTAKFlXJ1kGQNn8ZV1EFAXL
KI5vieVBI71fc0Olr6w+vXuyX5HlyRL6Yvku0y6XQ3O3Bu/B930PJk92QReyl2smqG27rcPYCm2N
8M9DyrTcjONuZeiYh4D8Fz8wcFBK44ECoWxzkXbu2GE9S5zg5TjaEEK+7NrzizVq4TF0mPPCQ0tS
5lSzs0J4I86WSMwNnpmn2CgghASCeAEreBuT+zd7sGnYi3BgCeWr+n4ZOokOqyVxa7R8NBXDxVoa
4w2e0B9RM7t06eRpkm+4pqTdqrZ1D2PG/m0AB8VYODCOC2Mll6Ev6bsg7U4Ce0U88xP0GMVmH745
mv4jzpfLw+jbRpe4gEI+t4UrvKJ4xrc3Mpg5Asr7hbxvKVM108B46qrSjy+ApQt068w37JVXEPeN
Xzbvdt/59wp2Kyiogs913A3h9Cm6pN47zG4EH1TpuOYrM808ooHGc16phCLpTy+rXKdwmXcCbaoo
HuO63okijnjMMIub9k60oz3lymChB0eOEHCDxkvv46McyrjBmQ7gGmTs0NDZNeTQDliXcKId9G9V
DBr8XiZInwb2ZqNeQYcYMwbFnwLwYCXrJ7n5Wt7cN8B0Q1FfcjRNkONZWqL4jW0zI2QwJ5MPYQ9S
iyJfZYsPn4P2kun35xnNxS860D37W3VQZ5rt+7rqCzyV06QFZSNdiGwp5X08KZhKKDcK9EkqJFZU
vLXVkDTGOWa4nYz77sESiDnqP3fl8Ukf2UpAiz2CtTAa6H6QRPcYUIZTyRf/s2u5aiRSZXxOtJfs
2fqC4aRACybJpzl+2M1m0+NnPYenqVKvUl8kPC8iM36X2/OL+zO/Gs+QVq9Q8dSZMXmvjqyfYp8H
/w5TsrRQVxltUgfVt10ZU+dFhk/Fxn9thhutSeND7MxnFquom+YmJbILLJ5jevZ8kT59Xi3ni01p
oSCRJBjH373uRAHSq2mh0+rGmbH8p9bE8ew/luheI9m260DD5BUwCdWJaSYACsWOQlD0gnzpo2Rz
XVtPPxs225b2r/r6f7DM4WPCvaZvaDoMSFzUONq215DXK1F20jw2ij3JPAfrUqahLPZh6Sn0wY8H
AlJcwSpnJ6Er7sgk1G+9QOFGK47k+6yddDjssBoQY9whRjntygEQ2relDTs5cr6PKnk6cmUq2meT
VvTY0IagYzEjZT9lwUoYpSozfaHeXdsMAE1VBbxJmPy4M8bnUNZPFEN2T18eA/KRtqMGOF2t1BiV
pFWgHRvtPWS0+p5ElYQ79G0WMhK19gKSB6vUOjoTGKiALn2pc94smG9DkTleY07KNeRYPcmBmifc
Pcggj256yZcQ6X3MY2Z+M6hcfvcIwO4809XQZ6FcfLZ3ZWYdBWq/zNnDMLCqSxRFuXV/K1nC9pVW
oU8JpbLzjdQNWb9tftnq6M6iCA5qArl2e3WOo0Q/ZkfWB3b+5rlu9z+SlprC9JK8puIsKU8paIMs
U7KsTTOprmWjgxAoSuUj88m0dd/iiGMRFlH2OjvLaR0ZM5UvOSwLrAHtxmRG9hkizMoA1V3mlJgy
usML3US/Cu+pAwsuz0LQtaauT/vPRZv1UlP7ex9BZh1uEvisiRAu7x24N6TmGnbx5z2jyZCuzKc2
nx71V2J73iQcFjN0U4QTd5WVhCOuqQ5Qa/fgiA2d3LwR1twxvPNzzE9xGD8f9yrcr1lNeV8K8hkQ
O9aXjhD6pCUwkelooFRu289hoLM3nRCoNcnms/NLQpFx9qRY2KNddkLb2m5O18a+JkoN16lj7yFc
DdQIMGPYslN7xf8Be5H41ne1iT6pWm7/qik5yBOco80B69lccPBkNPGNO9S3Z+gG/JlS8gIvE0qD
3LRAbTZm+tqPZHrFAxOUp9TSed4nWT/9fWlXTJyu/Xcxihx2LoFR7qguLLx/dGAl4kB6MeAl5OXq
FFYYSfeFTW9IcpjmA6E0aA3N1lseKYvS+zJukyLZtM/Z+jeELPEpsqjFIuDsN4LB12uYBpGLKFLE
j5qhcMsVCr1ZZace8mr5mWGAd7Rd2bPf9VQR9AhqB0rXTd9J+27HE89qfQb04dWKz21ylcHSprJY
3qfkvXaMZ9VH+ayuzld5IpOGDB/UqrIz/L0/D6s8xYjiqjuC2HUpuT7RClxGF6MtrpP/ntj+5uxH
5hSdgD0PVo9uDb22rifn8kbgNEsisnIUyNEJFphPjsB0JqFvKALHA5WxK/E+YtTyApS3qafOU8S6
UVjpF3Y2u4V9cBK0fQkBfsGYNIuuHkMVJpI+4+c1MOFbi+sg1M/aEGJ3/rI31dq14HchOk3cokX5
RxO2pVWOWfBJm98f2zHNERk9yojwPy+JbIwRZ+EaXqnfjyc2ppS6Vs9MNIMWyzJrJygpXx7YS/LM
vrRim4OJRReN3/pLZ4rbTYs0eJpvBixHeLnPCvLiTH7j4NpFeDKpSrOq1x9i/eB8CIeTmDBJMkMj
HQP/mlcrAFU3g4D1KfC4E0W5kMiGBrfaagy2vaIsPTHyVELgO8XUwm21nwdLbvxHJpvu9DAvNpu+
FzFLLBle5EDeZg6JO6SLyMXO9fpDUzYSWPA3IKY+VS1LPsfJYv8LeLk5Wo7ACEdwdpfDfxDZU1k0
LW3PwM2djD19NbEQ2YgLVrs8w2ZsIz/sxBPu5FwmDcBko2FRSPLsl7iUsoA/cAxFqGvgObXTGPKT
TAZ1b4vYsmhdVrSLDZ8cpSm47BvhZ2npbAo/efem9CBK3fSfcsc3yLsWwcIemQP63QkUbkq81KjT
gelJPtUux0aXMWMrj9fabBKDFa2N1QPZhmbCRQZwN8tat+EWmGA+8iTchDPkVUpH3VvazZ1g8QAa
qdg71kV491CKCRAYXIB/nxgtcR7o+hMeIJ+NYFrm5ZQ7nKmNMbuaKSFQQBnnb/FpZ+IXGp0k0qjs
H3MsV969L8HLR9GbE8vHGOsOyU+97JQiRMZB+vs2MccK1MXdYlGOQlOSsuMFchy52zr2XavZvX0f
40oCysjzB1DP+ZTkaudh6+mQJygquVv8oE7AP2yJ/u9/7wMeb3kP/wKMaalgfvamvhNh3MoBRmeM
M2qMfyhzf189DiNi2QgB4rwEbkxLrGboAcs9hVunuRCCvZytuoI3U4RTHqoESsV/PTqxOrnxrpDn
FnViEQm8PwV331CsOm6s0oPUpIImjMoJQ2VnuRKwTAsedaU7pqVohEjjIQ+2UeT6YI17YZJn3cfc
tutGTMPgYmMIj0GatgD9uUVZgHV9fh2zPfWSPkmzuW+RmtJ7nVP9k6MlDpGgKTL5jhjShiDIITWj
lBRufcNIXfyqdFv2vj2g7eLXVk9gkkDa7W2aziaDLOI2WZ8Jx9Xd7rIek1L61cy+RepZj/somN0u
Ih9eSDSmYL2qGzdDIg7nF4fcWIaIXgoaSbRMh9O5pRz8NZPRniCx1Y0qaOCAYRZiim6rzaA9ktw8
kxczvsGzHkUUUj6fG0KmhprBqxr8cnFD92k3f2qa6Os/wZOhW6MOhQ2gyno6bjIx56lFHA/A6ZVJ
RI0+Sytjx424mVyTqh8MImf4TjKCJds+b8J8NUV+VJ+p5LL81LYAVAsLhhstRAX2N3yiVbP5WJwR
1hJbANr0QdA/zVWOEemzS2uH7Y4tlvRRgxP4UcmrFKgYVCA+f2HsRkpdRxg+Jy5AzEMdDclZ52Kh
OyeVuRO6SF8xOVD3foHIDnY/qoX8pI6EZpstXlF7v0Ca9hZ0qer/8zIZX8nXxmzc95zFZsAxlXad
O0jVFRPXRZTMm72f6kMYPmI+sN8gA2QnqmBZEJAvsAIjd+EXbhKRixL5vszNR/A1lRw3V8t14j7F
IWfIUubWwiizELLtaBZKUccLFWp9IDUZVtYVo9rMVbx+Nu9Fzng2/hiosxwcum++pPGfw9OoChBO
M3Un5df2WEnl7KjvnUjr3NniRdWPpW6FnsszTINYYBEv7Q0d3h5Ho48RnDc8J8kTvr/F2KS7bgc/
oOBuX5NLCa3IlKC9eJ7jSobJbGCs7+fGXpskGRk/45ya0VA8+iqPXUwIS7NVUuVybDgHYb9SdYtg
d4tkrl9VM5rdFi5opJLrOBpr4zx6XDLVwN7Rbh/t9Ar+tEWF5a2ZFGHXXY/3lBKi4wkG2VjeGOAs
p+N/4rfx8GhJlbzEM9nd669Kfb8bl0a/XowA5FiRfbj/7qT8JVn4R9f4W66OEasLXv7HU/VLFikY
Cp0mi43tByAh7v1WWA956ca9kdSJxyCpxLWo/fu4UaJeyq1wvLD6tye7ukW7AuccBDFyYbMSAi4I
s25t9sxQBFAcFRMSRW1GZyIEdqBcMqJXXBS8p4CQB8oGNvGL9v3HGTqWUiKwRrpg8iZL35bhvLcv
FhM0jJ7bMBEte0cHxS5Oo44K3dbIG4o3VijLi3BCijzNQnsbCbln4zRGavNeOp642gTy2/G0Yoj7
VDebhe/fjz6E0TFiDP9Er5JW+kV17m5KVA/tp/m/B7Sd1x6F1RA/Uq9y3ssL4pDzJJ8lqegJkyTw
2cWo5m+kYHn+ZAYRqasno2+dGzbGxa6h61UdB3wzVkl+iWUldW4QcOdUBADbfOv9LijCOHLY4xvC
U40xDNoZTdzHcByEMCBCiA5NrkAeHDzbd99eUcT/aMMtpLNoF3nPLrZGuTNJuQeKP9lkwe4hUlhK
beW/ENIJkty2nF5i2kDvY8e3/ZdgHVcBxXDhsMaovGWHu+PbykdaMUQ2oLi0w76N3nXWXkV7u2KL
aRLivPiTnmRqaBF7PJqWFpJQJ7OF6OISZRgLWN/qkMtnnUni11y/2hjdGeg0bzjQMNEcyOiV6ozb
HAvJIP0w+FfUX2xYCJcQGi7jhIY3I2c+O4LDm/QFks+0nC+o4EJuE2Xr2IEzO7j4wKPtbLuwnqys
rCsLUDT/n6WpmdU8godqfYSY0ILHCUxayhk1byqFu1Z2kcJUDa89lKlBYpM7KtmzTu40zXuEgnk/
xCCkaqeHCjj+eI4yYW1kO43QMfGTgYZAf4qBrfIeGzPkK3GReNyhpLrJh77DNWdyvlYiMICBp5Wc
AmHzcHEG0tJ39QfOvGDy/vOg8D1Nan2bsXFWAog09UoyEW5cxqF1CglN5BQ/YHDvTMUT293MdTiV
cz8TzUzauLWlhlAXvS0snOboe1dHGydbdLwPuyrhh/JiI6J4OfFiIARguKSMbld3sxXMuOS7BG0f
URWS9rmj/cFYlEE13FbdGyG0b+cLjveoEpY2GgFX2zMkNygCsjCaF6YCl3eTvuyVZprJBHKLVAS3
MCpCrmmrOo1wzNes5nuZIf7yC+U3luc4I8p5fvo9gWFDHUAF2RNzmZR2VFCOiyL6PcsGDH2tckJD
lOd35fxJdFEynISApEeCXcZyG6v3KeC7yJG0+LpHUESw6VHqZkc5i3gjoGhOcKgHNKJJPpm4TuHx
0eh883wCI6v7zWG2gS2WtLQQaPE03AGqhFpNdRZrccfdYhaQMxim6nUhyyYiXOVVwpHJ4pD/4sln
1XvvIsTuWQMHUQJxK7iJ6ivnmyzyVcx4hs11XLeUiwbwH46HyFCPtYTwA+5rm6+DB6Hnbt3m2dPL
w2YfLaML+16nXQW41YUwrB5uRTmfs59Tfks4f/t+TIrkBYNocn9eNwy1CeOWq4w8J6qoi7AJQGe1
CL9EDPRbFNZWBO318PREcSQZH+mOFMOe20BwT/T0nUvCvu+EFy6ho+++gG3W08DADAlet3G1C9vS
sFIEv9dXlEva6bqaU1P3ToX4zsmmlwJAlcdT/XObUarB8FnMQc7g76/xTy9QNe1MqtQW70+POJGc
v8JukiMFNE0WKFdrMp884JzcYODxjNj1MgG4MK5PGofidnPjQCwRyYZv70mWgr8O2vXTKiSHZ1FX
67pc+kI9cOoc9VZ2mNo7FrhaJUIrMLe/jgwVwUbrABTNoS4kzpfccTsXZ8TgRzALvPSso/DeGcrN
oshx2q7iYu0qkNJQpQskJx1OHz2WDXMgg+1083cmIu09q+25zQQ+B2cJozNeiAVviPv9mQynRDAR
Yd8clzLrVODtbCQpWYZVhjBBuBqN7HEbBKxIXGsC4APaIuXx5FXy/qxDeqyVRkXp12iFRw6crGhG
YKc3k9A9PoInTvX90h6sC8W2jLgIVQVfLAxPgVyYoDwyjthcBJHKwo4LuPXUlkpMOGTglY8dGzFY
AHtVuJYVd/6HvWlEcXxckVVcfgyy4/9azYgC6Reavd3af2apXnjAVpG9FQ3igMnLSCs35/Zz/N6t
oei2QYpJw/blgB3g2ARBpN/ZGffC3osWjYRnA9tgo11MG4m7tgMSz48i+zNFYj0guJTRj1/+Z7pV
pCgooUQeKFyeq1mGQEMQtb4PsMBSFAThrGE8r8xRfPyHD3ny7JBM23du/56fguJ654Gmmk+hmuGq
fn+msddPpfe6132LFGeYWSGFvYbo47Q36cRngpxJnNWtnr+ShTC1YTKewj68ncmgdnpzjvIlK9JU
RlTqPxyySZjjmPTuWJFmg76lNRjLl8WHA6UpdLAd/l/OGBa+QS2DGi76DxdvWODS2Y1WFVv0S/RC
vmYoTL/sDlUjhCfPU3x7Cq3Nw2ZrcCvGa2UVHnZCkCrKSHXZLBtdSMRivTNlSeC7MNwq1htYpmP0
rh0TlicSpGuEEE+pkhDMBxGHQgr8z3xb93qe6NP0EPWJzhbjudjkoGevfP/dQO7bKSMv41+aDiLv
/daTH8tmiNFI5FdTC7OjS4W0Vh9/jOX+8E+m/ebjNYVy3qm1xRAh6D4Alk7e51O0ouEMaB/e01HO
nmO/XZBmhVSbJdZUzs0v9kJY8cO3AcPU+xAMgQMnlH1CNRtAnnUyUNtzzngFD6OGwbfnM7F9xYQP
p4m6philobVR7GMr3EXFUSjdlP9xDI42bThZQQ5L8bZaHd3phgPZrFLTacxzco5JDxGqefVKDW3d
lw6rb1lhm85yz7X8sG3ezQHeB5P7nAKakAnDrG1F+8FecaG50qsqUJomShQy/RMxd1jpBrKWzSOg
q43kYBXubdJPiW2AjhuerUXmPyvzM9RRq9ygs+2GN8ApEDzmjE5565ca4l8sVdTUKpYe7mb+ixbH
q7EnGyt/HRHC57oYTSjs7j0LNZlDmkaBQgo3SoyYYhWLFglCQu01xr3oSeKZyqu0Ahl3xHxO6UBV
OkzfQYqLu9CSEsGae/YGcey2rlS4W3/cJ75rFswHHbTG9oT5fUvrSn+F0QB3LBnShW+ercQfNY8i
33eDnd+d/Q+CdjjYIn1vVkTXgpRAq29JX/xziYqawFC4QO5FmnA8MaOvi94xX3E+yvLCYVHLPqlx
Ma/+eUqNAuWKGGwd+TeccB8eztG36Rll9Afq3ZVA+CSg0dMb9e3kbBxmVd2vBPdxyYg6f3Y0BLGx
LwzyxcYAVW0ieYfmS2bF3B2bNAulnPBk/p0hIpRemSOO2VcFQTDyvBnXrqI8iRk9zAFIWISrvpo5
/Z8/baxWbkKi0gtksTt6v50uihCgXmnFyc0ClmC/4K8qBJ8dhrr14BGGfpxTLu6tNZwyJRzybd7q
3GrRgb94g9kvge45zbC2a4AL+OoyC5WzZzrQwa7YBbirCgc9MK190aSG/3rMotSWyKGVU3lksTrD
ZwekGGTPu4QaHPtKh5eB8q/aSL0nawpGk9U6PmV6szg1IdPv0hpla7sc9EkyCrb84w/P0MqSk+mN
XYxv85xxHexQeFUInI3IZp3ggzbmpAl3q58zD6oKpZHpCciHEPoHSF/KRaX2lVPmnLGqmlb7xqkO
jYE9Lu7jGnTca+b4m4P6XvEccSTf+PyrPRzlK4BmSV/pb9ZfURB+RlkLiLBySqxqJbBlhJK0V8tl
HEt/OiZbxRANtSr6nbQN5FgCUExeEpf6iFFoG3oSAlRMSW2C7CW+lwtyLGno0rI+a8Et0Em5Tp6t
uoCXaVeh8VDKEtEgzf45F0ODCjR77mnh1y49v+tlqQggj0J73wwg2Pc9nAmUSM/Y2vRgzdsHK5xp
5oGAEzVy/ezL+LJ/UDYqvuhFMkFCcLc+2F55EoPOIP61x60m+c/JSbBowwi2XL/2raKxM7N12Xom
Fk2kDiK3RWIxV3BLkVP/WG9XF8kCpAle0YJ1wtI//nXFh+GjbjddsXrxaEcwwSEKbOTtuR4nsfOT
jPSJ19phC0LuqtdicOGubYHt4TXx1P/jCrei39myjKG6zpCJMGXu1cUklvcBsS5byEbIC3O+PYi3
JRxYvUoOHcPY76PKVClM79n9G1nO0nbYvEEXvcK8VaQVpfWCu1aiY8T6YvLHoOXG03nOe2H1+TU9
ZsDyg6EdDDpQMXLKkkSU19iMjvvNvIKWaWiBKYEWcZBK9JBf+/RmtYtTD+FAzD+T6vgv2C5AURUL
XSFZAfIDLUkYTOUVC3nov6zZxGVym0tdOoyN8iB6KsNHCR4juh1WfCITg4w6lMRHvxyVXmvy9+II
uJcDnlt/4ysPJumscgBV7G5Mv+Ll1uK1qsRJABL/ca0wvwzWCmmf1n+mh46v4OWT7PlUa5DOgfzJ
k2MAqYAT5opSSrNOVpmvieXoaCTzUgJ7bb9LOQfeweZWutSrfu8FYQ0nUZdzRUwcvJXn797uCIb/
qTztizbUMj0rNAX2mV+p0ltshnGOh795cR9ZP7fSWmhv2PPEPtBv/puA9wWehq8FYWNg7LimJd37
++rLoYSXBKw/CgHcpI+JitwdxGhCBnRbCN/wKTjl7CTeCk4qL0ajK28qpErgMnzNQgxEJt2CQjHU
Lbhd71r+79/KWxqmm41zHU5ZPsvb6OQEVkeiJbJR78Bnqz2mxf8cHdKyMjBuaJoY1FaoXbP01vDx
AIt+v+WkvlBQBUYYHo3q0g2dTCqDm1IjHyv816y4jq5sdbloHZuvBuMfiarZ8p9r7GBO0Ax2v+a7
UG81i6OB9s8eDAN0/5Br6rKYLoaoP6fBNdbU2e2Hl2FJgbmMm0j8XRHLVgQ+7Z5sz6hInpUVChFg
CrsF3RrO8mbz9+aR1KbREANWrAHUS0eEvFNWsUuZVRcpuvCneewb+WqoftOPv0fLxfmWzkChJouI
Y97MuSptC2xMu8r5zHnvxs73Y2xPgo7udUnykxKLypJhJ01458c8D+VLagCW2YBXCHZIE8yh4GWv
rNHyVaHFb+ooF0nNlFGDzMz2LQeIptKds5mTv6A8X15NHKDTBOB7XB5iaKJfgNLxbM3zX1ESF4za
n0IB2x5Wj+hAv83dJmA6dPzP7kBJID4Up8qG9icbzcUJIgylUzxxHB/vmTOVZWFz7adDjrvqJ3Sb
pTzsBscjwoNiT4fgQajSC5wgRlXaUjL1Qrpp5tvNtvE7V3xGg10O12r0iHSwPFl2pevPnFj4QVK3
fmOP9WUE22aRNIaMcMhTAUwyNL+KkygzGPCnlV/BCX3mlYi0s9YQl14ZZ41O8zBrIkfHSAmCaPKB
i4ZTM0MTpH43FiPT9LkUvV5vKl17nwsii1a3dVZZBdIDVTcxcjMFYRKoklctyZQ7vU1jKKMWUuyw
Jx7kV/ArVYbrUGj2Rl6KHYkk1Z+aQMML8QEMLKGqo7jZu+XFs93QmEL6OKS5kqD4lv73P7CduVyg
YfxpJJoNl1EFOz01qcr0I85vDfkM2GMi9mAdDLOAsEeaSRPGNI6gi5AD7WeswGnMDb0MPs+EBLZq
hi0FYz3m4aydoUToZTPxfZbfb6dXsSMPev71ex8Fw0LZybhPMXnDeVJw/NYLYJ8zW4zRmaxEI+/p
FlQMLH/P+F1zYmBq1bUgAl9L+cvl4aHBdspOCnjPyijtMyLETjRhaL9SMZz9jQ8wXgl8qtycDfEy
S47ATjss1vKM2hj4DuRIq3uGnGlq/AGonDV2pq3XN1BCkoTRuOlDZoG+h6/MimejFGL2cxNE433s
2Yk3CnCdtX5RE9OwHlguUBRaF5GFXstnNsqESXvONZPoJwYsOnW4gK7mQ3S7rYncdJ2IPKQThDeD
LEFCk3mSYlqCGEm2gKRpNhY7Hmq+7LkaRUD6VwSxCvInZZmrZSoZtk8o3f0oTtJxb2m2H+mmqgib
5uJLAfx8SK1V4NcaWqYYw6UWuNnMDjHdsRpmro0R+5oUm16LYKmnSqnC+hYAD0HJ+5qe6r4b8lsY
XSDd8vbpd3FsUkvN49RKE4+IKCaSQmZatwh8VERr3Cjvs1FD1VE1Y1Op7kC4KxN4qCWBG1xMXI9z
pTBeqw781N5UF4MmUaKmE1Ml/pxwQ57HB1ojmNqsmzpoUzUmwNhk901aKjP64U7PAG4DXqxS16hr
f4Fp2kwndMUSwqNPlqYygePuO7otFSHGyg94a5ZNh3B9mklYC3trZeaI0DEB5Ko5j4syAw4k7rev
cc8pacnTRLFd4Lhuma6Z0Tp/6ZGLn33gK1fREmDpAYnuuyDjcFlLoBRXRUg6A+hhSwKQRqTGv2YP
E0AYnmWav2AXhQzdyzfUvoEHlgVDJ2tkirqCujmnj/u+/IPrqBn4lV55E2Jq53PHscHszLi6glXv
8+qld2YGd3qUXaD8/rRJCKoxoBgV70hc6f2mha53sem7mDRhgOHuxh9C87me//bxWb4FDl0j4eiO
sKGWKsIX6SYq75HaRo3kZNiB2zhp6MHPaRAas88nntMORoHlaWnnd/3ZLVkZLwEHxg8fQG1/4VPx
rKxUejvLw4zRrOJ9EqpGdOjXYmariAJhZtVZN5IZX9pJ3zu7277j0u0et5X8Hnjt4GBIkSOEHzce
3sI7La0qNYrZ71X5JpFvs9DSMDLMsWFi0yEcdQi4S7yM5TKI+TYgX4kX4DcEnUrBhsyC5fcuDP8M
mj4nTdWCug8KzA72q+tL5F0mXCIjWZQoZFgkvbTZjhUd+LR9M9/WigIUDRpZ/VNsxw3NRlI7sW3Q
PHImBY/fHalEHM04o4XEU1EOnn0G+gFEjet8tnNaw2WWj9r0vjX4l3czCHeq9/qrwLWOgZcG1zsZ
3vA8FiDtbwohmTkvcxH0Y58D1eYW3Xg1Es/S8Z5BOmKMd23H/NNSS8J0nRRdHKMgg1Si6yPNUw6t
/+bxCG7NpK5wpw11jyddNoIxo0nzbtt2yNMgUHhhZdGcBdnY8bw0qbjI3HvC7+e6LTYdjjdnZ4Oh
ANW/AbwomlXNLfTwA3ZOp9K01iUmpcFRKjHb1vGuG59C2o4arJqfS9R+oytuqeUrvvlPeu9/9PAj
uA5fj25xxFcvG10GuTZXWVpTrXmIWCqqm4ltHMObg7t1Rqcx2amyfRJgUf3t16VtFo5xsO7VO6yI
YFlEjBR8hh/1LOoqVfp9iD5guuXKWb1oSsMAb14rXCNXRZg0/v3Q0TeCYhCxWHtKcAS74AIoRxZm
gbNV8a2U+f8C8+QBunRZa8D1+4u7ZBPdqzEXQesZsSmkt20l3i4wXiXmZHIlIih9cPWaVTctAidW
ps0IQvEAq+gpmipA1Q5/RkgwKw5nEUDTlLKbcTPukXr2yzpcFdUAQvyhGPbZRpsaalpSJyAwinVV
8Jsggdk1iGar5IMadDh45MA3UNTNKHqyqwZPvEDWi++4FlplE2srXyOEzrDQH3jgHzVmDtF1QcBo
OvBTSm9YHbS/a6Gy3aBBXfiiJZ8FAdh/X37WW0zDALWyzy0dz5rN56dwnnhiBpeOqBi7rH4O9jGW
KQQYGHYB7sJlT+kEbLKK3sYL41016DN7lJ3fTB7+ZMhgQQdkndpxXSHI5C+XptTsQmWAOpY60iQl
OWIE9L8CoRZk8ulRtG10MnOmAddkzw8rR6jU7JRC2RP/o0triAdj3w0fKgfEzrKj+iPg/+UnjqML
UKddpIdXcgGhNQXyE0hPDgrVLYNPInh4naA/betR4le5IaXt2Mjt42Um/RefVd3PfFOIEBkyuIXw
jWnf7gkoMuKBDv9HflSd7xIE8jpCGsRTpsYBGAOJj823tvPLYz9lBmoXMGHVYCX98lNVsi6soNXs
UZIBej+GTmjpFtv7OLkeq0qyZjWLjli6A8fi4PwgbmE3/T2gElqhgOn51LMrEaZ2s3IshFK+T0KP
Sl9f6HEeodstniRtHxmQH+ukjR5Aotq7mfzPdWxs/bvEV/QoYe7KR/g2M+O6WyRE6S7/8NeWcWWy
a78kQpEgGiCQTTmqFeSff6ukpJlBFN2W9C/1D6ktAjdxyQtjOlmv1S6Zu25kB5Z6UJkD6UJReLVp
RZ1IYwJwwn34RJ1CYkh4vldlvX3eVvXapbbAO0K0KYW9KIfqEfJj/MlRdzXSNAtvI9XipUizF3I3
09+BGo4lZSX+sez0+fiyCONN0lHlDLywfVqqOaNUj8/hoNyr7cxRvAsL9WHa0YkD5/PQfgyBaPoy
deh8iQNN6L8tbBlPvX1FIspnCT47I1lzVTKqgkW30kfJEd8G4RQLIIr/WCBZYAdOIQOCx+Xz/EMI
Z9NZ2bQ7CJ/YQ9GctK3ENNfs9ugDr2y5NvhrPV6BGlKc7BvYm2xmJdqOhyqgH+hDSA3LzQnSwmQI
MOdaS4wctVt0w+zvrcljkJMiCDnMXqk3G+3gKQGspsKuBinM6d6LB2WLMb4f2loIR8mAG9EGo6zF
mmtOg3hYEyD4R1bXdxiLSwFHS5z5dE/EV4fpWuA/DZr2S13nuCgELzB9B/ArRgFJngL5ynJt4ZWg
82cRR61Uw3GRghrGJ9MdLsk2s8hzv7E+D7jQ1b0M1NDRVbjpw1B0xOgQBpE1v99JZRR3t0qrC6h2
gfTJQaJ3Egwxc2gf1e0v3ktvrSzgBkZ6PeT8Zq5W+8nNL/2e+3O0Rp9Gh0yigbNrsFcMB424ZA8F
9SH/soiWZOSZsxGcV2tuTsOlCDm7N4KMx8i5GyLsJ8jd/a9/TifzD+WVfHbKcb8z920+lZFBXGxS
Ok8v17LVq5J7p6WNX4hlR+7RwCo//bu1Zd1IQnNcXnKMtmyeESIfp+hNsaEGAebxF9JDG40FeK7n
GwD92zEbB4GEdH4vl8DLrhbL16YzeE0RCW+lQaHZrACh99M9PApkHBq/wu5DwR09DnXnQRvGro4m
WNAy/XUOknTu73tWqxtarHOeUM+NM+/U3X5tSSOVNUx+V5BUaJOb7Aq2HcoBflaZEvhCg3Ixr86e
fn+FKQqw+IOdEZLEohsCb/a5aq2ZTyZaXqeBC1tD22piZ35dmNG79M7aWbbzr33cZbMWnR3zOcfF
L325DvbmUZJSE0pncH/Vax1tXf/vGjQLzj2SECijSu6BiGEfX8mpgbt9vUMN1LnEVdBiIcuD5Y5X
VqwL4+3J7/z1tfWKuMFSmI4XsVIUb0Y0+KH6PBGdTMqlihPhYkIgOPlInfRSjgP6W2Z+Z+Rg9yP6
+N1+Y7vnKXl5V/wuUgASxgXkYdGU4Xq96+OjsXJMCgC+ESP+lPnUxG4ivjoqw9uUhvlav6A5Y+RV
rsSjYqm305Cku5K5vmOMyAhwXaAeX3fYcVydvCMAbSfNBabm3pBNlY65OFiUPsvMGnRPIwU7zXi5
rHktCsPO9M0M1sebd6t4+TOET0iA57nzLoNMsD/C/5Z29FMJH2CrAem3vVSudW9ySHHh/xbXqTDy
GiGMiliaD/5ZvdVq+15fp6yt96aq1TIR555+kNPN4LyELLV1Z/V0kvGKuGpTLamD5u29mCAqBgJV
rN7TOi6OZBJx6IPC/H6CYwnF5u01Re3/7yqjHaWkS3ZPPfvnAAxnJWPzbuJL4rrS1SBTT6mE5XlB
veWoX8fvRQkei0H6kFky82o0mgvdSMXYH3S8088xk70cFGTg9zAxY2vVWae4VdYP1w8iY282TQeo
NOoE8j5SzqzOgDEzw5jqo77B8fCxcAON3auORwYkCLFPY3GXzvueMchqiVOvXa27AczaOduZUuMT
KrPYIOfpBkx2L6oYZUDQS8mX5w6aYEgIUH6peo4xD21p3ZRF9ja/S3n09x5EtgR+mygzuu+2MdUC
jL/0m1YtmC94UODISBum1hkxkg+Xz2YdjPgvnStMoWl95sIXrqf4mWgcJg3CvL5lrzElmKS7akT9
6R40U1pUTSkkE0J3zmhvo7ef5QyYP0/TOrddCY7JCEqCJC2VNb9ZnEigVJjW4BREULtQS0jvi4F/
+c3LTdOIABqNj2q9OtMITYWhrDys7l3aPIuj+fnhTs+aLYNkIfhNcUK8t/H8MP1vkejOLzP78l9P
Xgns8zXwiSYUIA6bCg53bGTUholtFQuzlB1QKnqivijMvNsSDSzmtuWRbrV5yqa2BGAHaPizh0AR
DTZ/NdN5qDhLNKqTaRQ5HZn53zq0UeAi9byo/T6WfVJMzJ+arb/RQyf5c2s/b2SDAYnkmbAbpyZm
NngcU6G3bQSB0oV/5vjJfO6VT6QmkknsvJoQKIrrVY57htPB1KlLNDTz9S1h3Tt/0Gun6uG+48yg
JasMygXekIdnSMTAF/z1/+AyFu/2oNG/qhGy6kH9w6fIJsBr5DkJciuxRgI7MzmVzrQN8IDy6eqa
54XCh7iN3x+j7Bt/ycp0CBbHcOtDbYHKHXql+AXsTqh3E0Go8TL7sMkPIMepD6rKeuFu/VAe9cgZ
I1panbC7GZlIOXS9acxJbTo9yWlNqdhuz+mwHPkYMfAmw8NGNeJzVgPCUqPf9XEIyezndGxp2nxH
lpUjROSOH+h6FEtCfsaEEF/LWSGLz490rEnappMGr5IvqalJOl/A0pnKBqnKkzeAjftk6uszRlkp
ZX0EH1O/R1cRz5hBDFq6T34O7OAJ6SsuwIQYiFBfCMM8fbcIkPJCyXLfNUADJpf+DBK0arpL5UKp
w6lVVpNc2DRMTAcvVhpV7O72ZH+b+N/khtbHPYcmesuDq63dbrHAQFkIoMxMcty8SQi80tnAZ1Pe
HOzRIzkfvZHrML6RPGx4fIITPJqUjtBUcWr6Zs66ufiN8BphL9Cvr/Jog8KW0eSz11PAnP+F20Oi
OCGkPFVH4KRY5gSIboGplSBOOC/UBLUhD9cgqu5OzgeTLwqwdS3vJbffZZ4Bf1l8X1uqzsq0fWPE
2hICCRzXPzaGn9ohDtDABd5Jru/8x1NxHZRO9QNKkkLqzoW+JQ/muXI/vGE13Y+rRMOxNNA1rOxC
tudYteMfmyOKe3aqUaOVpBr6GEYlrDwnxxBNNgOdvBv8ighoW5h9mUS/DC7lSlpuLn7VebBuZ7W/
4zrfEWDMGPL/Ki6hnXFdu9iFjswJYzvURy8T8liDIlyec5iMKf4LZ/y7UDr8qJONLxkOIg+a9m/h
bC2fzjSb1wKOmCWGBtOIO3CP81o61uR0iZ3lv9GZqnn08Fp6xZw2aRpkjUkw483WNfcumjQBTqUO
4Q6woY38HwpfRIj8EecXxlGOsP0YjyGFSXpgigfq7YVWKhIu3N4NQ83FzL9pqVr1YZnVGDloLtFs
YV9k5pr0nQwuUJWoKJ2Avr1cWWO3inX+ireJSqQfsP0ls5yHdUOEYcQrMRfFIPNFnVsG8ZAt3f4w
Y1orCYV8j31Zq5KeqGFcZtcwjHjPQz/HvrAerKrtKd8iADRxoc5A8lNjAscMlc7SVapho9DIni/S
opNHZnRNYdraXt3uza7cspisT7eTpcr7UZvkN0em33NGWtGVynDpa1xqfHQLenr8H/l1PpmTJL7A
SlwqOp59BMpIwJV+kxlEsYGXjNU1QEykk3dwV0j79pJ+agYUlQa0bL7dxEUeBARGO+gTL6owvsRF
yAGY8gbPyWTS0n78EwS6IpjvRgb5E21Bi692GVE+HwKlEU9eFejTuw==
`protect end_protected
