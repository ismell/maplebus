`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ndF4Sgjn/aBs/bMvOIOY2UTDvGjiasz2t31uIAkqiqfO+iGbki6xxzfe3Z8KQxcf/tAXlLydXEEm
GQ4LdpvG+g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TJ+8FmtdrnqqsUVH8/Gib1x0AxdeGJ11gYSRoXsgZhlf81WgEitSWstSGkghryxxzvW8VOalTVx9
fEUfffCnwm6+hcLM9rFJutwSIy8jKJmN9CnDBtpJapYwzEGqkQAalfJO9ZE/aNJLoeW2gs0aq8u6
Y3KvfKpbK+8O9MapATQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UjMfQCHBwoc/r1HqR6nGojh2Gko/ZKWwaAWv9g+eIhlDsgOuTJUQZc7UFXCeSqZaIPrmotN5HGB2
12Fath4GWa+RzB56xyjUBS9wZfc64uhn+Z9lOZYHEz2pMKuo+FavKt2SzSFnJwzy7hu8BDg+0km6
ZWWSocEkQNkUPhwQLGgj7WtffCXOCK4ClV/dO8YVh0I9th7hDsdkLsckCfQahcgzlRO6pMp5zJNn
0LB9323hFRi6xYmxOsCHi92TW0qvo4/7y1B/Db3DlIpOlTa2o66IGUhMoZU5z6CwDjo44QFagDdk
sSmGFt/Iqnv6P2vUkpdCm3jFfdUoG9Mh9JFY/g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TJMHDoDHEF0AWHNCVAW3R7dBYh5NcBEQ10y89tzHGMohL+72pZLr0EaNDsjREvb+m49cN8IS9wBj
4EolS78D5cUwgPOVO09RIDVkS7eUCjW+gq9WbOGm3MlHDJAwNZBKXUqPqW52Uc7WsHSp6Umow9VI
As+/OLGXZxEqoRHYCmY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gv/XnBdJ1POda3u/pUUZ7PGn5FdnU9sZZ9mHMdPPxeeJexzMUP1dOGeK/DaLuqHyMbWbLtzhpfhD
TWfGS+H2s5hN5ORG4A2Tue4gVMEQmhb/m/8RjKPJLmcNlSQD33g0O3KLLh6t4QjzG1f5O2jpjSOa
9CQps8dFM9GqxSw0nSyFz12+CxQ3zulCt5nJ1hXZ7nhREEH70bZkVPBizPrWs30FoMBpX/d9ahZo
8iAkpA/HV6W+9UT95I4x/eHNQqFp059dg3HT4qhqZCwLNKxm56YbqfBQc1Mdx4oaw/GmleMoTq7Q
iWr4QP8mJbFb7SCm6bulLlIRGrFnoRcwQWrybA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31280)
`protect data_block
mwGioMqrESAIwZzKAFli5j8momvRwBEwpq83w8JSM8Vgch0yJnoSi9uvFJUKoSMAkF3OAgEdTQJk
fC/V5ydQnAvMX2rt9+DaYXuk3GWiw5quKtMyUyyDjS4PzuxLxafwJV+DmAQuUuesJYHjGM6snHkC
kZV7cOVKuta2dGY2klxq0yK+GdzYydrVTY1L2Mf4v0EmR3uDSU17+xoknt/dBbwq5l+VLUkQEgMX
OiCtSRKrm/n6Rs2M0/QED/ksQTbTwcqzX3bwdA1jGOI/DPoImIW3LfG+vsAUXhEzF/gkNrMU2LVc
HuiXlSO+MW8jb09eii1MYGXDI3xz6xfvQ4ZjCTKYrLXjZp25JlOT+rnlTQq42r7xfY/zsoLdzYjI
onekFgldOyWavEjvS8lwQ9p1wNzAtSG4L9jU7HELmHfZCEQETTUssEl12KGuG2aTTIbD8fK+C6tH
0GCjqVD3qEbEIk/rrtGpEw9Uir7oP6BmMD92rTUOsPt9LcvGBqw/dereFtdSJIuvImHfzhljv+RA
6XU8fLSdbFOKoBowWa5pNwMlyXIqthqjCfxH/GBmZck6EERwtJThIIIch75vyobpcCtRIWlDXBV6
8Mt2Iiprf9R09w9XdZNtgcv7CGdBlOZFHkbgW80M+8Cg8w0mUU2JGjOKjz8r1oe1dYQ4k4RsBbxT
KxcllBF/IJ010vEH+GESEJv8q/gAvJSBY1XC2/tIgND7UDS+Awr7/GvByQQBdDe2Tmg2lsTLZbLO
3PgxMqchp7gnIJcn05+cSOalU4VJr102wDBxsa7tOE3pv0MkX9B+LnY5Wk2+yd4Qzw1ihtku4puR
FkGS8AXBbnWJ8Nfymq+Tz8aaSdDR2LLiof23GPJdgQP5duN9clbeKSAd+4oVo4DhS9fWVXjtggFw
5Cfwc2tldB3gVC+AVUOr8DonDPivPAW1DAqQYhI+KIu5mJeiwkwmTgymn77srq20Cz+EnbTAbQK9
sJrBd2Pr/2+SDbU+aQA0OkHPdHj5CJeCBkeaRD5FBbjPYJsep+K9Fpncoqt/ct60NZ4uWmDzvl3p
kp/X8/F0adAzqWoq8o7hfftuF5YWAe007J+i/eUdS6jM4IRxSnF9FyI6kqKyP6bZVby9sKH2Bb82
B4exHiWK9GuVjVV1XM/1eiFCwH2NahIZ9/5YeRKuqR1E2Bxvd6R47tRh/k9/6sCysKxWTWVeQ9RF
BpScP68oWfRmv71fnwR2QRzK+YiipcYfNL9Ab/9s932P6e+RoPTNOor9BlFO0jHEBuGDeRxCctyF
aeAHF7D3JURjMCGKDjFRwZnADF5kY4A068lzE8sRd3yIz+9be2Rl14nugUZzf6YbtwAngvJSz1vv
lcIuO9y1EIoG7o/7fVglBLMUrMRmiUK36RYS6Qn7rvZhkdaswVYdhtlxic/fOyHIlDJEsFDRoVAu
OWDZpfQ19XvXjAcuqsRteTg5xHI2CwgvqgKQsCdIdzHCTBZPA4QIcY1IaFci/gHO8nePin6JSmtJ
G7dEwToCAHQWhKkNTbsnhqxtyNg+etNz7PbR8sAuK4+sBaC+Rs/4eRZS+rxc/AmXz9GfjaSYpkWp
zCX561vPY6uB7YSfnFDMIZ6IeIqJ2S4uE5zHxq5h4I6ToN5knqQR/WLwNyBnvVzdUCQFPBSZMHxu
gEPvZvO68qBF6F1VsNowxhxrBMhpFRES7jROIjS0hBKy29VTthdRhBurlmyasP3FS8GZeT+ZuzVT
Dbbsmwe9U764fVyxPDV+SG0MA0mW2re/Kig/CE1sm3tIJRJyPf5YSg12wYuvKspD21q3d5qx5dja
hWNq4iaUkn4zEXFXNYLux8csG2hFQi5XANctDZhAbtPovrmmvLzQd9iir93OVGklgPwTfhPzi1ig
kN53k6oYyZeX0NahnZacZc6EDItImQLz0124I+WN9vrMBeTACIrT3TmmrSiZsBt0ygmyfeLvrcUi
CY0jB/67rbmS8EztpsXDr97J/tGlieC8cWvmoyeZL72ZnQOOwsiJhf2hccJULLBSlwWYtD0CzRUl
MI8h4NgzLB1sWpQOs+bU32LhGjy1zg0krkLfmVYi6Kp1mrucrobcnV3oz4c0HJkYCcLdfndPxJ1i
BHK1jaGadHbjen/WQskpuIbLbN5V4InKzTBgSZvWxmFtUH70hnEc7Spv7nrGVsj2qfnfuhTpQnf0
wk+YpAP6WX29s9sUhtAVeyuVD34gCYCLGLWAKqI6vCADhpyWFPBBaEMqGNynHmDWBsuJZ9yphopL
H9p+3HbgeOnCsse+i62jQhjhJ8s7nsWmv7pSaCjtU/HRHT5s8Qz7etF40smzvyUxrvmdsc0J64HQ
yleW3uk1UesXSElU/bZ7dT9OF+ItrxqHAoxZ1UUY+Huw4MBfpAxBnqYBdq/H4UYPW94l5ycPx1sK
m+dhlsjyDQbkNT9G8tUz4KCEf5DWEcNLblvYm5U3V/oUOpS7JDnxga+dJYIKo23GOPJQDuVfKFRM
DlpEODkSpr0LN8M0c2vlA8Ii87t5HXSV+ToiVAnrpdQOEsHlsGekLcW3aQono7BD5oVdsrNT137a
8ruxEij483HA5DJ6CAmG2/5TsdySfIWR5yuUD2h2VJg46jX9AoIG2hUCoSRUv+wS7bxm1LCt7W1K
7RxgDlPj+mv4BSsW1uQFW3cclccvYrtBQT0cqOb8o7zCXs8xFwhbWngAoHUZRQg7AyLnhnn54SK3
rgu6F+zia6G6w6Mdmegz4ROmMVvyhaqSBgfdFJtHDA6gwhAPIzozX39A+aFMXXrEyJV4lHczRIZT
tBGOhZ6Q/LDV6lh9Td9h7wB5XimIBz4jNBBvCMk4pgA1TfWeqchHVzqk1Py0c5eSc+cS9BUpOfqp
5G22BCWHRk0A0UZaCCMVGF7pMHYotlkQ3RrQNdow9YQKR3TMQvC2x7Sry4KYS0Aq8pBMKYk761BK
YrhT7rTHXK5uJ0e0hq8R73sNUXWZ1YqrqNnDFPLEsaJ+yWQ2EMVBOsbDNOUcmwjCo8gszmjFmXzr
b4ew13lKY+IHPj1BVeqz7Hk/45qAfbkRVtKHHYprC5bvUMI7ejJoxoeo2sXoKQ5xp5vXyCNYa4cA
JXFsBG1wYIw9ydd1gbOMhmHGRMPeYnCWEeEPOi6Ciyhck3GpFavqBAKhp18EUiKhQrTxdZw4U/lU
dBf2ckMawEVBZ61KANjB4nuE+wFUN23h9Cog1b/GDtyg3J1vLXrpj/dQotNZVoV3Jh19rAxfLyTf
ZBJ3RaHOJGvLb8g/eVifYY2CQU4mYodpJy7U9VA2OLRDXr51GprquKO12RnRY3LN6WMSDdUP3UnB
QeIwNUzQtrppIhS47XmWdy5UIs73/YU4XNX3ghgm0+F5NCrNzIGvKBG/KQd1Bo8DKkLEIsFW06yg
RZmU7+OWgPt9u26Kzle1VdWKGdiJpEfSwkzTgleenFqWSDTiD1yjybdN8H632ZxP54LzoZtSS476
bLBlUGROhSQ4b3RL/T5b6OlmEQ6ReDyKSwjkgFV3VrK0ZqhQ4L6AhKI5AVig0NeDUbIjJtHVnXtR
LazwLsOfSvkXunL8mPfA4GO0IEF5RH9TqMYfMHKU9lD/gXNcTEpNIF/5FZeelImcox+E4ZjCfezL
87AoSsZtYMz7R4crY3Nb6hzIt0MSmgG5G4FMOdaa2hRLWLtD8PREXXUxCetquqZysVkpUvknZy8a
/wQJoyVMoAP9L5MHRuttYQDIO701F3RuBs/Z+KxtYPfwc0h3iKolq7HEOYryvCEwDNhaV3QbCNq9
S4cphQggALgIRYF2x4YyBT/xXrvz5GWvq29nHIwjEHKD43kIGS3x8K+DJ5Xh9KIRKf4cmb/V0T8S
3D4OGa3IgleFHlSPm5MnYNReN0FX3K+D9Nmy7OQZl5qfL9m8cRLkPmvbHWl8JBgJrCgDuVTa060V
ega9ForakFKi78FkOOR9P0EOVGvfnq0tRVGXex3TDg1QtTAiVoAJjD5GJjkU81i6FUymrAaBUTjW
B9/npo4/ACu116NaGAQAe/wNSQtKNR0Dwk0j+zvQuao9m8gFCazQwOYASUj0XZ6FA/CTkl04z47m
h9x/SmBpMjCJbgND6M2WktUHxaKSK54LzkLvL1JS29/tj3ytLd9sN6UwErh9/9bu1+IshTOoVIt6
GZze6dNxET0Puyhj13ZXxmG1aKGlBiZ/vjOFVcDIYENWghB3JaI7mbiovK1mEahra95H5UNnqsoT
PGG4pWZKHPp7uwMM6ip2CQaf8vyl8MUlSDrjG4fDuCrqhcrsJExoJ2X7LZEgJIMsHAx0zR5LWfiM
tHmNu3jK92AorTZ9ZciWQrdG1K74NCVg9FlLRctmFOIqSnNk6zA22p6siC//l2eo4EJyG652Fo0K
JRmX5T2m73/I3rhCpQGzG86X4WUm7ipNCEjSV6W4ob8Gbc6QV6edX9b37siimv/wqD/rTV8sMmBA
VfXWRW+zm3vk6OC60jJPs9bw8aEqkwz31IDniRYP+XKbR8spHmCkD7rjUDYsbODi+jqYhJ1rQ/MI
rtr4No+hQrXqLavEmYur14gjJQSOacgq8fMimFOY7F9/frCp/gm5k/dUHZeedkTLsxFXL1Voba0k
VL1bhdD35rGmsvtW0WR7/nmzCWXu0olsGZGBLa+rMHZi3hXZIQRwVgIMX2CkZtqPOt9KQsYgWru0
kNuSlGeyhAD5DTx0TYddL2GveIUixxqam2wy4IQWsjJO5ihu670nWCROcGGkO1sgCk3hfw1/jnOz
p0aiI8jeYiUrd6KUWvfoHK2PJtYVuNV2jB37ydfGbacogNdoYLWXFGxZYyr/MWVTTYY2SUiniUb9
H0dYujH4jViGie+qHNM6DMlUtMjF6vMwfnsJZMpxPIr4ZYUE02xCSv+PcNGx9xNYuDigqRb7UsHu
Y0f5Ee7TbTgcB/qyAtAchGNGaGRZ+IRz0iiNgD2Lim90/x2/817+VhC5dukCvCthN7Wb1v0LEYyR
FeOpSdiP8yxaRTidcCuqXBMeR2nUJB4F9uJJZdlymjlYtzI9dD2lK/cdVIUFiwwOKjWJatHzKG0O
wp96OBcG21Xib7+aBV7TLEsqxCvVajD7gswxTYAL8xtjNSzLQXkvofh4W0sRaao4cxpE7KXTbZlk
TWncrprUqh09blkCc2Lu8MjA6nh6jt1qiIAqjM3UdEbo02ufOBwrHNHpByQOLV56iLjq9eHw3a1S
4iM0UYwzDimGHUTybr9daihU5rMewYCNGaroEGwwVIF2FFr+2975bZZ76UeM0wLwCr7tfL6/OA6l
i4bvYWB9T3fu7R2eaDhtQjnEBGBJRjjvImVaMP3XZF7kjy9POsF2S+QhxsX9XpIkTdMVu76se7CH
Agp/MsD4bSuiTgcv+zY1VQRqu8HrvvQaZes6YGCHtdXM2dzqv2OALms7+fZH97aGAlUHXx/Re4o4
n6m1N/zsV9/s7gI156CmT9+p625dv43OyRk21195uStsILMV1tIiF0T3O9F52C7O/HhK1BCgta7w
g37Gyf5wI+kDJo/7pqEWc331EpaEEe+HRAEhWiykrOYLSfswjIWuHYjkiJhpwwWFORTF56S1uBer
RgQQ/5RFZfillMtb2dQY9vXkh2mon42CwJkd3cRcr370u+i3LCZ7Xz1dSJjzMM2lnWIrbqNKYC61
IFw0PT0xuZi8WGny4gtFEW09ZEj7XDpgEOim2cO62wminOdzXwMD8g2e132UU2rhlsmrUqebnSeu
LZsJ77gh9dzy7umEQj9R93JZSSnf4EBXEfnpRCxj2CaXZCEjf+nAf2j55S7odsd6ubVPUybVpGGL
faEh6wpALWCGEWwKDvOGt4Vc72QsMZLxh/+2x6boZxiYXVWtcdGLy2E23SNQcjutHJOaj4ADBySh
ylGuGadcyXCys/OvXOu1wtcPQFgqpEFhySbvwwF661ZClVWftgLAkzWwBqdMO8RaQdxhvErYsAQG
CcnWkZOvXWu6UAqQmzjlXGK0vmpdw+7vB7YLgaFotXAstwBU3bco6FVSdXt5+KbV5qPiJ2RP6WBa
sAKEMKOg8yqt6Qr99NAQSb5VsrqLmYBcwlW+AW3mIsUUiT2vUUVK1PbxP7c2BabFTZS7/eSGsEaI
qUmxXSQ1Djw1qn5qfFctkYJa3IzwrNq5cesLTJOUgTT69GsLBlOns0CvI8VS3eidtiJqM0A4Zmo0
Wk28h+BBvPYPr0w1HWghXMPxgTABKxfEesQCt1qIRBnbBvh1q/OuqMsmaXEwTdtFmtSs/nP3iOMO
aPwpemk4IEWuB08vy3bNAy71VNHjrg/JEtn9E6IpMaU+UkFeD82F6Zhg7OEYN2dYdq3VHiL5ZRTH
FWpPMm0kODOJY0vhTKZf02evw4Z1KLvJH9qD072vcb3vu+I82iXQp+QQbM8a8IIluXy4BpPg/Rf+
PrRMNLhAEwmnQozDmaT8woMgEyG6RX3/SrSD/ZZH0psCajZyC1Ib+N1rpv4SDrQLCK2nommJndVW
uH+yYZBW8/25r2NgYPvaJVddq2/GdM60i7A1mpVgHUj94AXkDbRQ9WrSekLY3+TY/p52MNqGrjwY
UqfmruwPj6ilTZ/rIHLT/UMd8W36hw2nTcFmNGGtTL8uiS/jNm0MvxeJ+XGZZzTyqjulIp3uwbfA
byIz1kMy9dHGLRmeQNUbMScYQJlxWK1xRf9/kHywwnTyDPhav9VbA3VVTDB9rSEaWyYyw3jIqo5p
5kRql+Eqfb5Si365nAcVueNde48aZXVxas+Ir7xEcZc1S9ruR+A159v+A2ZM596E7WHJa4X5FVWs
Do0tIBqyPkEj4LBSkTSggdIIpppsngVLjmXPrYRYSz96r5Ws8bakrDCzNSB/BBPRprHSmcNDISM6
M/yt6idGTz942B1fv0frQSMewzHYXmD4oMTGnhgE42zCoFq1ghq+DrgyngcGDstsYeGKkKSvxOlN
E9KaDHQeN5XNdbMf1HvR4gpYwDRdAOHxzeVKWpeRX23mihqk4S4FgFqIlUkyGONICaZFiCZ7CjkW
3aGexPC7S06Ue/UDfBc1VNaB1V18AtYDgeq5doz9MewpzxZvO4pVGX8Y69DCAV57sMhoNveW3Cf5
u9qQfAzUqwucQWPkkNpB6sIE+UL1cPPCqbilw13ANciiiLQlqb9LDeSFYufYzZYUA20UwNKLq0sv
/bB3FBLJT6KOp0FzZ3id3GtbykdCyiK/Ef7Q2chAYe3j6mAgW2Tj+SfhOHvcYGsnZFn5caY1+rNi
Ha1LTwVxDjJr76qDeZKjVA/kFgIWscGrX2fcfzmXA9JMNR6z6YtqjkwyCf0tw0JG3YmZHZPCTWCg
BIE8+b+InA8AmvCUctEEQ6ko+x8i7kMWkIl7MgoBlXhMKMq4cikyZHa0VXwtpIt4O/z3qYDNG3+p
QBJ7OjXxuyHzSDLZ9li9t6/YJT+GEGHOI6GQvK2gNTVfBqkN0/Gk6UK8F98hDc6jKmdqUL3M561p
/mfv9ZX/vvx1O8o3unJev7aLUHE8sHs+88PDkE9Mp+rq2XTgD1L5sRW+mW5KLKy87mZUde49N198
9AvYmQnmQjKDLkeroAiYs+kHY7qnRsq1thl1Zism1ayj9Y4stCiaYqlJL2MB43g/ihOQlxBXLWDm
JxG/Hls+zuoue2PAkjHikbNhajSJ91jC2qE5U7bVRB/l/ma+xEqMtNP1nX00FqzPW0zjabISU34X
6cMZ19yDw7VCHLD4hR93cJqDq2jy5OO4pcFpsAFu1VWGn937WVaCAM2OnFXcqMaaQn+NwZnsEM33
7n/EBNjDcXSODlOe379ZZxbSo4mppVXBIct5J0mBk70iIln3vG8KCsdnY1mkTkTxunOTcbjMoox9
aGisguYGXjwNiZRX9dOUfAcQYybQEyjsvPPpOuTUkXb9U6YSuq2jT0RSKmEBC4mj8fw4DHbBq2Jc
MtnZp5G0fIz2dZQN40fpjraGOxAru/doCTpoW20LEWRBh9wzrXHF1bQan+zbkVu3hyeEIRsCFd7o
TA2JN/ZxJZ2XZh6n/rVKzrI+9ABgUXVDnX9qhmWzUYOPCEvw5Jjn1v9VwDR7Zf4ER6iYercuIStJ
Qf3ucji/0iXU90/R9Epuo5dnKByiJFjy8P/WRdY9pvGt64Pa3vW3nAFMeNrJeucdePdsKSxhEbHO
ftsnjjl8LeoufAOE584VWZOGhhpCZ2I9nMNRzN2+lz3SkMRGhHCgNEya8iV4KsND8wwdwufqrjMS
AtJ8BUM4+U+1/dczSI194XzJGuY+Ul2fU47M50Vyi+nTOY5l/8S676ZgokoMjKxWXWXB2DCtIg+q
u6gVQMJN9oHgbL1Lf1ULXSITfoCYFCmfd8oxUULxKGbChXaKUnCZVDU44AukXNIeNKfyyXj2xRwZ
rooFAqCggn613j7t+Kmov729ebPdbSTrFdc95ASwlGgN7V5Hq3f9OKxj/33ULPwS/4w67c0+QUaT
lX/D/58sZt4Btdhgq/6zRI/4kU0quTTg3i8dAjfXNydC8yKHXw++cyjFnGHiGCuNAGGNs9OS6/k2
o3VZqg0k85bHFSZQVBgvpA87nA1M56WFyc06Rnt71b0FbHEUDen3My1IOs/Px3Fmu3i9fp8aYZ35
jayv/5IE9274TbdJjtALS5VYziA1pNNtm0hnF7F7oZJysObi0fTrE5LY9xU5Plu6eCztsj187FWW
d0o53IBQfqSj6ev4UDGPMoaTMv75YqY98j3GD+Q+gBu+Tu2gR5au//Jv3Q8ZBgNjP4UNLcWO4rfv
iNDuo3TvU1WJwZOxjHibchpE66/1vM1j4EgiVqOZsSkXR3G0zeQzEbg1yyKpgZlMlt4LptqjH3B5
kr7eawjZGsiagysf3dMNHsyhcruZrVvEeV67Uj0167WQo0NtDR3doNYlJ2FBMjJW7rSLPQGODFoj
BVt5DgS1JxoHaxnd3BLbp46Sr0xyj1jqzUB+6IMpUrvqWUA4ZebK0KEWrzzDX/824DoudVof8dMX
H87r+sjGzRmj6gwvwMeOdokyBsj3yYBRVQsdjVufhjfOwWrTH/fftVnda6+Ip6W4grqc3EoOM/gJ
xXoJ4irdmgDEbAu9zKIHdiwm4gh3Nl8/AJN9W0LkKZvDX5uU1bZauXuLo3udKZrMCNhGn3Byo6Zu
Uy/3oQD+BFuSpnTXK1Hdr9BBhTVv4M5DQkPpFT76aivfZg1740kEO4qYhoc4yQoiafnFDqN8js2W
8UGD3AkvjcvQYrAoPC6wh3sCBPdXMFD+9nf0Qv+TNyxC6sJQwZcK3DOL2S32VQvxa6wm6zysty3u
Umcqe9HrVDXkFGSYNlI0qsGIhfiwL4Q4UMKK3d/upj1SgG5YGOzDSrv6FMFFb8L5O3vDQylRkoyn
1HZEeye+Qy1GeWcK2ttSyIZI0qT4sIWGnMqfQQ+sYlgFJTLebsjXq1IvzZQkIfTbazJUiiCNoASe
NJQ6W13qTZHbxJKFVjJG9IGg+WgcSjLvzE51iJ843nxPUQDguNEGpWGfbwHTlqWpbLTpyJCXfk92
Zx8bDBknWROKqzIr3bAzm/2KUrKBDFfh15sS6CZIG0RcpIcIdwM5V51cXf83GcbNQ7whKikGQQK2
4/Fa1P3vN9KVfmYsqhVlDKIh/YtcwNf3bt87tefkMfoY3+kLzI+KRi4B3Bq9cMq5tlnORLNN2U3h
g1U087n7HQESUUPxThHVlX0IuRkoDAWfZS+ILKzmEbhTHnc3Nrm5VEdnsyaRHno483qJYLc76ADP
+9IKhdvJAn8EXrL1ywXd5PBhKv+91QOKAuEyjw/V5UfZy33EYRY21Bx8lRWqvaMw7c274mcZRVd/
PwlBZy2A93WJhsfCrn0/TkB4d1hIKKJf9lvCmJ48tXR0Yws2ZAG19Q8YmKkQy+k+Lo8GMlb2RzLZ
7xFZPGbzO0FqYBxBUIg7l2yb3z6ob3LQtKt8AiAWocWWunjZWD7rPRVXYWaRw2/DA/qHH64DCsD3
rhVivENsKpQklDOZIFKUxX8K6KpXg4ImIZD4ptUbRepUg9ZaYnbZ2+zvTJRpTpNg20DU+3d5dksC
0xGI6iUKjozThEj0pUuzIwCUU9xWAiqM+dv78gvfdWrNB50XqLXo2iYf/Q2Bw3SMJ0IN6MzZ8CU4
hzj5iOviKaitfTUjrKZ28bKmqVf43zVwV1dKcpnFuoUgxXtaBPkcWA6MUtooU5Lrl5lIYOKt68ny
czAIrjhW+5ICXL06++jehwiRNovyYmMrROhfHkuNs4mAD0dLxsEMnmUHbR4hodRvklwLm3jBB/Kg
ScF0tECF5jXu7vqKAYlaoDkjpKhbtPZszZ9n2sm5H1h5xNrDSXWMN1LZtreRHr0zrGbEeBhrDvb6
eJY8ZyUOCjS9Svn+y0032MUDqt/RZAVjywkf/VAsBTjlbb7cQwdlwOt3Kh/oGYYHYh/zig2UufCb
nD6IbCjZY2EWpOZuIrFEZZ1xzYWhnpyrovorsPcBlO8R948rE8BOPQ8rKmVfG2EnWsqmW21Jtend
I/iAnIZ1fM34tLdqJjpMKAcW+4GQyJ4V/Nduw+8ELO0TiEXWViQe7cSmaF3LsH6Q+/am8mOqKgSv
lOAfiLZoaMqHmR1BGzY/NG7yalNSksDJT+W+tIJ9pzeONhvpbdWd3N2TWIY3XqYsvBxdtVSGiwpr
Wkr7LW4cBdwu+DFA7u1bw1Wo1cLAE8MHQMT/90m7+4rrTVqQ+b4D/zyJrvzmQLyLbZF9bH2p9+3Y
ZrVmPMfwQOgJspQIk7hRKMwXh5kILPcgWExE9LOkXX8uWAR/YJYcttbY8nCCrpx3MnzBF8NN91rg
G4hjU42RHubPvidx4cVMwp2eUci1Rptg70k2AmBlFnPuCKsQrakes3IS4qmbd42923vrAyKJ28XS
e+4a56oCi05WHekjFQJUvSZ1LKEQ30qh9UkhLUTyMU/z+QDFpb2Lb+U32NFe76E1hgTnsY+Xbi/m
pN82cjL1gjqZKO2dcKHPRwQr4Jmb2RYOe+sytq2+pNuBjz8bAbI5gUQ7/878zc+NxTalv/ZpA4JV
IhLlCziDDjiAhEQ5boD+zqnpMLTRu5PuJlMtw9vPCVepeOaXmEpNooM88trzZ02gbYtzQwubzPeC
drN2Imxpv4xX13VCj8zfxsW8uPghY1St3yfklx/oDYM+G/FhD8bbsovQ6tFI7AZ91hiXWfOtS4lk
SQAjcFALrmUTQB83lC4JgyTh0tAOlw2IjEv9qh0b5Z3381vD8P4QZ0S4/pHQ8UCsO2cXjp+Q9eo0
EzCmpdIiJViJ2BamBzI/M/giYECAzXHgiCvVWNCn3MAglGcFWLasaDlKopvHrivi3ON4UydAW8qF
RyIxNObeJFLfe7dC+3kKN6BJcKk7IHyptt5GbfEcSxoewR9aZ4+R/pJyxgweP2kP3Qmebl6DKqHG
oIXZCGbq05Pmh4GQUNA+cNfeJcsfQPB/6VR/roxcGAwOt//nBr63iijs38/GJuMwu8qtZnXftCiM
UeFWuIHFWbWDQBekOzvl9BHlDueb4NCKtEtwUJynlPdzaqUfSWg0eHTOCTFBaTrm5lfj/R3ud6b4
0Vg//5k0C5vta++ySoFGVVS81D6ePgdp8QkGNe0BUuDm4PAMjmrfujsR6w9JyQBD+bOY+z7VHm25
MTvOQCHcwnzhRwLzxYzbTnomhmiG/uKSnTTA48R51ruVKOtny0RYmjrPSgjr81AiW8ZRYO+QbrLL
nMeyRPBoF+l79UsURKCPbUhrPP0m+Iyew+mXRJ2+F+xXxELjB816TIPRnzISEG9eC9AnIa+3fhtF
9PeLmlZb6kfMtSfkyq3jYDN/WpcdZD2jC9ynjSdDKrGXjhGi1Q8kBRRJkwop4meBRQHnyKgKRGBB
XGhyhUwYQbDRYh0n/fymtEe4mM5wVAOO1koSTO/mvJmP8Ds8RfqprCHu6r6L8RSzsmLrXFOnBBVi
6gyxs60R3erL6aL5yU65NZh5UsPV+gEnRKBMl9dKOqHeE7440kB2E9O7fNfoWpoB+XaerhAaIByD
rKxjoXH0l3DbkJ2/dKEsEfDKabhg/RdZLvJ4l/0K+46KNavQOG/spIuZRawJRCgMzqNV2Vp4YZrx
XQ7EzmY0nk2stqzi7ZpByhdkwCZCjqXstRWivfCPUsN6zofGifvq5fM3W4eAs2/fO4p1JO8/9jF6
c3Jx2dCi3Pw9hrpdytEa6xUEo6l3VMtmfIFgXBKuH9uJrfDYhgBgs+iomLf/m9K3pXr5768EoXhj
44m4xyacGu3WVpdv+mOUoWq0wz/LZmW8chxXg5T5HwRYBDEdFHlZ+o+TWNQoisjt1iGZIdw4ameZ
ooIhFHraxHrqWICHRC5HH5ryr5ra8OlJP/q1tJ7b5oM2GfMhXWRQ7FPpOfvrMifXwXjHPSULkQuo
/bec5PRw5tm+Q7Vx0v3dNKS4SxQkuJSCI/x/kArDaBPq6G4CYJdYQC7MNIZ2R5R3U/gV2KSy/oh5
HH9KyptOTFfwkPtTnoDmzsDXcp86Ox2MYHCfTo7j66DsNigEns1K7h5nFB36mSaKpv75/yf/+fG+
xUiRYgHgtxeCE/NMX80HdJv2ClF3M/EMj0yaQSHPeYI7+zQ5AF9rltQC87hUhu17MStl6iks1xB4
sM354Nyd5EcFGbZCz+1Y/hJXxDbjl5WFEahJgger4bD3cUcjgAL+NyKpaOHookoVw8+fi0CpB4Qz
bK7y3iR7WXfzjFQJ/J4qPQ4cX2NV19I4nRI+CldS0h7Yf/r6mcofgTG3POcZWKGSkb98y6VuozfR
3vVoPR1Uy5gDSrqIWOINGfDA7ZtYF/2IAIdb8qIM9OdpAxOR1Vmp9VO7a86J3s+38S2wAyvEprnL
MPrLsCskFcwIHLyh7+vrC6MBpnWdj5AdmpdeCIUwND7442tSs4Nch84pGP/8Iso3TlHBJCQh+RWa
DY3XbgJidcIfnw4GXxtW89+Q+KKexP4RsaTc7j5g7w74b71dl9ahIbq+/OA0goGNnXPxRNsPkSiO
a2NUqPibydzlBZuNfwjd904OV7dyhR8Jjifj6fGcjR53VQB4YxSJ1tKNhZUtEeCsf1P6y2+ijGPf
u+62vqGW8H5LdVHFdudJHSdIwLRg5/sBWtakDFgv63BqxZYR/utAg/VsXQ50cz6yhe0g25N07+HZ
Md00okY6dA4QncxTXgFbuLcFkFI9Nv7/vAew4gkuaAaM++PiIHCLJUeYJylB3KpggNyTFn92WYFw
2TPGhKxGlX3wu8PED1OGhGhzo8+1LZTNr09yAPpzs2FnFFbeVMSUrwpPdYr02zAX58Bxkx2J2s6n
Umf86QtloZh7M+pn4QWoZ1/lNeAhSPB6mt5wM/OZNLFcLrxZSuA9xQywUmNDbKFq9/gc88I6PTnO
Pv7QdASVGRlhr/7pUAIZo+IgTqGXqEdRaqamWyMRK5bHOqym5DNgzWkzSl3FaL6OGWtBHB1yovER
Ode8qxrR6AO2bPtZ72WGf6kX+4e62kIReNTS/N23rod4FAccETiEi42YlS/2FVrdLS1jjHI+BLXy
8fRrw1pBdZ7WxdOZiPx+yqN4AK+3nR7wOeN4zFfoH1N5L4i7dGf7pULWT6RfI1hxLl9lT60/q/Sc
Pf9Mfg+hwIHaM3jOv1oPuRKrySOVzHGcxTPHpFvESDNBGfOpUng6838BuGR069dqqTX1WKlC6owx
HFwmb+8unvh4oR+oejt7+O67qk1lQ8UOK8ULZRpKoXtVmk9Bxwh793/5mxeJsj24giC/Qg1DxCdR
KYVV5AiKPr5edVCdtFLm/FC32xEQwI8bHaIpdkyNmh2gDeWIhISWkZplScTAI6+3+6S8Cw8Cfd5U
dsw6QKYTSSAlCU3q9ak1g1N1veGKTgdn+e1EcKd/cJvuNpF/bh7Zy884se/VNEetGrM2EJvzdMIU
HpGD02XvYmyFEoNsxi/fQ5q8Xjb3fnbuoR0YhK9bHO1vwxPJDI2PBlQIob6CBu4LEDQkm7IFSFaB
0FqprPw7MIn4Py4+kFZ/PpM/777zcHCqXW3MfxlchooVsFmMKUSPL4g/QgxwXt/CpvURkghZrvFx
uyMfM74SO+fLU2wmX4oe3Tf4lEIB6XddA4pXYTuAs6bgTh8K+tSeRIUwv1t6bxGo5KFx/da2m5iv
2m3qFO0Pgf/CbO9odq99whM4LVJcR/zsEew5rhc3ONWbiNa1XzPNn1Aj90dzoU07ViSd+nRL1LIj
ljDTk9dXl+MMY8DU2I7F+9lQqcggjZ05QIelwxC+J7g8WqvAafX0nQGVgw3cflyyvTQJhD+CcV2a
jPBm4MNE2uAXnusP48DCam7cs4cJEFBnysypz++sSY1Mc6xoBWTUwj22tqlAHm+1qpGZO151ASZo
moaw2pdPWnRYFmJxKZ+uiGHXMRr9rRA6rotzFP6uRDC3itipOTXn6AFm9b9g7NU3hi2/EkAd0Ql1
HNGsRNn/QLL0cfLCex9T+txkkz9EbD53nBWnMTYBaPNKCdbs56XpXHvy7b5bGfPNohlT3QrQQZAY
7tclbxeUIAKrc95EMcmfb1N4ABF4tl12JxdmXOCmh1dhgRoTE4YbEMy+c6gZh/JLYHdLgh7D0CDT
n0jKZ7t61nDhPF9O2Vp2qKgtqxOtF+XUzxhRlx8KsmFqQamGKNnqojqnwFl7OUpUUZ01LhjsKHvU
E4SNo1gNsnHrecHHUakzlkovQ/oGc2kiBq4ryUPKkvOc7ysluSjk/1S9Bihoexs7D/DLeF0f10Df
BBB4Iz1ZUXrbisr2lBmG7HLaQaS1a6N5qfwxRPrC6brtogXslKIwkqMZKhI0pDoDcUk774GOfLb0
nnl48aPNYTLd6eypQrdlt2GvGzf5FxMwd6sxxaLhd/GOa7IzETQXqdR4PeMYTHaqPkGehdEgqrMc
NFargJeCq+vqjfPjQ5V0QmAyYm2PTAdVNdc3wbRokhKS89/O2GcbIJ16erOIHdyLgnaJLOuZDCJe
PxsQZ9xdAEoILUXon5UBvox8MIThsPHfj9+58ioueoLrj3vRCzwCHqRiBgCsZVdaS0eFltUcKe49
DLhvA2v6peBUjv/UiLyoZSdoBlG/Q5CfoHFsmeeQhTTOl5pTjH+YhN3Ol6fEXp+axJ72MreNaho4
R8lVEzt9ON0ggKucfZVOOMQspyFiNy5RVK906rHoIsbB+Fr88jqovmlYxe9D6xEfBwsjqzjVP4Ho
Qg12ubFLgNLQ/7VnRIfUFae/lwv32D2Ta8nRWrZ4siXfdv0tD7QIMs77BCVmVVx5sFvf9U/qPiVI
3drEZ5CVTCPZD06vHbRW40HeWZ1qHLK9gTftNTHNRHLRdSEGSPTUUNYQyiqnmrPwZhQ5ZBmBCccA
4cqravCeA8D+13ic1XPzwUWrDWDl6jvqi3/bk59UTPt2zjSgL+2WLHd0n887Rm6GgVMNLIBvry6H
k6v5p7ikVv8tYEkOUUCC6Kv6MuWM1b4w5w8e4mT0O3oWUf6fb+VrAUPk5+rhxZ504+u9wZ/KuYaB
e32i8fKiniWXKuiYkA6fF7UxZu4ruc/vicKMz4l2rTRrxQrvEq62CLX1u6Qqx9IAYt1L/lfyHwr4
N9JTFd2ouQvxZDW1lfTqUB76XKAw1Oh3aYPkaoUFJ84QfU2Sz0Gvf8WVIp3KnfSmFoBtdYnx/HfF
88x94mWgjSuEwajonvZ9NV+e4v4iyPPvczdJlfESKUBwlU1SACTgfWH433Kezyam6/PTzt0OTbTT
ZO8jHSTySCcF9/Vf4ZvNhAClpwqdUQTCRcg8pD2YPVyZTGHfFRvTqPKRGJkLlqXxL/X2kdYhjhzg
idyzgkwljbmzuS8nNlBmOdG3e5dC37ONv/eOp0zKUO4VhMYGYfIEPIrvH8g2BNUu2XuvIgnWbDm3
mttAIWBBj4iFfjflgWdPFBbF88zXigAmUWjusCGRicJj2mnZZXmnMkOeQbS8U0lUk+Zh0HF5F1/2
TFAiXkj1IHUU6ZgFug2nMAG6jSgtU/KJ46xymg4BJ4l8m6zS4Lzo2CxTnHgrfTgWUzaqk35MWHsl
dDpVBGAx10/hmdmNWtZO2wDXQ2M1R76UaSBigDPmTy4LP61hy99HM4NEPYTrxy939D/UzgqpjtP3
CvfD36c6TWGanMJvoT9FXSyZQts06ouI0zAkkOT6Q2r50Ma/kAFML6WRpA20ctPT2WGVTEXOQ1zE
O+OGradCHzo54rfWfZh1ksuZZBBE4VWgip7Y3yTcvY/NOXlUEhghZrFM3si8rkAT06mm7ifM/URv
sadvLhCfEHPmbEL968q5R1RHCTzRDLloJD63wMr03Otd9KAsK+UJwc1MUdXGB02nUcBzfZxa5pHl
NxOJ+Rbjlt+mX6ZBcb0ZTIcpAomGeS010AcMbRrCl+i345Noy5Ula9F06q5x6plT46Yi1s4752CN
RHVeIAnxIYYyr2Yhx9+vv62tQ7ewj0kgaMXjMQ+qyRKPtw/8vsisIUMThb8Wo5YakV5xssW+ti5G
QmE1y0uduy9mOwvkLPft/D2AKXg+n329hI3sSuhO67dHlVkOfPCuAYaetUe33LhjRmA34LjY05DJ
7857hLmWLTBM0bW5Or/rcB7CKeIkP8zgSw6tgYIge9w9mdTdSAQqbSnf4Mn/K0J6vWlCF/OWIi4x
Vd/k8+jDXQGUUijM2POTjdBkP4vnX/luMAHmysPQZL5DyGnFUK4KzRklPVN3jZzeDBnLfVSBfCCM
Ct7sOZqrz9aTQWguSkNnBOLd/ibXP7zzpJW4Z+nFQ9f1b/WdMCITqIHULOKg05MAW9qPnf3/aJ0f
6ZGIcONkSjo/ZUdes01U1jEHeByQyknuUdG4uXoA08C1qATfcQphvFlP7IXe3HGia0WQPbQH+RRO
tDJw2xsDgPqIrEFyUbEuTAqDoc0Bu5OSId8+hVM/qhy22PziCvwVAbXSQ8EQpVe1SrNtuIwu0Mba
uGvyzhQO3lk/phxWj/Dyxjqbmivb1sI80e8ww2gpLtRWq8E57q7zkMNsdDcOYGR1WZSv60BJ8nrS
3QjqvSjbwSs31IfBdhCgMhhYaM/QdtsaiHvBLrnQtP9ovE9HSsRV8e22jNjoz4KO05kGv+mTmyhU
ft5IisLAHYCl9AB+8cUSrzsP0bFupEahmj6Q+HeBrfGlJtwE4CylEfMG3T8m2v3lBgAdbjnzUpwg
97NyVEbk3ncbk1+jA9SKQ5qMuCzHmqGlcjrqswLygaDlBN5LDoLCW0FCoenC9iKfhIhGQ/CiDd3H
WbyspYSeerxmoXEEvTj/YrYytPDj5rzT3dN8ZjDtw2Au6dhVpr+d9/j2Hs19EnCvSwm6c3ST96Qq
tGg1MdCToLkz9DHIz8h0p0A5f5Sjko5Z9STeAnrePIahteG9PzlEdONkmkV1zuNHt61PA5Iv4iyH
H4grUsqcSBa6k60OOEKgpf3Lms0C0u7TDS+JdnZ1mKVPZZIglkgtfJ2oDk8fqgrm3bpJchrts+hT
BVFMAa7yj43m9pIm3rCvzu6KvqG3kQEt1OGhOc8CZ6hvmlA8k/Kmf7JOXLXmI9grQN1NkIeHu6Ql
HSatwFXSe5D14g0B6tvZIZCrer+90xmH+cugKqLU1yNZ2DFFbwX/6lDI0+xx/uS9DdtV0eQqb3BR
EB0ALMwtb3n8cUQ4L7Q/N6ODaGIRQQWX+co+XBbYOgIHWYII2FrZK8ROEQ2ImSQUkA4lydHl98vd
+9RSI6vcWa7gWryygOHOuwKK2lNJNuMqH1eZIYHyiwS4a1m4Sy3/ZnsMFuSzP2gzXx3gZymB2fWc
CWYM+H6r9aHWYYNB7NlGoFUwSI9XaQvH+t3gIbbmLbded/Nn6s9XWtaMHf/ZA6c7H42QQRDV0iX/
vbDMwHN2dGmWcmgxXNkflcZF8P4FtetOX8P5RRurizgg6O6PHajtHvgjfEl1MrWQQjVEEhAEj8Dt
uFuJ47jfMWuoEmciouGNrrSTGw6LU7xddkm9FSE3o21WQJnR+M4KTVgdMo6QNVoUajLvvNq/rVZh
KYDtXC6fXaM8pghu9L3X6h+TaCoaEOchvwhgzK4AxiQOW+KCyaOc2hR+PwUEZ+QDTFxnhPENLZjd
X20SbwMM3DbG8clsj36yNzYo609zLwVbgEqaVgjTepQ6eBHi3EwhBuU20YE3tESFSVfiK7s7j2BT
9/UOWUvPAd0EOWP/GqM94TdNxl1/DWV0Ss6OzEoq14sSQXIDzP7a4XaQSmagSWKXbQ3PUeHzZ/wL
vYpYI5MzYyu8NbB5++64WAKmZ9m05tKb9R9nMEB6kfxjc9H0krKk7uBOdbxqSTKy4bZn5SucgWQf
4uxZir1kkW+SsFROmPpdYuQdvRDcrBAjngaozOCdUa7juHsiVYGoajZgxxL72CY26a3/xm367y29
zUJPOiZ1NdQkxizBJs0W4xJKn7xPOESuz+IOhXEvog+rPbCq7+d6iEKfg69RutJGx/w3c3aDHeQc
gRh4qUUxATEL3ZFMEUN+cpIJrGxbWCTtWj2sDCi4msss5cVJ1stWAybrHhGcjOClgchCcc3JRaDg
HIh8rWUX6zZxAXYxRFg8ANlIfdjWpvujxTV4DCCA2iqfWQ0qjleA9hxstNLhyBe8pVcC27hUUlKV
g3p8DhYVZJ3ujTTH76qxWXvuSj9YVYjd2nDWyvm88BuBSWxEQK0IHD9j9PiMKYwOSAUhEoM9AIbK
ZitHZ9J8nVWsyoJOOMtcQYV7r8pIuRtOm/f+Z+c7lN4k3hb34PPpvVh+nD7vaGdFL4qAh+WND5TK
Ww4fRpDBFtCcqbkVKtdJV9ZDh4mfFq91VOsFbDvzD68AnjNa5pkUosW3hoHPKFDLJEd7/A4j6Xbl
eZSLDRWiwkKo/MmVzCwVJ7bXzeEib5+tSOA0FPugBFkj5h0FOwpu84e6cBikzzVggUQOV6nqZAe3
0ypNdqOwacQnd12/1eVaC3/WOiSFo15iMqNH/04PMwqy249Cn8HxMf2Vja+8DBjOYvfMvJHjZHvK
crdUm5I2A6E8wEuQtuLzO3RpsIiEc50dICY7/OxDWO5u4Hfw4tQNZ3Hkl2ZvEPZO6NcrGmUzkP4e
xbT8mf3Kgu/8lR1nMYWGRiP8kCGPZSUahqOB4YAleOwER9wPAaJvVWo6dM5NKowWHE7TNQvvqcy4
gDgozezO9EZ6wZAssgYFKxSre0JfYWigQjt/LGX66HTzvw6+8l5+h5IQnTonIm9jgsY78nmAElgU
l9uE/fA2qjb385P4ljoIJH6uV0VQPdKOMIkptzBT/7k6lafsqkO2lMRbu4uCgmKBfVFSOr6EUTe3
+aF55HnGjLIQJUWznDFprHu6ZZI2Bf5HA/aUJ8rbxeuL+5kSHLW90rzzuDz0ZcpEHSWRY6yHCl6g
zUJ7oi+iXHInHX0QbHmzx6xUs9XKMnKEsOZp6WyRbOjL0kxHPUhItuAFkgnXtZr9BeLhqSlQsHXj
9wwdx8bLAdxoXBH9f0uyejARRObIhBV+NAYbKkyTJIb7Qz4kAqu63DzAVjv/g3ElCGAyin40hIYY
5GnEIisEb128+CFOm1WKMGzRHBz+gU10s8PtlhZlcOyqNrxChsfUjq5A8CKyemOqC28VH/VOCtYh
xZy/j2p+SGa6lhtMnVIgLypw4wJvtlWnpkOryXhsnfVs2/qtG6e6dSi9VoM0nPMkof5VWUlhmntv
eSDk+zztzu+9+Wk3NiWyYU0msodEjdjxw/PtXVkparWqdTNQGq6QuUktGlkRDW1TewHasvOfuBDD
02ahxMH+zm8IZubslPvOoi7rlm9wwP6hRN0N0DEfHf1E7gNA0yAAuN8fcXqBI6gUOjrHt97X3X3r
vh27yYRyBvJ8Vl7XIZRuPmanhyQ/ZsEMFXjdObtZOUKvSmeFmFW3jg2XsViaxpdjvcRACUTWnPCL
KWbnEFJbpja+93Xus04JfJqb9YQTuN05khO3M9ywcOybRmjC9D0yOxiSVT7W9DwfBWHKiG5RHx7k
v1jNqoQIweJ9A8WLS2yTQl7nPlmCdfHel1+A8uOTfzfecBgEARVABBb3Vrj0E1zarsfsUztITh1Z
vjGJ9V+jF4/7nAEzRokol4U4+QQp9xa8cACNWNuXkOFxy9g7IIuZcVK7XONgOgpAsmZHkujrJtRJ
zEuNbCNR3MtFt4rLVCliloWippRQhAUCCoI/eW7zeFyX7AqVuf/q+vCvxFrIxJsWw8QBS+X+Irkm
I4Tv2cYbBqYRHtjA0x9BYffI6Czq5dddegdNxj+UWVDyk9tUgcxpjcwIcaYMKamxoYiipxRzaKkm
Qk6kMFBJkZesC5LRgkcbgjZkGP+EjyWjLW/vavs1tGrF7r2TYWeUXfamKzMXpoi4bVgYRbrL8Z6Y
VUThCEUJZOSMyQBBklpnr/VaJeBgwCimeVdECKLCjEWHUnKP0vnpwlG6Z7yZIjXwpKTf0wIb4AC0
rL+R/HXTA9zP7/5UwXnTMlxzLi04e+OGcHkJzzmS8aKsPkUffUp/f2mfkzNK16KvqZBNPGFHa0K7
L/HMjOQWYLMp9lCFpY75qb6/Ub5IFL2CYTO+m1H/pJBYmGNV6OFFFt/noyHWNPp3Z0tEDT4JdJXh
wvNLIQW/s3NdE+2MkHpWIUryeDj0X+QlczgLKkZCliboCMWYoLvdjX93ZdTR5KGZMqK2vXkQHg9A
rArz5VyckGhHsbVxNjdi06+XDN3p8t2HU87Q5Sdcc7TI2SyFHcvsWdfNPl8x0Cvd7b5mXWYK87uT
1/RIhYctGHsog0Scv3/FUbRxN/iNQoFmhzHnhubRR8D8u5Uj7hs0o5c3qA1adxy1TfNoMQKOqxY+
ex0Tzi0bN31VgRlIn8ltc9GBCP16VKnmXPmHu0z5aMLVBSvLBALjgvlIsVDacaqr3lt/BJ1ELO0i
f6iELlhgplL54zwcx3jPJmP2Z2tL9KaxbvZg8pmzQoPm4Jca7tQMG9Ysd6VhOSyxD7QTYqvKkIdr
wdiIoliIVCBdk2DQrvcvkDEy1LnZ+qkfaqT7EMWvEFdCBfg34DxhG0w7zG/XrlqIljL8eXMocyJD
cEVQyMSYL0/Jt1f3yQu0SMFsYCG2e2iO+GO4uSHYHuxhDBjdtssFl9cfhU/rilZWTyeON1ANfsiQ
5/JREtpn5008LVJFBCzBNvaf6Zr/+0i0VT305kj3MKYTOHAXh1u0D5ehxwYZ9+QZYoBxEfV9cOss
qUjh049yTw6/po1yNokGLoDhxU7/kGLmlTnrtSLeDj6O9RAebnAAMHlbvNUxpfqbtpGk6pS/dCVv
LWT0iUsEHEB8gnuKvZX11u6uRudgGQtTwQrhzrtYj/asL47Ws2vQ9IRVm3hyZVbYFP7wKr9x5uN7
CIyQSS5k0J2dZNo4wUuvkHKClNDhwNzpayi5pkpKuNWIU7brkBsAf6OcoI+YfBYV4Msg0pNr89QL
IxqDBAa+0AO2xQZgq6/1PxbAc3tE4rClFVhRyAASDz7sJDMCVxOnKmMAoOsAODEPZm/NB9Ej5e2L
CLfxkm+BHUZBskZ+JUVOm94tGcggwRBYPxAfqyrs7u4MSIsXdH8YY7EuOc++3CkWhQKkZIbN/BhM
JGZYJY/I83NybxuoTcpShRZtnqM//GWwemj54kjjIb5z1ML7IPoCJcm40R7je552h3ssGMr/vCtp
MPRy/BT2w/kCIuP6Q0iSXfM7P8Ub9ljCJRLKzuFVflFmOunHgc+X6JJTA7HQ+sDkbqKfz+inXCbk
4MLilNGI52zmfZodp5lZ1ZpuXt/OLhhRYhuQY5KXokB5/XSCKyJMX8m/6Dh/JJNm5xeGb3N66SK/
h5quCU27p7hnX6q1TfNkaJzUTNdkhLUKqlmv/0zW5/pZJiavM1OOQyCg8uVvsJCn2qzzptomaGUU
e9H/ms8b+K3+anXiXgDT1GBbA1IO/4R0tLSQ53HsH4NsjTRgXD9CoL1U9RE0XeZV7bUEKAL63I1J
GFnpJ8s4DRDYx/NMwmW6V/PVVs/aVKJp+agxVuag6XiMQoAB82QtVhEt3IEnEJFIervkaCAxqgo3
jhFiQyMkmp1MIFhrH5t9K5B+Dte9OA4Sk4YKkZ8RAlxgWp97jiBc7u+m08OoCGpeTuCrstfUbTjk
Fs6T22Wcv8HJRw1mJ3zBPBLErK83GY9t8qylqPZc13Za0UPsCwa/ha3i9yNM42YqH1HGPs3qQNW8
61nZ8Vdz6zlBK4J2xg7P/yRZRyGM8Hfs45aBSvyE1e0C/0AApV87CtAgYZ6+mDB04D2hiYTbSGiW
D/H3FqPlI5EUrxu3bIKgIA0XcinCjado6mIKtPLS88sI9vOAgGy7g0h2J06IXKqjiKfwF/i7nk/s
hmYiOtsByOmM5s4nhktfuA/bU5O8LvzjzirW5t1sYYwrB5f1vQT9+xvFhSjlLrEmQ9KjEfdCOq9T
fKwB6MMg6PZs1gVnW3kZTed+CR7BQ7qgAyeE7KKXoqq6RbiDQpXs0sKMSd9DUFVaftlZy8HugGzV
4gK4L8JXL2KTeSaOggIJtjghVu1SQqWwXHjssF8teH1ZjLUgDOc6ssNYTgIw+GuqJmDOOZvHL0cD
bp0VAGFvcB7PBCN3l+El/zycl0tVlkV2KNIyR8i0wNaTlDZG4iKyIDWkJDBuuxDnWFhzjOrzpns9
8cC8lFsVdls3xMnxMP+b9nbNuYI9WRrtB9p1+mi7mKZd1++ykmCDGUDziK5llCjYO9GPMdL7hic7
MIcj2ibCpbRbRpxAfXgCMgAb6Nc9YQWsE6LYTWK8Rkq+RaCyYkkEQyMjfmRzFmeBIOGsafpZgCvg
GBN4VUm8Z94g7y7pWYifeO7DzpZY1pleI+DSqrXGuE+MFjAzf0pnGF6nKLsCx6cbzLNkRHtcYx/z
FjLh8ihunyAvgE606b2MEIo/GrItwlT/ciBR4aoGy/tIbQStTmLjQxTCWorfPcZqmL+UelsIxBK+
GUfN6GkCb1HzWN7pIoDwQ5g4IT6qpmOuaGywPeHRnSNA6DIJitUJArvPxN+TecPEqxsB4jAh+QOp
pEBi6b7Drihnx3wKIzB191qPwUPwxu+MSzmMy9kobZr6862FA2omcqI4uySpbOoqBbrgLynJzijF
RAUtAffhAvB64JzhvaRHpDy4x9cfk68+aeUHVVAfgyb5yUfu34I+Wc0+k/hnkDd9YjkKM9VFfSDO
rMZ7UBN71Qaa9ttlMWtGihOgEEhNeBIMWS9Cy4Tcf31Gpq5vfBEXNyUId/QP9a36JsRsBNZdResr
x665fEnxhYynlGY3XBm/n7MQPrmpjA5VATg8bgXGAzJhKZ7aWto+Q8uLHk1qjUqowKmtxz/Mg0kV
HRVXYJw14b8HXPd+IVqcmse76nHGEvBbX9Mckt0KkGOIUPtRWvOQsYieFi8TKZzlPGWAr0eqIazg
lYKSGTuihzvH6Y0YsmsGx3eDVWRhI4b/WweYZERX9KQKF5hzVWm+XVEyY/ZoH41JGsXo973bW8nL
yglk1XqUr0DRr7AVNFEIBK/FoaF5TJsgl6NBXj2n8slRANsSWrhE4an5No6jOHDGF1QdWZaO7Abx
u/l0GAaQbS8p8+bSC35SopXdc1KrgvwT7L3ihyDliwoNd81Q4/dlikXfdTXsTPxUksDo59rScZP0
N/r32I2lFHsvIAJwaULXlAhu7P2/uFGrVf5ccEiOVOFztzaJBVZuPfHcVN31sQpZr9vHZjbWVmAy
WCeFrS+3A5v3MfhXbiRv8xJGfIHokG3la0i5bAp998f4JJqnAavgD6+EWddxeMMrelBUN3RFJQ9o
dVI/UE7/lu2HQRzOUso84f0WeIAzClaCoX1y7hrsUNA+fVXqgggXhHoZfoj2Ty6u1QPNnYVgEQIw
rCGAdEyHif1bXtpSn0zZHZ6oba9s5gTv+A4KKawMebs3sMunBEqbKQ7990aJn1ZRPsou/i7Po7LG
BBaNVNO7z6qI4hkUaB7faV+PgWXfK3xbwxXW5KMLdNQ/D7Ovk1hDqv8+BYLsN7f2ul8B0Niaacls
a+D7iXzxiJANw1MMa4f/r9IHxWGSKWiBrMVlK+8Xiu4bCYqSUYC/dUpKIoO+7rSM2ByTA1JNHxcg
KH0e7X88fDYkANzX+Sem+DzrZW4F44OjvbXsBKRZQ3GdFTAJPesqA0oymoeF5mXMzkhyhTWBRwVN
r6NDDf9ndK2e4Ga2kfSo4gxBMSyf8zsf0qnaQ6LTP0RnRRHsUU0lyp+NeoP25gSCjsLMvfjcm3Ke
6noUSR18wF4RjP4EEGePBAqq2y6s0/9+NUfOgmif8fPv82XIwN763MkHLnCTS1WZM6DS9qft4XqZ
oc5ceyF6wuf7ibCuGcAtSyQmUzR7XIQI/B/WPJhr4mnu1lry1HXuyHR4XfhO0DKaiK4H/iAfyl/N
myikkV0y3OYmcLjCEb6ewS52cVBgDFUZ6sqHz5NUDzDjzvZ7MwyFTIG3egc2RmBOr7zx1OjiHwWQ
t6U97MEYMCpMFprNf9UMfQtZHFRIIpobUhZmWoprE9ZQxqm5GizNV1hzLXxWl28hFrFJW8JyABYl
Mrc4kgJznXRDdZ4TT4rCt1VEyYkfUhJODdUE3NNERvOwVf4LyePLOnSQ7ohc97JYp3X7gloSv26r
bralO2quSpCtqg8ozL7zPK/TqQsf3nzlNVNbJTD/UMbdfOhn8pQdvjnAyKNTy5gSw5LSF1WkzJy8
tYUK0em+YvbHOWlQZjVbt5LivE5+E+OWvpDlhg1wdp1QwrRAxqsaecY8yYZi8wNBkWDDEZhNm3GW
DXJy1oY2qWyNY9FY3VxhjvtVN7tMYvJPXTCFWW8v0Luhr05AO4JCF/zLHyDaYyRqybjuIjwhYszz
DS1D/l6Qjnj/Fuw3MNBj4q/rKHoSuMw8I60LnzzPJvnIDGwrJOj7r8nPxmMKH5zxtxT3eXFmE5v5
2Y3VTllL1Sovbez2bUMAJeoi6hWQmI/yxaIZOJ+cmj0y+weP39OdMaOEZPQLxgHLoS8MjEQkSJOS
btKCZ+bb/BCUB1FG/b86FRH7KulW/3Py+FHDR8tCDNtIIs/dhCHVDegK7ikC7A6diE0LSQcP5t3w
Y18NlVD3DIVGL+/YoPRydkXrScJy3KQ5BeO6YY5e5MA331UiMdCAL3hLQiZvsvDEN3Qlk3rO4shI
doqaTyzFfqQdkJGC6EME+N0wYV2nWL+4DUVsNFXzFm+Z3quLvDThYPJwGTQTjjmDbDUoqX4QG5NL
kLmFYKO+SDzrIyMhokuolOlUfCAnehHmLOfbhrELfB7N5xNJSnO5iBMtyZneEbygSVxdlRwQn2sK
GiPPOUFQ98WlLWg5ffObSD6TO1BzN6L+CHtisu/9pSGHL5nLKK2KtQ2UFUVajvBT4C3/mS5c7D1B
DUiPrzhLiOiJzU5/pakf3UYx8WvFqMbCXX956czRTZJ+LmlwIxfrHKxMm+spY2fotAQfnv7HhAz+
+/yJ4/5t0JstPKkvMivzsopltIUX4btPtefBw+cyZhicG8alNNkOD4BCscLFy9s3XfwbqWiUjN6M
QIb0xbi35y0h60R0/09S2Iv91D72Iqadw1YaYsKErCmTghbgs5LiTJvL3ryrWrxZpp9xli/qKQoz
cc9MoDivCFCVQk1s/9iXUnyLX+pigBeothf0RjrqKWpSsh6GjskNJ4m/ql19xs83xLivEGNHoQB8
KKIuoTlvQusHwVBv9RfXEwBlV7lal5WIoHubIBCYFGl8fOAwTBMYfoOUgJTfmdKzU/xdQh76x150
1a3d3M/1G+sF96fvsrIoCzxIA2x6q+3/OAdpSOxGCG8KsWG4NAp1C0/myyKOgSKhSho9IoGyZLfn
wxN9dGJduOkHjpqGUkBaoEK6i9SlokAOlTtE7sJoyx6mqqZjKBUCcL5AgZ8zV1Fl167lR/qyirq9
Aq0tloeDivpsGT8LM0wv36IPLmAJ5pb4mgYnEZ3QfSiV9GAdO1e02So6AqqFbGTdGjFQyf7yD1ld
kJx0WVCT9P0P1kpRozI77cdYNW1bZij+rbt/XS0obtxXFa/xCGQPD1c24NbbCQCWanYgp+rZbfCB
rZ/9IPvzVo/BWyvZP5+yVId3wCww85B2ZC4FrOoUbzNm2hFTyoadIRj0f4rFIHMgSvpg/3ZG4jeL
cxNvuXe7YobhlMYXZ46XPbXLLie5r2SWCk5y+w7jej85XFey8Tv9RxRwzTvh3/97mtwzjIUXBvxz
vjTj1o4eZwe6XzpTTLJ+HM263SpVM7OfqhEYAAeA0s8LZbgM1ORDHf71iv5MkO79VVqzWKv+kG6E
Rotpy3DnK6vnNoOrBBnsAE8A4WsV3cGOusQGehxVpbypbJzu/o7pd1R6HXIs5CVIqiXqsN3Vww66
n25qa+Dc0duKVsm9wiApv8jJa0qdNTQNvjBSb4roCjmLBxdTdLHlQMYHEfSCdvUJuP6K51lsH7Qm
oEVojcUgHZ7kVdX1msOCSpzRkt4OyZxNM+AJbTyG8XVKVGE5i8gGVybDAC1XeY88n6nGGAJAAsqu
Cuwap9VRnHQqAXDEWP63ImV9e5idnMzc+KiMZUcdOj7WKCIT7UEGuUBcl77AiE12g1xSyX8nn3FD
bO3Vz5oVlWhFlAHMX7i9029LzopFiJTNa+MOjcSQnRouiHOnQi4qg2AOxlxtwFCKx7t3LiFbv8Z1
OgTNVywNGa390YnMIchm6EPt6X1e3KF058gj2atQe489DLdc8b198mpN7to0/Rn/5oeaZRQrCIaY
8mFTnpS89E257oUhBiu2TNeYyF2sMup9eUYlEsXGeMtBJOY/MWexNoOfdEhNWjM9hScGtSiF782b
fGvKiZW5orpXYP0OzjNUk4OH+5qaMuStyLGSqpwnj+vZ3AlueYTLdVm5RN/Cx+XdVPf8KuMF9hks
hqJz5G9Nu3GpjL2QxQp3621LpZWTvu8KCnAS1SNUsWAKckRBI8Jl//3NIeqE1pcO1JgiOvV8Y+Gj
apdQcknl/TtouxMbjJzXTEhUiaCGLoSxFTI8NHDsJkTGwRnFzUtlr16fRUSHIeRy3h8JlUuGVSv/
jwxJp4u59qSGR9cdPEqRn/EvSQ1135nPSHfifZ2zCDPHWvodG1kn16GS+EgM2Nr4bopPsW1QqJAv
pMzafDor+LnQ/vH6a9wuafSxGGxGKKe33orug0xbEPaf6+JcGL9WBKpoP43izVs62bzb8pFUMQ0Q
ODMHpL/rbesW0H9/UeqnUFlXtJ60Mc3PAP0x4LDgmJM1cUeHx+HS9U3kQYy/Deqcmh8iNYoUT0yn
ZBWVh1Tq+5ztkpU4rwCxU5wscBjbKtlZy7ecJ8Qcxsqhw29tvf16+AV2fGrMi8fHOfXr5PI5mun9
h1avDJqQkKnGwrPIqqQhtd+xoLoELH4FHGIZjUdoB3l/39JbUJ+dFf7TmwpwL+/+ES9d+9vlN8OK
1tDkAEFGo//xr5xWcGvwZ2SS+f0/PaN9XpOvk3LdGqE6WNplAncTD+afcCzQsEhro7zDH77VaJrT
++7IMcOLE0cYW7ZhrBlS9Wt29F7RSdwLULDzG8mI7ZyGUjgXvOH8QC5/imhKOasjKK6x1acOqkEO
L/xA15gvdw2UM4ywlp9+8NlZxw2Ek2A76XhxUEDhcUSW19WzHk68ULDM6ZeAZ6oeVPqsEoxUZqmI
zK/l9yfpI1oH8/ecMf1BGsUordQpBN5Vc9genUvpvxuhAaV3lPNyest82PibsfBAP82dNLde4boz
dyN5p0x/Hsa52MvbwIWrqTQ73JQhABPp5R4koYP2Kk7VWmFHb5MCCTmxrMZed8AwA7I3O2lNwtd0
DAb0G0GxNLdmHfW/Y4JMiYK70+ZtBadg4nNEqWbpMzIvJ7nCQzVqu3VfLLeGHiW1fw4Ik43QpecR
ixSbCQ42yeD9hhBLlY5jbVXWyepiwwCIl32b7RyoVw4/1MRhV1PWCqj+FiJ3eHt4J/Z77AT4PrMo
UOOcD6E1nK/bZeFtUpkvtMrw6joPRuhlQY7FAzkLCttLrjwSBK/RkpMm1utGPn937BKhPwf9TKmN
VkaxjLC7Pc/91x0dgf+couRg6j3V19MJM32BVljGPY6XUqeaSmIhOyp5U+AYlufCpXAJFBa1Uuuy
zQnN0CdHUwhUQM3TVfo+u5qDyyfMcsUv+nzV9HE0RX+MBrS8d2cjmGoX9UUXCeR2eDdOVEapRPO6
LuPXryy5hi33QBaptqetsQsQzrGoJvv+aERVGG/UA3mXBbj8rHZITpGQI1Kg8SwBD4hduPTMRpVZ
BEwvyPadRcHsYE4qvY4mKJNit/rNuhgn6IpbTINEl3H6NCxKdnYR8VZT1sHyHVO1g/6LCxd6JLRW
B4RfC666dqZntDXfIboLK/aY87Y4nQa+x4XOUkWrZhAYIPdc4qMEdMawx5Axcm2/KAT/xULwfUWp
RINvjScmaFZBk4YSAiufvhAxvx1CORNmDemdlVICvLSvskw5pzBFNGoOAwXbbbe1FB0hS2PophIY
ubn4+jcjM7tqlqORH6n1lj8nmv5wZp54bWgRLdQ9CWQm9zoGGBa020KthmMMceGVkuqvhVTEUBah
pK/eK047J+7+a4Lt35JHrbgTgLew6m71715mcqbaYpLxCltBjADz9iVolr/fS8aEpxsKuNz6a5w1
3hk0dkxuqhbASmj9Pkn2+xDdvU+XemVtTHfguX5/skWjVPAKy9NyH6qk2oAw8MsfKuooYbL1Xv9F
a3mjhGSg83r7rO3oOWtC1uU7ZgtV2bkIgL2IN54CpCq1jXvXOQ5/1gKnJynaLsW3i9cfJUxdMVMt
tr/EopnsHNVcIzRm7epXviD48AfG4D/9Xl+DFF44e7u3dxkVLkmAKeOTBo3veKA7u3SZLPrHoIRK
hKQzaRI21q2NM9DDsdWKIKxthstg/aaT+FmTduMCa0fTSYCff2UvrOGexW30LNlh9ryVK+2LgnjW
kqVdRKuDa48/kdLoDLe2VNh49TU+UnAMwqD+9yoadjy+erl0f5iLgvvjgGhjg5HZf3/toktbqSAy
YaSYu+9lwfBoW9uAtOZGNEC8fAlvp9gNaN5P9ji0IgXk0iJyf40zL5GvWSj/K6ku0GbjXSparxDZ
Oj87sTzDJyEau7taOENI6ul5ZjOcYbW798I1y1j1I2IHlEgSRXKz4M1jAAxyFPOAxq9MDgpb4orm
EIFy2/Abx02zAV4ryQPdwhRaaeswiRTvwcSTud0u5y1x3Y/DOhMLa3J+Cw6jsj38Y2vHT7zycLHJ
mQkAbHb+d6q/mYyuOo+8D41qx0NWWQBeI/4A9zvAAhnFvOK3+dPrFYXaZznQrOw6/oxGQgJzyWOC
/VqZ+c4+3p5BD7X+2JiBZjuq9YQIwCWFm2XW/2Cir1k66QuS24qKwfWsfA4KZ7NvQ+6DttpL2PrQ
W/NPQkauAFqOr74ORaNwHq20yatDo4N471HgmdL2uRdMM7CHTqh+shyqFFPJ/Ejtx9ILPXsdL6Qi
xs2eHqvDTkVt37h+bKD3kuwgNUJ/cmRILvwwUaI6gcPbFEJrA8nR3c0rH81X6FumaW00yrGPKlYP
EWKpefpz4tdSwrSScE/h2vMSgaP6W/hIk4gZkkUBJyDSlwR6kH6DtOWOE/QEAp0QPxCEaHOyFKKU
XojZKT55z1439/YWGaSLmachXdx+UVJyzoDV4EKuH4WmRWhon7rFjjIlW37IegVacdqdfcbA17Mc
ARwGhr7wj5J/Q/nYYSjtkay2yl1Lik6dDNx+I588X96MTBE5FDZPNqjg8FRVwodLL+m6gSPbev6r
jLJbMwNkHLEWU4GlMKLS1v1h59ejUXHGyTN0ZkUVXN1DqBLLNtqGO7JwXpraFSGOMhQyIyfDkKgq
o7nJjatbCQnkH6n1MdYVebzNorfzMFWiBuOKo/v38x+soa5wWJArfok3Sh1+vsBy9jcL7u8V8qzw
ZBwGzhoecXHYYxXlEMU/4VQSIwDi8jPOfHgVFw2XoGFuqPwtI5SEp3xWi+B6JBcnAQ+lMe65FA7g
Y9+WA5CDzcpRXk51JJ/5GuOA5eK12/IV9rZpcuUe2pkxy4lEyhJH+VtkBC8h3Hjm2V1UaAMeJUJ2
l3Jjf21Hw/y8NUw54fTMI7b62T7NhzOj3Uj2H3DXPU/xzGo2qypr+PM83eAUGXGiV/ZDHsP7RhoP
7H+NwXs/RDuyVCIFaj51XdPxdiBt6zVkKurNfsctf2pNMI6vB0eGv/RPrLEhUvcwapQpylVkYu5H
UIJ9ATgw06aFDf0PFf0wDRq2SoArD9RRXQv5x723oF+K9PmK6l4cO6FaXfj0sdcKIdhDr/ck7liN
gmwCeE4NJ5G38lx8AvMGpAAGVWEpm/+bScpWnA1JZdOyVXsKJdX7LwCMhQTe1YpSlQf+wkiCX3Te
e7aRiNOXkC+VC3cQ5yKWn99sp2JOirJOoeJ1ZYBDc5iu/B+oW55bMRpsgAStr3NTpGNbuagKVoAe
GAgNZG1N4a49HCMhOMPb41eFs00Sy5tBZPjpcTTgZompzwQXihHeqdLgbtSG6mfmv7+v3zNdmeqX
YVDJsa+leVD8tre/k3jXS5YePyXviCCUeLyx8ksGnqh/UZWMFgY/fdNlgJEU4ibbiM9ZtDEo78dv
Y6srG3xHdk5ngoxBkVX5CS3hXMdOmFwGmmfv3uN/NtcM20vanj5/FUL82R9k5hnVKQDM+Z2hji+M
Qp3I3JrNOrh7cRZRJqki0cmP5f8JgSiasyDV+12zRSSSWG/m2sH99xN+1uyuqrCmL0ZSsaopVHTM
jx3JArKty2xKzjoy0/kuqZnXk0pv5lQ9jiP5oBLSjtDsMIJ6Ojjy0cNNDRNdCxYvpykCv4zVGwDc
thnuvMEn4qNNaM+5VpWSCVJttZ17qQbLeWbGR+dlNc7M1kD/bJSA9fU1SeX1mmsmUxzsCHaYYIXs
AU+S1bmnuNpn3axg8+OUbPtwpEJkYDPxZmIQ7y/JL0+mKOopGkGSQuwixHnsf857ba1XC03r+9rb
RIoTfuYxaqFCTStBNnHWL9dD2QjjfhfivfD39YH0TsnVDRNdWi8AQ9Dl2s55pcD8qzBsYpRwMDbA
UokTSrTUEvapyZsnrm1zO2HtvaQpLN35W4nxImjEvk7hNRVY/xCg7eO8avMFYenMxt4O6ssa+eUV
zErZj01ORLMuv8rAjJysJ42Z0nUC7SqHoLtTQpWtH65anIOoy8P+Lp4X1xJ/q3XenBhQ86YfKZD+
JiwnK8W3wkKjc+lQ3LtW/d4xJq3Co0dx48q/MC0nnJV4FqcvgRRcic+JZVZl15asBzieuN4YruuZ
NmlILSnSA6K6IW5899DPSNDut4tpBiNmEglE09kLrSEBeOsFQ1uobQW5EAQ+0a/5/JCj33NNtEi9
pGwGvlhL/DbYFYX7udnfo1ylNLbDC3yKlABGj4zY1xrOUI4ocS1k0IbaEFLLgVyL910yPjMYNGwF
9M2s6Hz8gj3QBU6NSzNpMWFzuSem5f0Gb2pQPjLodgWecY//CpLuNj4y8Wa6KtMDe7CLYmHpst6a
BMm1kFLhtpyiq5JV4/KZ8mrhjZD6ysmnkZpF2UdN7oOpziqOBeUoPHo2yEQ9/tBqdq4KAlxE8mE9
t/ZceWim+R/WWSYQqnMiPSeASG0yIAL60BRPIfWhUl/4REEn02SMGSKXYZSXWIPEJdkwu7LMXyIQ
JCvVK/Kwgk6vrDw5edqweiLjfWFoaH8qfClG4KQMnMPRIYh95PIHv7PjjDDwV1LbXDqdsJupwAxE
9lLOFdno2du/qrs324LmDQrKudsMlnzeYeN/1sm1W/4VbGcXwC4FuuN8Gq8wnmdmNiVa7LfX1jg1
hmGIll0NYitC0dKQnS4+b8rBq9e0Rz5zY+08zewzQJwHU9C9YfnWYjAr8uVTGS0q/7ChjdCbhvO9
tZZViHPjd0b1i3zJnCbvd5lrNEZN/MMWssjreyw5arLV1UuY670GPmMq9BgdJOqv3xj5KE8DxPEg
eEMHqsw2CffoBJMlSNmvbQEri1En3MXiu3TEKiei0ZfsisVAPfeWNr08lGvkF0Z1DcYivHyO/KUs
1OdjQ6f1K3kq/whl2zaC0+Hs2EKQ/TeUvlmfM5fpgXZ9OagogGx3MRZq4ZUrVhz5UAP0+5wD52N+
UYmIi4jeyUAAnvHkl2ZzwZ8gV20CLZNTPx58HHYnYJez3SeViK0m+DgRq6ZyHsoIuY89n4AHSQuB
TIAtUG2/9J1zdwU8zaD0Jw6Bd6WaoJAZalnttzfgodJ93Vl/FfK6lAJ0t0w5bV1b2x9YXGzLgOWB
k+/mUmocwl49Xi5IX++82bPnDS0Jyg19vPpS3amLz199K/9s3W56xCrwLe35rSZz6MlWncpefwuK
tYrvDHUiufqB8HqxuPu2w8/qODzp6RKWWilGREaHaVcvd66DSM/NfD66zrXVO8P0Hsx9cgYRBzzD
Jb877KmE3/pNdJTfXQ8m9tIwtlOGUx2CLC9KFNFZ8ARMOnqbe+Qs4BATRarWouvksa9MED6ohaqD
lON9YxCszUhk5P/Xz2k+lFTlsw+yt3eqBSPmYHE4h9QKjAlMr/b/IrNuojuezoRX1RCIe6D4Hh5N
+kum366anWnFnP7pny+M3wBufijtKIUe6j3bbGKgJbWPsfkDIW8yGK39sqCryWyIQlt4ItR0tI5P
VGj1XaasxMLuYgTUhjPNa8vmJYGdF/Hiviui3RfnF8oryad5tYGyFFrtgHJ/XHmVBND0d65O+91+
dIQvmyi4BD5gfpgAmcHtu5KzuRBGGX8Zy1IibN1oxzFyaMaAkGOh8GkGAFEvBy+yumeZFk6P4fuj
1VUpLlvpDOtolan3dKrs6JrEa48B5fxxo804SwWbwOJKqkw5UUlsMMKV4l/lkQLBFIEPVLvsrNMP
G38vblmfD92B/j1/HdX7N8lcNgsHNX0nwPBgif9CytN+zDfjAmgakB+IlxMev09ntfQwqSEh1MSC
QrzK/Ba8yh009c9csRBrotBoSQ6nAubr/k0gjzaJNkE8WSyBCP7VpWDMjdITmZ91ku23h7F6tPsw
fKXaYxuQxe5X+IDrENw9ShVv0nnM6JiG8pcXBnaSI0FQ8OiFrgcRPiawk2c9GdU7kmFH/evHwwpy
s9HsxjSkEzQ2AjbUhvv+kZ+GOlD8GRlAOXw0Su8Z+wC+IFkJuGamcTHmBi3fMvajpbe3J2fZuJrP
sLbENkVt98IMjdtaCOqmbeC6RR1SfKiTPrmaaw5IzMQ9MZrBOea9iaIvj18OecXIOosbnXwW3Ia/
qt7zQu7WWy0BRWJYONOQVsAgHIesCGbLhmg8ePzuZeh3yuvLR9ZP4vvvS2kt2cjcersuOSYQZKwa
XnucEL4e0+uW3Fqt1lv8F/wSOyIaub8fFyDhTa0Ckbx+iSwLVsdXW5gJqKzSE753x6QFbIc27qyV
S1aMdoorMJRLa3O5EWQD1UGQ3yftozTnodAhkANzOgDZ5wNqFTcjEQH+3lUsN1gRgKFf0e7vfUia
BfgplOBz75p5eAl8BslE4SoZvrZUM+aGi4JuzGpqIu2iQAg+QaP5Q+7psqy6Kuxo+o5s2fs6qJMj
xSYDWK+/iCKoBkuuF8rSiioCICNXgYWHouKwPxRyVHItB4GCrE8CdOr1a/iLCmhmaOFrkXQ+FmMf
MKsmzq4C47Shr0eKFlIYvgKa9mUfP54XWpg984Zk4j44tMZwD687qB9kJ1xQUX4KSvhclxjfW7dY
kfzTPaUfDSczkQ7Qzjcr9+RCh+NRB4QN//bXlefqMArkpjmOkhXvfwqF0+RCYvC0t9vQoOFdSF+F
d3qfR9BTs5Ob+Xuxfku4BnUZxB4UTzfUuWhTo+3FTfFRL/jF3y1yGmpXLBZLlHSYnLeMWP7LEIp1
S4tpd04/PVow7qR0CqGfESASTWb0Q2d2SZlQ8no1P2vkLq1elQHXZT77ETI/8iSM5HGeeI0kIb8u
Ba+PZBCDzk7Tm3jhCNBal2Mf+RbpA8BuZ1hz/5HIKarVWixQBy5NSQhIyLdQCMonj5wzYLoG8bAg
GTjf1yXYqj/NWcF8aJkhVdyBl+mFfsh3vn0ixlxI2dKKXftLmJBMMC/udlIeyEs4C+bQbS9v//FA
ohId7kH40Bgrakq+EQNrgOVET4O39DsLfuNe1a9R96ahJLnm1jRjQOqmjOuYxfduFSz4sb5KIdlj
4upr1NoV3/SlGgS5r2LyHFfdie78acYmYbBaSea7A3nRS2GdTjaybD2C08jr7qGrMLvm/PjtpZ5a
3X3QplZ/MmFXFAK1lr5cl1Z0ai1cFC15AL1LxuJuMIwMfduGfmowufKS8+ZjZVwhO5M2yY5/Qj6D
k0Lrup51xbVXmTrWBh5K58XEdS7FgxBW4I6vY/CRXF4yoa6Fvg3sLuO1/IuCEffi/zSteRkRPIlE
IQlABdduYqaFFzywWff5S9+Ev5wY+1kmHC0RkBDGqvBb0TpWUjR7EG3iM6R029RRXel40B2kY2JQ
K06R1LhxuHPVMMxTBd+q1DN40rMyJ1ElthYHpDGn5qwP7SLNQgPLBxj2CZe7s8LEDgyaQh5aIBPK
2lQhjGh7HT1NcXdOTuZ59hozfWo5PnP9mVG/+ToYb1epJszMQxe3Jp6hZ4A0GgY43K84YkkbPz5B
Z19XfqNw3RBf8Vv4aX90Penoajqf9oNZ6eoGMzIjkbQONgVo2zRlB0XzUVrV5OdLViShv936+sos
l/golGNrIzen/DEdpMt8yS+6WWs5cH40FepgV3yQwZvck0ZZ98XJDHsoyq5LQyl5OFAl9zlyM4i0
zaW6VZC0gtmOnibu7RUzlZND9UZjV8sQveY0psTVEgQPWLbqpiwVMjiFR8/Bx1NKFnAnPEa/rHIK
5d9yqYjAAAe40A7Vx3rzbP7Qiic5elOHUAp4oN9C5z/UHjkRDie2lVI2B4w2VXnqvufi6gE4Dwcm
cksQzPtQ2p2hBwJhvOfJ4cI9CzjIpMzZdA9e1UjBDMR96hPJaTJlSGNoxetQhVdjeK7mDTMMm3S+
tckXVlAjCYw8mpjoTMhukH/PbwqJvnfnfYLcuptHvhck/GhEC6Cln/nXnxhwuT6/06kr5N8nzidQ
f421T6ltoF2w+Xy9CAvzvf/tTU43Fr6XiCqDd8u5AOZkJ8EIOO9NUNrbZY9/Stre8400Kew3z5U6
ozUOw4M5Xk+F7ZKILAGunJ4lX841+qcyzVhBV0vFZpD9pN+0UJ5HLCDiitoSWdCqiWBlhvC9shFq
c7ZLL2QcuGv3v7N/VR7SrMzyvdcQv5NLIhLoKlCv7034bOSNDjnnUh2sIBqeHYFH7UMmRMPupHGX
VEw1rwzKddrr5Eg1fMPScsK7IORGysaA2wwoHi5Ssh4HUYsAMpW5spNSGVvGT2eUp7JYJ2vc/pC2
lX3uwhZspfP2mSzUbPpzx3jRbVD1WesaKcmz+1pkXfbl5qIHP1AJesYQNt2y8UfhLr4FES6i5mbQ
kodGsugZmSy+9nF7/jiLEmmXYuHO4x5VIXkbaJlckssQg+pv6Fj7URF6GK4/GMOIsiTZtmPpNv9F
A3brqs0IOvx8MHa2k7e/iPRPvrbgn4iyuGouc5dUedPN1cuonJN2/BYC/JgaGuWraeqS0h47gry8
tyfLpkwIjjOjccNIfY8w7omIvgp2ozvVVgRh/yMYp9biY7MoVQjyhhYiNvvc7Vv+h7iw+kRm1SR+
yzgBeyu0sMEqjEP9wqQjfMP4oQW7vqnJXDzYKW4Ft9zCmRoMp/91mb3+jo2GwJfRc97KX1GxBlmj
qRY0SWAhy0sshkLZatv5OX1nBykHxJHEvjmyfcsk1mk6gzOWSIWTXywDLzcMFgw+sVU/F7XR8FBQ
1+FDtLSC79CKAbiJsUKuQF6OVbDOWmHEHqqWLoJmNcuG8Ro7xaJCfNEg4ycbgCBZKwirBgAOO0l6
AniEvpIkOptp6YxT5DfoORcwAcNcusu0gixP74ZLTgLpwKt/Sm22X3Sx8drNyqmSsxvVTLJJ/VRV
GUi8opMSyX9yq9g+BFUmJFxH9cXNs4TyghalJsCo2TXdcJTrS/6jfF3J6BpvRkriOG9SHWe0s/+s
Pee9Z0+hrnYnRVxMidrxgYBvWKihT0zXz1Lwsoy0hLOORJBXetSTm2qHp/u7x/F0Pf7Pkgzt1Mh8
aqagMULmTOZvZR/kafJ69Bp9m8xy4Oa5bh5ogFg9OuNiihI6cIZQYo9UYfsx8+vgm8Gi9UFVYGE6
ESTH34fzIF/cUuerjslxOY7ho65rA/K79AdTSCkSeivSq/k5LHSAkqGcH/6OeFMn37hOcN58xvUF
nvf14EE0ooZ+tOLDx2yl/hzIMwXvvrR25Hgg5xhZUvFCBb2bqfr/IPu4fRqTpVLBU5qPYJhPpUAe
Psnq72r+e5qXzAy8T2zWXGIcr82ldQjIeWlIe2UUePnK3dBzyQh+BBDpQLXU4sZTOW78uCBIHK6f
s2yKf7yRHG8fxqvTg+cVKC/HhmSgYCUxcLveur41o6HGnM0A5s0D/qkUpo1mX3TkmzOOrg2+sq1s
O97HmNEd3agQqSIVx0PXP8I9sBsfNAQ+keeQ6uNYuNmSPOqCwhYpZzBYLKktvOLmJF2mqsHrcXXr
hfc2euUok2WJSJutbI0uoEKGiriIYFp+6GxXm8BVXJJFX31ZnUveGw5ouEECnKdS3/3THCB/idDm
KNdLdbhycagrn/EUK/PPkkXyOyX1eJ2OxmCmzIoC3zQuWhyaea5be+BPxUcDw/k7Zz++FNowa007
wDwFNCJmwoXsmbXLw6SOwSsTT9Hxx3jpyUgWxast9ZSFbJhyKXUeEgBsFmV6mkyeQJ1+iH6GJijQ
PznNWoBviy6mYdpg+gvSPDzIyTF6p2B6wifdl8zN0IewRhE6tOAyox1mzK8abKEFiNbbze616VNC
LqXGmlyRhlacAvCzrl5ZDnnlb7tz4mNsViNpuoa1PPW0TfcKb3O1Ym2yiGVwfxZmKsgT7UaPhxEb
6RTwYwMygiE9TZ3g4LXT1oNqhxvnRCrIlVguIta2tCy3eaBDD0l0iUL31SmYhrYeCI/YzuSaViiJ
vF/6nBbo3oK0HlWVda+HdZmUzU9BvecE0yIBSmRmiq2cSxuzFS6ku2NO+BssBKasNIYTHCCWj4Vx
Sk3b0KLEvE6ELRARIru399Dc29ZIQDKxGxU/GgJYNr5T++NFPS+clgXH2Y/uw0SqiwtRpt3gA/Zt
eDdIDw5wVlUdSKD5noqLRv2QoWJSIGbEI7UPjYfHUtq7evpSU1/c5IdXvSXzdtgzoO/FVuiNb01C
SRuo1DEUTgKdVlMnblvReCIcJCBoTIjz57u6RTk1GfV6CDYo59roIpXojbDGcnAJEQTglxWZKUJ2
YKC0ZOZ0HMbAgu70EnYL6vOPMcDe+mWPzL3zmfaw9NaCt1/RydwWjWKycVV2bSRabz3Rz+P2x4rd
CFuyUpJ5sIrNK+kzyO0IXo00JKEdKXnmm9/fZBblszUqFliE9K9IJq79v6BESs7QuyfPz71h6Rf5
0YwdvrsSq/TaucPz7ZTctWybyjtFokU/BYv178cxbkuB+BKlnrOw0GIG5z7z2mdeU/bxa1CaOTBJ
uXIHnNMFUi08RU08RMICxfiDvL1uKU03D0PdZb+0upFj6bWm/0/r0+QzdLSU1Esi5r+lRGwxrWQb
FhdqtUoqym/JYnGOUOEr5LFnHqnHAiatZMZKyMhcyInYOsG9j0908pXuyzTlxqxpvTTqm2lP7w0t
tuc/zEPUxllSayUDpjiu8Dk4Pv560oU26mmEwE39GuUb8BIsuuEePwRXWTRP2yC2Th4+rj/etNVW
KxO2eBz8ZgoMZS8vCjlBVBOeL2LxOJYPovT2xTEcezcNR3+OGicJ4jNAp6Z6NMdRTzW8Oqda2vtv
PMWA7o55PK7q5GGad7LDAGCPeQFaOK25q9vz6UtYvYA7DEzDmgsuRacNpsLQydRKdPBDGL/IdNxw
VkTZuE3UbT0Y+ynBcweFObKw/rOaFO9610UcKBMtlGXAyvD46QZu7ZodA38yX3dB+uXUCYtS753k
j1aiY7WyXLbJaAKw5/HFgRUX/tWZIScpoqbGV+OokEVKRFt1Luf98D3/kwRoZh45Ghg/RBJTEP2J
6Y1ojx8sePaqE9E+TpC4uKikWmNiSV3zp6rhv1DrdImrmhzCtoHG3/tk9w8Vn14nbV3Nj45vk7gX
zhyEYd6Zc636quxZaFWvEn6KAQ2c1vMqewulhplJMfUQ8Xy3TBaEyl3j2wlNiO2nNskBlR7wfVBc
ddai4lfwSksqRXCllb9ak7bnWA8APVtismxrFsefnW0U/AWgyQY2gzSwidz48VeS/BistFB49s+P
Q+k8pgbJwv29iiVZJAh8vQnfmnx9Lo0XXs3GHJVXTVaBu3L1fI1T6SdmHEgi52W84NZ1xHjpQE10
v66jJP+hA5dLUdewnQc9smEtq1PX3PuHXR21D7B0iiAm/jUAjjaWRn071kuNkD9+ubgKMCvi5YaG
e4ZeIyYC98np6Bh7uGGOT+RO6axpy6lQ4F9iFpBJdO9k00RgxGL4rmfkAgcNzggEl66qA0ap+fxl
a1tGPEdQSQxa7YH419AaukgbIbo6WE0x5iEJTTIFPQ6uVBsNnBKfH11pNoe2AIBpvoe2nge6hDax
x1Rs5ICLX4z1wPK72iiQ2NdMXmdxMc/f4KI3MbFR3elqT7CWyb+r7wtVE8vZiZxb+w56cjazr2XY
3tmWF9BTd/qB5Lq9ew3KhWMyVCPTTeoYP5KXZwgJlllMQFbPc3Lgm/GeGdCKYR2WRGez/uWmXOVY
q+wxZKPUzx9OWfyeynHO3rvY3fz+XkLoHcn4ESnkxGWBBgL9F/u3ytsNXdOea1Ww0Ufh9mXLTGbV
oeaGNfeAEqa1YWuGRHvhFyT6tfoK92NdSZxAEkIHi0xPDv1bTkTV/ti4ZN+Pdva7mCXCO+X/rCpG
kL/IqykozSd//YsYWGCwEE089NiLaNLXuAwRWmys+avOHbPIQK6pprE0ZLYgHXzdNHHJb1knhWr5
KzYKngxLYE3mfCZPs4I4YUT3fk9chRQmryVjNxM87gvLps191IiiNWpdZjGXgl1b340IRYDE0TJx
gmOfpmreO/u9PZMy8DAkHNcga6p7ZuDqrASvgFO3GbpaoHPxxUbnLOPKARUjCCEebuahv6EkSvrq
AgBdK7199I1gw4iwTb2qZ8b4Pbx3i7l5+4lgwdmcKzrxyBk98VkzxmzSfkonRuOIWJOthgY/HcBk
rzLoAAtqmpmzLZzwLHzHRzYWtDSffR+rg/YVsdL+zSeVcyFFTE5BslpuhMmnIeebQ5hBnIUBwc/K
4hO5I1d3DlOLnu+VoTQ/Rh/tV1uRf7+WOqD7YHXEK4QFFYOPUuC5LGyqEtPnmzzgeNSykvcQUdjz
g26XObD2qy+ua/O2RfmoE88/LQoIjJQvr4ARIFEFUZoMwcLJ4ydTI2lty0k+JseH/jyqnmqZKk5E
EBt6V/tRax4BkQHak0SFQUTmTPh/sKgHuNg6Ziy86rAeFvys5KuSZhe2kpfbnXvZwQcBzAzkTVql
fBMmZB7ohR4OYRJo9Jq5JtA389QKC4gqAMwMkj330U849PH81tRgeiR/RJRT4PiB4y6YeJRF0c9L
HHfqIrxr+/MgeAT4vDkGFPy3i2oRADIpG2Xld7QHeI7aiwYEwHBLYPJ/WiHUIlXhPdfJFFZzlsbH
OvsFAkLMzrcU3cBRQMO+N8aNjwVmlajCv/eSt1OXf7+evtdbSsxHwc0dOtsJ0UKFkgwz8wt20hmp
dXqfxIKvoX5osNJo9LTxYaOOsPjpwonvoMTXI4FNoNugkRB1Kc4AquRk1Pxe4pcFWp+/gvSPowMv
ri4ezzzrk7n4Fl3GMYRkS2qlrKsPxA0u6Kx7rd/WXWkR1pT9pzdoGZF2GOtJHGx7wZyWmhPgrpND
nVwTwhfwYYD/jF+HAuUXi4pqwuROGTWKmLex+35b7fdaYT+5Ho73jR8JI/L5lOXjvLEAd+EfIlsX
cYFQpRO4pulBde3QEFn7ScNbeIegz6MMs1Ji4sEPD2jxaDdHHqfgLuaT0TSise5mInH9o3MK2hld
2BQiZDtlaSAI3m3OjY0ukPvjIuMAEVlPE/ZqcM2Znwg8KClIOGNexXh5wxe/pwm8C6G9/eMCq/M4
B830MqjSFlJn1q5cGmAnLlhpaXQFFVx1+fEnqzyAbAE4+o3EhwazwxakXk0S4aHjLP1gq8koj1q8
+c3yM1/Ewb21NzlU6o5buHgIpVyOt0ieWeN3hJb4yd3JmLIHQXBcJIyC3NfyEQtGMBwRqtnKyN9X
4joUBIRtxcwcJZaq3mRhE3NkBHm6bzzSKiigsb1Tw055S+ZFIHcqL6znE/KETwlFWLyx2UFCL8Y9
7uDlMxmyNE+OCSKU3hNYu1BQXHpnv8irUEsTdQoG6QCireYTok0EsQEx8/i2j8O+M0oiC6G9Og2e
XyghK0JIlNHpOw7YZXD9yu4klHqmaeAZFkKFFaHvizRtYC8IEnZAY4Fv6p/aFI1Zcr9BT5RW/bvJ
vSYCq2Ol7pwZJF51lKKsoFgOXxf/+HYUaS9ars1gWyfCIRA3NlnRsE56l4pcEntXuztz96sIBRqO
/PautMkjgWtQTHDcgcEHsH9jwlAqmOjjZ7dO4HNM0vgjjPA6QQxktUiAnnCp7wXiJhc0Kx2Z7ACJ
FC4oMS/KPEydmZSysMhRHzmCl2HQP+ZHbDBvtw6WW3KTel111ptuPWXae85kKFbBm/7PTzVx/Hoj
qIJXwa7tmjcro/cp4e/0nDoJmrF5Bs5nX0TQ7Ryyk336fDB0t5iy2xNjnCYweHMl1/Uj+CRUNmcl
7rNnTk0HmnMPdfvvGaolSODAarysaapXnjZ+QUXabofMVwphxDowACc5lmBa3I+RApE88rFhFWX/
uK2rmTn52yYnWRS+9TDtdKKD5VrMaEQZThuqBM3ffuJw2ooQ8v+yuFEn60iF5mKTSHUDg29eqb9z
KLyLRrDOwGf52v85Lyv1at7b+kKZd4RuHFQpQL5Jn4I9Xtt5TTPyVesQ7YQzQgaSCiLjc/Zq0cW7
taQ/t9J4qKFovGtjoJ72DHzv4vRY8aOmVKc/KZVJPLy22DBaZYSJpGZBuO2Irqn/cbH0vUMMvaNr
OxzQ34P4Ipk+oiSOVzJj7EEfNXyCG6rtlH2/tyOuJNykwI/P6e9XmsFhmb01grVRcs9sGpjYRKeg
BanIN0g9ZuYCKJ6u5aiqUZEwUOMETfM4mjS56mozuIMCJzs75CaVfjd3/X8V5qZiBOxXkBlW1wtG
NKzk8n8pH9GL1L9B2BUT52wq04mtWfaXaW/NUe4yWHnj8BKBj9QpOb/fTvekMQJrLDETsHAUonoS
982BRnOCmAtSkCeCNPGlmzBcfDNPLzLJ5Qa9fV9E8YEWWberoBcJa8aSet3kKXv0EFAfc5vLEais
s4GD+AqjqJKorKsqF11D+Fy/6TuAbKjqjBJGbT/PyNxAfLA4tjrbW0yRhVbQpl2wpmGZqb5jQ+lc
VPN7wfJXEu3clWfkN+O1RaduzONTdpTfH9pOknFjMIHhEboGlokDBzdiGiQ=
`protect end_protected
