`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iV9RScEojiIYavQLdmhYeWlVCnGFhhcYHmKUz5KTBhhW0LvpekokIlUr7cgvImmWPpJiEPECt2sX
qiIhhZUyjg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hAEiizvT6gbTVOuCKPqs8e9iJKr7DE6v1Yswz0NfOd1f78QdTFAquwZhRRVpTKc55oCyF1cmsJgi
484toQVbDo5rsG2FItfuRPaMP5uiWApMZkjGECC93QdNHOiavmGKwehQmIifadpdw8cu8MTU8oVx
rvv6XrKpyyHjLnGIh+k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hEgx8LhPoov+7F2TsULzociaL8fj7xI+oMiG0ZCm5ZmcJYJ4/TNy9JtpgVN2IH9Yl1Q0crglW30w
mQjbBqDAbngJqlTDxTiedOofunRFFeyuz3X6QQ+9+wXP8Pb5m9lVWxgA+GUJWcZA2PXqW4IKUh0x
DJ46hTmthnM3XfDSrxz6txi0pg8x2Kv30ya9ntDIto6+F9M4T160lpoqdlLfKR5XV3XnjxkFBSA/
t7G/vJGIYmH/woQNzlQ4lAJRL0ElxgbDDloK8iot0fmVC3Wojw3cHgmFeiRKKO2Ozq0qQK9leiIL
1lkJoPRthX9WG48VBedqbZvc/VYtQFsWj2J3Yw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cC1wfYe5/aqnYJTZsrfGoSYlzsRhNYd32nBp7LOqgXSUBSxmLg+VrFQhSHLMLXFYjuHzM7Nrp89o
n9HTRIExQuCoxsfblEDOzzeySwZtf/dFHCh17c/0LvZ7GuFRxfpfI2oAF2Dh7h0e9g46egBIabo/
evmlJqQeQ/NWwsqak0Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OaPvfBhqSU+PUXK0gGD7gvz4oJN5TvNleV/oyc9QYEuG7LIEC++cRcPnxfQTbiXDXErneTL3Gr27
SsfvQ2YfbE7Fg2eqPxseRbZM8UW3u/YMxesWIOs41v2XX4dWAuJUg7x+SUqVYmD2jJ4WfpPQjXRI
NczDE2hiJ5JDP8JV/VRe/FT5DLk6GAgZunNse10+LkAb638rVuCQTmwWzvySs33zly6a5vPyDCIv
w5lMEWAJP3MRvl02c25vQzJQwRpt0xNsBqnbIaCMsBSxi1b2vvhw+w8OT2XpJyUjdk+siyVkJVXd
pkxaIy3mtqpzXAJ5ypV2/qxhRLyzAMMRUVDiwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53792)
`protect data_block
rhl49Fj4syyBUBi2k/XhVSgSUnmuZi0Ix3t6qWaAw7c911DCyEiJhGKrM82DjF0TQg6XYK3q8w1/
zz1VGdntSJAU1cpTX408H6T/m7L6O17sAQmP93WCWl2VC+zjrCUpPqCJIBMrjfjCQUWJLd9UyHTB
d3kcT3Wd1g2yrgLPjbhi1vFUu7jx3apGtsDeiKvKQS7VboQIlQYOX5ZrBrOQrpalmIfj+V+DH+Ii
Fik1rfYl3o2XX2Kmax+DQDVpL8fQcCwmtlqy3jPICqiP/tPlkdYT+VReD9gxtEi/aXGLO9/EhUGf
sKGuLBMU+hIHwvTnM5Mf7l8os8kYVykYVrPOEMno5HOHXIbuShJwNgHay5Z7uA/m9JEHERx5v42g
19n9ZC+NTFpBi8LWX8YpryG8g1kh26NvNux8p+Bbgl2w7Nbrdl8bGldMEleir4lw1TUzhDIdWGyn
SNffx1Wz/Y7csWbpSWTlitaF8lckNwjSHXShXd5HqrrbiP+A6dRVgoBuzXGjjooP2JU07njVKkgT
dCa6HgDXsEz6J4Pfy3TSPZ1cbM4mJSSlRlpOPVd6h8CFSb9AkzLY+QhZ76hHB3iGKuZH73tkFSNf
o9uD+ge5urWpfqu/qYMIOwabmWNiAjPIXCs8m4DiFlI8FWcN53PvLvMX250Pf+9//Gsc+XNjIrrs
H5kiq6HtHKJ7N4qZZX2b0NypeWyjl1mlMjks7PvYwwgxV2U8WyeAKoWOFkfRXuMQ2KVRE6qy+ZM7
+kJDeyR2FAwOFHKOr3IbAfg7UcjvIGt/Qfn4HXEswHewFSIT1kTabicGSeLaheTLTb5TCCTxAV2S
QN6TdM8dSt8cyOhBfZHN1KWA/VMM1H3HvJmwIw+h/xdAFZNbp4vlrOg08W3V39bo6OI0xtudLzut
7O3f/Eu5ZCNwXLfycuMllkglPZVJLJHLa1ROXmoWCc/Xv6VXJELpld7vbk5V+oAvNHq1zIYoazEX
lKQDyXSrFxzE/omt7VOllJs/kuFjctErXPJrdnm/5/1gsYZHmPnAbVDcOibE1fcaSIbcgt2t4JBR
fGppKv8cykf7BYcxvD5zipr6Wqct9MsQbPdLP6a9TbJlho1fi0F5UmzmWawY251ofmvpFUSwMmC+
s8qB5ghqYygw3Yma31cicj1xyubMdmUtgpxTHcGq2DVz1njJ24xy2qOrxPCv4jrSImmnn3dpvE20
3rSNeq+Qr7CSwN6OzGzszqEr4gquBB4cW/RZH4ZDKHj8wbDFSiQbVleeeN53PQOFOha631tfyxX6
tcpAz7ZtNqvzJkxw+Sk0i2nUnV5A3kKEWZELpoayRTXH3cMsPSXRIfAaJpu0GdRq3w26uoj/Rd4M
ofFdFYt/6Yi5yOZzTyHVZqqxZYYkTiqVUezG9HrPIp6TYONRRvisOW0HuRz6h1sV2/tJwO/qjqq/
DiQdekcbTsaXdvCGBjoVdL8boKRyYpmLHuz+8zDAYZwtZIDEMLJi9GkoKp5Y0smkNJkYi30W0mE8
iqohiEDKtIad70k2aybjDU8xlrUDy4LszFHcerADD4XVmSa5sccNk/YIolEKWv3ZIfpPvdRxy3rq
dDRUWJhk18RQbXLUO9pnLxaJACHFZuNKJAsI0I6GumcRztbvs2okiMJh1Be9crE4MnJwloOZ7Bj4
Um2Xn+wBPoA7jzE2EpesnDVHwpfDyurYRPPEmt9SCnq7ZTckBqcFTOVc7B2HcVmiAOklTwDwZ8oa
+Ka8CaLWbUJfV+a0Dl6PIri8G3p5Z59Qw0QE5zYZCHdOKgvQRTreKXDjISGDNVcGjqXLAQsUvPkG
9ytlBWngt2qJ0Lk6qvMqKIA6Uf8moN9SerpXavDosNk+2dkQ2bLTIaXjc3ru1qN6LP6bwvO9wd2J
0pb6LrE9YJ7ydOnqiFEk/17ObGXGVsfCWVkW3wBdbepbzTKFS2pqw+lKcBuiIKoP1Yf7b3DaKjVw
6PRh9Hs++gnTm6nk+/ZHZcXbT1SKOLzGxL8SYlxQYj/y79PvyiATe6jlo1JV8bPmBTO9FCa4FFwF
VoXnWAEi96Fh52mNihMF8fw+sFpQErBDDBzQFmeCWOrq7/mRy1zH5I9DTZLZRNMsLvT1KGb0qioT
g3vTBBhp3Oz35uBShrFEoO6kRHJtuAXVGMpGMSLmcFMjOlpo//iv4We/AKVoDkk/4VzpXo20gafA
xoXitZD2U+SfiEO+ZsLEobtRtcxIIQEUMH8Nu6jl3G0tn6iogJNdJmeNYcRBElePuEg5/Kgtcxob
bo5FX+h0P/ZKhH21U7+qn2L5k/fe0hRSd+mTa2HV4ptk4mRqOFSWH3aon245DRU+Da1Mq1JiWdLn
4MndgaZguRRg2IeeDHWsXMqD5kdiXGJtoiSiA+wTduEGv8wJ1tXzr0KSusaMWdyGeTxRVbdkT7aC
Xr8c8WMWeZMhtfGktucm0cI34gbi8AgYEmrBaysZTgfJ40+gRIUMojoyszir4reXAgu85CBtFmq6
DKdJttdtdoWL0pkWAR4j94pVPoPchxFbi6QieyWt0of+tXUY+elTSasSFGw4swqBLZkZggZoUyxN
jVR14MDtTqaJrXChefo0jnVQyVQ7fuDIYkvQCyLgL6VXCe24XTWU+M88ZIUFiQ2SyrheBYhUhuKA
Nt7o6DLCycHOmB9ulM9THnrKsigOl+ntEQOiwIGooppiqdtlfjk2vSEviWj6D9JIW3DQea6VXKX+
V8SMq9YByzN3RfjDwj9epmdgy8nOMum/1qtDcy+ud50Ia9/znz3zJ30ADYqg++peCtuDQCHd0P1P
bSfRAKRojaFeScjkisR4L6CO6D4s1JnUyy7YxAEiqtgw45xgURfRsNVEGHKxoGyMVwTQKgzDtX3q
xQfzOMqqbElcA340T2KJxBLTKcBy8Jw98/1yEOBI3oNPhPZUWgSzh9F7zwwz1Up8XTyTYRjZODhH
hcvPORjVSJJZvOj7VxferDXbVs2hEAbRZGJ9ZwFBorSacpMlOAFk0mdX0ErB4QK6Wu+XNhM0YIpt
lAQVz1fz61gD6VoCMwX6FvEZtaauDGGi4vngR3yCUDtSEtBM8ymveFzDBZwaXdsmfJUSxrOaAZBt
AagZAwHj8/TkaCfZdbxTBTuCjkXLF1oqLKAocMZOGf/ELJ/J7ky50LyPMRCbZecZbz3jfriU/DQ/
3lvTucwPa9PM+3jFVy5BTNNd8ugeglJ9xFEh4cEr2b3HIETSP0Y549oqXtvZDiPZHAzR0XFpm8LQ
iS6gvEEvTLOKruV79ABE/ezK/MyiZz0ab4aHq9ZYbxjoPt4m+tY0lJtAb3madADNkrDiTmbFpNCI
xl1Du2xKCd0s4DSXG2MKrp7ScemNLCUunyGEm/fy7mDPamxgdw+/bijWpRMBO/QJZMORU6vI/T/L
4gbXcaSe5Kprml35DUOvjuRyoKFYTEiI6V/M6R/MpMXVxmfBjjkKEqenSnvFn+AQmjhHBwJkOLmX
9ZHO3D9nsvkrdk1B5AFTx8iuaO9zN4CNIdVVprpHmtkp0nd9RtYuBV2J4BCS7kF04XIFAEn+kA6k
RVXuBNAMTzPZPZ/eM5YBTkI3AuYslKnGuv2tC7/FPhi9Z2s7F8Sh1dK4Hzb/L2ZmZCIalLzoXDKn
klqeANLIly6x6yKYBZQVgT3HkiDakPt7dL5wjSEr4FvYuWa/Nt0dq0dHhe6ZWSVzq6Qs4fHXZPY/
+aebnE8mCabPpIy02EXmakbU8iWM02Sxl157NezGTC339ChQ75W12IosHfCmzlwoPml15FfLL7CW
aGSVEJXbFvNKYeBY55l8dhPApveHTpwAJGgQBLwHVLeUF1j+2QURQ472xwENEUw49pxfMKceqqcL
WejOdVf8wxe5LQZb7vk6yEI0KwkuLnqgX/1m8vVcpZJObcrlVPlYYhYxbFxkD+23QV4frqLuYRoo
5PSswFox0aaZi0sh/jeIBgewCxh1TIlxs99rRFKn5UETbf/2GLoP5X/sShNnbew0kYboRGyGpFYH
eXdQQ6iObVjPQsNkOmienCJedIjQe1CySlubRG2jusm2Cr8UuUKphJpu2mHnp9iTxxIRH0KlpwW+
fB+8mxUBNAtdLFduqQb88df04jgwiAkPvJqyJsYQlT/+M8v1ZRiQ/qXyUCfAf1ZRlZQ4SHTRuTuj
cWtEnK7QCGPG+22oybYoMoVq/ZxbPLn6/TrHWKg2pBFUZqo3YI6pbmbnXQM0Gr0SxBm9kNxHUYHO
U+2SsEe8yWNfwH6hOCI0fO5bWNz1qELeKDEw+YNUzMazUUfDVdpZj7IsXrxOSfHf02l/CCtK20vo
PcdHKuElP5oheyB2YP30ipvx3C7ovHfrk1uQxcUgR3NvJKA3JPa1o7IILSIc83diOpLGXxTnLtbM
QhAAV+I3QgBM7NvvEjBNp7qX0/7TKAywY1zGsYzYadeFpJEcgKl+2b71PMVmtXQFvhVzVASrdZdo
W1CYkkLKARl1Rge8Aw/qvYIxCqUiaqDkcA/dzguG9GxNjJuC8eP93UP620OCjfZRWczB1JwRaHXk
oZjtaUHdGkLk158VPvdm1bZ3iMzFGhMRD8voODmeHRoxsZql2oGXRGRQCqTUMcFYS1LsmdeYixcV
1ODvU3G1W9jNw4Uei7XiZISPDsVGJkf+bRXhlZJCbIi0hUaGb5Y37XoXxDFPf5QdRt2v1cxsLHeu
dMp5yO+HECjCFt1o0mA8LPFrDy4UHxOqUqgGlqh9m7AGoPHQe8nUKybaoGPl3fAcK66/mFqLiKXO
83yDtPs9Vk/FAMl++kGE7eqOlIM6x8c9PT17M/8Yp2iWyaDim5fgD1efXRgvVQ0eTpax8Li9I/XT
2vBDKIMhbP5OKtxaigdziYC4hcqYuNDiy9id2NtZ5fNEWIkOgmUl7n4YqE2U+UQl8q+GSL+MmbVg
vbX+Jut1S8gmOWtGVH8ATjjD847/vOxOuhOGazqSQOLgP6vrlZygGt4BU5ACKZibmSVt4wss1HLn
4p1PT2VOZvW7/anNO2rVm5oKdiGM+WEksSq63cJUhT18cJ5CQu39iWLgCf701sbvh4U3S83fGFMv
QDJFXHnpCfyK0i8LJLbfZeKvza+MhBVfwlqqTrGBOSLgAyXFwlby1P4HxgmV0UnccghAjKVWdOtT
XPsnXU27Rx2VOukNfFBS6aa9ioAB2U/8nSde5jfOPkSVLSu5YvponaCy1KS9X49w4bU7L0n7RHfA
npXVJT8gQ7bPQUlFNTmQ4ZjHqmwNNbzOM7saJsrolDp32wppQiaZmGlVLT/69MRscN/ghc5Wrrzr
TIuKGiXsxkan6lQnTKgvrbmrdulXKESawxnsq4TAmNOiZXlgIkEv8q8JUdbSGyE2E/6JY8Pm8iQx
jBKVL+Wc5IPlYvvnPSf01CR8dGRATHp3XcHtNmpo8VUombqd5Sioi+NSUAT2okcdNGgV1wYhlpQZ
BC6vIT8T7QB4/VtG8Li1V6OFwu2xbKygBB/4hZl3ntAA3x3lEjXIkbFt+4yvF/6izn2ZxfC7IF/k
YePJwnJSF63oFojdb/8O3QS2TXJv0ONCWDi2mNg9vFhpR+AvpKavgqHeBRi4M172YIrq86lUl+kZ
34Rl0oeDOd5tUzc5o4SX7gaFyJ4y7XizddzuWShpIwItljEMaRwGsxQn3ybYlWlXN5FtRyraZ7Sb
RHsk5lFMx8oWWi1MNz488HRODCsT7J9HRwGkGmZsRS6lDTND+A9AyZOPu/AY0N7khy7de40yFmIW
Vchybh2CGIUY25P3G7jfL2s4VdcOHkha3KEYJZx7x234nv1H0UHyovc3gHUGA8gOqUD/nPuLHuU1
N5yJRVkBfhwRMtounhEteZWib8Pqcxnl2mfZ+XKJPB9+1XdnQj1vtMwwYz7L+F08I7hcT2Z1TnfF
p3/kP0YYLeINsiJPVTG4T51Vs9XwNNNf13Pdh1ieQ0tSAyVipudliRt/oz7ti5ShLU6TU3clb622
uJkRkDw7fCoix/VMeRk9nbLnjsoNC/I4vpqBD+lPhkWab/unTmn5bxZG0UOgMJYvfUfBe2cJMJIn
OcrR0SliXrC2JEyEW2r9YGEHht+JgJ/LLbgbhL/vTNXHwZFbFqy1UgJ+iK3vVP7hpiM+9BbdwBwk
4dPkkKBF7rWtPMrZAcPaQQNdIuVRajVrotDrElA9DKTkWTDEFXzz3lgGz+jtQrgxIjRVg6hjodl9
Cu2yYlboBd3iIgdp/P9yfvoV45c3pmESD6GNb3lK+vO6bipMWwbJ1WsmCHV6LnzezMdPPKAvJ/3B
SuTvAMnA0X378YZzeqdCOMPgpKq+MJmYP2aGHCdKxnAvsyr1sj3jhaXo7wB8Q+go0XCut5OzhrNE
2SRWWZSAW/g4dIabNl0dGIGiFDmoTT0tu8zy5AmEZlepb0sqq4mxEgVimY5X4JRkaYaKQD3MDXxD
//QE/1azo63gf5wxqVIW3B/FtIwnz8aqXzhEJf5sJMNFGCl2D/FkJMIfnMlWG6rX2hEfDc/RGMAM
HEi9tasNsS7/+OIFNRFU2mm89JJcBTRFM/E1LcNrYdQEaWN09qYe7TgMbWHvo7800kdMNxpslnLR
VkfXgbdgP0WAwDUFoGmoMBrEQHhiRFIddmrcDfdWXEy1FOxnv2QPbIzghh8yhvFHJjZ/Y+Zw+sYr
DY/ydPp3wzk0LWppax+GXmsDmPkffQZ7B8qIsxFli2DsS7WYdzOMo88AG1lx8/yUHxZMEz4QkFdI
d7T5VilZ6fjpK1h2/D0a+vXs17RAGZUkjRlFX+2s/Ads0V9TZz5XU4OlpmwwzC+F9HilbuBmWzp7
jhpxGnU/UyC93o35mBFavP6snoTgMo8ryN9KMQF1EMCAM/rbUardoIrqlqqiiLUyroMdKAfbynvO
9jpQiKOhipD/OHJviTvzTy7K3v6+l9n44s0kdR3Y88Rm/lNdsC11rfknysPbkLQGkpsaV6VSu8hW
6fnuSbNpWrCh1cZcXAaHt8+5j1UrAc9dpJ/2ZInTHPFQf57FJpOhwNzdOeiIlt7Ro3nrxlW82Imn
p2biammdDhaS8tc4rliQYsEkMbPWvOW92o0NxObEKH2rxV9zuuraYjhGJ2d5Ru4Q4LLValoaVaar
fvl/HVHxjEP/81XTnYdZrLrTUB5Di6X6wMbZm3Ss3j9TP8XHAKwmE6HgOYUF2wSXNIAWLUgEzYTQ
7MeNYbx/Jrsn3oV+NklTcdRRISsDfl9KxckAdd/D46fM68nJ3d29av2c69dkjKZJamsbTqty/QPk
ado+9W+VBcKDTmAVzkyobQzNHZ//c+ufpGkzDeTLSfumdnd24/BQckzBeOCsAlYayGB7uny28Sl+
j2z4KZyoqL6KkdJVPcbh4eJSux1BZoromTIKNwVKPOjy4Z9qAAWJF7W5XcRnmuFfd1tdIVjMDA2o
lpPDZ4ArHOH3KHEUFlzBU5/T36QHnzfryv9mR62sGCxeIaZRPwsn65UA+roP6azeo7FTNWz+Jpnf
qQlmKrE+k7HYkIxEeB5CEduJeOAjm6U88k+KFIemj74lwMCj0gLJ2ImM0BSRabkJXNoIVDt28Uew
5D1pzCwZgVSpcFL0Ypko5WozjV6yypk91sa6lmXRZ7nepWCg+dDthI3+ng4i9V9JD8MKKDbNLdbK
dvK5jJFlEKl9/lJdBxJX46nR/SunzDG/LrWbGB59Uf6U4bFSO/ROXXwMVDSYeHDQFBRw1bwdDi1s
Ixl3UOvpgMPFzy20WwQSY88loErACsRLS3AFcDbtBQBZsdxp+kdYGwD3RjT1+16trLDDtVyEHk+Q
dLI+/gSu++zeprVHGoskC1zGFlXnF077ncKmD+b+4dGZA40U/O3hmWVEWKdISaPvbGtqfqv8YsVf
zIXEVIvrKZzUw93mABaonYIIgZvZz7AQpdRkaFdXH9hSNA1EnBgrKZdfZK881AsCCfRc/kw5Y+1E
ROeTGt6SrmmQbCvf2FQVerMvr8mxgUS2e1AmG1aB3pIFqbQyocpYL0aHuBcSItXotwfE7SCPwOFf
mKTiqkOOpH1DRm52uAEUHukISDr9j7O9RPQ2Nl8AITcu2wiMs7jwbWOoCUpAuA4OGsK2agftEPOq
6xejrDiwJeH55B3ubCmOaMTIOnR28DWqQN1jF6aUGnNIMd0tj7671htzjoHvPbETu3GqvHWcO5VL
IJWBAOrXZX+O79tPoEwheWsxmw/LfJG0VWH2aud1QofLqqsvMHxY6yLqe3VdS+MTHxCyA412nawo
lYs58fffVvIIRuBQJqCINIfaH4itkfyXFdQE6lfQd0qPchX473jencMtkJqMP+LiTgVy+FJIaoAU
HhuGksYE4ngwRfaFBLS5Wpr8THWFNptMJW9ojKm1LFsbCKB5idlYhe8WxvSYFMQpyb7RjBiU+Z0n
ki5np1sjjmx3wHxANPb5eB/9Cr057TF0Khppy3he5arg2VCAdS/tLOIj2+41vNeQ1Infzx8JqmIq
zNs0F6HlOLHi8Zz9eO3ov7vaqHbCtFKT80ZlHC4olA7NtCwlH7hrQqv1QKg6MXV1K9INo7ei2Qcp
9IH3HqGysE+S+texj3VxAulaboTk6wXMLbPuR8EZhUcXtVmqdqkWp39brGENR2CilD46RmvqFdVF
o4oy+iDONoh+0xIQHz4yWK0mPi0j6Sem3dduP0QtePfDgxHSb7TDPESn2kO5hMeNQ5l8TM8PfqgE
SqUzWgWllzB2wYF9jRy68kL3Hen7pXqodBapsw2TP512sT2WZpvpFWd02tWGvP6DYc1EfGqZsLUn
cxsF9v+Z8ComsbEldm3wukN/oyXaepUQZXaibhimDrLq1MIpQDzJOWgrS5Ycotu/dFyJriThyBeU
EwdevdRtgfWztSj4d/Ts6GTTecHnPSO1SdbI1sKshnCuvyhltQrBq1cn6/Pi0dUDXK4f9m1Vkb6J
k3D+x+n11h6IsaWvONxtXfSMH9D3Vik2/Ct0DHmGOJTKcOK9uXI3FxZHHXdPPBBZuuyjupxoUbHx
hXpfYHJbmpFl0laR4eHFpQz2xDqPf3g8qUAbZvMgjGzTaUgiIdAojk7ydwQ2L3+SU6GCG/70hEvr
XEcd/AWurEEbgrKJtP8dUSaboL2novVeWKimWs0M8gq7v0NTYYDwP+GPAlJvavTpM6qQdcpd8k1B
f9t8tVlM/y9kjMl6KBHaJWaTtljKu7XxkJbNkZGyE0VjhVLgEG8toopuJxCFsEdWhLScDqoz4WeP
ytnTCG4OmuG3jezDHgo6UM7J89q//7vELV9fvUD8p7nZ8AtyanXeSI1fenhOOjfHzkz2GjWHdsMH
q2aR8PqRtxlTTzQCoII58JgTXXBq1ej+6d5KZ95IyQ/06lEXYtkqwMjs05818cTwRo87qdnJpbWT
0NHOQ3RyiHAApYl3wP8cs/jO38yCUcS29nvX1jsj9a3UcJJSjMwwrYoEqTY2j2RI70sN/juBbsLj
5+G9SFO2OaVO/5Ro09QfqO9/eATL7zSq/T/AIctc3ClNKic24rcsjDTVL740KKuQilo2YfDi9j+9
tZpvbSU3qAeyV/kdQnvd6aWyasNync9Xmu/C0OwSyVYJMYSZu31y10AU4fmnUxOMQD0fBuaA55cK
TPT4urKIJUiyd+FiweSDpaX26tp1plqnQmzcLSypUvGB8ROVKFgdDO8lXd5Rm5hhjyeNhzWF8RhP
a2Iw1gJWiWnB94KAKNWRKB5r8nAo/eRL5GHA82k8hoCLQH9gO6fU0FLV6oYrKkqfuQOitZN+7x6R
joww0lonq7VH7S/kzTu0u7tfAu9Y6+eZaNfLpaqNBEtJhHVa86UTUeU/R2URiHn4Bx1WrePrnJ15
NmycpNcMkRv7tu6WkxPaoY6WmMk4jcjvFEQq3dJF81dM77+yA5zL/DBrW7WO8dhiJSbLfNjDK2Kh
a6QnuYpejxd9eKbN4+aoMocg3of/jeRnfmX1wWjASguLUbOvwHS7JToXOqaddrL24g7F2hLEUMFW
o3eTAyteXhy+ljt3YJLrEBaIZrMPET0Jgo7deUBO7GZZkTwXnXhLwbBz5R1kvq49punnhnepcCnh
r6vktRkqIdtXnuWVWd0eVs3W1qs3xNvKBrnEGXnsFjznlczMMlIJgf/KDQdH/b7CpJ/5GH0JL/5T
cmsGjFe8WibLi7fjD9m5Lap15BOZZmRYgbRPItEo6LaQ8mTqyErAzU4IWynLVlaT6rMkozRTe2is
6Jpi7lrkzgJosqQeiS0lFRYuYurV82+9XRJnBPV23V/+SVvukPmfYKh65L/JyiP5zwLr9/tzLdGF
RR4OOsN5yuU4ca9poaR+0YGDauoJ+wRH/0tV/FPTLWkEnm3ueknMhEMS5U7CFcJpFfCWo5RYfxnp
OOS5JO2nbLhWwZxpMsbXqvr45EVQ9l7wKVL/Xlp6Scpq8FNZJ+Y5X/qVFIQRAvMkQsQpJ9971c0h
H7QPxx1MzZhSKetu8OTk6u7vO28CEuku6lW9VUSLDEDQTRFzYhEPcdbapQoSdAdoTq5K8GLimcCZ
7bw5Hv3rpSOgjzSdWiolYkW0mISovFJ7UyvJgE44XJjYS7oOITyZlz/zrkXHodCAtSDnYFz4pRN+
auqS/9JFptDiZ4rlVgEPEc8mPfCCOMKx5PdyJZjc9QdiIE1IgcxtH4pQJW6LwIJzwBS/34dVqgWw
nlBc5NGapk5Dg+fL+lZwdDAWPLt/inRraTsBDH7UTJVcT3LXLbbU4OL0/7yxNFnzAcw+YtcCoFsd
jZPH9YJoD02T8XYQ7Uc2djiAjd1Kl6TaBCoycA77TRMb4oWYEGL9ygFCJoMGcbF3ykRYTrk9+EYR
pty618eGgFOP5fpsPBt54LFiO4oaHEeL3xGdCKFAPBJjzi35P5LF3T/mevdCq1Ag+mC90hjMbjc9
XhLUXKwcTaZRs78BBp2HiGID8i+0Y7jchLcb9TO/iTWwMbWXuowUix2HBoBmJwFPg9Fp462WtIS/
APEykUkeHn3N1dgbM87Qsd6a/D/ROQmVqR4VeNBmSrR99WctVCSq5rOcsPT8eip6/5orCwb6PW4i
Y9lgbCcHQml/a86BAaCHEGFIl7m9UDg1wSbLsMVMDU5dc/UGyAcj11WCVRMRfWHm3EmpvjpJFxcZ
OEf6ZptbjhfMfj4adyhp+NSZPi+fP73GWbOiGvffhlVYE/UHrWJVFjryxN712zAVVdGvPmC4q530
XXqHtJPkXLB5IkgfmP3Xr8rda2hb3Mx3IpSVNHKiBhJF1JgyRE30Sk0K0bLYplQBgi6w09itvrx0
k3erA8VvCWxYzv8kmSN6aoYnD+NTYoemlz5WbNkjL9ysW5GOtyuXACVt167/k80e7QpHnZZSjwQo
6VZgt6lM2XxuKx3gnSg+XVOrEw5jSddUAtZNAIQiZ7ocptwvI7XuZNo4U0LnOM+cJHndWxVS/0GO
YSdwd/xHu2YCmSccaKYLm9pic9CzZ3nvD6LWAKkf0iROb2SJ7FbOhG/WSmv6MoaODci7EVXJ4f1a
qqbEIJITDW4B38YzLNUL7ua9qpIndSYVnQbbKWEcP058deZzuLFx81Tck2pPvyw36vve/0JA0u8U
7a1mXCe1Qy80anBsYZqcnMuFhoAoMgLJ2Ot6ZyMWJrZSRY4MksXtxXofGjVKCNJXSLYCOQ6njCdi
fSSSjkvRYZ+3j1P+YPFYYsN/t49LmjKh/H5LeIhKXBVZKcQy+meb7X+LMAbgfxr+Ee73zUS/heMK
Zro8Srm5NoOGWeS3sY4zBjGTFSrlQlEMk5CQ/7mppEQfuWwvdoXgtPcZDOCYcPda4BATO64jrLJC
UwUxuS1pXCQ8URtyYZh9DN/ha2pcaimR65DsFiBBWW8sZqfbKzLRZbnyPPWGfIw9kAr/47Wv1vxx
UJ2Q2F25FP5kE9U7+rhruLjpLzyfs0Pvn9aY29LYAg178kig5lFAmKzeyST/mRkyCsgHMPfae4Iw
IxXc2CpW67YRXJu73RDaMyFngf5gVvFfHsHAbnwS9o+fF9nsb899RV+1cgbArNV3X5un8RSUw3aU
i8LAsdRZurKKc4QTzd/alT3NHa08DrHIaYFgxCgNQKTwnEmHmF+sxVjFgumThUpwkM0o7s9W2xJE
oqDfiZFHEbZbANF1+MzlhsIrZKA72P3bUuI+BCkYhxkwZ/opWGRK4ivXGg5D6orvZ25kjbv5aGhi
W6hljx5I+PIZ6a0aYtJlgzPyqDSMl9WCxKrn6AB74hBwEkV1b1AicYNx7ntmtyYhnSWb3x54sH50
pqPUuUNQNR4W5BQGiX+zZJuY09dQH9tWBUnQoRg5NGqi8AysO3cucEG/2KZLjZC4SXfjjjc7AheS
U1Ha02/AEBP8SfQUYQmVJn3ek3mI8h8Dyk00qnfB2nhXbOFqF8LJH0OWHcDkkeFbjyQHyeIcF0Km
dwN5Qcpl75H14pMv+NwWNmZVcO+Q913xtOtd2T6CC6IeVYTexeT0fOLQ9PeDuzRq+AwSP5PRB37b
I37f/0K0vneddSQhz77gJTPtgUh+35gKD/Hrx16QDZQXC3zBbHLhSQFBF3noZ+8zrXjQL8ZeZeeX
7spBuvxkkP8wTwNlS0MAwhT/4KWAdmWIkfA62a1LdjXO/J9e8m0+lOXzd+ttweiEr4KcZtV1mb/s
EaiNgmFYyjejx6to+5B6y6LhxhOpXzLD1gM6Ybn0Ux6pRPVKR/nJEELKwfr50rpr1PgF6mxvAqSM
X5VvwjF8IprnUOwUwbLMdgXP/YwcHnFwcVbVEnsvwiYgg+yqGu4DLNzYCJfAVFNNbJFYTK4SiZ9l
YC6XQFlJ0vW1Sl8ZFOI5nUhfIGQVvtDr4dPivcGu2Udvz3SZ8uwdi+9+jx7egsjGj9Wl3aP96rnO
WwFFN0dqvqcWyFMkBK6NTzkJK1ko1SSiwlG8C0CHMh3TyJUnczpLgq0B9WesIxvGKTq3TjWWA1Q9
rzVjOZOOX3mzBNvd8F/HeJ70AoMIGFBUiL3+zckB8tM780vK7sYlbFv7D8ONnY4kJuxU3qxEvCjv
TSZHC2O6L2ELMqrJ408rF9ElmdqLzxEyCUDQmm8PYVbIrJf2G8N7sbf9JaKZ7Kr6LDwZ0H++YyrW
XnA+sl2O7Lb6XVGRwPw7vHFeABUtwEGo9WnWd4Sxd8QB5pcNJXKeNba2DYup8M8zAe0/C7EvMObr
NIAFmYOea3VSMJMG/jdlOIDYx317gQ1DxnXECCzuwIJ/qwF+XC/D5C9WkIv3ywo3Ok7vY3WEytqP
j5QSjRXi8ewY+xtig9XYTkhljekVD47Bz1tGqMhJy/ZK6sMg64O+gKP3HxJHrFh2oIp3ehvzyO7H
6rn945N7NZhLPlfa126pcOOjyYo7b4Nnj92RCO3O4P+UWxCNQuRk1c6naBOvvUIG9cGlYVu5J7Bs
2mkiv4LKH+aWHLvjOB54dMMuCjT7xHWrK/r0vWQIYQeWPjgJXFFLTYEBKcZPBKalcb7OYAza2eF+
QVqRyba37Jze4FcR18VlqXDZ4HKD8b2+bBIitxh6eRVWFhNDPNo0JS0ptRicyoSbQlsyTwLoujw3
R/FdcIZXAorjDnf2qxpcRKwr3hr3IGK9s2oL1IOpXxm2E8XGfWRVVq61Ey76uZWqZiOIyJLHeb8s
M7xg0nnGNummWlpZZf0GSuMcF0uG4/eRAu3IBII0uYKkaqLnsaIEycxF5vPxFhPuNXRVUhI0V6Yz
6N0tC0qf5TKpBkY5opVG8Fa2JX8kwThd2srFqljffpiDmxxQgR9K1/Bk0aOCzGbdnyuInUPVLb8Q
2lVynnuwIddLBz14/QWvtnjVJN1pkAJsVQlkFwmGIuqkv7NWYXOnx7UhZRwSBtVQtdzyd0wdhW2J
X4H71VAHXbLrbABSdYGixeJlvJ2jVR6gfSUsoMB1c9tIHaKhe1hEuDX6gSABIJ/9o4sw0/7iU2+R
Y9VMIHfIIA+gFJxorFPNQOsgrpkdlkD3Zara+wzAYOdu5D9Ggd2xciXChkbckqd19MHf3mZ7w/v9
lxw6oO2gqGhnjeRmeT84vN3UhPK2e/arrtrkkaCVAr9RK5eB6H3Chk4HeVeUtpIV/sCne/NB54pO
iT/WYuB4XKHw2BHLpdKaPbMG675aLKBfmOg3gsotUHJj9LkzoB9BaXtSu9ybHCF1JFlQqCQIRpdV
WA4IYQsC4EKU0fKMcQ125cLgXQ4V4J8tvaE6xU15vksLE3kpMHpsGoZacl4/WN/FrhQWLcb9fFA2
1gP3HI/ahLvj89f6ipCWrC29eEljBltztHJWzjBVDPNjVO4FzGGu2RnUj5OUo8EX3o6Kj4KOnknc
IkNAm+IEd68IYh7FGhd423Fx/VjWZ2ve0P+NAFxb1ZXiwwPtEEI9zOR2w+DLiZ0fGAAClewrQqW4
lBBW5xYE67j7Ckj5Ksspm3N9bgpSYJb1vlGbX7BJaJiTFKUoSNx0MV5UOANkVSYdSBhMTMAxwToc
CkzEfs7fuNX2hcaPrZo1dMtcZpBWEJZwJI5YKeuh+73kHVJRkk//EFX8n19c4Cw87Cwx+H2ji+aP
3lfLBkHgH61Zca5YKxkFSPT7QtACOcF5wggTuaPv1tZEp5Lc3piWA+q0MPqrmVTlfpm9bC6cnyfS
3asM1OEupvWKiy8sPlU9pTCr8f4kzyrHmiCTQaLZuQhq35nf7w/2rBvK2Xj/m2G3wFr0V6lcgI7v
EeSBBWO5nKys9j9GFWYfWR9ifbjQGz8MfwLQeygTHdfYNidDuJNNO++bq/CSPmPqTzO6eKSLetcf
TRFnXEDrk2TvwHnIo6k2HiRBqo7eOGV3/4s9Q2KMy5/50a6o9xxjgqShjjg8pA5I6CE5GDPNv+fU
b3u0u2BACqjSS5IvIxvQOSCz6PZJpplBo31axaVAuiwv0Kuw68w2UCndlFgSR4oeMrLyrhkBaM4d
yulX9CYOoeIKax/lAEawQ+c4e5uIR5m7/9EYPFF7WSO4fWrP0aPhOhmOXTXkqbw1vJQa1bOPG8lT
jsXWFIfWxvXPlNdLe1QcL49T0UtxJKtBQPnmnXhtCtr55/P1QLdTGr519kxjR74jJ4AmznfizfNV
HYnnGSVVin9d7KpF3O6p5nSNd+iqWgEI+RYuc3iz+k6MiU8oUhDY6atdcLGO3sddJdLWWVjXEed0
xAmJ9VEfK+PdhZLxkBsL7LYpGUEvvTnYLjSsUrRUFWcW3SpICJ4MFhkB7LYyWkOUMjNuU73qsFVv
pFTLaSdLcMxxbJ6f/vu8Jjh2Lo3XZkMVSONukWe5c4rfzgenyToR6JqL9QJdXH0XhpC6JdwcyOKh
/3o+EcZ2uajIqCoJ3XwOTPvHf4Hovk+dhCO4Ex8QiLcXT6TdyMEl7QJYgQFhSEOW0b71VqU1rpa7
8KV/99+bUxdOnQSfsAkIfisWedFmRGgU98gpVQvk5t6Kq4ihYhIv1eNiSsF3EgCZzkKUQ5wj8WY9
vv3TcS/b3Ama8ku/6bopnSd5Alfrku8Wreoq7Y51Z5p2SGkExjHLugdA4HgznFnOSbYlar63fX/n
uda7GrV4RZmSL2Szz6Sen15FC9wt9n0qWhJaoXLgUAOzHoA+MN7nd3AQ6RnHBSbHQ9fQB3+iOVkF
yiRlBCzNPzPwEitJ0X8DdJS4epwS0r93GkjtH6uHLNiSms0ZQCiWcwc3EURfr79ZKzDF5nwC3WD3
uMOYmttNHry7Ea1GWhKCubeDRhrjXsVOn/1kqVkVsQcfso0S7aMeVvR+Dyv2Umnjilnp5CBRJ7MB
MWVPUN4XrOx2gO4RYu8aRR8a/MxfXXywIERa3dhDcWFVRWr4GkGJv1WDIUF38MFiDTzUsaNp9Ax7
d1EZiIa6YwjHsij3gwYs06B9QnNS9C65b7d5dfCMGwzTRLCtTwsVAc4aDTm0mUmSP4w2Wyei53wv
B9iCovgDH90t1APEvcO+jjRs3N7W/GvYz5E04+0+6JGZRQfwXCyCKu6FuYAwKp3d09vLyiwR16+G
gC5HpLmIUyMxsqtcwtOqphIY6b38dczjpLksIt4QMH4Hz2aQuFP1fAsTcRhKRd1NwPEMRCQrgJT+
grzt+F+MkoUEgA+Xeaaln6Tm1SsTjEVR8wanLmfCj5yA9bPAunjax049jJ6lkYDXI8JTE2YyQ8UV
RPQYtH2CofagQgtLBZBgKs3Q6RlkvH8ARxxylAtayugPB4NY1HMKeF/66H41EnMy05LUALKiRPCx
rrElM7eOHFzDE+lPRY266KuC/2MVANHGyiMutx9Y/ThdsLb37eTqgCKr7I3kzcpJS64hZ1Cc+OUS
uzK4cMA3lPU0w/9b3JxiepJMsRiDolTOqy0f27plzF2UdIyx8FRO4ASk6ltVOxIASGNkm/PgD1KU
HBEhCr+OwsPMvHanAzhwVQqC8VdwJW26YeRmyEqirrfm5cfJ4ZtRSTc9MVLGpfpCESc0eHRPXjh7
Hdzxk7/XRLDIKV24vtfpDjM8WE/UYrhNP2C8ZE4vgUGbSQEB6W8EsIHtFgeeTtqqzSH1vJKbgQ+B
jFZFAwYMxKsKhexyjtZL4k5EN2cmH2FBSWJ7v0KIUSMh7I0MJKsDXgUOMZUeHdPOA7eQR81n9jlX
P8E5k/2mBRt45UTmX86O8JeUPzxz8lRjodGaceIEoDu5WiqUySCMUDwoOi/MJttM3aH5zdjnVoS2
XPTLNj/40OivlRlYWlpE7KbXsyU0VE3qqDORvj4oLUcPwSUyacqvtEdsmwDRa7lU9BQjrU1/WFY+
OKz+qgr4sLqIsl+2JRN/p+dmsddqWd2oL48AEvd8uFHH3VS9v9q65c2igU7pnz7O8vLE6839a9GV
GItvS7EM9xqnGXU3jl+z395l3vLP2QglAqKftQg8YaDKksdg6LkxwpYBk5SFY85EbspLhmIOhu2V
8f7pKtwPhLYZCcfNCZ4+Yj+B0gVmkUXxHn08+jt5CFYA4zstRjhUYPrxkyLAukPRQ/RACf6otU0l
uDJPEDcDp2XorhahFeBV/Psi+k6Z8mk7K1zzL8IyAxT25xgXkdZRNnZUjyM4ahdSVzRT8e5nuK9l
/COKBwym3nTacH6xj3wE66RIEn0A1hT+v0PJ8sMtrHNUmQouydIqVKIp77iFYkls261YK6erfkx8
zhwP7dUvzBCwWC4cCRzPiKidfiJNM3szbhkHN59gc3fJ/CXH+S7sTvJ+4s5IJhf19d4MSBJPnUiC
GOPXlwvnEo9PDOYRfde+1kjFIULaca9AuNcLjbX3WOcljVhr+W3yQLnv9G8yUa5A+eMxnp6+9qb3
F28FGgqEBOQLRfPLJaRKB4k5zA3UOcj9f1wLeTZ0kQ/He1880LEPD4Us8dLRHaqcdLau4dZbCsEw
zCDzM7CY7AUmrNO+v1ZnYrg8si3gO+K+i+DatvArIUelF827BL13H/BTb5OYygxMhhp0Phugo6kC
Hj0it57RJo7ZuAuKtIEsDy+dLfPI22MrXVxc6r0qykSBiIZQCpEk3aNjki+befBAXFJLl808DDjb
x7SCbPhh+Mg4Lpr6c7EQO59tFTirmXTG1UHcdVEtD8i8DPNv6cbkDvp1Ws7e8i0zcExcjr+ZatDP
ESZ4ALBpvrAqdGDmtOkuY98PTffq/nz9s7vfkizI8DhzErsJRA0pXRyBnrUKM0oh+c5LxEELpgnI
P+umdfVDyetJnI1lLB5zx/bLJAqzqUKnq3TzkqZIaNr57zBhVHnkZt57zSVgidH+BDYKizMZ8ja3
YSIm4pQW3EZffYZL8XwUXIdg5VsPkn3RTcwE89XZjTumuMuJr3oVEEHMd4QO8NLf51dIfn7f8Xrx
ci3E6rfRbgmqHxFUPUzCw2KQMMVHBQRonvgTul8EhQbsUm9DAkDzVxHXQEhHu/5NjOEMcJduHX3U
hVQ4ibTmCtf/DvabO740BlRYzAubmPPXEGmz4w9dwtHAYu1uiiGqExl2/+ortkpTaWc5SaDWVzYl
jZS0fYd2VFH7Vqq1feTVWFh6+3e5CkDyAlvrfdzgOuOISYRpmsTsbhRVEbAoCoDDku83NUWChnYI
H1s5egPlKCaAetv9t1w8auE6y5fWqMaIoueHhIJj2k5FbD1kI/iq9VqoC3/U5gsUOVdjrR2XGs6F
GXJJ1Pz6+hVJIMXng93igiqBfgOvRWOWi1VbUwMk+AlUzLlXYSeTM4yiOxGdwuoD9qsjM5EsNGbH
1r8F9vmyM1FbEb/QtiRVnyd2TlD9Hg8l9hPjmXsjSZH/cy1atiUMlqRGC58O78zUHjxJs0kVAyVy
+9De2+9L6zWno/UykJ1kzhK3aMYzh70Fa2O67a8tEDgJoYe038b3kf0lIX/KAkI4g79ZIChhe/e2
PkjMQEzn8qjD//rAjoahsUzD9f5YuKrUYkj3K9zOBwPNAE8PRkEEBQXqUeC0aEfpK4C0Bmy+vn5x
dZrAJQf3tD9u+7QvSvRvmqPT3jPjR6Y9n8gU6v7zDDpnZKP5NkIc2jNeo+JjN1MChpVOcOGFK5If
aV5E0UchIE/ocncwJXcpZ825d8d6e4R2Fal8vy5JnjO5AUEqMFSURDeUtrD3cOZl466U1aVx0IM0
RPMRQ4N7rNv128IFiG1bmMTJkcr90mwpkQ3uffTKCjOxje/XHPTzZmivJhVoYbbSFc47fol4vNaD
gEEbILAu/mKwns9tAW9SoyOP9cGcga45xwJgKIIGMHkzhTmRjoF4RnwwmfjjZS7WeP12DMnz4QpQ
tNzxcCbNoi397gTzBp9riDPBolyqQQncMmYTPmhIFbYk0cGqpZeDod5D4gjDuEVXaut8ypWkkiSu
4mspYHuldCRnf/ZeWsgDMxiyaDchnLuVxnkNeW9xGr3quwz95G77T3YYNbMGbmWdQknVn732118Q
8CbbKdc6yeUmCj+dNeTZLT0gIZBju1Y2Njpk+xbwwO/ZFwg4WwmO+UPKxkfP7iYYGRTaSPtNzwL/
wvYAtUpoh8wM3btQCSKsWiW3EQnG5k0We4t4jpTnykLGX6xDoyqsblOWp7fhB/8Oc8bArgRRyfuL
OgIslhoysVuJ9NeR53eh8K4cL5ewk62nFMDAqI5YJVu7G5lP05WB6rWzQhEsCOYLUahHtk7w8wZ9
5EV8o7EJ3lwlU5nmmfmcnq9+bAQRq62xxaH/7z3Nxn9sgzw7tpWxPAoFbRq7NQ3SvYN+dFzSQ1Ph
TtE56WC/jjCuKO8eM7kaDgtDp0DAJa8dhLyXM75Kt+kYOtdmizKIwCUach0ikKhuR6roP0RU80WE
i9RL6sEymjfS6TTLbkBP61Mx+LNXBhVdcxX2FD6+h4GUDiOGs3jgwd3flrAwIM1f1EYByCKOQRwo
M0mtcCd4XIHfgaPbhwrZZ5nNAuKlhZhgniv1oFVhkboR52xhhp0t5m0ndyfxDhOO80KKesQ+y/wF
G//8n3DNBZdxUa06eXq+7/0WTitgVGUfr9hqNxQxxSmWTXNyUnd5Yochw936N76S9zj+/9ITnYa1
oDtC0YJb1NSQqbL/R08XjbNkLn1pMeq2/J5qTwtmI/UufY1BLaSKbrVWmprC4Xk/j5SI8X5Qa2Au
WcpdTPAr6RdH2ptAEqmZW8uek9RACCek1uq3HaP4ruJtbLY5FU8nAiJxP3ZCD3PCCHFQ1QZ+KOv4
YqBwTu/Leuoc4TPUi7DF5/mQ9pKsuTjmx79irB7c92JRPe9miYkzW8xxDEuGD/7R0qXRIFXYIiJ+
OlaYLbrtmu50fO1oUbujG4rleT9L34QGYQYu867LFMMYZ/LZgOxKTMtfDFwb2PqOs1q9IGtXTG8t
sGGHXow1xN9UGOmI8IEGLX9TtZA0fwJfKjU/bYXlmosiRoVtHxHQUcc6+j1HSB7wXF/4sDAZIc4W
6cdVFCNlROiVl8m7UfadpdzeFoNuIu1zsAVNU9+qVIDt1RhHc5jlmASklQ8OTn6DlFGwUBaN46k8
W6jyp68P115EAlEHboXTFx0mUZBy1PWI9FU0MHKx0z6pJwZJtxxYpjtv+UTgdSydM4q/3WJT+1s/
Ct5ydt1n++F0kvB0/bItP4uvm8zzsaFkRPJkGTiSb8J+ESpHP0wzYJsR9i07Acq3M2mNo4s/mHz1
ArB6JgnTXmxFbQR72Ckk34BLED9Y0D9ESlZbsWSuIW29WyvzZ8s67tPBnrMVzjVihLLPG7QoIGO0
fmCYsXP1n1juRhbooDEL4Vh1Xgw9mVsXI+sNs7kEyId7JdbyNwcmtxm4m3XpnxUn1wu1TOFjpKf4
YW8PaLPJ3GOnXVhGlPnd72TYogyB5m9xQSJVpQSOQTuDy3S18jmLZ3yarDH2RyWGlxkmkHv/FYAo
b5KtFfmCh2eY3Sq05CpkRa938gP25Ydg9H8HRPPRtZ5rlCmPPSf1maBGabLrRMz9a4XU/unjlNMQ
F59BgT1SqG568+7YTeLux3vfi82YD30Puiwfy7HUIhOg1Kur+4LnPEDeVBWkeS6aOmMYSyB3afrS
pgBdwIeSYO9Z+s00xD3dSvVtMdjNshKp5JX4xoMoP+IA4cLzcb4B6i0sGLPCKLL27dvhCAmOc8jJ
SAlui/pa59NynquzKLaUUBQatgGOGyHvK248/TOCd7V+t2Nw/ySYLrfEtiTAUWzDN0w9GNv4C+kR
gkoF/bF8TGK10XHdvhr9dS+w8Xg30y8HQiTZ+3/xy33DqSRa3ZUs4lLnYIp7kllAWYgwhNh3W7Si
t+JaCr78nEfwkNrFsVRlbFdCFcxrAUhha9gd4QGlPP+uSRfkQQJz4grnUK8es5GH5OidIsWrWL63
ppndBkbXAClLxLD2PxHRh7Yc9kLQOC1J1U9cso8eCUp3gSoJTTyKDQNMtw/NIvmEiNnHE+koS81R
UuRIHtcbyTWfHd6ZRY7yUQ3uG5Bt71R66WxODmMV8ai9sNj6mFeWiLN6dv/sn/05m0fAHvlnCQvd
tvkfXZK0Vs4Sn5c5KGlD70BJtVOyn6Viz6KfFcOXWftJLwBfgsEkAqHi8E0GWfJ713j4UZF9lH6Q
F/WU15koHizJ6qXhn9R54VBtagE2pM6UOsnngeQ8gYeFX/k15ZM8EJKyJQKgdErwSMetRIgpUcHr
uE/u5hkt0z+nEZizwY+tpKGZPBX9SJDpAODk32FjrqGwnv9EJEyLZzZbqemLV+yCZUwN9FDAWAfr
u3aAFvE5MPaIAn4LkUI7NOMgP2VvrmAiWzIh1cJbEGIXrEa0DoLTse7B9WYJ8MstQkaiJCe7O1NP
eZZGyUQR9C8FqeJRhqX9OVIILq3aKJ/CjNjWhuWRv5dyzEgNATGdh/HHk/mm+3xPSS0FqxKQZhLC
jWESXdNVAYtcSpFFRBCJIIv6fuNcUYhFfo6i0KTlrwkqW2VGGv+O5Dc0iXGhn7RunpVGL2Hkk09n
gAZ8m3p1YsMcj9LJJ0zr4UDMgBwb249lD64SHASaScM2qkc4/55JX8moWXutMZkBcLp0h2d0gkfA
0eAMfRQFS+/hjtXpcVbjV2PMpv7GEofQ7Po6nVO/2JOXH/Gb0emepYQGXCuSjA7C1FnNOj5duKYW
PJ3wzSbvpArVieHHS5o6ZLFMUzii7NLyIvpiJSJ8IKCUHuvJX1coKq2IoKJBIpPJnXaXlvAoSsV7
8hSs+Ap+T8iIZwtlyjg8slzWCkuAOKq4zHhqjlm+TPT0AEiOPx8+JLvZxGZoVPKlB9Lx5Hkktpgz
TULfuX0y+vpMW3nhTyOQkwsN83DDOlXiWV1qfB5TrORToVWGKbSb5XLRfCpFq5B2NZYoNoyAa0TT
OkJYRr50ledwfOY1hiRGTRXjxTHQaeMe+18qrZobva+BenmSiZvacMKmXCNG5lfn63CwrUqtiWqH
Jvn+yWA2Kj1GXwmEqeEMg2ZA7GqP+D1HGlMzySvv1XJY4wwI3Y4Kp19RMGy4p1T4rE3TWgrTt1gp
PCC/ikLTrDvaeIquM734pIMRc8g7CU8Pqr7QRIFCguSjhqzboGQjvC6/DEkyMueIoOshXWjSUswH
HxYvji66XUg+Wj54d3iJZz+M3f7tMkCTePnhQNxtrTId5qRzdnrp8txOd5c4/ahwVNHjcNP/tGvr
zeioAX/fXsyRDkUC+tkLXz7z1UId3OiRrauNim98ljuS5kLhtKsoIJL15piK2CfdnMbvYBKGr9l2
NH3kQS7zizcYwum4YxSLYRDUQ1kH+zJ46dB6JgV5fG9xJdOMsCI+0OP1cqhioT/h1fWe9DczcNEN
1uJX/xl4dMCLvCTxMq5ogqLB2OLECAVCFCFKOBQmnA8amWgogbiAQDSB+sENucVYO/PH9pUtEGks
kaB7WCyzNbZyJVYWJ0LIwlrXj1pls7WHl7GWvbH5E/rvqq8zf+C+9URGgo8zF3ndoHpU7BFZw34S
/CJeYfkIq9YgUQ7UMKEjFYoDRvfO8t5yha+GAX4SoZBg76bURu2wdlyPUf6Hkun2naeSuvFBsRL+
r+btFJBK0CPhWFFx1Y8W1YgcTsTSgYzAlBvRfbByg2DgpXoBsxHciJjA1R2nn2t2lDATMed2LdiM
+FqWmSgV4rEAToJVIGf83vuZ8e0Bd5aWRq2eEJ8jWetwQIwRy/GVR+5i59RpDkJKEJMrEBH02cFS
Rps8R1TPQzj99iQA+gjsJ0A55fs09c4NKZoXi0ztpXIzOvl9IVtpebW5RoNQFzA4K1rkcVoGYSM2
876n07+sgak1DgmDz+mDxbpll19b4P3cXjS5Hq37Pl7KPeMx6k9UqI/1H2xHNH34BakeWel0kBlm
7EbTdX0mnyPlCMp3obRlI2HC5fFTJXqoscG2a8A2IyMnwS7Jo9flvnnaICv1kuB21EOV5gXdmQnp
6YPOBAPc1mSfttf/oopIR5UwXpCCHgR2P9JBeIIoDd5LGpZn7/9TynvU9LW+4AZfN8YPlH32ZtMZ
+ZYpWn5AUdMeXuW0qTLbxH1UkQWPy+2paSXwR9pJ4QadxUr9QFI4bmFjPHSr4+XF2HUwV/jRU6kk
iEVo0Ol6v8ziYyMMSfE1TqFpm5Wdp3S9NqPoLN3nC0+rjWqBHA+r4IQu2ywBJDkbw+1XScd6/cwq
IGNWYFz5E3IqcD1wk14G4h4+U4RdplVlaSrHVsuOC6FWX70cK36MMUd8ry7oPpjB2ucwpD++G/sv
1B4YelZcD1Xf1ignMkx/jT1+vt6XTqMUjYqwi6v+qGkoQ86hYxOU2ki1SYFDa8CdGIV1v4JsnQDn
qYjSs6wNu3WVt4xIQSFbNltZsqJLsUlxlsVeg7++8/+Gus3mG3U6Tf/yiT7APFU8i6vbpOYOUJGQ
adRtPJPq18h4DsZn5IE0Mg3BLd6rr6jAe62XRUL+Hp6XpnEzzdJGaOi+RcxMzgh0MXLE6/YxtBKx
7Vhjroby+6TCNOZYJJvzM/74jmvCqJRAxXmihJUq5MSU6ba4mwdlvKqY4sFwO9WlrA5OnBeNT0+i
vJKcR0I6gWUPvgM6qzmptIuCfbQ/zrYCqFsNOaxXkMiOAgDFJzBgwAM3NVrTbRaaLZM4p5Pd00/z
pwlaK8lh+VBwHbH8yrez4B2TaLTyEsNCYMWz9lEhJFmNekfAHUQh5bqj4R4erm59eLOUoHpK9/Ef
WsHryHcwSbvuzKR1YlHRwOeKVeC4YwTJ/txJ19uJE9bHBR2HbheohtKcETcK0HZk5/SOxLnEUWyi
pVj58umFL1GIYH9TSROEpy1lvO9XRBd1iO2kt/hqzxPnQdC99T90zIIt9RybENGPeo/1ODKBpVxO
YfSTi0RJ9+/3kPsoJZSrfxBqrQLOJO3nvcRVfdSWx8GAJajHmeEMxYCliV/vRWcVTXCTVdt8okgR
kQSiK7Amnhbaa0QqvK+tivL8khxcyI1WQc9zfIsqbO6k8qUF+DSnO5FWX9qpvPLjnA2qwW7f0OOu
P8bubA+HkPOj4HSPAxWZZWsLXKrSZRdghZbFUjtHOi4gUni2tY8gW2zlZB1c2zdO66FTQaU5rXJR
dULzlHF4xmHHrKWyEC2V351yUlovs1ELBwtZp773L6wDR+c4s5uOk5IEdHe8jdgdhzj9PftDaTon
wH0O5+o95WFZCRDvY68jkizxd2obeZx/o1rGyEQDti0fdL8YEGktNrc0/AGSlt8tM+wiqXpAzqoe
iS5Ic4rg569maSSV/HuotzaUZgtIHahPj+HDV4rGtrdlIAnMKBKT9aSUVTcCuo/aV+WVGu9bPqDH
42Xp06IF5aZR7/G0//OqWAyGDlKczyApY30O8akOC8JNhWGTnA5bOi6WLwgZQid0dJk9uVGKkfew
EWjSSj31OE5pOUxhR66s9EyMZzW5NSKErlhsf1QYKnSDGoNpFFEkYm/VpHRIJql1oPzlopNrI4IZ
KmEk7Kbrg7nvU7WQ2x9MAXY+RkBwgsSPgLdqov5WIvqIZAfLRcfTVSD5EqNsoJS2kuhaDuXyRmmo
EXy/3Y5966BhmNBEWMIlQ0Fi2Y9EVHchqCYmUpL9iXH1Af2SMEV5n/zF7YFpxaU0pytNouQKidqk
TQFYm7t/L33rYFo2EndQsrAyyQI3pSqax4Vm7z89eX6XlbuAO6veNjDh6AjMwTVaGgnSoxtZpLKd
Q5OA03rcjquAJ0G/q5WI0JtYPkDF6Zu0JTq74Pkusqx37k91slMhPFtjdf2YtECwlLQKBn7j9SwD
E+Ziv+PGGKAde4q/NFPv+9aVo4ABkPxRJCPbA3Jvu1v8Yq9hr/DS6s9+2aAxYCnZrONFHD78c1n+
garJn9RFtm70knT+xZxuzNul7Z50FX1PSrleq5s6LCo4Em9hWtr77YQnghRNj01zaXJTumFInnaO
9CdaM5RDrunX0olxLsg/zqdq1l/LgUgl4JoUe24ubwq49O5nur06eMTf+nwJL+XW3HWyW8rpF6ML
ZULRshHghXLLOY06hjvEhY6ZKBttWoxGATQcoiZrcsZHC3qCBDkON05He1C8qYdgtYkrfvCbNhLj
Kb4YBEX2c//Mlb/CzJ9xcqQR9/80TmiD8QF8G8wTB/i0M54hYsNufnRpJ2frVKYuxBdm+1E645a4
Yd/oh82M2KLlrMSQ/Z42RrAdSrOgxLxZ1wcxQbGrZxG31YYdn1LPy3tgkJhHci6vfWb0v3cXHzWb
47pXbmmW3+zzWew7/FBVg8hLZpasxbUCawvaZqen9FjZKbWwbS9lEwLN6VUhKAhO1dP1ibNb8IEk
+121QwsZ3YJlSlCIpvg0FA5QTjnwwB4x9oy5aq3pzzYwV9nuJZQd9NLOcfDEUvhewzjBISHJna+/
pOquFnuIlymQZ/JJZ6FixnbfvcjWs4sgi9FlLU94xNxLzWWQiYySx0jrdysrWX58wfYf959elLlz
dGNWIp8/EKpmM9S6VHZq/5vST+hGnYcv0x5vHJDYA7wflj/vgPVXlBkemACEW0OOVeElDZFS5xbh
12QY1ntHbhieHl0eWrR5jpnBTmkj4TITZIEqg8SW/nAM3lMKLFEYxUtRyHVBR6GhMP4iysEXIznJ
jX3m68MLOb0iAtBTrYjlxtGNX4/ZuwIc6t0QoJZegS0Gk4S+EQVW2QnD47pN2ZsSepX6Hz6Yu2Ad
+g6s4W1e/6E6BJYokeeN8JKRnxItq7wuyLFGi9//aV+nOgN81YuZw68Z/XiRNPxIB9XJYVzyUuJ4
YLJEsjSrEdzvm2CpvJp/bb4GpZvfvv84pRKUfSRAPAqxQe+gnzWc+2qUnGN8dU8xbz77xi8rh1vs
70HdlUrxCPn8DzKyDNYjrAkLciq4BZwSlN8GejCNHs+rvWr+Lx5rlOjriEUM+4QmAG2+iVLdW1Ls
Dr6omia1uBv5qqOwBK3VjYfhDgip03VXzofwV0BUsJZktbHv/vSiNKePs6prWi//m2bX5miMHG4D
AEzZpTItE2iJPsnn+5EmMSzD0WF1sUchEXpui8BmSmZo35eDLN8d/NS7FG3lSGI6aHz94CEnSf3S
Xx87qQGATyrDyS1HEeRP4oMqA7XLcecU00ryANFlZQ8mmkN7wivU5XXCTsXvlyrFFma2c8FlRN4N
Ya9fFQcNQQGBr5n4ZWoBVbNKYDqHWwDGqUNgoKey/rzQ8rD3XSw5LvNFQCuuyOlKV/g4Z+m7CnDX
YAs86agLwrn4AD6bZpqxMf997hC7V6xBWrK8yFu7wvxuxRzOutIassTI45dgUZlOrhYM00aOrEuX
r31nHUKp8nUmXEevgl/SZQZsizr121jwW1ps0N8YvrfLusKwoAyiwgt0y7Gc6VBx43Ly/7Mw3It3
TdJjFFC+OBpAcSYnQWAUUIZ9ccbT6vInsvwLDN86XWRLcCits4Btroh6McSN7t84bNeLRfNBfeV0
Z17bk2W/5PR+TdSBbNpcvvAPLL8Vsw3MZy6vHd4EIT3lgN9EukRCn41Pv7hhLLqGHGlFvGtJBGy5
bREj7YBAXzfmyV4mB2X5y+HQ83NEXAt9nGnfsq6MEkk9FHewuNEz3gCwjYchbug0O7pgIrztIQYT
idqaWU8h0bRdtBOUZfFq1Vk6KZjJIdusucr0mg6udpDQdLD6iuYsIiTcjw3QkU3Kla3jFQqbxsZl
wgC+/NXNCwp/+D/vDuxt/oWn/APBoO8iJylHX42ELi4l/dQ4SheqCjgy55L7UHO10dlR6tN3JdB8
ELzxaX5cSpHvQA44XgDUTlSlq51oKd2fCyV18yW+T4n96L+6oexf6ghYBhr3q9yfMghR5FzWLZGa
VcxPKK1oixNqRGF6D2lcHgpuZiZhFkJopY/b6e+dWEXiOor0dWnqf+IKoUQolDXyjRTmcpiBXdVU
aWgm8rjynHVuU6LcGCCR0HPQsdQ139L9AxR/O19VEpMsBXwmZ75ssvVQhekfvOvYJjErHOYKNlbC
NCHIppdRIXXTnH2KNa4tpxjgnw1vnCar4pRxtBLpFeBfoPcd4tE04/0nv6eKdR6jLBkUEueBm3Ol
Pn1w/zUihu8v/BUjfXEcKV96F9j9S+22l0riCqwxXZTSXoUxuzwY8T5QzD6oOwqJX4dZNAG3LyPo
CzumCeuaEaaweu2H08ytKCsJ9hNIvdNZ1fBXZZRPo9F9ICpb06SEtpuAS8cI+BsgzM7W0sKq9wlo
LxkKTAEtQSOiOsJLu2uE8oLTcB06lILuvgwg0X0IybxPXX4bEfne0oD/SV/jAi76hdJgLTz3OWNO
C5n4UVpx5Tet93Io05gNAZZ4A4AvtDhfW6BIu/YgPZYivvY7bogPwjTjpQlI5ATfBShj4Fb7Ou1h
noy5CuRHEqqcPSB5PzJ3MROEJtl7EMrQVePY8/23q1hh1E5+dK2pj/ZLq8ef6PpoJxepiOr+jCYE
n+/mYq8Vy1m2zsMVZXDxytoFY/obehfECaZGGuIVpYMEslaQzUTvCL/4QyJmwdNQXIOjvHNCLRLy
WAQNWqlV9jPhWgkUWN4H2B2+J+ACv9O1I83E/zrKd5ya7/DWZ3KAXNLeNcof6SL1Ho9hpg788Iwf
Qc/KZdLAMwT/ezplKz7f6QAAwcNmAUFe96QqeLVHn2OM9DTXuPh0m6sVl1Hm7+Zgyz15yyLBwX/E
FHPeabYaWJuleh4femzy9t0YteK+i1FBtsMa7mIMUyZN0zJII2p/RLD5IgcFgqZQ5Y77EM8cYxoW
IYnRXfFL+lU7NZqoJxbzKVklPA2k4oZ+GDyBLEQ6WjQQx9a/SbP32T+AOirG6P+oaJkGgU7Oe3F3
YztgTI5sfth751F+5YHXfTLANx69dlDyUZV48idsNiBRwTEJVKkOd91VedQzRVZ4dZYBi2Iu3HCy
USU98MYLxDZ0VuAE31rgLooDZUDfOXYfP45f/izMCnrMeBNWgXW0iMvoVLYHgITiwE3+rDL+16MZ
thZ0fP+x+87+9/6wEc0gQ/mqaw2bAIRxGqWl/lMuLK78b2qyDLTMPreWwhUJtUX5gen8FswKtjIh
sHtBY4tA1o/sK/9vSf4SUCWkeSFHFDF6DupjDN1KnpVyu9ANQEjNELCCygMiOBUQR5j1fAEG9peb
l4QCD7S5q93xk4+N1uU43xml40TTuU5Kq32pbzqxCf/cQs4ZEbUGFCv9tEbOWij15cBKewIcBUCO
HOMrUmX9XQRxoXNJKk7xyLXir8fML4ZCmrHJmEpjbikqmmlRCNyyt3JzztRc18VhAeMylo0MM5Vx
7OQnSKCzNdWCu1dUr7UgsD2Q8X7Uvo+gotM24jkGM4w2MpsKMMZkDYvHVmtPx+vTRQBzqZEH1EQa
iA63jo9rKFm6N9nHuiqsXMZDBNvX4elHzD5+DQQ0SiqCL1qYvhUahM2cVN95veFSO7HJojoDo2mI
BJkewsPU209b0NYEkORIOrODe7us2cUsDyRGO/ycuVxdfdDTRIKjnv0/JosarMHmhxfXeBmElQTE
LOcCjky1lInRK3Eu1DmfUuOLcibxvExhfYklpK2Xdc6R+rSx1qgHF+k1SNmgs/Y64pVzOLPMQbD5
Q75j8sIzSVaXuYX4+RjFs1/4N3EvBKms1TegEaPsUIaj/h3po5LLWBQAuF/S3rECLxv6MMGaHKWL
nGHgfkz2jNd5TeAYxH6ta8I/vUUXn2g4h9xe+kHrbho0/1FDHgnZApIZMSV/nD6C/MH0iIpYHIqV
Mwa0cy1wgQ3waYUn7sIyA9kMeJPri18rhhdYR27JLAw8roRiQPugrKSHoaY4cBrc2Ll7ZsXqM1zA
O1FOFnpxGoLxUF1gqSWCxXKVL3VYEWwqhKtbolNTWzhhtuCsSPIR2msK0dTj598Q+TlmoC/tXEtx
LD+9RboSJA2XJSS1/5UjyDWTZ5y6Mzzx6WjDqz/4Mnn6BmNWTpqXSHXK87FF/eb3EMGT8sYxF6hN
ueP34iakG3popKyLObFhGpsA7zHmDRt8GpaJ7nCY6F7j6LJ9Mvqzk6H1j7Q9b0aq43fGpW5mlnqk
obbtUJtrqSL+Aybd1xVl4i1Uhz3yJt3IzLx5Nb0Mnzlx8Bui/DY0wr34tfD4QIJMe57+Ya1u1ydU
mAZoDGR17IEptyI0uYq6PMCxXiBVIPyhSw8xJACAg7+vfeKZaCfJSEM7oMaR9lbjveE0bu3MxSSt
N0/HvlKJ3HU3zMfwDqmiq3FZrNIFt+zcth2jIOswtzZWcPslCDNL+Gi1DrsAmLE1fqtP/stug6I9
JncwvevcBPp1lsu4mATWs7cfm/40/QSfybXimyIRBcRykANW9JuJXOQ5iCPc5fRPn92Goknr1p5H
dsUqfElhKUP9nACJUWBdRY5T8h65Ekvbr66iKGYQ4RchmAf8pZ4cvWdhKqnKyvWtSU9+q/xWJabP
ymYGZUZQ89OIhKNmM/AGH+peveVGAibi490CpTcFytVwp97cb02EnOe1ASWhxrUEV6XuByiCWeEZ
MWKDFo3INPKQ1iLofJQKsDcybn26egfY/T05zMiX2EPxlQinySBFZL4LhIy2q28DJ3JsgHcnOnzE
nNN7dwSA7ONbxkxXagZSDS9IVWdHI7i2Z498r598z2IOAn3v1JQohC1b2HXF3/jRz106ZRjdwciv
yhCQV8nGzGqNUeeD5s8DGF4frqqahUUx0n1YWEvnXhQze2Lq7KFq9xfM8azFzkiAO4s21YOdtXUe
t1nM33lW4finrbunxkQ/vMO1BhtLEjiCc22zN7/aK6yqwtXxweb6pYQyrRUMyisxrPmgDTE5FDGo
HIsE5PVG9fYMSTjrntPIT38ceWp2kAYT6i4QVVxfOVHGFNAc4DN47MXoEz7ZU1DRY7+6iphc9x6y
TDc2FedU+Yy4ZqfU/T9yaJBDmU68kiJEitEUnr5XJJy+dSuP2C51l1uZe5yLapASaMFQ7gxYJvBB
ovDmyo9fx/PfqzqMzQLApEmAljdYDONBbI1Oy1pXkTltqTmJ7v1Ts+9DcX2ZLv/xreck63QbjY/+
oarvFRTXwhhc75XB9wCyipdSdObaEN3aZgdzHGnzcrAo6r2Wjoqpms2pEBFuHOudLU/oQxfi+p9Z
hTJvyra/GsKMl46txHZoqnCoR/JPsQDNSr5BhB1b0+hE7shzifJ91ecs1fUYAq5uc6d+HxERVFNs
lU/eM9XmLPAu/8SBxZRZF+yetkSgvW6jgnM+xO3AfrNfKH6bhHlQWsAFVb+8AmHQJ2bfY/6WPNZM
fGO82x3l+/7hUM+iq2PYV06lt7SAhUKmKTLYuSMm1rRvg/29kWbmkxHuQ6AbK7F7njOdV/Z7UkAL
jDwjtVcTdYJDkkIDxg3ute0SUl4T9eiZUuSk33n3T68keZy44+H8elocrVJNEOvFOwqAKvuA2CfO
4/wa8hnZoRT+VzC5r7RxbQyQqRk+EnRDnivfDA4FaE735SxM3Piq3ISJUTw6QVr5iVIHc/KgElVg
PGzgkgSs+RNbmIyPT+J9I4y6YMcAjYklbsajPaaEAEsc6T7mxaUuY+39oaWZ4/odd4V9/In9JElw
1VvXebokO5jsdGrFyh2Yue8rLu04uvRoxsQNZni532tS/MLi/sVUwnsDeSOUqfiFRRjJoKGVtTxX
oZH3MM+b/nYdLMzl4KNWTkRAJUYXLuXR1fLJ7bvVnXfhwgf9zjLlgo5t1Wb2rSXhRBO15tHN345W
UDcdVscIUZzCGmI5+N7a4zdjKhZ1dZK7KQE/iCVJp+O9UFv4QxRXGQnjha0aPmyu8yA0H0cpjknm
1sabbgd2ynYc4Th/FUn867bzQpU3PUpaTTKXTCSAkv8V3Pkqt4+l94P1hKaTrDKYTYJ/TGWmG/8f
GHs6fJ5QRYDzszxhTkoc96VI12SmEt73ys3+efQvKewwvSBHFvjzMdNTgsq2/pAYt/eFmhv3U8y0
D5inQnjVlQ4rt8JMPm1Lu4z9jqMUzTMsaYW+ZgVCQ4uorpTOW3uPDB5XmtXXvHP1Gdbl4j3z3wPD
Zwap0HFMvVsXaa0M3w/juzl0512DbWdl0roQ92Gjv9uCRUKvaDDzqUzdoiWW9M2hYEkqdO2goeMr
9wfoZ52BFb0sx7Tilx8KqmvG03ZzujyJsslnYCHuXkyEDYyLQx5Ado3gt7ylktdjDsWBv3Z7Mbbi
j7pJjmQc+nm4CVvpGPegDGn1w4anauSeUKBRbytUi0OPYwgCE9uGAASBiQEBkaK2a4DWBu32Ha0S
MS+2C65J8GXGyw0gVY0Tu+YYURB9tYbH+FRXXfayoqJau3jwUx8lpp3kTu7nxvjCZV+wUEVFNMBy
fieIkmGFSOBHFmlq6rC4fMwkS9lMC65ZYUdLUBUgjKHSbleVmYu+kszQdSgnnOXjZLkcWj0no2Ru
2XXzYlGxfffOc9r6CmNH3q/WV7aWwYoo8d4Wvzs55XYRVvup3wnJlXCrdBv4Fd7u023EN/D2PQWK
9upEdfcXgka6pukkZjmYA8WOUg8MZZhDfMULt824UMx8QAobBhfWZdV8hJuH0+oDpNfvgmmiyrp9
lONuA7939bVQkZNtJk6SvFI/hb/izYHiMAXBDeTO1A8o3436qw/YOMYPOznOUwaIssj8gBCUO0Eu
8W3ra4EQZxcdc0ez3evxbI/4TI9IRnMMgaq3xkIbkEqYpP8/Ee9V3G6V32qe/R8JxSG8H0dN+gLt
cOIU5/XNaV4FpOTKm5fLRkYB5RbmjWV1k2EILG3T+kkIka6+g0C6FXXmzjnGvQGMcXZ+EavCcDxa
IHQYiWeTjd1nXLIGhos/5c1jFyyQR8+ESkVh2wdFnZXSIqJvopax2E/12z5+J2399+wihQkF500v
iqnDTMJPkOhj/MKkZljjLUTEaS6NGWQCC/JnNEDPrG+W3nWumv1csnPEzi4wrQ046HUmq6giQ0ME
U/mB3DQLwfT6ZP4TSTshHms1FHy2LC4/iVzoDqw45GWA6F19d3d8x3H7aAY4tB9m9TADiIx/lZrx
yOYjLwIWxivqKvyKNCseaRqFew0AEXkI4pc62jyVWRhnXuWRk9FjHsveSWPdyZSrV0N3rUX7P8AP
k9C4IWsomug1+aWQ968UOj3DWLE7XzSWxCMiul9+MFd1kzf07nKWa0ezIlunr1Nh8JF7BB71TQZr
2ukOKB4PLztORFdzKfFmPSqbJ0jDN9ZarEMWHXFlP0L4/ZcqZdGSySaZ1AyZ8JbhdPBZJMk+ZJXY
TcT9tY+fHl+p36u9i2+z0CcZWgjdDli+z3Ohi9szT1iTp+vmM6d1pktu0H6QKgpImTd4MTjpHamq
XR8npCOys3qsADxURcteFAsqw677DjCyZRBl6CJlhzwAp6xUbT6YDer/Q8748ZgYSfitR+pWqIgC
FznnuwBqqXlaDy40hDBP61dege7jYGfHVZx/ZqRres3+Y4FIy4c4qOWjg7RRXu5ggV830i7sOtYv
w5bZzgxFWVHRv0UP5HFRXj7OwfyUf4JaPBKrPEg0Yk55ZN3znycnrb7/cyv8yr02a+ugKxgs2SEU
isTJVXGhgMEjeDkPy+bkIEH3DgHm5bc/zmvWBhCkgFDYDhRbupxMsvertYiD/yGaLDgPvMosJUYW
zqxdvziPzD3rOUynBY1XhbLTk7nsk47f95dgjGJZv9k8Be0ZL5EodwgHbBzMflk6YNF8kFLbcLOs
qU8OpV2TSrSTp1q2QTf5h5fhfKXjHLygtTYu/n13CvJaRVaPEBu+9fH6m77n/JJ12ZISsiwrgyZ0
tfyuOVCnehxVkz/cU4mBmBr7t8vuHBQH1cSez225C7UhqUgdkNbzwHW7T604ubrlwUBakEPSpxE4
u1/g6ujYauAKug+kDP33Jpm45W0jnH6qEohKulk1o2QUA7BW+nNgcXa3cjJmSZJvgvJGD3Uc2xHU
oaF+2bOsmmslUijYe+SUAvVFyTaK+cBV7Uu7bNxH0mDt1y5HBEutcs3+gaa7PHwxWGbwguUW2XjF
l2vIUfVCYPLkx3+tsz/2lRfAoK//XkfyvGDczMt8YZ6D8+w47ETwRZtJbEvkPn2vf9kK9sBixaOK
hfkG7k1onDCGbfE+TDcNGu0c8jtCah3zC8aGPN2Al59Ed9hmkVsAZBfuTPOugpJv5DI/P7bm1neH
NiI3P36AXKh99IyWOf12e3+bwLhgWAL9ZrbpMOszaKZJyemv7iCfOIo8lqkgrXX/UJ60Zw3k+nzi
Je+Xhf27WbN+yhevfe+bHhjviV5MGtCuAK2TPUTNvBwieC+ByielMxjP2UTueD3DYJ7TWpw3/DHw
eVk/rdNCcS8ZODEaf+Zm3YzcvR0kemcpwyhp6hyBhmd4PWEjbDpb0tbcHVJGEL/wZAHnZLWP4+yf
ZaGg8laW0injbr/uoU+Nr+6VW/GVQQYieIVvrvnA3PB0DmoGfQQOCUq81f68NWRtAOSkP7fB7RFn
mljrfSQJeqf8N3wTNjJXTFnz8I9fYJD4CCb1SYnD1n9U4Knw5GUp0hwSV7NJIL5ReV6YjYttsvei
xovrzewSCg2AgrQBXBtyDkhNg1nss86OSsayMjSP1n7/cF/6jJ+Y5afSSZeCyva0uWkXycAm5UlO
JDNMsU7L1SXZ48A6LXmmAszZZoYkGVwze09E15TPOPhaMptiosp8MHGfpuXiyHY/6PNixvChpc9Q
8ftrM4oNySsJXxiscR//wPunBSM60nNhN+fHWAfyLtZGsDyWb6IXCd9qo7NDgOwJvvheQYyGoPiK
sXk/MaxGO8CY+eGW4sZreyRh4F8h9fNOXETHpYfG4zuRqQpqESpIwFzkug9tkOJhLITSqu4SavD7
cKjOY0Fbx+EfB3Z76vVI1fPRZLVir+8ayZN2YzAfR0mN2bVgEgNnEtPtXEPvPzO8Rt2bX5zYifGd
peOQd8uyy9/phAMpocfEuBRqGZq9+Rx/2qHUsdbAKgZHeL5IerQOuegomATbUZaOcbpEv/W+p5os
t3K6PW/WG/Up7cHySKOY8EaTdiQnOw3pWxBXV8xTz1OWPQ3LIRxbBv0eK5gzxGcu4qMl/uEzhWsJ
XNRvdWhG1GBQOgz0NlTsvTMpWjik7tRSNicXijfZ/LmHVzU7uGt6Ott1eDZXs90dhqma2wPC/XMh
C/eOoM5bAmvFEh+lfgXZvmyGeuLNnV6fKPWxrMZ0ixJX0y1GYjBW6axOef15v/ndt91Cd0C4bTS+
6lcKKzfLtBlu3bM0oPhTQQYQH+VF3N08m/k6yjkXgIVuY4OPWr9ZjSNCRoI30gPqoilzo1dORag3
TUPd1nYBhQG0/zrQqWd8vdd4UYktgM5Xrr8a+QsNLHfRuczc9VxU4Hw2rfkB5MqxOKpJ/uj048YY
tBqSZ6F1YM22xO/Qzm8UCTmIxr4gnr1emj9/kVbrkbaej3RIco4Vs83FKuIkwdprwUNnaObyCAvV
Dvz38CxvZeQhlQE1RQbRqjHx7TZl8z34v04ZLd2Yo1phAmMC6M1dhtC93Kx02JujddGQzDSXUrLM
2L4Bnd4//sNZVCv5B9mv71GKiKjurOnquSPDNqo050yN1LwMWgmnrKqpKRyiGu63EejxhDFhetde
rp3pu0Tfaql9vy+tnZvhUY56hVnWQY4znfq5KeqEkr27q7E7YBlKDNX37lDtAiBPsUDDJLARLfun
pREqRzE4KcbOdiFgjv3ReWO+XS9BzM2t89CrEF2dtB+Eq4BVAHnHyoyhXjTC45al1LbvaGXCxJy7
2IifCRDL97nSJHQSUFr3qqS6F0zTuTH0ysuGoZOUweFWA9jqui2018eu/ye+teJhWu0E9BAMCt9D
lJ8iPdK6yFk+76IYLnhUgDGdKHbG/2DZkpuqQvyllX/b4mJTf5EtMP8QS4jBS4I95+zCwCa2QIA3
//yBHrjlB8S25mbUeD1XI99t3JtPWHyCZM4riOQfV9Q9m0L2Ql9wBH2LcvAjgE54J/maZZIiaDsx
rkNbUlpefFQzQcAaO4LoMARe8D1GuOBFo7iGt0+Pay/0xz7SkyLWuDgOIil80WSUrWfRmScvOGmc
ZmcWODU/3fT+h+zKoX6ASfVzrcG7/9ueADBZ2++R3E1g8n5eTtqP1NKfOlFSkxeBuo0799wrXdCj
4gwpazKvR16RexBd7L0bBR0JpeQO5sfMYS8GOdN2dCgqv/V2RTy7VCy0kcny3ZT7eRBgGpdfW/GJ
a0o06yDNwgYv/KQSGs3NObAYrePzjL/gOGHccnamOzBpx1bxguDg7iDXB5LoCQkHDgodsrTQkSbn
TrpgY+jmhTIAl26K+KOeFkvNa6otROHio2z0Uk6sHElrRdAnrpuDmzz0f7dO4ekEVM4TqoARkXbQ
/eG/Bvyb58A6XZcVjXTmVrlR4yeD79APLHKkxQ/bdLzd8iRCF00aIdPQxTM/Ql8J62n8Ms7Zyqt1
2cO3ZfD3LW1EpeSHDm43Tva4g84Dy2l/fZ3E8YvkjNrr6r9pfhRDYohWiqfBaefGCRtwmU0ixnyx
cBl1Oq2y1btQJfhYH/DoschePg3E7z5P3fsdRLOSjAzJOpdkvJZLZkUwzAX0O6I3M66DoEBqOVRI
096/DnA5s8QsUm8jyrhrP7717DJRVxeV07sxWwwLZM9CKPRYtdGjKEWstVywszbAK2hbZbduHYxY
9jATX5kfxJVKc4GlfbW0KOtVkKDRTM14xTxeYoG73twtSEIzrwVM6d/NL03GpmJjz/nC8cubVZQ2
Yrvyrqm/fXAzrjSS9WZrfppkjZvWYdO4AptJwJ5ZNmUXlDE99Uf6LwJzgSPvu/18gXztoMzbwD/v
uFC/cEbZZu7RwamCkFoJh5NqgVMfIJv1LF/W+xUaSSnXrqXusif5wncmQkoY69T7P80AgvvycJLH
a/ou+S0C35+u2iqvpDGtKuGfDDZKyOtIgskcmk+6EATGe60EkzyoWQAsCrnOBaWZoLTP6ibkv37d
5YPQoZexFxAzbk1T6pz09Z4CelaT070VvLWp4ioFnPA1F7RlT6Avl5SHB1Oza2gmtRCyvGUq5YWx
DYuYs4xZfJQ3lgPTl+ACWjmcEX/2M72M9RWvA4T6EjgHHYRIKJ2hXesnrXAlV1B5FlihaUiVZXiM
NzGGiqSmZyw6P3j1+QwzvgPJvRLQ9bxrFafbM8zIa0upKEVCVNelHl52xVsmGZTK0aqduWVxmUXr
s5gQ0P8kvblEnBAfq7dcUVFlNXc2SunSU/02nIROSofh+I/biFGoSMgZEoAr8GFJlxy5pZewXK2F
8q50ea8q6FTc3Yqh2xZRm7wduXT6U8hZOKDHVCvZixztdkGIGgl3JyejKtMF6l5OqCMq06c+/mU9
HtAVg9bwumHmW55TVMyd6SNo4/DKJTjyEPkBIL+OIKTOdKZY/e7aieI22K7RkBBjHVxiNvs/IwiW
LeXIHy8Vh71OTPiWHu51Cb5ycv2XYDxJRipcY8eeOduvYaKipeGIb3OlagrK+Y9Q2qka64ScCFQ5
EdWRqUtn+3aRYJYiKBcMqvXBiawh1L9WxrigdPf1jux84S9vS3Gz14K2Aizwg1JRisWtrmzX90YI
7EC4A6KmzHKG71M7BX0x6NxLyu/2rL1EnLGkR3FUPOj6oTjp1C4nO6TpXZpHtxKWmcNLeTMpPg6k
c4YU/PTweTYJmifsA5/kiylJl+Da7PV6SBbNZZlDOylKcq5gWIuJTW3QbD3qZkGB9047f2xyIwJ8
d4hl8Bu9eOOXK2TBnjSs6vanPji8WtW4c4FODqh+lnA9eKBf6+yh73B7IOz8QYI4Ut8Q9wyG/ldZ
tIO2o/j6xWezjQRsgY9yYOKz18p3VIpW8eB7x4tbSiQG2uXU9CBJdR7Gvv52nXF1m4Zlq4xIZ+Va
guVg4Jafjsbu+zL69PRiFkz6P6cZKn+WItNnu1WvebqMYON7zpeNIawV1Srcz1MBF6KQOnXZJDl7
p+gyQGirqi3YsXT//L0VhMEsAm34cv/7Vw5Xb7be5vqDdCsD4mt+HMo3irehga07awjv4nqgOL4/
u9PYgeAFkaVf/WR8G1NHmzg4xXO7SoZL7/YhUaM6KFF/s5HOVGKx+BhPO3T4rzNoMmY5mYl1lShY
bSnFlvMA/hPA+Op0EpBz4sE6b/Y7W1OwVXdYJ/LXxAIu5/ZBnPUawlgGVGIPO6cWpKwUdR3KNQfu
6rHALn8Qa2PZMrGoYqD8YZ12t2Fg8GTpity6gWOY9VMYhNV8Lrk8t7l+INXJGC6UacZYQLo/jsgi
7BXrAEOP/+sy+3qCG7NzJvL62E/bXKmVPbmNGwWHIRZoqp5cjRPQrK/uWtd1EnrbNml+DbJeJQxM
VHx/Lq3CUnI35ofprldRQunRgK27vrzxkyCnOXvSiA5oFUVHC9nGVcSzzlLF0OrG8wT+eqvMdDpW
v3Lt1cMGstB8akx3vqVBGjY+TDAXeWRhhiffVOI/KkCKl/tZiCCXhV7QmQQvvqRrd/za3/WmZDES
1s149ezGoA/sULdiahaOfhNmzY5/xla3jlBXM1w5QLaWBQqYdUelNsUhWY/8SmKzOWAa3N4fo27f
rofBqjWYaBhxETNGl4/BkbMzraBfBJqJ+qXI2GExwSu0S3aQAZSSJq2PdRJDrXu5gff/3+ObS4BU
skkk6IbtV4dFsnlDIQ4SCUv+Fdf75c0RB4GpHMt2z02ueChX6nZ6joJbFaAlFJNhpKDFJgqEcbu+
yncI0Tca4r3L7QhoI1+5pjkY0yxfuhaqeBqNB439rLn2TKLs6LkvwkLx3boLA2eMfqN632KlCC29
AqjoDg2c4iayoZilgDvfCfMKkpc5dPF7eKVHdkFTXxuNxP38FSvywO7LqHcfbmqSu/LLal8XjLdn
I+AyErIsLxvGUb4Buq0GIuauogLU5qKlbE5kyG/pw6hcPnulzMDnTxBsR0xk1cORsXS2p3NAylgd
C16GFUiIEONs2R2Cfuo+NQPUL0UovkKru9bVapWL4lU/ukXqkLYeZE0/doGNKpD+IKN1iEWKkU6+
+eseaQ3rEENtGzCjjmwFt4KNGrUYNRNyOV7o20nYlA8h4EHpGCsoXsu/RuDB45vDA3yHxXfLBAKh
qMbq4vLdCUjPBrw8rOCCcbK0sLojDTDZ+8GCOXasG3ZbjdlHve+G287fyLZoYjbvJnT1IY/Lsevd
M1lpqQvZ3UeRQMC/ys8fMrxjptzZ4TKfseIp53h/WcUvdT91Vp0wb4+MYa6ssBtv2Ra6BhiAK2iz
UhcGLo1AlB8Z0DxyQPwY6YRQJdB3+lFFo7wxuBrd9sANPOjzMGJu79LYYiTUOkK7aDi15rQyuh/q
oJUdv4EtRYgiHCajdy3i++HXoatsCVodDEaJIj98Rs6kk9OAr/3SaUYWPNqFuLsk7D6YZ3m7OeNg
+4/CeDDkGMjfnMsbdXhncJ+4uKYjiXKdeXhI3u6tDM4isv2W6G17QVEbZtV9wGn2b10BpOZbhyxg
Cf2rN7CwQ+CvjH9h5wfKIRKBDMVboprQzoCJhMHzbXKzA2mynrEt33+4lygXb/nw8KG0RxdTV4Gh
s0TeCDq96Ks5iWR+NU1Cjj96NAVoSdxpxaPXyoQX/mo28fhPoRQOB3anOaN/HccfJL1DnFoZ2pzQ
MNg3lFw6RAhldIOj4ZIglQhJEQgSai1S+N7baJffSZjA02SbCdCHUJiQRYwuVaWDCXIbEpCfqU/R
ZmIBywN8kx8TPc2R05tSXXJlcM4Rymzs2XfX2/asuk5rybzE2AsjUGlFu/+mWaBARiC0U+yioM3I
m2ONh4f1KxiW7PwW0iWYPdwdAkxyVx1SvUFPB8en49NtMA5xo5CL3/klTQNJfESWnXRe4lE99Ijx
mht6phglJnzL8F+RmIDSayMkYYMgvRngG7nWe2YX3f0DVVagALxcE4H9lKGpVj32YclShtNIkZ0u
HfhPthRpQ20rJ3moCH7xH8VJ6j4k6jJy95LSfEfeKQrPAo/OIHfPhVK8stH644jIlIZN7+iUHYpW
U+iGbPQUXqfgAhYfZTgon9W/IB1YPuO1SXIysSro/U6k+tcksWUDIRDAHjS5/qVts5n1cW+83R/2
ehKxeTihJyAAZOtC62XW6hmrPnSVPFgcTp4B2L+98BSErF/JNe7BB9rK0VRIKXCcCEwzo2+sELJx
UmLJdv52oMmQwBRTmusM4xyqokOjilyaGms+NpcmQwiqXvzPkrkpdxaeqhB6xbKyiUCAgxsTICzo
jClY0qPM4TCeHgc3HF4kW41CQA4ir67+2JVKEQ+NSLXMC/h52D3HmrDek6ZQlVrQpr5hIC8evff7
Y67/iLoxdQqlmQWzJGskixFRbcKfS6z6zzcrkGp1EPvrIfTg8N1cJACBbYorN7x7CihNKbkHwLgx
yAunVxA36Hqn1DyhqlkOXdYX1q8MSzhacnZ3Hd6FryX/mjTJM8HSqRmTdq34kFZ42iC60ZDcJs42
Z+PHfnFsF/sqtCS2ojbnGdB1JoPKQ7zGFLqpnhlEeCZW1Ky9Iv0FDfO/zpwts++F9AZs/e8wd+qG
Ob6VUXwphF5tZUiMs7NGKsdPvtqvSvKDpC5lch70m+Oq0wWH6tSshI8y4wwrtiviCBAibWdWuGjY
rK8qlazrmGzX+P4NvrnYN79M6+2/YUUGpVdoT7GMkMDLREWhDJTdn9EAa3iqp9mpFdPQlGbyIdSv
oWCmO21VcqJ92R5Ivfeha3NYyF9RX2cCQjbUjba85cT/iwucNpPIWhTqVYzDp3GfUzTSgSBLrQsX
/i7gDY3LIl1UsihIbjHl38VKDTJIP02EM/+i1nb3iidFxOCSGWOPEETNKQm77sDFu6jwydsoQmp1
1xNYjCa1vJsYsgGdhl3ihh3vogENSqqUYPG5PwjgOliYNJJan8YLw80LKSj1jZwY3KJj1KAsQPPz
ZErM8gHSpEd3xIDhAilR9aM3JaLPy2n4aahANGJ9A6kFMKFYUx1xBemkEi4+4Hq8DSk9IOfNAc//
taoF/vXA0TPELGco26igCKOlu9TmLmk6TGcSPrl54COSsAgKCsbBlCkUh4jb+xUUkEvp3dL3RlrJ
MkjU+qh4YoDBPdwCZS24gU0xDBlrIFiMscSWVxsvyGgvMUbOUV4PY47wufffnRDCcjZZVIsziOmU
FN/UGlzmM59tKKn34xiTCeDiNa87h0aosyL5I4EI5X40ZG4fE+bGUQoxIF85q6hGNyIJOynC4hIu
Rqvx5TaKdRRN6iFdcG2qz5hEOA7BF1nZaCPoTJ9f6aQQuOAO2Zc02qItxnakH0GNFMh0S/Alx0q/
eVFpMQeqWjnkSlrXFizp6FOt1vsmrvq4O4o8Ed/KXt+JMnsizKfAwPpWEB0n92J+kvCiYs5kWQGM
fQuZyklFihFxxOqvvfZWzeb+MB6fBH/NxlWQ/X3MJGpkML5hfgdEYQNl6ow52SWJBG3ORnnxg0fO
44jXGyGbSh09/6Mdtxr2fbjsgRjgWGBfhIkxLJeDhnUWg894BT5DYuvQ8cMdDIBTbI4Bi/ER0UUj
msfos+Ynjm5uKBtiMq3/98BC67XuGpcAOVLq6cRZeo8jO+EA/a6JBJlafqQZaiH7Sw2tyn3rFgoN
VGtm2rJPr7mCsPTQXBdcSfYEbYxDywRcCZg+NKhlGGo6LXhFVqyhSSclGfXVWLBNwwWTxeG67HdJ
EzA0r4Eq/mk6QiWKV9g8vd+n5ys5VTQfklXy4kUa9G/Q6T2MqNYTbvTBfFJwar/HF8i5KheVgNRL
ShEO+LZAuL1WEsVZsfsHDFxrgeRWHnEtQhTyAFQPy+4sBFKdn5xdEaulfWws9vlrHJ5QSEGcV8E+
F5cHbWT8mMdpPSA8Vxn2nEc0CrkcsWTveyNCTutfZQtMs6M2Tr9UprVFSHIQT3m+Hrnmp4s1WxTd
V+VwKUE8Zt0vdWzpna0DjdUQoCWcLLGlugiKGKahI0Ml6GsKeShh5tB+Bm/2J7fj85vIwAbRPUGT
t6EWe4OOECHt1+Plljz4+hfrCdlJG8/H4DWVZ4uYCxpZxOJ42J8EsYNrqaiCvO1/wXjSFxjsUj/A
x33XB/0t7AJ9q0KHaiwSZopnd3YvCTN+gYc6d1q6fsnRooRTl++5LwqRYidvAeimRETeg8hWB9M2
la+7EXFZ/PSbJidmAalSujZCq6R2Edztt/GJY0ao36Ngj9DjhpXNA8Yt4oo9mOzefbU1H/HxDOJQ
EFppZCH7uPIJg1nB5fkF26gceqmI6JanjD6E6VzlUB8aCVKl1AvobxOdHGus8NFNXT6nmHIqkPEp
hUoGmz64U6WYPOwqgL8wZiUxI8U8OPD/mytsU/cAXVFo21J5PJ35QnB3wsucwaxnRkPKU79vRcKL
6mQ3+uPwRAc/Fld3lT/z8Sj0hdxIMAWYehEnnWuCSATn9AWuryArAwsth96L+6w7fSzPrbVSGxi7
1kk/wE1ejiKBY9IST3FXEFLoCnbvsP4AMu10y7G+LWYAotzmWGEcJ2tMA/H8MUyLNTWahpVH6fdw
rVdv3+wBvD5B8SbQpMdZmRUtuOc6i0oi9lL+udopYlkgYD/ADSR0oBkjpAaWMAU/nsDla2izROch
5bqRefGFfQQAHiDCMZYHJvvTNUayMhikmRXaRfkkmIRiuVBGQov9UgfX+OrTWHdqFJmWqhCf5sKe
Q9QSxuoPE3Yfhhk3WaVbu5Y4Wskr6flhT0HskiBSm6geLop9Fg/42G0igGfPZCRJsM0sliYe23zw
4blfal9gv4Wql2TPIa5/QuVkSwSq8KZn9X1rEZ/PqnTKDJ75yiLnNT8uZ8/ZkeI5iIUvH4OjyIue
aRundKiSc/p2nnR739o95jvJni83P0yDfvyAqozYdBwjRI69U4/vnq70KFAMTQf0dbBS8Xxwqeq5
TjbR+PiggBiWDcVQ/U3gEginCpW5fB0wvHmib40LTYc3UnW/x5Xz2K/uw3fAAtu5pxHvlgzCQU7W
re9A+xTxJ1i50dcOHy3aDMuwWrpkq2V/aE2k6Edqk8RCOu6Kaix0nkTj0xqHtzcvl8DUyxKEoVFD
gtGHCzv5eXMIsk/rvXovwf3v7CmiLIX/HBYIhwBvzOIIDTccGVqI1rMiOqb87pdlSQvulH+2H4hs
nQHakq2qB0JUnn761fVYWHXBiX/uiFJy/ZPoYPDgZyhIGX/W4lOSFrio2+hVcykfAUTqbeFVWhkv
IFUycVxkSmwfrkyO1UPsNWIcot9D5EAEm14d+NHt+DvMqSB735RLAf76cyUDC/7u/zKtWd3EzSg4
6gfLC8MiW3YZFV7niRFn3KjNg9bXjilArq8sngXNkbBRMXd/FknXnd40L6YySSs1mC/uWOrg27VU
PohftAxUHUoesl0nUX64rcJBPttgNIxbiNsnQMlCunnblzkaAuDBXPE6K8hQDfi4JalhQlIK7llY
eDcCaAikOBhSkmA+jdn4WTzEOWT17YOUl+zxwW7Up1coFWWcdG20+W+GPPYEJ4a//tpeP1eveww2
psqCOgdT/dceEW3rYj0NrYyXaagSToJyp/50xHXvo573rW4Zq0oeh9CEr8YAN73dydcL+/1YaYal
oc10lc6JJPNRfjDdIq8He2ShFPgPxi+ion6Q6Fv+KCx6yHwLSF54HQd+PYj5gA+dofvLpiyuuLUt
/89/OWPGG5k/3NSUKneatat/s7+wCkzSONw1p/gmSQW500csScY08230M/+tZYYpZIbX4S17zQND
C4dFFOvEC3JdmHfA5nHdOp2HrM5SkjdXksP8tFNMSZ4G6MnfxVgJPBCbBMSxSEXs6BMU30M8DeXZ
dJAI95Fg3vN+os07xSeWUsH7MJgIZp6EsKg8j54xzbzLWKFGKoK3b/nYAmRS9DRgaQWyzwg/8F4u
fZPb+63NQ5plRHFM9ncrPiyPxDZsXStdGEsTK75JwcO6hngIdn9ggWpK536mcLWux3qCPK7YCK/n
1+X2UxKAgRGygWkbbXZfaDkgIBJiPc+ScY1x0T21/yqYovbsWdfY9YgbCCmrC/2FtFXhh73RqNsM
/51X6wgmSg9+OW5okxOrrwwv3pEb9ipO5DO4O2UJJwB7ol+NNtBZJzTQ7+tpykq7v54fuSpEHKfp
Rr691dkGPFEoDAjXkrMCPCAA+sVPP0Rr970F2g4IQXuSRrw1vvrAgdZ97eajpd98CQi1LsbEAEu0
Rv0WVGxN9Ldz+qCxrKOZo8p6nFzAhYL/gLU1xG0XjQ+ZItJiUXvGWN2dd9UMQZ7dFzeF+FQDdZka
hzy3g92t4+ohXrwGxaGtur5YoqqHcEM/uMeQoekInZs/yXjbkeqAmet8yZKDeiiHfvAjCcuTvKRW
4T4P1JzxuRDpQ2MS760R/5M4D+wjf55/E13lbK1v8zuGAkNmyslWtzccZmC2lqhE/7+R2JPmrmV5
3vl6Q0YlH9tBuYWz4nfwDVq8nts+RT2nDYJws+GO5dh7nhNKlxWGg4KqZVYU1bQGe9jDbhdGWrSQ
oD6YUVGN+8Wij65ej8/n3abaWHjFYL4zFMQBqus11waWftJEpOBgZFvX1GZ4FyODcgMFX8W3YtwG
XBYrvVbSW+lQXQNXyQvsoG506PYTofxjaPhZGQPrz9uJXgW23SriffTmlK3csUjql2bUi39dtMgF
GNvruUisG9InkFsEUHZnQNELE9JXF2Wgi4opwZDBw7tJhKMQDglotZ+ti6V14uY8EqDftLjpt3uZ
08jQV8qLe6ItdvW/qbVf6It6BS92n600Z+dw1YoG3eFC7VUbqlDDFUGSSKdvXJHhczPNmuUQY8bE
VszpmPfcCGU5eigdeDeDGv5OqlX9yQSeb1Q07K0NRtDF8AOkDf80aHnNsKddK7/3zXMAMtICRhXd
TSX7a6NY23jgZqnHxyoqdQqqLvoeZYzlgrv6e3XmZUCVfOy5JjW4pJQMlY/5RXg7tkwt3pihKLH3
iLVNTNLtJ/vhzKLbUp+M18QxhF9mrOeXzaMQWN4c3cTEl/vrxjxxzQgxKOyKvVzfnOG9lTqHoKam
FD/FhaAslqkHI3Agui5b25WYozToEKukyrKKK+1WsY+HoMRRi9dtCiVOKpff7FnwjDq+oy//Iomn
TJIU5uKgCVk3L5q28lDgIUiu6nz92bWhge0JGoHEsXjI2tj81KRylUD+Pf153CJYm06NO8LTbJOj
/io7tlDOCTg1ricZrE+tbE0UhB8KZCUUD7pshZCxd4ufkrkAIYkmMJpnt3dZmAXAe9Kfz6n0r0fI
zxbRRruRkcTMvTXLgmtRAhMYt/sy8Kw+mxWxbXtl7rRoKd0JxlByhEKegNyBCJ0jb0unadMEkTF8
437Kv5qVRpaVvUDeBMM8u+bc5xaIlqEKh1L0T3XEttAGv8hm07EjUm2YoRr7Jb1oNHlT1DGGi/KF
epeWLt1v4Q9d81kk9SU8R51y+gjE0jXaKcv4y09wC5WGyyOaJsMNHOkE8IBTulz035ZZWbGcDTK/
ZyP/SCBJnUPKTYQBNGsnJPu+ozgOOanRyTFmzC7gMPuaVeK4Lvy2BWEwbKpjDX1CEdh/SsZZW+D5
1JzMO9M+ZMZ1fGg4DESueWtVfnHUOvAz1qyB48qSn1+soZ2Dr5G4RHpnKFE+kFAIMTBFgt2DEqWs
I3PfDbSKAAk75hZdBqvwPRWATUE1gu/hWafecUlcXSclNk1w1O/n0dZsCMBTADppTga/BBXsm1rs
cq84ezWvQRSo/wqTrzrSN9K6ZTiuBZJF9mWAU2SaoXA0G1Z8QIr/wrM1etzzsd3XGIMeCj+SlfMm
beTuFWRTe8+NN5iVom/Htwn0ks7YL1mndR5cUi62xJAlDF1w129msVPMFr/kNLzziVRGZFTBpWCh
DAWf1IHMiMR1QJW+GisMJe+dLMXjTydra/PeF5o/609Jf12xvzUMQe9HT0+g2DG9kvepMNwuJead
7zecfM69OaOYWlcT9m6AouKxmNVHWILOAIcPA4W5PXmJDKtjCurpch8u2bAt7j08BXYklHK/VveG
xluZ2Uq23xkX5LDd2p04aBg6DHDJmF3PYjVpEqmOr46zTGkb0VJzx+gfXcu0t4gTwtAdFQylnKZ2
art7NMHM9scGtt2r2ENrkgBbM3pcC0Utx2ngFtQUuTnca1T1yGcMu8rn4PAkAUTvIU9QuYhYaNmi
0fdGO0IwjC5zDHuA87sAGYIOeReOtVTCynzLo61kHMY3zbZBpphQNU/gS1KpUBJVpRxeW2r5wOlL
lTmUQqVpy8K7dLTo5v+ksRqRrr4qEEavfbqBtp/XwpqFg98MEjTdfSQMw6RDk17Up5NGGECT1tF7
RzQxNDVAWzAvLM8AxA08gLK6IDHBOPTHq2trJg/7/o3W1GHsai/BjjW+fob3MvffWgct5BawUZH5
X1TOwXFO8/wonIx5FxlC9eckmNPlyK2QzU/30hFeC7+uIwJqy8kb7Q/eLifiDX52PINXSJ/AV6Sf
mrQaGXBk6FrebxcfD6DLcNRO/LR1dI2wIOgxlvWb121esEfhHt6htD27l732N+q34jkTR8PJajsi
AwkzHTwujJUWDvG7JVJZdvyoYugM0yUPoZEmhovUWebrEu57g+jw2t71+G3Kt8KQY5zQLT9HH1rY
xQA4oEmClaKza56+/JDgn8xwxLeEN/W9UedEgxs8JArAX58QyaualPjpyPeI+4K+eeJGealgWIGh
1C1YdtCmNB8CENCr4X+xaoJPOy5BxtWUDfaEpB1IvCefPyXg0daLAKintOtVhAMolUH5Yx6I2AYe
p7PNTPltEN/JIEPhse368wB0N6j1hQpqSuBAGMnZQG02SzPu0QCfyqA+e/nUtObUhwNWnEEmKT9T
OP2e2IeorDj8fDFwn0w65WW7Di0b5I0Sb1OJjZPd8V/JtNhkojGRMTu2301J4W84RDXEtvw7qRLK
brVVfzDLx3tRRXhr5nY8BPlss2Gwkl3PWUTNIO8awKVTGVxUHMZY85qDdvpVM8OlumrAoDeJLKwl
zyHFzjAcYccl/gYLI7C+2nkCNiKqOPyOROrCyQ0HqYwnTMXAxEGCVkbduhKWPfFV73QmuFiTxtEi
SjofaFuwOK/tHLUiemOz4mom4ihZvqytkgXjKvnUZFae1TTbTOPCJkjCETP0VcRKEfpwahgyDjMT
8XU8VI5y5TA+OsiTbJWGLaGS2bEjNXdB3chrEgwdGLQwHnsGffCACjWFXbsWB6H04h7+U8RxD64b
Z9IyvbB6e10sXq4J8BDBToeuJsBE7COtZmNUB29Zasl9XMQOkd7qcJpmlWGq0RBwZDfxzoggSVXb
WEpETYI0TdAd28yt9Nlilnu3sYOch4o0uGVWMc1OLUENO5DosKs6I6Bk/+DZ3yyE26ZGkFyBm266
NcNzMFrX+j38QP9uT+nc0wEN019WT7/Z/5dLL+08VfldgRWahiESF+O7CLYvMzsIVpYLfvVBFb37
/J5wGT2KlhWF98UyebgGS9acyavxHZMJX9NkLq2bz66NThbJ/wHCGXo63s3FrJjoZ6x85aHkJ2f5
u/wQDWjl8W8rGdPutq6gZlzAvrMLt3T4iZ/EgF2JOG1MZKQ7wMbcZFsL+P6puE9V+736C+Qi4CQK
EmjeOKYNiYnjFOE0qH2unNozco2qmR9HsJ1iBJbaXXPSZhwqckB19MPMBCYWzitK0TEkR+qCFM3b
2dJDromkELr5SI8JCkOTZvpdKAo0X0h5dglCjdPc4imRcFIzBh2d+y9gmUPLcKBc5XJeQxu+cXM4
olseddrEpugL4qINEFN2QJdBu297dYntSDCM2njr4R7yW5enUOGQBUfaY6vbUsKFhaAEfl4Tb3yQ
J7ihO89kBTHCkHdc94Z+G9ohlSiVBbA8IHxI5zt82wVOf60VRBeA9JLnkU430Yj31Y7tsYDXE3+H
urT8Gvjcf03mxMOG3cEs4gkvvI/plMNbXsCPt1cEw+dw6yMPn/eTQwGSP0fm8hD+7po5IqrMuZWh
JgpKcmlP0Wd3aqKyu1uuH1y0TjTaEUHTCVHsMc5HgOY+fhGluXKDK8xKwzWo/qDoPXb+zZ+AvPIn
fa/I7+yPNycYggge08Bgr1fgOYv6et3IUZDOehRbVvopz8iJ+ehNVmPxy5Im3Q1Mvh6k3hoohDbO
vnYqoOdXNJ3pTGAGtdtMFemFDirzbkwepYC5WmGiOVpzocR6h39DBjt+Zhx4TaRFJ0femmc0LYtA
1Y+ghC6lK6Ztt+Wh2dLVvamhFXkdRvYaQSzuXQPop53gqxezBkxApLKlqdRP7GexJIDGKQ70BKZf
0Hbf1UDe8EzPhMiPOExSyXc1Fjydpiirnm5JUogrzHkzKSLI4lCU39qjSRBrpNVdg4ThCydzK5nx
gJbt7Skrgh/ubW1kmuUh899tkAeDl9ptPJOvUPzGxQGsm4FUSFoJORKnK8bGq/FzDxF7n7CoOwD/
g/3XKoLsiTtckjdoVG1gnGRFynfXR7Rzw3ffiIm4+aRHr5qstgwl22DUh9kgmbGGDsWVsXbhD1Vg
3fbTCErz1NOdGHqxk+z1dbMovxwxXX1YdgN6+QqAKlsuPJJ2DRiObn3hzRAdG+TygwONO6Dp3dyf
K2WH94ABfA0r1RK0MtkjanEoHWr2OOq3f145e0FdKuaN2B7SmYfHiqWpqXha09osrkaWJC4iFfzS
EzjVJYl2JhveDehqv7HTxT2b90PVnFc4KrFmPNh5Jl3CN9zVpsPcgoFIqymjtpGBgroftB4NMHWe
gktX6Y40tzDCI5pWxPBQ0et0xbREybdjH4AfSL6JLCsSlmCW7X9YRehu8K/MqM0qSRQQWC6gX/5u
L9xkW2wan2Ar/bQl0uBDP+ZYFndVM2cSv/94aPG5JWFGBp0Ts8Rx5BI7Nf7Oh8Quu8xgol+ZbWRu
rmqHlZsuURV77bAF9++Op377YA197MFQt9u1qvftv0d2fsAJsPoVRxZhdbwh4DtCbWyTSD957sI8
dkTHplQBM9cyqhONQ9sP3GirsQWfjcKX4RdmguHlowg6Jbpd0WzKeEPxZQDX6pG/IvfkR3xpf93N
yWFJOGChydSWm4hRthXS4tkkf7ksNeTay3m4CwF0iwgyWl4Xv27DfcLyn5fTIOeD0i2TGMnnhMEe
oXxP/9LHJB5PxzjiiK9DEfze8TtRfPi9wk0h2XkYvE25NFJzVyXforlz5LJOf7YVEuskDZjro92c
0l6MyHYNgfw/6stOY91ucJDQBhoKpNYYumvtvnrW9bZi9eojgQtbdqm5ES1dsjpfgw1oD0ckxjIa
QeUxjflrISwcb/LXYid7hxwvHPLdlUb8f5wjWtEIxn4a/sHUoygI309sKM4SgR6KXjEdLFO6lQ1l
jq0MN3HkU/nC0LSRpEkZmWX4srnN+vd235ZnhKhWVU2PEQ3GcQxdOguISh9aJ6Rp0QyQfh81K3di
BPiueuRAUKhm5TeLukyVo+IH9oh0zgAsR3e8kr2ixD/5d62TqsekmvKBEoF20YzZraIQq1Pr/kEl
ZfXD6dZAqfPOo4ui+MyOlwUiWETPid/3tkpskcy1bymwridhzPbit052RJUQoKWJEtkITtiG7D5A
IozeyRS0XYEHBGVEa3TyGqeWjhT2yMU8a4IDqoMvXtm1idN/9rBXpmSYVWSEBV4I8QQRZGgcr2FX
c5y8qDG0PkEk0/5v4zlSjcRaualsG31i4S34UToHb9Pm0vPsG/7Q1KZrS0GP453XaBC8nsUlZ9Vr
yv50r79SNNAcy2whD+I90OKgnJWtJUsfWke2b41ZFggt6K6S49G6p07M/sR1bZ7Q/+UezbmqyLEA
e1xRHWLqq6eKo/8SwxdSKiRCyzxkACB3nUlOsQaLu8JTyGycxtraHENt6DEWyBN/0ZxSVJGxcJ3M
wPTJq21cdiZHC393gk5ZqHsHxzNK013nWxCN2X+q1H521yTbLNho6DL5RJiLNjv02TYZnSuCUTFR
zFgD7LxtHU8+gWAJMRh9O3kjlsk9krVRKIRh8BXpdpTY7S2a5CJjl/q1e54D/2u3Q3CpPnfSP2ed
3r3O/OVQiYQTu/TqO6N8XgCrIrLdDwKyN3UmXIONcaz+dh0Kgkv1toYUyEh4GYo9TcPhmFM0HSkg
vwEtU4+bwpr6L8i0FlHEjMxnaTQ7s0SGIoumv6V6NLsZVsFikaErMAf2Q6DPQm7JKTJj2wgCrTng
EzJTv5tdbqecVobr+0zQjlfpS0DDPHk9glqdbLlsB0g9PsTR52obFijRSh3BcOLLbnPA3NlCNy/w
Q65nTL0uryDM+zfu+CdCOP8j7k0b1sVgB5RP+1qUNjItLe6W2fX7y2l55WVlMOGS2MHbKFyc6ZaP
tXcyZk4jd1mePtpy4IW56Kdp9uhiEwpEMZrmNpbNz9DIXE3wmg2SNDq9GmCk7iYm0woPsR82r01L
0+mNpJEEhVpFDbTz1G3QEdQzbAETJEgXMhh3gH+rcDjzkencMMf2KjVvYPYbs6PAz2FPsNRa0Sgy
ik74jQiqejSoSR5MzZ6KtdLtfTOT6/jRrCE9ghiMxtzFYMC6vrFo+dlbMEa1oL8E1DJTa9FcE8OZ
AoB+rrPGktrR5QF3AAc124ywZqZhk3dOFunv5s2kMZknShNpfQTTX9kCaUm9EJNHiCrVXsV0QR1U
uP6pF6bMsq9AsY8UGqs7rOJeZKB5NJGsP1/vIT2bvVtrturCRXeBxuCDJ4dCA01pObvQD2BtXK/l
aytoDXax8l2s+k5g8fJ5dschqvJ4s1Pu1vS/B3hZulE0q1rONq6WjMSifA+o96CkQkOeI7Egarpu
b7Y0fB/j9a7WDlq3fmk7VZqGuzZphxNhz6ZlOf6D0+3YzfA4EKkNdLuRX0aN6VBpGlsXQSPxIwXw
AkZePyjWZj/Y7GJxxfIff4LU8Z58T2DLjngvNhwcMTRhUiVuN8m6tlA4tnx3AqDi1DdmSYe9Bkde
McRraTEWzzC/rZrRtUNbRj6oX7He8iZSkehxRIKk5hVuRLNvfF2F6tJfG0YamtNI5q4g/HYiMZ5i
uF3aXZJMxDNnso9Jh1eHlpuS3UoIqJS276xm50BZw+REZ/wbvmw0JRq1tqfZGErOoGRzhtsc57C9
LWT/nAJFfREGw++jFvXNpPPCfc/ME+wMxh4LRL21DYHFgor3XTevAjvrRzAUF02E74x2BpBmxqOK
2ZGdHSXVr8pDLjEmnuPkSHxRvtNI6HiTrTEUhqU6nAEQJ9qGmwtc/4YYr/N0hcpeBzkVXkahaax6
UIki7g7E1VylyPfZWEPvN3EHkSy86CjjyokEVnWNP4Kb5uzNHlj+5JPgBywZuxTEGouYNYm7nZfp
Seq0gFrhTIn6lHviBXiB6JYMax3IyV25GsDj/PUbYEy+wLqYFWXEuYRrHYSuWbxI5ah992lgC4fu
A98ogmO3DuvQFAyDru1G29VUtntPDijQriJ7LIJD7avcrp2HnvhHGSZgcSDU9O5nhmHACYODRZJD
0Yu+s27nTHGBmTfz04n2yMRQCGYCPdgQojXH7qNi1zzNHz7ibQyOd44Q2gQfQakEIZklDnQ91cXf
GnxFlp4wyekTYFGKpa3ExEXh8d+IvP8GHiLwNFr28AbdUXbmXwmYV7gfmrmfsaoktQ1UT3P+jSoY
xSw8PhQt0fVbnaUKS7RFZQ+dH4zoryvphEpBhBc7gbcZ/UcqlWyq0ksJCAux4kqrzWAIn7DwHUkB
V6kGtL/gd73wOL4kB40ZTYl60x4L7UlgQZIxndLBjSHn+H+wp3iU0Hz6Bu+OldB90us2aqIwe8Bq
lG3BqrfoUWTdewLg2SrP/EoVJdfB0QqeUDA3igTl5m/Qm7Q61AP10g9lKfk30WCR0cnePItBkSVk
iTo7vR6uuYO7BHLLbxuhKEt2R2+CYjBAxUu5Jq25KvJ9uOigGBTbQpBJKs4+JF7dVsdzMEvR/7os
Mwdu/QPqy/tt5xBBRm1c9Umvp9yywGn+q0+Ys6iN2a4CcNWSxogP3Ene8v8LeNSH0c8bPacjh7a1
5VnKcg6QTLKNLiKPdpdTXLy99f6VdEm7T773CAXb86QGXiNc7F68CoZ2R1ilFd4aMRr3joOm2DK6
ikYfa634Cwxy38aQ6rdKNzYokoxqTWS4hNKFBQ/4t6kopiCLePZTiHn0XRfDK11jL9muQeRN+Crl
42zPrriUAhoXMrcYa2OXZM7geOuGAQPqnyxSHtRz38QY6eXVbiRsn0ZxYd0VjEXtWjhmNW7xykhr
PZGKBwiX15x2PmQ67QO4oU/DtzLeLJNoVT+SAxY7n6v4qNCDLjHBJiyICwjP2T0og+NTWZncP+p5
VsZ35dMJp3yeQ+8HkD/g+WUjT+LAgvtS/R183OxsoP7PdPHFzz7X79mMmcO5nr+SrrtdvWbzTwZV
jxw8u6oFCxx1Q7v8JsAXAG9iqFM8CM0GrR+6wMExaLEjuEZw4daI+tvNCUB0WCPU3FMa64QgbdF+
qet5yfWl5uUJt4v29fpV2O9UtiiotxmM0v5c2WLO74ynEHdixE0ULdhhiR694q0chVKB8rwTeGdZ
GF00+VUpYJf+cSjSjZ5GLmF0748Cs8lIOdNeMUNT7VZPCW5pxZjQcYe1vL/xiKhAGr4/cNPud+8S
zYBYUCwaAoHVlDxQ5b++3dERcNz3s/7RFWBE/48gLSLbujQOqs3V8BMhEG8y/AzvFvcBovn0R0ev
K07yDvi4djWqY9fAifIcU94NvsaPAYAWaLFZO3ikW25elBvXjzKN+az0tKnTUu9YOAIRIC51xGeA
tC5KqVDYmSigw+1JMpTWxzrB6vAiRw7ysgbs5mHnQ8WumDSloc6sERhNanUFMLNtbf4ZEqGIwotx
bZP2lhY+3g9Yy6ahUQbVzQrBRctB7lowzl1n72JoEc4JUtmkeSsazhE8J1kiqgr6iBtEDaHkDIkL
/vPbgdc9FW9L9PMYHlYkzdWPCbTNr0qA7AZufJgbAaSFWZdQuu35QORjiyV1WfhXnL9QZBA9tKr1
kT7dLVi5CxDakya7kArrUUVaGCqb8zm+fjGZUAICBDULXLOKIfXvSZR97k/IJ1WY7IPvbI6VyeUX
AkiaQPAU5mIN98mhX0ZOYkwJAHwpJsA4Y9Sf4DxwC5NF7h39l4TQLzwXdpUJN5hoacnnFC+RZyhl
UkoQ7aQGL3UDjCutUlq5BB2PqmHq7xkGgbep9o5Cf24JbMEq1dctkhq+OgYbC7CLAb21gDhVt3kD
l3XboxZqTpn7wOkx3z1lolAwcDNnIwY0fZI0crg2mZcRZSWYoRf5u7iM5cVlXR/mRabhGVHYbkUx
hgxEtyHOi6aTQJ0ECbkgExwmCij803MG61iAR2RcxjxdS6Cf3Rf/a+xFPOlFlDGUEL74t0YajAiI
KWgZPGwILkLFsATnnD8Xc9x/fN1oab09WHyi8L66BanCo9xRmo1ZzwCd/QSuG9XWK4s3B/k9l6s0
yNc0VE9nYv+/raJnVVL+Kp7E2atcWMqjf8r6BW464BaSa885HHJ/jvtYsiGjoCMDYMtZYmIAg5UQ
RhpYGBXTsEOq3VoInAnXu5mu/SZ9gnYuGbLl1boqV7RN4vBk/KzWAs/+gfDZxmeXvd8eRpWpkkP1
xGJyoFPsS8CkLJ5apUFYCiEhKeA5GPJcU59cbL0Xjzo+VCnYljNpcT5q8bNqlw2nyQjEQGHx/mLh
fY17o3OmvFK9pfNBzxOIAgAWWbBGCLJQBhYiWwraxFmOHBa99ZAB5Z0g6qmvtMstzQg5C+ZZng/C
jjmcPYW9B2D79fOuBA6GzXKSPlMlXt+tCqCKCpC1qol/zUqmcZbxG4NgYeh54C9ebd9+arLYn9/h
1NgdOHQK4l45F7oF9GCt670TlmLq462hn0b/aKLPOTx+g4oJ+57O10PKTiUqmcVLR41gYl73Bu1Q
znkqZE8MDBKmi6xCmQtt2+IE9l4lrYdEXIwBISZclJZs9tCINMZGAmLiu2jA5CaUqJqjheJPJ9wP
QZbF8AGoGU8knjEBhZ71t1dBGIJMzxRVy3WsI5zq9exDOdzvKSaMPDbYnCV9TAOx7Uz0Pz5cv+YK
sGYii3X8FASqO7aBdXiXWjRJoRj87OMc2v+3LZy5Ub9hBFucaC6bpFDvE0Q6UIGKk1MXzC78KsNT
x6AvWZzlM77qbDHiqHfeyr+V5Qf6t94D2bbTxS+6jlKHlj7Aq+ObVcpzqAIuVPLjRergiIMFD8An
p/4IQPAiv43aPXpGd5k3yr97fHBcqhv9HlXXysEb3A/Bu1XY+qaQ3ArUI128XtxtlqAkiAPIfebT
5rpVVB3dIGzQrCrjuzfklAcggEe69FCtixVFtFgNzeORE4GM/BmiQVHzr2BuBx19ggOROaJCIf9b
snJrbvakYqLAV7sha5Yr4QJ3TPB9fY76gIjzn/SHC9+A7Ap3A+bD1mlkmSWsprJ647UioT1rEnyz
Un7OYhlibwYQ0ZlI6oas3+dJfeP8VMrsDadf80hhlU3pewp50Elo0fxv1Aedrz/sGB/YTJ3/ZYPY
fAgxjwu/wbIhny3+eYttw9WgH3Q+RdURtItNrdrBfSF1FKHcnZD4KdqKJXViXJ4gDstLOi2iFx5f
faDdidZ8eH45WFq1jg8NopxYkhpHi28d/eGt8LH8hoMT8XHVAsvYr3Ko/pl2vrZ+5IuuoX14bi3H
S+Y/LnBvewPr+CgQIFDlVUbU4Q8U6mCFWLtYOmE3+htRxG3BaCHowQxhyKGxMxlzYWYB0cN+Kx7X
61k0wAKLJsWLjFl9mgIAYTYzCr5Kw5u69q3q6Absn3a+7vqLKwj6EJE9xgrqKev1KyuzUPlkNKf6
jXNPXRg4KjQwI81QgCOFSW5BH8OFJvDSsxNcSn/gLFbDu3j+g2itPGt5QupKcfoWSYmRSJsWrMEl
xvWLQkV8xUbo3NQRx6kKnsZ2gs7+r8RK3R6LirPKZTc5ss42pLarIgNF7UfmrZINEr6uSg6E6R85
RZ3BPUEtZuhSKcsKvo3olqpROqZGy1Ts1uDkq+X9thQ0iCoVMkEEV2mjGHX3Tlw0XYsk6f6KdeDZ
2kTutxnEnF9cS45sFbrViGkMZALY5glVgp0+07Hlao+UoEKE3xybXiIo2sb6D8JZBQmqR+JqxQ8n
I4QD0dy/FKS4/De6lCUq0zxz8M4u7qBLuFBv0Ay9NHvwC1wj4QK5skMbTAEfL4UvBfFp2nuZd+l2
ppkhXq3cytf+1MNDG4cJIm7Ehiv3SiaQC5CP+Vfgf1Y3A8GAtF/Pr08XFH8XD/5kZG5lOG5Z+QXY
RBoAL2Yf659bhPUELEcXmSQtNMRC1P4iQEouIJl/7crBz2hxGL/fLAKMYXbae3T1wZmpXnRdseEb
o5lyhvBmndDDV8Vu/bqvgxoGv/UQv00ER5U1HcwsFbGrZUqxb1mZQcl3MhsoXEHVOxRqVFfnFd2b
C3Jewuuf2CR2NFpLji/Nb75BEFzYulFNH3WNv3r6aBSF/wxu8kADczjNwwtv7IuvVmmSHvwqfull
1U+EljBeB/a15DvP2hxANnRqShgiPiHvZAcjHX0oqe6cv0FJn+F/tsNBJB9oVGu3kXMq+ftjfMky
hsnOr4god6+hnozrQt7JiJwE45/FWpwyrN7AC8Bb898W4SjR1f54228TVmNUhQFvZB/GrWZM9obQ
qMoXYHbx4j9ApR9d1xK9pFDNXOhKlqscE38l4FLQsAGoZeRVQVItRJZjIUejf3mbroJmVL768mk6
NJ2LWsSGR1n4KLo3Oqa9RTWocJ8/FBne2XF6G1gxxYMPe7Lh0rxfPNECyDnrlmQYgPaEclwqBerb
wzE5bTpL+psAsp7jgLnzHhbdCOZMgQjBf1niZoISo0hpLYIueq9cHfldOWRiuHYDjyLl4qALG8F9
ZZeipQfnIdz2sR/Ap//ayvTezZ4FMtwKv0qKy4c4jNE1lHSFktXRPPpZS+3PcXwtclEaU2A4O9LU
BJSqptTmht3vlxOs6QoqozVzQ5m9qDRapzwG9eDL2dyZMXIhfYczD30W23w1JFsEboOg6XC6H9xI
rNT3qdQV2I2qco3pSsKtsNCmzqyNaKAebBQnbIkh4v5sjNc9O3EdmLFsUtu8T6/G4lZI6OOi4whU
abxDcA9PhCpUsQmb/NqCM3TYyT+HWSEqkCHVw2ZmHTrah9daZxJH4phHIOQv5OqTyossG98d8bJo
NX1492IJFC6NYrWvWn19xkdQq/b2GA6DgD4LreMrNW8S205ZLw2jI/sS0yLc53NDtV/hw7EMytw4
9bDrt2Kw/5ii365nRWicnmHFObUEDfFWmx/5pmQHr9rRZmgPYssMHNwSUuU9SxioSpZCRRxml2cZ
smQTm1bLtA4p1rDTS10iF5zqdYns3v68eX6691sN57LEReSY7vZ1RFa8PjFAjSWKl30XcCnXdolN
sHdYFJD8V3rdsg5iSmYCI9Sy1e9bf+cMMOdngrXl5SUH4X0P1//a8CKUb9wxRYE9Z6sATUXp0yD/
WqGGSuE1OO0WAviT+5wh6Su9gUrHuzgEA164Y1OCkAu7KBpeum56IYr/889hubd48XSBKbJ7K567
YEDTQY4i1fQeH/o6aPFMFb6Om5DBWmdcmQ6Oz/ikrGIO3SxBPG225N3unyxaj0O8BBXqibWKH8Zb
dTs0HDltrOveb9UbabFSb+A2z6fO0ES4YQ3pU3DXcgD/PSIVBJfiuX2EyXfUakLg3DiD2dL8IRPq
XhNo7oofHiC37zNkBbyE97sG9GmOxswrgOAdCmoEXYf+F+6KtVsZuMBvdRU+YD4QmXNOo7XWLiaw
ZDTV4aGcd3FJUn+3qCaB0/7VqfOHsAPSwaOgO4gpUNYdllutaQE8hNNWFcU+BQaUUBLbk+l8GHw/
S+F74t8gKp+GmP0E02Y37ppFgD01Z8f+4sjVo2RLp+/CfrH0aB7wSqnIA4jTEFuK+6FcmDK88Xdl
ZIvsXluD+dYomzsYYcwgokD8sH9S4Ts137NE0tft/9gyEj4UZr7DWVcDn5r0egt7kfLk1UYaZdvN
W/sMAXLM4dqXtE7vP8wWL3hkyC/gdUQuHzty/EZtZu60M2ftLAWfNSFiIqBTxWb7RotfMW9o6Qso
9LnqzFq6b1LiGy5aMzajzcF2n9Zka6QmQwvp4SdrHjm8hhqz0WQuFkv2gFUAeJpNIGREsau6Tcud
S4AgL8lLMRpGoGjrV7fSZWrUw3BtLv+CeNEEDuwJG7knTQZN9eqSnk645a7HsA1rBmyjg3mBCeAo
On00WiJVfLScLn/VaiP2mxWSrsw+dXXyeQNqT/vEI6Aef9Og4U6UVXS5lIZGM/2e9/n/rs2RFU0s
zxnNhKbYmhUu6qwsyvBqqd64VqFcsshDNrD5DsXSs5efDvKuKHfWeEqh5m+ih+ymSyeltQplJayz
UPHGhpqgJDHj4IW9061fbRVNeAua8B9WbYneaYFtjHmlxp65BjnArulFrCX4E9Ou5wg+PYqjx6l0
5uVZO6+X9XwP72kYPHag9OUJE9oY9QuA/z6x/Z0etz4UQI/9bDtGQkzei3o/l5KgRXmhQMO1iAc2
EaZ6+O+YNM/o1TPXcLx1qR86c6zExdvsAUZhiJr05Im5DI/LaKeay2VNJSFK87SyO7hyKTnnNSBC
yZOe+FC6O5lYsZ783vF8lGFUsSbLcMvbXVDWyOqhYjjgqpLrOwmncOy0Gj0LxJT2I1W5uX/WqgSo
bmQYyZsdto/Qw3NVZlfCizvM4kh0grydvhrxyPZLMfk+bhjgGEYLI+qtyxzy3I0XVhWw1RbfMnqm
0ive2ydz0OAsHECLBPuVOAI/8V6tEKhL1DlgTpuDwsGcepLKLauQrnuiBrj45ailFCxpyBm8sNbY
9u/3ZyZBWqdhR8h3zE8p5dJVk2UoCKT6sBFFws13vkK7bM/WpVavWEmoTVLCwZy4Hw56GLw8dDHD
AlvLO6wvzukzXPz+KwVbxdD4wf8ZXY9Y8o3HNAXN1naBEeiQycLPCOYcnKEdZi77PlZvuXHvNP/h
1FZ+MMeCvpNv9xsoMBhQCWtgE8qhOK1fap6/RoGyXWbMg6k8e5BGJqLbVHzWx/Ku6JEmpL7p6aEw
DlZNMMzK/tFN3BpZ9jIuB6D5V3efG/pDMCsSfNhsv6OzynV9YxIpnKcTGWNLSj4IAZXKKQAByk/Y
XX0NGhb2v1NSXyaa8RvykXvWxQZQRkdq8YNR4SF3NFmkRchx5bqG6g+SW/rC8iqfoiQ6cWrhPIvp
Us4U/Jyvs7zQbcq/Hp6grTP09sQpyCp5m8xiW+91a/LWOjwo7JkBHgio4+riBRNRxlXoDh0GosdF
njrW7jJmdPyjV3QftlOPnserGjkhTw32r2fM9q0vhQ63WfSqohdVZTmFuymis1S+uZIUFdwTF+Tg
vu7btOxge75XhkHdzzDkDEcxurAfUuy6GIz6gfHoX5oiKW/TwEJmDqeQ/o3ln27N6Rz0dQ2wfhf1
GuSlGMrbY2TRtzk7TmAoySjbn4kSLLvQVT8SXRgO3ypKLOsQpNYCGEageCRVFb14o6v9GmItTmyk
CUJKmcI8FPTVeBjyA13hrRaEe79bW33w4PC+sCu+0JqYtLHhMnUM5YiGQQA2Nmok6Nt/+2k659lF
+YpagcN+JT/9H4A4PixpXJTpk6ndwdKLZSQ18S3MRxV967FzYXejj0cSyic1KqC7pLxELP2jfMHR
0FtcAHiH/kC153pL7KzzmKtjFkU+PmJ1kCt1ps3sWO07b5l5s8DOG3wJxXEQT7mojr/whyMyHY7F
TuSfUCdvBDltkyB2WppNTY1MgBgRC78fCMnRxERtV06WsXt6eKn3jdyQXDW255PuavF8jn80IFhQ
it0WUoCSBjfW7Kir6fxdR4Ta1PpJ0V3V4vc1gbkFrcCfMnd3OyCwyUYo8nfpTsvSDN/OMTVqJSwY
LfIo+vOuVAhjpwr9REsr0SAVl3DEgoO2XCWZxCHDVJQga7LNcomim4YHGCo2pqj5tZXgZ7RpfVh8
UvAoTpuffxXVxdjguyV72biCcBVWbTfJQtkCYttIdtzyz5DW7+U2WqocDcINvFYPTDAM3bxNNnTa
LSrO22dxh/oVo2SnLWSP7QquLbJ868K3k4T7lmbLHOOGy7lcNWOnIXfzBn2orwH/7lqwx+pnPC8m
farf/Md2fFuSv8BnGzi/WGhDkUnqDvWucKuH1Gy31nP9CTYuwV5EJKRmcTObwn3soOE4dAOodO5z
L85nLAcxuMmA7jzxehA+xh6h2G6jPs4xjcegD0HXLJQ65R/Rph614AMqlBGcL0LD0o4WbnAJT18Y
kteKC27Dp4VkClwkQkWyVyIVOYaBsn/ueXTE0YoqHvWQNdbkD70I+1w4VXF8jWY4cSBQdb96+/Q8
8Sy9h8v5ZX5WIxie5W2okcqiuCNNtFP0J05hqPSQgGscsjbVZcjnUqjSn5M1kLsDN50rwZzlHI+c
JmyNWJu8k88B8yD6KVxW0PicxHUhrLwLEpjvCN1I2Z+YjPV8DB3FSP29bH14bGoFZ/H4dVmgdo57
F8n66IMIhYmVJLF8bUwW7Zsc8X338AcUQ+4OxwoUn4qVVwJUHQ7bleQW8Xp5L5mGNUCcKctf1r/P
/s7dY5NvPSqC+t6P4OeZdLzSYLoqOx45Ko09xKC+YO2fp1dey0eIGuRgHThtlFnf7PdBP8Arhn7Y
8jLXCUbqRQcXVA8jWqcoJ5VvMtlcWiitBeJO0nWBk67V2PBO+4ZhRn9TXf71krmfREiyfUGwIZt8
LYryYPj/tkC9p2NG04v/jksu1ZW1lwXwDgiGfXCumEmIYQSktwaSCNZP7KJfMypmATmaYlK7oyH8
QEFjdwyAiWSa/uRcn3L5X65C69ohjM6wXMDIB67isr19Ip/7m22dfYy23l23HozLSKASyJ1Y1IeE
v/kq16WkfJs/GPNYU03SoyRuBrS7giiZSz3D8cNlxzkRQM1evaks2Sq1rMbcU4GrZg75NJp0RJg6
oDuPyZ5DEX2WUPME2i0IOk/ohFgGxC5TTEsS7Q1xHsS1aNFreWH6guz+nW15x3fz89o07AgjsLVA
bnkRSb3dNhcbrpbspb1iYU1nKAeXLk/sQZT9o9lJPM+1f1mXoMRSi8ZM5y/3OSKKNWGRQQB4GAeR
BcAFER6AGdP9w6HShFcSquLMfL2cvKL0JYNOlZjFfCGcQwIVSDfHE6gP4+dgFWvpSRj05RhrXg/t
fLpZaLtTp+/lsPfKoz69zlIAP7lz59ty8TwThsT8K0/JRhqNOTOInZBMXnxxa5ZUiiwcS1TAxhUU
Ln8K3ad7cEzL0272pQYBX5Ef7xzBM2ffHaD3bsdXiMg0e8Lzy+UhB0TtW3vEiKO1NYSIYTx1hZ+j
TMjDNjUF66+CO6O+UnARq3B1zujUq2BjRLECZiFPSub+egST3FgLSgx/ZXpq6eUd3GYuovNLVVC/
7FbPU7Leq4vB7tg477OFBa7V7hwJT47cQxEwzrEIL08obNVcnhpuSFTlLTYTgVsliVufbMulESKp
x+RqrrylUHZCQ4D8X9dE0Ajxy/l0jFUcHlBKsf205CHPF8zbE6QYUc2Yq6DiwTvPdz6Hi7iIAx1j
xZllxPpVG8sptB2Qmx39Dbrj9zrz/u/0EPCprvuGKos7yzm9EgjSa+c6LoZK9FtcgaV6KJSt2UsD
AHtbI48QDFVT9rscvK8bbK2S1AvsfyjBzvu8Tjr34O1s4FeemRs5EQfks5g3KhC8oGEvTD1slhAG
9EwG6GTtVm+pyWfOacLMOiIDZdtNE8lCT/KkTIdyr59GjKP+eJDjjBagGwssqERJ/6t2yPYDTqCn
H2nXjdc3FHfnioHBEWNAEKfcjXdljUvXmKz8YshYwbWZ4JFiNOxil57DgVQpShZWjF6YeIglwv4S
/5EkJ/Efb3LBgeTP4+3lL5xaJZm+NWyEV7KMq1kQGfMX80gVQDqoQbwi5ES/KsuEMVefsyC9FfQa
DxHFatnDXsob3jyxH4SfFCMjLxIU9rEOxFRp9BgFwm14xH/wX9DWjpQWfaPfLT2eEg6GvoP1yUUH
FbtMm9WbaQYtileOCH8YQgoTcKfZfd3Mcb8lyvOoVwl5+DcEwN1iOaLzap66hpfuoVW5ozKluJbX
/BvelJU1Imk+fc0gzdN1t6kXHeKI3CIfacEMx1StZwO4eyZFQ8aH6CM2MhBV2bz/OxtYjE7OiFz1
SdveXs202H8j5QSG3d65geaWAhfb/rJ6aTNtYDKXSf20DPdozdAjmsWo4ylcHmb3HyWnRbP7hwrg
+u/fNCzFvBXG/XkY6f+SCZjllPbUIkqOaPj/4DuIWNp2tRM2FkvLlgZ2aeb1LKDzXdSvKuyqt/qA
+0FXytVXe8vesAKZiPG76vnmIG7Tk6+boCNI4NVvhi2QBZDFUbVqONgrNWc66RDwp8l21+ABrmrN
09Cyp7qO2XelbkDuwT3G3z0l068xjgI+kd8Bk+YyQbt/hE5ad+flEo3pYBean/n8P9qOwjfkvd7I
xEK5x7w1sGKuoN8CBVeITuJdg3LRe79sjsQ0Bqp7NK12jlujmmzN2AT0yDLArH0FH4yiO3tSu1Lw
KYU4+YqUtAVIVvL6KwVgf9tsXIzNOdAc0qx5MUYiEUA+1HqGuJwfgK3G1o9u/Ml2aFOPouNTC15u
cftRd/zyBQg9sRjomNQnrqKFT00WRcaik1L2cQIAiCEBy1OZG1KjeH7P7lG0zLnsQvvZmVnJSYwo
gLhWIJPm/heol7VsV436v7o1t4EnyQiR/4vlQTjEsu/XvJjDuETGfrfmjq4F84NfWLjpkjpdZQ2u
GlKjiAcnSbV+w4i85PDOCA2nN3XlKzV8DmOpONXEDjlMVjsN4NWHKi1X6Wngg+T7kS4LHQPzRkI+
3wX6Ksjynd1kZSTP6jkPVvTqVMV1sWmgLZ+SEvqXOJnCDT7Ix+UiXXdGXfp0/RVbeVAN5O+YLanQ
5uTDiuQQ/2vcABmmX/djzEQnddnaswlfMXw7mvt8wqa4Cn+wq6uXGawVEluHKsZfuo5r8/11V9+N
z7oPUJP5YiSA5MijARIqSgVg506zlYNpl4CuRXlvVve69QTyjO/58Meghf2Wm+99HLlsPT4TaNiV
419TVx0l2anN4FkWtfNaE29+GwP/bTYXv5aZNsv12dXR4JFSNZLqijSs9dHtDBOTTwzYdSuvoWPK
6prWJcyYqoDbRe1T2TrgBY0R3aqc5Cytu6SVmYnSjQKr8M08BGusg7EltD4WZDNvm0OQgRnzEUyZ
6kU1iqnzOSoEA8hsKtuNUXLOolQJFuyG99+zCQkXxWmBgZXSyD24ta3rJC1tWM/53BvO1NPvK7Zq
4ML8z4fjV64iU72ebby3BLZm5XKKmg1IutSbGa8WNtMBWhatogOfLd9h4whcSgYdRueLJFiBWB8h
I8Fn3mdz2GaZcMVlAcGAmLM7gXebjxGnXvFduAJD+nglKfx08UDoGOuqNk701hzdhju+m9vsd68x
ogV3u663ks+FFWqyvrgDuT455u7AoVV8IgVjLGYK9qWbyLxGG/48pkRrlxGOaegfs2bY0B3bUV3b
YgixugA658Ot1he9sUBFR8P/OB+Jl9OM6F5OZNflqpiTbNAxiPFIo1LWlS2Vs5gUb42NV0Kz1+Bo
Ldij1VEcfmm+oBpgIXJEqEFEq6Gk81umA22GrGbYIfTWnwavna42l8LUc+9ynPU60p1CDLi/b3aW
IB0eHSq6WHHuzBq1aOKmsWOMxeFJoHK7apoR4QEzp6vT4VwaxxWN4b4vL6tN0OuhO1xkY8D/2ju3
xBiexmXMiXqmj5x6z58PErTK+dSkVPHXRnngF5V8Wy+pr4jv62xwH1kKy9SoitjuqS5+thqlEBFY
NzwPbiVX+dZ4hSzSk9hzN5TIyENqjSH1GMedQlcSvSpZdUq/4D8iMGPl/xp2OXA0AS4gLrjZWP9m
VNOrSpLIZhiNbjEm/rwCUpC5J490rJqeqFDoKyUWIYNmUYg7Qi4vetTK8Vz72fAPcjwgd/mERjhE
M4VFkD5jN1KfSx9Ye+hCAVb1Bb/xP3+vTB1q/Rmdzg3P+m1JxriKcq7Loz9gOEC5XXz9iKvMLXgN
Di41OUnX6HqG1v7NTthnYaC/+ygzNKZiQqXuklBCFbTC9berN8UY8SxYh26NqxGW6DnH8K8fNxLE
wdufjcctfQwQPMMozppTeAe4NE3jIq8XE+lkmRPlGiOI2WUeGhbpQeAJc0w0oLpTNu/LiA/GULmk
ZH8Q91JZbLBzzNWihAgBYHcixiar2wY99l32mfJg3NPiWRaZEUKvfoeO5EH9amCxuzhuCtuVSIY4
5KzRYyow5KR0lpUuRZQHlxlQeCU8pkbe1nFv/EJq4JciIBYHVV4r3DaPwgVEoWB9eWaUGho/GSph
4RlidwNDmMQESSUIu2ImXXn2j0ygHq+qgNQTISpnn5OLClGvRWP500gJSOULDxZAdHrJImeYBJYL
O+8biRYdfy9OBZo3+B8iTlI1eBVgUhy861gNCF9h9PDSU1/2vUIYkMqD2bM3HKfjDrQg3gzAl769
88l3rof2C6qmYdGIrjNzdvEQcH8rJajwwArIf3ITe2dN4c8dC2alYwNQEQpcqI55Z4Y/GoknYK4r
h6cOIUUBgML5gF82R8L4j5hyCRJFsvtNfsSGv77aiagxtzTVV4sp52fi6WX2kazBW+EPkJSKR5y4
5L7gPLdt+HgFhSMCT1ANClCY1xDHE2eKcT1QFSxZV8jSUL3hFJ82mgDGW2heqfTEy4utYI+LcXgF
mK8GHVhD9bxAfcbckYQbAunOmVJbmVqVfWQ/JRfblh6j+/S5xNoGyEoae06aEMgMFqHy4nItDsfr
K9aUWQ8QS5Suvh1/xCj6q1woqLo/NLxjqNjakz6m58NlCtRvheRv3hzI8U/tP9bWoYFSWEXB4Dti
ZX1hlk49LH0xZjvS2UbprYltHGncYtFmvF3Y6U4Ow5OZT9XNM//yPPuzEkCveG2Qls4pkTsLy2F+
OCd7bvVsNTMtgvPghU4h0m2Hiz0jf0ADizBmEDckXFGHKLtGNyWE3YFMDhRSjcMTvYZ4ubUS4/f1
tT0nkrP3ljlKdglwE0mOshwEWQ9AlT1AF6l2hnP5538LxqMJsoXf3SdAnlr2SVC4Dx2yWmZkSM8j
B7ORbQAp3nGwq0lCtmh5SCdOqOfiV8v6a8/sNy8RuaySEKNlDYlgO9fdRz0peSQA8Ty1pqaQ+CgP
uRnONMmxpvr8Buo2R1Wq97r/l7va0tKUp9lS51/DJTNT/W0X/9b6cA06PwX4CxWMfHkd2irufzDR
Mjd6q9EIE0FsYY/5Nd61BaKTDmJNuhN45iWkhwROkF9FMfC2wUodXbS6DZ/R+KexzLpp8v9Q4krL
euB87VTJlpn3TOihfBd/PxHh6285d8SeOv5zqfOiB0uPtcJs2JHA9PHTsdg1d1ExYxiQcr8/qvjf
YMhbXB8isUBSrigBlRFe0CX2sJsZIp8j8Fzlooue8TCY26t/c4D1twS9d7qo50UHcYIYd4guzITA
zM0P6r2cj7H3vcV4UdyfHRrDtrzIL+32wjazKNWrVqeeQ5p/E+9nDTCMmrUGpheNUpz1s3YAqxdT
iniqsDEd5kjN0zcBx4ABw35IcW78cUecYqa6UuG7/5EgAggCpHA+8kzOassRx1/idDaaEWzCKTVv
X7gXNklIEmy8/Y+vecCoh3H0Ur+bOxxXnsGL/8ZBCiOs3orOJ6I17+zJ/M4Mnhb4DIgab3YoRpVK
AArdFJnl78bjhjuO9mgdhkWO+dXTvrQsS8JVKEBstkHzsaQuGhECvr4vH4OJJMyluZ1brepxvSFr
4bh/d1X44zOT7AQEdpxbXIjfToini+nsSPbLTAov/UMSdXUnB+r6rm3sk4qAPQzClCodioSzIOXS
DbP7u0xgakMQngmhs4LQeQgMI3hpRqh0jblHQ/DzCgc3aiR3wbVXZItWHTSGhqquff+cb8UXkw+z
Cj0bCSu+fc8fOCgNUJf1fok3+zsKg/V9g4LR/RG0AAWQx2U8jBvpbV5oJI0kvD27GpX8nSMOugYu
su/kNN9StPmFPnvma/IDjIBBlzpylazcbB1hcUR5Ugm4R5A24iV149DknSyLa4we78ehUy5g3fPr
GgqSLIsxGST6JH3uZDX7KUDKe+7cG7KA1wo9RaKd9PUmdMtOh54iT/OSN/MzfaITvHPmOBcBkW0z
U1fl8wp2h3bmG9+U293T0I4Han0LhOL+KEo5lByno0sUmFF2zSQEHQ8WXnuI2icBKod200bGtTi0
YMWzgcTMmtCfQz3dSQslmy6VwQvbrKPu27+m6VwIc9A6I3Ye9NHypqTMQ64itYeo/N6Q/gVpGgd9
Xo7S4tH6kyxEENBG3lLyyTVaYAt2My7rmS66zKwa7pRMH7aTi4sfVGiBYxNYhKHHjipF57gD5VVn
+zKftOyDEpqlW/yhBJxMnXzYgkIcbo7VW2qN73KCV7Znq7fxIR5pVKalgXL9bvL8pfajOSGuHIE9
5T2u2Sena05imVKexukM0r9mgX4BJFrN0JvRtD4EkT2V5Od5vi3mAcBTTXaZIwcLT2zZLKm2hhHU
Jc7QHgAZccQvARw+QOsts+R2hRja20cIzIZN+rbNM6ZAxfUuXtKg57vOTRW2XYMg7wIwmJjQd/II
DnG1ATxTlnx9XMSFoBcIH1E5qh4+r9p/kJ21+HrAx2DSTSJmjDjIHCU5zDxXm4+XjZkOp2yalvag
E6koSPrV5hGG78P0Kj6qPnK0eR/BcEt6spbHU8k2+4lnNGnpWksYJKCmEFVhWy30s4eSliL+CCIb
Z/9gISya0hl7K4AyjjaMP/B2QVhU6EPkfjLOqekfomGy0gxsQvjmNE1jLsggJy9vGrjcNwnSO0ZV
cu9GVcsZy9GUzOikRbnujI8OixuwBw+z285UKKFh23mlg1sQdi4u8QCqXPm4qeyGCcyyTG/10vHu
6QOdGq5/ccpToCPI21194XFlAVKi4qJcu42HzrR8KtAVPSUBn0BmIyrZKWR2zkI6kc+GpvWbjVw1
Qy4411KrgUoIns+IodBE2frAV45samv92nPReQbyVV5THFxdCL1bhETUxRgsaTs/+pYleZmoyG6e
7pkSPbof8/qcphhJp5ZzfcvKixy8A+rsEtXi/BbTQCHykrZvdBpM6WAG/waAZVNXK0e2ZY9WVBL3
5rZPpIPe/RE+HB1A8FIku7YUc6WNLU368Mz4QoliXvKQo5Y9Wq9VWf46aO+p31R3zaXNG5wLNX8S
J/YDsSCEMuwvGoUEkfE0CIimhcECHgjNvzdG9Et122rI3/+JQK/b8ojR5mKMj0QyV6ptO3FSatBd
TVmiPxG3i6DG9Hx9eovhoXMkHzSo8CE7bsXXr17DHzmEK34dGdL9MdWIe8mv5dHog4x1rAhnRR4d
lskIiztkGNGFwZ2iiRC41W5vjBmPCYpCHDJXeJGaod+SahwUV7AzDGugSWE+ZWYHPoBLB+w1IQcT
GssPDUuZ5n+IiNYdNMG2YBubc3YE/gTnfwyyHLcvQjpFFO0twzO5cORr35ByFT+tz/kB5kaTK+KV
HjdzTncQGBHo8szyS+Dmy65o2sQGJa4sz0e1aiu74ZaMC483kBRnmLdIlaYTRdW96XZ3+oVtS8uq
PQn51zjNot6WWdotAXvzLlGCc48z+y1SoYkzjLejBF2P9wGm2exnOEc3FTECrycGrlTJeOCExnpW
t7JDtczA6hOL9Qk5fXLIMYo6SMXVLtXRNz/d6wEzUBVnVUfncWbTVaTsnAmb8/H2HMZoTD+4xqyp
CRcVhvrM7cpY7ikjh1/H9+H7wu/mvx+fvTqmiXxM8dpQsVo8EzgEpB+OwLRBkcoHS5yauNACnh/5
aU4IK1rNolVZ7zXMJ8jOMOv9R53b1MpR15QKeKr9P+G+FxxsLILySHnUW5eIy0zUaJRK6ahiYlg7
9y1Z0ZAZedgC5uHky8zMmdGAUK8PZlWht0bXdTwJyug0hWCMh5jrvDiN00IhOzkmkOsjw5mAWP/g
D5gQRhyGfAJX26qwv3UIY+i7vr2eLANs7V2GXyGAIbAOkHsZ1YUJD2UP2y1511IqpqYBWd2cGnM+
AAEJTe/kNPYoCLHKYe5fqW7B4qtSr4LHfa1vUoGL8+wov3pSLS+zW193A6u4bv8tFmX5xDZv50tO
TMKEO/hEgUkr0Y4g4MVW1FXvz54WJxeA2q1ehtRaH1vOWwOZgTo0uGmb+UtPlS2AndgQiDhGr0WP
PKyCHGUrxYVUqQvCqxwLRgbOXxI7Qv2CpqtH+AEOBy4ElcnYxrbmzNHdGDrb1JnwmJAkzIG6X9uR
UeOcPQhdgjW2zHDD8ezzpORQVO/5X+gXyUpVI5vhSbB1X1mi0AWspS43pusIuUOD6b9HgdIghTGt
ShRll1DyMgI9PFkgnT9UspTk2PwqO9TNVfvo51BlKlPOSCJcQIuXT6209jKGvQQmsxJBaGlFBjpX
d9GpXEuukhppe4vFh/lBqRpGxfrgSbOpAqxVr4zMibSjYBUS5MBWhgACVG8lrxXCIQ5Eodd141iR
NRig6cXovvoZ5KApH7wzR4NO5A3SSxdxLL+Qhe07yLqltMgM+gRmzWevacK9xv1myXZCayMPEQb5
sBiHxfzOOXQyrVLB/6Ls9QuP9/7G8QFkfjphEzOkWfJFhxkWh4VTPxB530lMdPUuqfiwI8PnAabT
pZSkjbfHQD+erSrbdwARGTcTEF6oH8UBzE0vmSoD10+60z3EvZ5Qfs9t09F0Nb4i49AniWd1Az5r
UN94FB2tbNofQriF2Cv061Is0QjeST1Ff4WRBj14iK+UjP5mNiItTkD6GkPyhIJEX1AwvwsXTpdv
+TUqVcp+16bYUEo591Hpmw2+iCsf8rWfTEzi1GbsT16KYgs/erHzJJp6XhmfDAcUM0H1fpRVkiVq
aZo4rh0H5a9/B7NonW68nzZFXCYXJRI/mNLimGBSmE3DLFNrv0PxUx3OuUXmcLIywqhJv5MdybDG
yvSxey9WV/d1+NRyOdT/NslRRZKZkXS8eHH0I+NE6DkUg+nSTPiHJcXyT8Krux3OtnmqJzg1geao
fmkqW2gQfXNBhsfwmADRHU3s8qkd3v4Djx0ymGcP6XT/gISBlsrYeIoPEXJFFAagt9s0vgHxj83a
FKZUO6ruSvZceViSK1tS20bph6iF0OwAN/StISt3BavH5CMG/rcKFayYw1G3kkgHXo/gXL8W1EYR
KERQ3KMsxr700OKdXbm8yrQ716keQi21ezOPhSvR/Nch7VW6JQCuRaWMsDzepbVwtZGWq0KhGe1F
pcE+JVVb8hnkBuIVS4hdGcsoHU+RTsay4cwo6/4MlopgP0NZmb1C5WeRr4RUlMy3q3h1Fs6j4UUj
zQijHnMGYyUuHczS/AafbVz5uLvJYCvWKbCtlGhLUAvQiX9tSX44w4BjIO3hQW+zN2wrndKTDZkf
tAFXE+6MWtOtZWZgjwabwONlOvHz2egzFfPNDg0d1qsbV34Ht6p8qs4SpxuYAnU6eVftZWeQl6+B
Pvkcq5qwAdijOuV8aCmt7FAVZI/y3YrjUpY00loTdV+yCCt6Kve3qGBXyqrDrzaPxfO/qv3mH3/k
JM62rHHVJ7519jPtIJpjHFxy0u9G8ENxGCRxhn107prj/5ZZqpDSQrigOv1AjtHKsznXRtVbymks
C7B7Uj6Se0rzZmQJMgjR0atMe+PDoCbmZykK2BmY1MAOhnbM8UharV/uOfgKeETUlVorNvSQeoab
5cKP3UT/i/pcNlMB4j75FElA486FCOLfzj/c4b8AD8Tjy6AoqdMFpsAVbUBf4bNO3xgOIWtuaDM0
tmP5BUMwQ3PXDrwwuI25sUe1rlT1zYWjQbXo/JxLYCiOknAxiibmrKbSlYM+dw5/6gO9kuHiwrwZ
BEIHXw1mw+u2K31N6k3SQ37zzix5HkmCjs/RifIV3bVQ9yc86wzjjDb1jCTxSeNCfJA9Hb5bz1B6
fFqO6m/+jFxY+4FToNDA/s9jeiCK2MigZDZPaZADv2VHsy3IpKE3meGAOG2K4oBm9SWE5IBTbNi+
h/1Fn+gKZ0vvCaG8izZIqG2OxvLPXgs7ZB34aiFO62xsHX64XrS14Ecm5Zkl5AXVJ+0Wq/pVQKPf
1i3a//CAMs3+1DWXqIC7UiyLr2QpGocPgAFjebOXxyoSvxhMTDeh9FZyCBW9r8JLthzxGV+RPcC7
qs6PlBxaVzAh1UUeUBql6uiE2KDij1cpWzZpjj33s1xpXsOIHEnbm7rx+dFgL/fHUmRv5x5sT94K
iX8FKI7xm+spUo6wOSfbOiU9q8qnmM+AJFdtdqgFeFUznu/qaZvCHWCVP2hY3zt4/C2IOLDJ4AI0
+Aiw0b8QQP2+FXqPyGjg9Luphqv91CInAEWH4DdLeVkjvIiQWHFWHSBbTNqIQSNifLwJJr9rbccB
tix392m94HNd1lnAScLodxsFQFkL14HwZ5dRON/o3+otMWi00PRNXNsT2q/kyvlZ1NP+QvH/7BNt
XHzZiDRl6bGLeLd3IQjnofpUsnVz7pbwEj3AeW/2HMvgBVPgTkOdxYp1pkespLOONoVSQ3namZHV
fK1tVa+s0vVWmAfH+jv35uW4T0jm9oeWQsGG8eCWg3urKhWLSTS7Y2mwNsYtAatzR6r23wu77CyZ
Pz2eUEMzqPvbOIyAriFNoIkSEPAQP15MAgUwh0a+VtcSk+vq5VniShE8kWAKCfS40I/UJ3Spityp
cHhkWiT69SyjbhQnUbSNrLtLiKI4GYiMwKAfpb/LrL3UFY9IF1G+8oUBTfx6BYeh1vuCr+972lvW
WOenssFnFSrNYM/gdxGoep5AUgd//B7c6UxrEXIE89ZeVfb4RvVVu0bqswIUEfnwbVrKitoviM1Z
jTw0hCTUm2ZV+rdY1c8nxo5rCo3A0D0DGhxQzblTTl9rfPL/83tEfjFX5HunLtuhmsC8kfNEs7js
qQFZtcPDih9NFMaUu30zXyrnkoRN3be5k7hIy57nXuKX+HQyyvm6M6Ds9si4lKycLFxeFogf9uKp
Un5yWiRT1G0tLBLaI5VWG08rOsKW/X+Th8VKYHgv9RZlbhZGKVilXVargcQEgX0Z4hv85liSFEfo
Wr+c8spoLjGG1UhJJ0fQhLkB+7or277fJLEzENvzbkaDm9zOWGPbeChPaPYkh/udb6Z9x4F0r/4j
gXsrjERNUHJfUMP4vkVEfZnUwEpMXbb0nFrJjf1ZNIPxQwgeiwevWZ7jlTc57M8B4LdjfP2Z5fpw
updMWQbH/L+JuaD8iP0zdMoHM4QlicUym76KcSQHBfzIDZBk9owcfC410iyOS6AzGbkFwkP70NhG
UGdfDaioBlQr2dJs/G+MblQgHMVmHUAy7KOoqflvF+BrJdEYPBv+jfvrlxMgMSQIWFzqROK8xYAj
ihk2vf5/OJ4R3OkrVOtef3lCYZaHCylDVf9GlrwGHstcDe/AM9ZwYsbhIkAqHfKvfetpkgw7PYoy
yrq4LI4Tn3/Vv3N5PdzaMFs1O++LLSejvQKjKmYpN1IT2KzyUnJ0TwfR4TXl7c3ISiFA8nuXlz9e
DXmfCbz36snmUsgr92m9wvf0LO6qydq3eFlXHQ0aw/RZWN/OMMxZDOnlblfkbuBFMAzBnmmN7zGk
x0tTpABoAau5OJklkgGllicsnMcnZhqh2BIzEgZ/LTegl/DePN98EODncnFlyp2Qvho049GxDxew
wwwpgRA4uwXaDk28yjRbZZgopWycawzK80znv0ukDPqG21irdzJM2aMYQSqRq5cX9HYHcViMe6oR
tjj5x7KsNWGg5gxZHLR6Rglp9sP9/P6TK6Snsxb0pierxOlCJ0Jd6EqbpF3w/AG/XKpEjFirNxCu
FoPcUNo5f1QZ7x/wtjxJSo/eagI/MnIejvvLZ2Kw2PPWl2ZnCRgk0eByy8wxPF0AsrI1fR5l5kNP
smr67pXEyKU4XK24tX9SxQds93lAgrIuEknn8AA8miPDwDXshTCx772YUtfyAPzH6g08zl3ex5a5
07XHRlNc2b3ez6n7nqcGXBp81+LsaOHhaKoIo/0sg0xaLodl0mAVOapx18uSytGTRcI5B62J7EB1
KgPGOvDjGwFzUOG2lp/sMyxPOqDZ4GGXcrqMAkP16PXoCWi/ZtxIX/S7R6eYbk3DtgBm5BnzKecA
U5yrA6OYNU837EGIvoTqGObpGSm3JZO1GZ1Y6DWPwYCOLt7MnmLLPDAi9v/Mjyj79nebenbX34cM
fYGMdm5e2Yt4gPUe1x2Q3//zl+cDYph27F7D6bRDdUsYlDeE6SGuZZImII0l8MUo8aPyAMHwKrYe
iVytUodi+XO7ni5oXY9+mJGj9YBzGTWfZRkhmIZSN499PkrZjI94imhAo6wcTs8VTe0J+Tw+RAIR
jYaFBlRH/5I9XSv8D9ejA4jBBOdWRzy7boJcjuEppMUYLqDWdXYcE3PBgIkELIFWQcvnPBlgLDq9
W0jWMqd3EVb4ro2JDaqM4jNZSQR4yq+sQqSYnuyCsACcIJVzvV53iBVEJutCxdo6W+e6Z8idmtjC
nwDWHAg1XlJMmW5Chg+Y0koNpPcPDqdR1lN9GSSCJmjUwNyliOePviBKaYabvedZxRa3ZNAxGgHW
pATd/oGVTW5CRq2ekhU8JNrcLFLwCcAzrUq6ZhYo7re+ki6lb1twYkHF7rQciZT3dc12BQVmOWgC
wcDWo3vNKXVNY6rukMr5sCB+dCrXmjReNN66KvJZ6uAROuar9fA41uGt/YafUS7NQhv6gwRYJoLF
+lmBK3KP/E+62RiavR/ggcjXEDhTvvxd/ZcVfUiHruqZzuen+yMGnS+a6pDGxnKlzl/W+u8IqMr6
lWq1en0IAc/kD3M2oEBIWUUvY1LzSb4/TVn5J9SyatgBTHX+GYZxtWK4AiR/fQIhA98AtxdBNkF+
PC5cae+zUPr4w1DlY42HEO0zjeEeBpVPb6JJ5r8eL1eAOIkpZvJ+lRGBG1gXoaYJPWe3CQ/sCYqD
ATWXa/DRcbRVbIq3v4Zv5yIVeEFNCKH6RF5ujXH1qYmUSzGKE1hSTtBjT2GiADzUWkPhSByR/pBk
MXNvWu+lC3IGXKpty/jgqtHPPDX3oJ2vY6aWi7+6TzS0U7UE90JSwNlZ/r+EuSFtmewyoIfJ1ccC
gVXA6QBd9LmyqJ5zrZopZb8yNxse0374WLILQKePNqwHhPlM9qW3Hmqoa9UMIs4dzrqfE1TeW7/a
Gi3NRKuHwTeLBxGXOAOEJ/s+DfXZWmSdGTf2+Sum22nK3X89ttQa660H7agsqmSWUgsUozdZi5ja
bEFEEMNljcDX5l8QOi9b8+jdCf9UKfHgPVt9uPHH1P5izMe9/SYaMOpbS3vwj7YpJgrb42yOWxXj
lnGr/coXKVp97GuKpkLWphpdbyMF/m1jZtDkt4g87A3PmNEZhEQ5AeqtKhVN5D42WtT+Gl6BKXIw
gpYC/S0FVG9dsc5JfWFNZ/OvAZnJx9sLPkwHSDIt0daoolXwFWVNRLgV+g7WuJRMTVtLcQvvXaSU
qoOBluaSsoWWP+6tlPbJwdD+19J9f/0G1Ww3B0G1HTy5TdJbBrBmDlvlxpT/dt121pUOdmz3EkaD
8dDSYDwWz6ytYpRZDbTAgiWU2NUqwLjJyTSmUhwJF3zhT0qXTDQmpEyXAJpZW0AEIDoTFe7yPJen
dAKVdMW5K3eNrbcmWfcmD01/avksElr+tJr4FTmTBoZlUbwJ854tAWw=
`protect end_protected
