`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HMtBu4FUyLzOdvXt8XhD8UkDVJGw2ywmMdYA9VEIa7qfttBQA4LzKjOcnIQxB2XlOCp6Sgmn4eUf
ZvWGjdLzNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oBWCdzLMDkwxP24pHggH/MdGM6OaZ2X+xNiyzZDYcuy1xhIuUsROmz7lguwjKKIoJZ2SKCtlOBky
sPiaX439nkETncTP0ztk2qIYugAYsiXErWAWg2KGb5pk2uxrGSbSSG6wwjVHDKGTS7GO0Qkq/VeF
M19woCOORe7vSS2bBu8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ykx5Zi9LWy14SITVFA1GVou21vCBp6Z4mp+JC7ZcURn4TC3dU0npNxKIujU9KLmWBmK+HMbxVzKg
RE7YM3bI+E1m2hLE/upWQWFovjnkAP0DtUF80qPA82NaPyEMEbXJMt2MvVTUWZoywvnVkCcMHVTc
SZ6FQyY3nh0xaC6V6inTc1akQ5pub8hoyryMuyt8F6JJtfU1JJVAijJGcPgYs8XvWnQV+pwcy3O6
DJK58pBg0KgPhB6COOiwbtTgs33CgJNK7uOLfduTFuw6pV2QnKK5lEG0rkzD6Ra0cUtAa0PbpBtL
4UkY+auKpxOCCQwa6CaSiXvLR0NBVa7WJkkUIQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jpJ9aLSNo+AY6AO+kzhV24u/NDhxjvQWp0l7CjPnGOqtuRqWMrvZJnKzDI/ektPMRCDMcNLVcOZh
OmDFqNES7PCyxJayIovb1sHL+5Fo2JbanmfppI5/HAHl2DbHn6Ta9egJ+dZ3DgxYvalh+M7Pw52t
d1+7UnNGeC9fshabcPk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MLiUrcsKmBFvNxNKSKHy/LFQt+IXSuCwj/MBJgcVntzVU+FTrasCY6ppQHQkDViDaWB78UWYvPD0
aHNdIxoHpK2PcWPjbHJ5l63CIkERjRhm4/Scf4M2mIeOkvFiA53nah5pzxpYyBZNuYvRY+sQkN8d
FnERQsuPhk9vfBQSx/ZlzI6g8yuM/VbbAeQM2kBSF+Ehbt+EaJvMyOgrSVLVIwuBfNNA+uKh5xtj
X0QrspcXIq/6V8t8N+rHQIlLLHGmUkh0ZdheJLGpyctVZ5c/HGBA4EyPrLokqw8ndDWj06ACfLWy
4CdGa/iqiOwDfHSGckQMNAeBrEQOvAWmQXTUpg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 44832)
`protect data_block
Vt0uEhUouCXoXvSKjd5LQt91x/HiJdCyTe2CarBGieoj6bozCZasQqWiByceTPyIrKg2xJBw62LM
Q8Whiu5JyCUQEUKW11lopZIJQ9uQ2HRGAu+5J1PAt/2wuBHgKtBREjrbF2+B5WHrSHynE5roYUrX
sKkqsMTof8ucIKnQivkmDSWkF4bNaDa6uPubsUgPN7DKUSeqG37V5+dDS5lHaYDes/mbCWDQY5ip
fSIWclq8OV1hy0KhynETpCuROsnL9CC+G7rRknFTMA8r1qzXi+4xpvb4DJwmhXtzu4878zkMmJ9I
COZ6LmdGrK508R8kHFdClALwBvXdU/AcA1XgQWqS2p9G6+esVlwiHi/AsQwnzBvw15TW/imgl9/N
gfrKAWZ3SDxC+JU+Gg1NUJQ5L1457jNEJPSwzChNHyiq5m0FZZVXNzlRUPGTMbqQiFdkzlj/nIi3
P3YymQ4VwYP3Jl1dITkajNR2294OA8Tiw3UWedzziN70VkibxBmRxpR22UxoUQcW1mxJVmyrQ1Tq
kZEgO0nNprjSp0q0j8lx3Txwinf2e+xAsYM6n0/VlrZBCHZGJ3Pb45GWmvjZE1Mm/cCrwj+iQG/7
/X+mCr2iuidZnpy/IqZdERCu4FoPjM3G3YyHjfV2lnj+YGd8iSgqcBkRdeDh4tN2+SUUjxsZz7qI
zB/MjGJRLT+cN4HQMkLxm4CCgBcN/yNyejaw7Maaf0U8X2K4W50PGoLkuxmGA5A7XrQ8Dzx5mCaI
8iODrMeR9tPKajVUEFwE6UCpAA2HVXhdwqWZvsS4KpxnjvNHY4Y4HJz61utla7WDQ8AHiGx0CA4J
TYpZkbYuHfL5hJSLvhp2o/jJNKc0Dfd1JwZK1XaDQWFwAlWFAKKZK4dZpeN1tM0JKVHpBmFDdt/3
Eoy6vZZNQXzDIDrIN0mGJBCzWGRZCGsKkCCd3Gw7qfdGXGWzq2ytaQFzh2sNoYl8bJW72U04Ja6K
UnKz0cuYBmbvmr+lr8PF02xrNZ/OvfMeNyS+sdU8sbqpQb+jOjzuP+J/4/v565F9Q5cZSWYGsVQ4
ODjwzi2a5YBc9pCexNmIg1n2JAyyHpli6BSKiF32TRqoyIVCoYx2zlPgiB1iCZP0Icc62tsmiNUH
cyZ7wu3rYILH+dYYewGx1Toe+zW2gdQ40m6s+Byqg+zEgG002cbsrktACzoBA66zz12+PfZBoEqS
NwN9XPnyyWLokyN/cpxnSILJIYW/B5UeqkolkDVyqj76Usk84o7p0EqKqtxSKZNRok/jh0c4TVAJ
DvhzzsuahPJewEuuLwAw7LBAeBstV2jsE/qrMmeEAB26wRvg4uQkiVvzcj8eN9moDNZMDw0picxa
7C3bgicpoXMJmr4OBeDQA3JUst0XOda8pcdFWvWSv0dWms37TeSKusNCDnLEJJbYVVkiFIbfDOL9
P+xkKseYee7Dj24Ue+8iQARqkO8RHgcuB0fZA6hQLuSDIsLEK4DoxJ1yhUtP9zd/xGmSxVEIF8Xo
Z5+wg81USjD+bNXYZne1CbK4D+ya2IPzHj4O85+qHH70omRk2/SeLvdv9rnkU5cx9CBsvT3SykJ4
roS1r2wrcTzKnQ8TBwMAloA9/cjA+A1pAXYRYw1OquM7FDIRMvpcBgwfss2ZptAMY+g19W8Gc+oM
q0K3QMJC63qYMeKg4nZ5HQ36qdrlGKacu7zpyGCT6s5zuZs3QAENeITiYfy2L6ZRQ4D+09XZnzWK
K5i2X7iGjFfKfTQQGBFJsMYG2Jd9av6KLwz9dm+oBCQxL1nY3zpPOy8PWNcxpnqkCZZj5HftzsJE
Uh/lCpo/T/It/7gH5DUiyJtodNwHQ/qSVn3nmNW8i3DSkDLpht1Zsek/DX/Lsh07aw3Lb0kXafm/
GjmAQIVcCN5UctwDcaTcHUyGL1crZI7NGYFjz6MDHagASTndCObZv5/dbI4VI304LILbu3UUqb0f
bjbld6EaGz3xAwuVAhr29lw0gwnBhi2Mjph1iwG7da1m7Er0s1ZT33+jTiVCFnrjSYyODyyZ72VV
GvW7Fp3i8cdu+uh0B5qYuhEYA4Ai35sMT1XDgCjSTQ67aK4G9xZdt/0AHkwFYScxIiE6qExYT10A
xGLoAYxwE3yBK8SFYHGLangDz82U0Q8VNmQ8Jc4+v2rhPtn9Cf7tvB1+CZBC6jOLkPmeVaQzDtT6
OMJJVolbmJuEZl+xZwA5uzOyG84tMjmt3NRLHUR2djRT4H5DL4J17FZHWbhTFOrsu09QR0xKa5B+
p1o4fwO6RZYn8PEPgLSrvG21LYlyXsevcCL8FZTEhH2fesQ8ZFOdBN9lqqXtBSkj47wbrXGJmgfy
ut0P6GQsMMWTUSy/UCvFrLYxb6eIMBFftyTtXDt+cIGgGi7N7MWIxtWXQ8q787Zxr1rwpxmsh7MQ
EoE7KAErrt4SSvvKO8Q1Vb6BMSow1HtyFc0brfI9GdvsQxfaLvwlEC0crUf4PzGo2SQroK1nfVsr
SdtgBh8rH4yP5Uh266KbFly0gfW3GI+g2V6ltAOTqeMMqccD+FkfilehdVBn2D+WVPgqD87Hn6gO
xmmh7plfkHTN+kwlO+cUkieB2nkszo2Wq5Vrg8RiIX3wK66C8d0SZm1yfCu/B6WDy/4xgymaUMZj
zsW/I/ZkwZ9Bda279a/C2FeK7zuJai9XaNMRMrgcFIB2kAq8XUjBLGqJsBThVEGveaVDkBDwW7vv
uNPz8oFJ4JHTU/CylHBsR5xa/tWVGeMteNJ6zWmZQAAy/dJA4OFC6/2ZlrxOYX8WK5dF08sS3IsX
9BwbQA+LainYGNPz21cGWF/OEQD/oaB4w7GWoTN+PY+AFXATlBfIXuF9laT10VSnJM17w3kqgxfH
GqjjLG2A0eLCH9mBIbjOP3pp7mGuZJjwC/tVfLC3CZAGgx/a5RPCegzpy3yCZLUvGTkpgRK2jdkU
iGLrk2zcUBpa57ivEycAg48wrOomHoyil5Mc3XlR+9or3njtn1lxL2eleZiq6bLTAhNB6gVCfVhr
9zJe7cgOjG6cZvREAGFZ/r3Rrwpxp8laeG3HwJqXmobBOk64c02KdO4/FEvd4D/2mpNsTN/Y+87i
5SimF3gQKVF5hJVG87ScgzWUfVAuQBDN2MuLTitY3APQ4F0FVemInP3jKIAQ6cbjKCAmUuASDNqP
O+IuRwKamNWxBrunOcgyuB8iZKaakAByCzHgHIY2pr9SA/2Mhg1XlhBU6wZLZK4zlXch6gMXboE8
yzcdn1reFJG1anSfFyAidNGDa9dUVsUg6zQUBeJh5F+UZ66IWqv/fTjnunQ67rsne74z0Vu0198u
3dkzg9oPxnkeoNPgZlFYTYJnUQlgty80Gc5jx1Sn1sO/5ykRH88akim7TsYT9nMP1nl6jhaubacd
aN/aAzTkCdkSWIjDVX25aqAKo5+eVJ5n+AI2waTnok3k03pdo6C4/8fiYTg//sE2V3Y783I5bv5Q
4ltTs9Ul10fqFCgLJpVmZ7All1j8CQ4ff+xILB1yq7ZlGjLMZg8u00/YX2Pgn4Q7wYyFAGMNdw+K
KyG3DZzQmoRN6rR4YlPri56FWwksc58zwv024Kg6VEB0t9pZdjzrcmWpq20X4jduSYcECaoPzcML
ArUJ8crvMzTVR1HEN2q4uh59T3v+dGGBTOwRx7JIubdJhTh9IxT8tTtbRjTg4yl+dmZjaXoQWDFu
YO2UADusEtfNSrtwmdC5K13tHLIt6Mx+rDghreAjfxkPuk/SFoNJu3Pk88ikP6mJm3tzpoNTGLCA
WzA7O7XgVqVP9EpRsWrNFxiPCTiQAnKjOsJjRx4cefoFK4k1Hsf5/RZGDcHUj/Z/TvsIRGrzZFxU
gkqA8FpxsNwlU+FDNY4Hr4joxHNiPTXPVGcZJbd0zZvnxkNfJkMLrk+jo1idVxXnvSTvoalnpUCz
dyDTfk1z7eRy08C/F9ixFnteibrqdKufreWZit0EIHARBkLJz7hOEZTyztacRysu9v4cRaSucHHN
xZ26QC/J7zinvlTgh+MYRiV/u1RW16Pzk4/igZs4KrFR+BbP0nnFA/X5mueLce6oktRfMSa34rni
m7NYFhfuab34XyEyIV+WVAVbrzIAgNvwTGRzAfKg9WDcvGBRmsRsdD1SBfS0T9JVXJh5mRMhNSlL
Y2T1SvoZ71u5Kk5zqNwW6b1JDWXv9bWHRnvOnDq8Hv3FaKKfVCASFgqvwhp8zwIkj5q3lbnxrttd
3RuPz8WCd1KooxCgBZzAxNuCm7GXTmItyzW48lDwYN/kDdaaUYE3Fltop0KivIfX6hBKpWZKz71z
O1e0Q++A2r/84+1cKMOYgmt2zrh1JPKJ3nycrIoy1zrCFfDmImjq2XOJU8tuJLG5hAN6UVJKE3FX
cnV8WIZ3OLIh1Yq+y+h7hx98fV9RlI4oNjpQcewmrAgjD78ph9BzlqWAdOWjXDOhsRA0nzGB7I7b
O6ShIqlidQdOi6/LcGD0kvtZscL3rYYdJWeyTTdPnkeTxnvXiTcfRojxnQd0WZbzEG+PSLtKG9T1
9VTpAtwamkXyAAC3ZMbMtVNenD4l1ULXK+vbHrAkAF8uIoqTWh625hFPgQu2aG2PeJ6D8efM5aLl
F56vYHXfXDdPiq2Ohj8I8ghb7ODMF6yAdu1WxDCnQ1ipcXqhCZf1uT8QZ2EvRhIxoiLSuUcutZRb
nCK1iU9J+YAZlsans8BA6ilGtkSBdUk+9wHNdXY00RExdkK5SwL1VYA+QL073EDobHs9D0ohe4Kn
SW7SH++tevSvSBzvUpUBnv7UlmKIccKL0ctbc32cJen73lscfJm4gkN49RxZ15Ozl+KyxURBSrtI
KYhviaa2wIWjvBEKCFrPDfOCqkr0Ag29X+Q8Z17NJdiqELYPFxV1fpX6bvYJ1NAU2x1aqHMViqFa
ewyBUeLaPY7nhR9tUNNV226mIPN6h/9GMhK1AqPaLdObTLCc6/vvcV9glN41HjGjpPbjv6CYO3Qu
aVy6dcwFb22EJ756eJ7/fcbxpKZ/jITHtfKg0Y1Ra+gn/zdPAVcf2LFQ7UmGsHhATiFAwXXVyJOg
3We2lAjiBpQWxDH3Bj7QPfgPp4Fcl5Qmu3EO2gGKVMxv3rDtALXv6CeOfdRw7NeGdETDG0Fb8ScW
p1zarC0iyfFiSBnjr5FzO+wjJyqbajtKqZ5In5qqacpdp7vIMsLiF/xW39DK37bO2xf+3Ls048/d
8h2e5BiVOfa7vjkOOiioajRbNPYVqoNpdkEhWcxgEBMtlPM3RGD7swnGXDdE9o/FPICuY42GnUNS
QOFgtil5LvJ+19UEZqEm3qEf89ieI/WA7qTPJ2CZgovO7dlJzq46ijFZAfDcrkFdtbFSF2eCzTff
FWF5VKKp+TjWt3SIvjrTFbOdpVIqgjBmwaPHp0XiFiITgjn1poEqCggvC0O3NwLm4v3sOa8zSmmN
U8J0BcH8UEhI8TUMduZXiyvK2fzpL6mOnILfU+Qdp7AIzDkg6VscTq3ZgHoBK68qqraE8jqrufuU
tFrevKPghMbi/Cd/ijj4Ip0/LeHaZJkryEyKaEc6b/tDPTzCEdK6Qn+TuVgEog31RPSoy/ZbctkH
XkQwT/QahDIbAdyuxEgEDu/28oEOOMpqcmgrpx17uPKGeUT3UoipVu+jXzpRohJUg4T5XJ+U+b2u
1u8T7sA9ZsMAwd4FCXR2MZWAVWE4Ku5jaBl/OxrEkVjkepBA31JpAacrj01bKzKY2wfArrsOjL3e
8spS4c6gCeqpVbJGwosUSJcFWMKJp6dkrfmFVVS5ZLXwbhIAhKcbwVmBP0UgzWe/WfpyZSi/077q
RQS8CnHGPp140v9adlJy+q1DH0Uq40+BqpgZeohkFOIulccfIYNwRGVRQwv7TwIoqKVLGFX9NOVr
HfUlC4qCi4pYgJf8D+RT4HNegIaJxt+OjWL1mHTCL1cIet792SbFSD6Gb1iAh3f6MBiT7qc9VZiD
PoUVNYSyiUp8qZVPceVVJfoz/fQkVgm89vDOHRMeIDF0qj9TPiavo+trf5Q6OaPxbfhVRx5ZyjeZ
atBABeNq4GkIDepghOrEk4izhBPJsIGZbBfKGLY2SczJWEl3Wco4tqJiM8t85NJ8A8fTZhQf0KuB
TrGtNcIVlIzoPDMm3q4vmWU5UqUeBXxd2CFdv+HqmrA/MTwvJ5L6J5DjtPc7rHzGGnxmGW/OqCUp
4K1YiLDzhzXJNrAz0QZnfTkk8Bp1YNcxWUIdOksE9gJTmMuxuwWr320tLLj4dNzDP8Gh/CcAvjxK
1VNvCCkdbm/i838yRtSEMcnP3JdQx5XO3i9a1qecW2/8/gPWLjgO6Nb04a6ZkP8Czx8t3wu6xJRP
isRXl92h+aWcS/yrezOvVtoHO4N5sL9W5ulOy81aYbgqbH4wmlK9hDMzbt4K4/VUEUVNiZ+Wr9xi
70aw51IvKZZGELXJE04rZKjpArVmvAJlzbnAgaO30iKiPR9J5tah1H/f7653jKSC+BcqrhsOFrs5
wMQ0Q3KBrnGCFh05NCsPirI8TKX2EHmwKeGG/nzSik0l5RgIH5+gBcVbKycwJS2HzNyv7t6B5e4Y
ePLUcYBbr3UPi810y1L0eNUis6zZ/H5KtDgQIqx3HAZcHcaF1wE7QgIYrNh353FEwqXBRQw10jwv
f5CxwLeNQXTj6waWkgKjIpA/D5kfQ7ThbPN3Y9yTlslEQ+K4tHjEUI5eHKd5ba9QekM+cX/iSt6X
cB2bwOgzb+7GOfsm6f51+7UxMoWTJdr2YlqmDgeKzF4/S+MR0k/YVnCX9B187gLLTT4tXUcTMDbY
e+Jvv7K9vC/L0uZeJNHMaz5JtTZ18Xx7idvDJcc/BfWTl8s1Ot6VcC6XYPVoVIMuKoYvp9L12YnS
G5gEGHPqNZCHr+nLw8hsZWjLSB8Pk2oIZcpJpRfvPIkz1fzckwLYbK2nohFUVAq/YMLTfzdN36ED
5NO0hCDLUcD/8Q2MGETPPYSg2+mUIp1qaVJ9ZVbj/YdWcGQ5+WSd3TUz1cQH3owDUGUMmKKdwueB
a8SrSbd1VSvfwPLSDIQI4Bv7zHYySRvoHXcYbmLNsmT8qhMoWvi49tuZAMdtjLPSs5SUeqRs8ZnG
iHKe8DTy1mdy4/2rYwU30hbp4fGWeYAFLrrTzrl+01CCXYmuzUhpO0S22alXe9mfQmAp8bEvKe5H
PBKmCvcgoIUDX3JOFE9s/B5ES7xvBgh+HHRiDniqANXfPsaJUT8LVO0Y2GG6F0zizYlDS9EG9Zwc
60nrslzplAShxzVWAbOlHM2Wh46lx3fs5fP90T6tZ08LEIebIevcv2wNLeL8Rl9tYrGHQ/atQ6VW
4a8bWFlxVTYnGeM6M9ym/bFT1MxufT/2NUUrmA/hrQ05emq+43iTPE5euKZXBai0G/ijIYp7u7Ks
bhroZ00hJgbOh+gYw9Ciknod1c6td/0cdoP27C9ZSZk/ck7ZKf/8wVnxF/spfgwGJ113U84DaAhP
3Z0ko/FTw1WAmaw9oMxdV8LEDSHYUMuZD5Pa6DOtGKE9AXk8NPBEBUH/ta91jen/RORts0VtaeRa
7l5/sMqp7rPPjRBikfcNKulcwJ6ER6YerUFSDqwn/C5TrGNTarGqbWK6IaMFiYLIEnqFg+1nYqQf
z2TIS48Gy+nV2kBK+horTurDo9hUwhLw5fKcv3KjcWuJja/EWEfw6J5MdGul4qqhT1JLPEY8E9LL
sBG21wFrEWzqsK9ESQLUMWLx7IOQbsOvbhth7zmjvOuWU/zVB84i2KOVLf254dx8eI/JWSDqinEc
4L3on6Ig/x0AVX7FX/e6GNuH4UDa7tfK+qt+hUt3xx5jiAXwfWu0FJGikiXqew7vqfLeLxwq3A57
qg/FWMp+3nceGhfHd23eoVNK79EhiAQ0GMIrTDh5bsQUuol/Hnr7AREaPN3MzUZ3jNRbg2Ap7s+k
wLYMHu90SZNfKyuM19lQLKwACv7vS8z3eVWU/Ns64Ohv5DwLkM4xKMOnEp3nR4pveqVtc0e5qW5q
zcdvHy67HVjXfFe4HcY9WTkvS2R0EmNh1KjCH7hnRz82OoNfgsejQUIpa6ionyYjwsi+UKTXP9KQ
ec4kS150UmspTm/lGutjer93C1pFt4ZriMBfqwnNqNXm/xojn48j0srD3iorcSkZTbdCj8BPJdqP
Ek2Ps0Sn1oPsYQ6kEkNiw/Qe17Vymoi2THoAZez+MfpkZWzqomOFsezyg/YNBPwUFH0ozma6+rvS
afGQLuqR74Jtry2WkLhabg4qWJ7W82T+jrGMKSI+hBi2YHtkYwO/ivlGLKRvtKvbHflULepgIINb
5Q/lb3HymoIHGRU9SLkZnqzMDoVfjlo3XYKAfQN0UmV/fN3JR0NgLif2tdYcdnNnbJLMn7flnj5W
dumgpco3CchLHctHvF732+rONqhaGMMpN+X42kHv5AnxEnWG57RvvMBLnkz9W9ZVv0o7kTGwYB1p
yIsz9JDuxvZEQGafaeyQCNm5AwJ0VIrTl8+YpmxOAqs0sXPCI1WY5t7K9DQi5WpmVhDIh0XZ2yK3
YtFm0JSSgUykBhj9pXnzcJFPmzLSDB/8sJ/hKEdfTG8Ez4ruX010PWHZMAyHenezzne9qN5ri3YE
ZVemJgt0YqtoDTTbE+AYs65AtB2YRWUZ5li/LB543vLRkJc6DGJgGsfX8UaP9Ulbip82kISTlS83
LSme694KziWpAcCXn4ed1ynIS4NA7x441eiI17AfUvU4E9v9Sa68UCwhKSbVNtKxksdiILSKFPY6
kZbBJl0TDSAbIkPOiBP9hTQVDGUn/zXqDX9ZUvkUunYhZ24HRJHkqM/PocCpGjaHYHhKWGBW2UQd
5OQ6pHJjUDeUXFJ78BCn9ghM1RToyquwbEvCBw1iTzqbOOuZK8HCPJiMBOU6tvPMsG7qU/pFJ4Qf
K0owOP+LLdMBC2OpWJXbLpgsqVYfBJy16euej+9LPaHvGYc4X1ffa9kr4fNVF6BDQ0WXwlpms9Da
aCBiA0B3VqqbQpqrg8FEWeBqOplqRhZ3p45F5d0VwuaURKiFUCxk4ppH67mxlKJYpnbyTfFj7v1F
p6R4+dg24891zPji1RyjCJDtTA5DciZZ+x7TRtIvCnSycXRYKrjpIMxlnB1JzrJTDm54bhfoDa9J
4KDlES4IAuFf1d6YcqjQYLNRiQFYnnygPrDInT6ZU/3xq6Q8LMmaG0Su9hTDuuM4m7Hp4R7D3E0G
+j7of1LyJQCGzC/u+OdI2FyCYEMPVxs6C1cGWzLdaqiudLk2v3gcbE/cXuLKupJBI1xTzThzxSHy
QZxY3W70pecvMF8j6XmD4otoBheEW8O7t18h3x2BiqhmOxG1nPFIk+v0xcMqMt5FMOx2eXOatt4+
cIjgzzLLa65otNHskVO6ePj8k8qKoLFOZtssmmpgewp3Ijvcj1JVZrY0EB47TGtbR5EeMQhuHfrj
BmHTDfSSygIUrP0tq8pzBlzlUx8ACHLYco4rsqVf1uGEzYY0JWlCHyaDkddxBHEzPQWQkhjPvjKD
AbZACMqua3/j9H1izfGLGE7CT1T5REAZqLyEKDU1nydyo7HqwhhFaiMj3EyoxJMW4vNpwiujbMtE
sOocD/Qdt1g5lfueTYBWZiWi6cF/lvNCQHmX8JrYKvtC5dtHHsip8brjBoLQysWdIa8QZAI7JsTl
ga4Zqsoirrm2SGbJiR4ETR0ml3BTqkeuqMhNs3F5c3cVpB6YuQ5Jk58VkREUIFN+SFccomMP1lKt
/HMVwwpWhpEswkX/E+81zpRspfocoZDIIZJ+h1TNlpChFI9xXsN30lfSl0DSJ1ALOMPhRNGSZu79
9wlbjH/4xH4O+/0AQQU6+XhrCRWsF5DT+ocPTd/v5v/5MHzmveS+ZWln8b6XaY1jjDI9zTQbsGs+
ABWkZIe5k5i1VPkehiLXxB5x6x6ZciJBvKnHAnafFIzu4uR15H+HqPapzG9uH8ls3nFqsPcvSLHb
OMelxDBzQufVWu11XRukW/z+HllOlWUMB7ZciVrSKszcJ1B6nu5pc7aLz5Y+/2q8oepYAGQ8Gwn8
UmzugrvCRY2ScvpGCO0derzynhbOLXC9bRvuqz/80w2QD2YYYTQfr7DS9qQ2E/1XR+qjst3TKtwb
HePImhps3sZ6Nh2N/DLqSSP3zCRbnOG9waucxmsYe1CjDMn3vql+kg0PyNVEdZXD+r9ArhVRSwXV
pb6gx6xlmJFvMMzMRQdS+u0g5Z/Kn0VUCtMP5HCGdv9TtKTBRllofDZ/wmAl0uRZif7qfhWL/uwe
Rzir6ZzmP9uakr9kLYdNhJRtAZuXxZdCiQ/s5lzZY7DhkloXe9SAaKRubZFX3zu9HFWFc5bo5acI
nzpxAj+Ovr3iRJqp8UIHAlHU9Y1v8e6zzb71/7z5n7jNlT4Va4GSKYd2xSdyZmhTi0V6SpLAtOqo
ytHmaRqTDAn7L+Kcu+rzmT8LurqqYblEB0TWad8y/qHj13zdm3d98KWY2PSjpAHueBroOdyAJEBX
NT2mqVQQiDMExfhBLadrfAeOQIuSbcZYpob3fNx6bjVwKvQEkFAQe/MExYpU5ZePFfwXoR0mh/LT
SKwjuHCankrrTPm0KYSKQzDz0y5NBVkAk3o60XaSwJy1n6FXnYuJ7GHK0saIvjtdRT+DgS9Si84h
N7Gx0wd7Qc9EiJBweUnfLfBJVzq5ryHxzqdeTKg95wylTCHALYx+NyrbBnl/NoTNefT+vqB9kzyk
NuL8ftHQXv4GZ495igcyigPtvgotS7UirY5K8S60VZE0iYSTLco/TY83HTD0R8H92+jGT7mMmLCh
BfVhXf+CloKm4IaUL6Dp/MVw7SOlyx08pTGHuqrOvEUnLXtx5++YwzhPx2smG9KLgaE06hNP0+KK
rV7BpTYdkeho51iWYQHFnoStvrh1j30etyKsz5oURF+zNpwsI4A1T5aObGxFbRIe8aDbhe5t91Bb
dh4yR63cl7Pw9gRe01y03k5KsmkPSlmLYrOQLAq5/PmCW/0tiD8R3aKjDbXHwSFZVF0eDps4aMLg
JxMOOzsK9cA8s6jqGawlkhKsPY77x2CVwZrCWhOV+uozYkYadardyVJ2fRB2SJ+UP0eISmvEvOOr
q0nmim/71kAf8oHvGBV5fcFh6CgSSc73UpIsCzHHON7ojjB/t2AqeT9uGmlIGOnzEFD+Rt45hTIE
7Ik4DoLsjQJ7pobd3Hf2f9cMZjuZGVUTC6wbgCJQ0HRnBLUXRMkD8bwQ9iEwndUy3VpZPKgQ6Iw2
tLd+aJDwA/oXTGwWneWIoQrOejzg7DfsEQ3ef95+516tW0NwI9FmznxkQe0i9pzaR457IIhiiRye
XAtYV3qjy08UMbjUHBT6aJOjOXNeM2tzFQ7AaR/qKbLcE14/RWkAThP1nYJg8M+i5vKvaLz7C2FL
fd92aqhv9sqihTMN68NaDCrBAHMUlfiKQu2IpT1JXxSMeFxCjnnqovpL+LfL1N3F2yWKlbbN3Lj9
aVeSjjwfZRk6JlIVHywaGzTDjWbJUe1eZRJfkrSsVapdiGOeh+L1h0CKNryXNykqz2SsJPtUaL9C
kZgOXI5HfGC8xX4e3871guivG1ZFyZwWbxlzFYRzLAXDrwPr25S2JujS7WbAqZ/wXCOMT2bgM3it
FqUPNJtoA/evTUjPAZFc4QY/ltcRixOhc7Tbjj8h7wT08fQxNzZrgfU0GYBKfLL/jFbrl2tP+QIr
CAfJ+BN1Y12e7vjgwPd9CYzt+p8EPC6TXOabg5Xg4osjphudnC8PEATTZ3PZj/EZihpRHesmFRmK
YYFO5q7DORaHIIxgp7fsihux/w3+tIrc+zSecUSQHaEFeg6t4ZkFiQ4ckZ7Xz7DWLWijTzdUlAKV
mfEQmTR9EPs7vuTngd7EiqHIsCzFAm2gPHF0uVx0bC5vfz/FfBBRnlEixnYBVha3/cH++P7awP8+
0hfwcAKVPYllDGz6VbJIHXgCy3AOBI4rp/AhmfoS3mS3sUNs6Lbq+3TiAlNGKCHx7smqj9zEOS4n
S/mE6QuHVX5TV72pUUxM1VNC0LgK6o/s4oF4LZeKw4q62XEZykpPlnXSOCjid5sUk8NRlopqS6+5
Y/+w9LRblWB2WJPnK2YPjn402ZPeM4U4mGOJIoaQQ0Bc7SWP9hov0G1tpWHrzbP2ehs9NtC16h5Z
E8+a63sKT+997E6cn341MI0yj9zm+MEgHMLfHwpQwYc0pwcHFy4mq/6q5EqJ7La4035aVhZHKiiX
QPajv8zfX0Wwm3a0RwKqG0/cqycgDchIWxFh3PkiCfi2Ou44EaYxOSOU53yJfcPPztX3qjRjEcIq
9K2XHb2K6Udj7I2zT0GmMNkGNHXYt/jSx56PtJ6TeSSdHuuc8v+jW92T7d9S8vYSAAv6wJhHal+N
DQcTV97ZSr7fduwWUr7rjwd8C5rnw/Qqd89Yxr6/fdOjYTRuobwRu+QTjzt6cWxZPYTJBZI/bqe8
yqlLtj/QM8Mj5Ww8BGSv8IHlNi1RKssVn9d4nGxlB0YU0NZ9ybH1ZFGq/563zLrq6V0M2ZOAGqBP
Aa2bxZpaaOWVIq+2EI7JcncEz/nWgWkXfZTJSOMq76RbwO2c6yPDTPrEyEaU9ONOqwqLfN4xySYz
BR0I+Hv60u5ORrMtr4BeBED79xOL6OX0AOmQDzxkLjzQoniwdacsXxwFwkzBWDF9I/Nzal2AvP9b
yN+dFewue8bS81PdY2GFFE0nomz2sJBsBXpOzvx9fjmfiydfRf5bqw2yrWhUqC4AWQT4PX/K+tOX
KiPpJjCSywDJs+MDvfZDz8c9kjhwLI59E5121iV0wRh4vSv5s82Fh2EJ0AWh9+ylTSdsMDBY4r9V
4NncJ2VPcO9xLjbyzEzR8BIZdQ5CbjgIFUt8DjAVtay9KrHIclXqADSIIcP74zPo/Yn4x7yr8x4q
SEdqn9S40/ofwDhbfBhdE5bf14+jtm81kM/98aS0fA+SWc9qkYHsgQDjN2ayvVFArTtRvgwlJeNL
+fyXeJpBIBzCWJuV75MX58ZjFuNVkK14YkSnPYmvT8jTJo7XNfh6chldd3baKSg4Kf3gu6I8sWiO
mJBGQTIvxaws8ao0V8bBbATxk3S+6sXzuDluAIB+IaXVvO5c+YkuUsbPBCMdRAYi9YOai/JXroi7
Tdv1IIw2vg22mXxBlRt2LdvqoEpAD6IpqXCd/Tk0/2qs38+l7oRBy3zGXt0N27EGHJAszk38FpvT
QTyXyYcjbAZHYcXelxOD+MB79/L18vIYKgdlEmCeoDYSo/hwDnSmV6tjZNuqtIXxDlXawGgJ9q7b
4CJuSjBs+i25C0P/DBLngZR2HeBFK+/QeqfQ3FQ5WxeXduFeHX8Cb209eQF7iLHoH404YRxpvg1c
8fwGogRFPqHqlpuqtlRvYM45eMYE3MPkVfJQpg2nn4j7c5yw51+HQfE73giGUyFml9+vOD6OzaVV
jbwywv3afXPBNebaBgFuGizAV/R2aprAJDGFQ+wpA2OxRDNmVEnmFd2uZvvf/J4LpP63BwS6eco6
uEXM4YSoB0AiJfmya9a7PERNqnQqohtsqR7g5hilw4lnqLdH+thZa9oR8J6q49Uu/6GUgwB0P7Nf
vu79PV95qlrvgaoSryX2eWvMeWKnG/OJtc+p/F1KnKKMkXWEKkgY8wVWr154VHlDBDVFeFtUrwHg
wkh231elKKXLCv/mLFJFjK4M8oTjRwvQEBSypziPNDkmtSX5z7+OVVQj/uzbw1evKsYS6Tzr7ooR
PpIVtqx00blDqFjRBOVfxikSXI+HJa2LxYBp2S3KkgsxcFfoncoi0IvkCqS32Nyo6UE4ItNsKAwE
r5BoNmYIvkqNEUSn/dfJfgQbwsHphUEhFSkXlbZeu9Xx6Wrs/8HQOJyDs/Hh584XuWgQVNEfxYAy
MtmhqKq+/BZtHgG4UAPRMxfSqUiUlcaXcf+oLH9kA7zbWVw/O43/RApIjomWs+bgFCRCfS0oN19s
IOZWofpsVavRRknipmYtzb8kYWmB6JQrIsPA+csNUwrYPJgRnRFaCJb9+jitNNfggV8CJQBDYquB
xUwroFWFT+FbsStUtiMN6Wmlf6jmU5rRqI4lvt49yZpelfiHBHBkRLeJtblIW+uxowzL16Am8sq8
st493VtOYYUyOoy/LcRYJEqLNzK3wU86wgZRAIk3zsuyzIoKMdLaZHic89kmXCxYqwaoBMYSkuOV
0p+c3YbYpTC/wRzK3Qx4sw8oSnh56B5fAvAihd4jOVWnQlvLl+oWuLTLp8GDGdPM5zJwS6MK3flP
LhyFmee9Nz7lWebrkEP5ax1m939zlJbDOWUqxSXZDwVf2tGpJPoc9z8nYSgBiZ/GrSiPdvlYI8+V
XviQNrCcRAa2laeor1XxBCbGvs0tLnzzWLhJpeHU6jO/E8aI1a9rD7xuO4MtBpUibZbUEemWiRtI
a44oZkuO/sqx0MlInQb3044MhPs6eziBJtr0pFnL3sEmB7Ky/hEbKqvCrPmOWDMV6JpP61DYNDp4
j4Gd20EPbrOzeuq1KD103JJczjWUuNi276ZWfO2rbaoVnEYRQogeqSmCBYaYgJRAGO2kjrSKxaNL
KPlasPGuvLNqVpSgEac07RaaVqtSRxOIhgig4JVxHLlmjw9m+qW9/NbW8ZHC1NJ3a73bCzKoxQMu
+MfrJYya4QKD6qOdayR6Tihlvt2vwr9FmGSLuQ/K0+AhT1yXTHNYtL0t21v/URoW/e016VmMorbB
1RGLcIu5ETCGfOuvux4TRfX/9GqxW5wrzaUmo2+w+sR+GykP8IlkrE0pdeT3qJl4EA/Wh8SrSvdK
vk/wO0X5b1vmAs/VgoR+7Ogk3MnYCstv1ubc6Jv1dSUo2u2rE4ZESAcJDOL2oVan9TBfEC0JtzSy
qky/vg3jGFCwYm2Di7QVMHDTHE31os8d725CmuDftnI9P01/BizkSTL2xoa0l1koDq3xSXwDfqu2
yRuG94umZiGW+w8lTJguKSykEsmfUMtBYUigjXkvU4J1s06uA03R0KKPMwekxkBqsO9p1OT654dN
M31rD3QxrNjKoTLiUZTsT36uK+ko+cjO4Sffid7xXdbpJgjqr3NXv2RcOBgt8p30p6D6KAqxRZH5
+rgklLDkajvHaxq5GLqinHHdjTxcKBTDc+B6rrqjwol6D/BZo+OzbRPsbVkdt4GK63vlOv0KfQmk
bf3n9McNrRlHrHAN7vkkgv7baAGOCCc7EdyOdaQKdW+5K9XeYqQuKmcGSW5FmGT32bK5yhTnJADj
yeePazObSXGzWsEsJgtBkRoo+YH+KG9uFB7v7tRZA1a18wq3oM1fji3BilIkIsPxlLD0xK3Sg2tF
DXKjD/2S9t9y6p9augWVoghWZTxEvEpbZW3Ik0g/MYCcgfVijiVlTDhW8xrGCJyF8oWK9el/+Amg
r4FR/O+3qVyC6y40YSIFC4k9dn4rCkaf4tFwXffzX21Rx3HCkJaJ9yiP8OrysRNkSB2+KB2OKTdW
1yu+cYLxNHST8lnFyZETfBiHFdxQekubsK5J2Y4ewn1CTU2AO1HsBev4/0AYWnKhb4uwv0ns6EnB
9E6vMd4aUNx52z2MTg7s0UOiOPb5fcCSdNUiQQLq2OhyuGgLuZobKSUQNJBYRu3DIZxlYC3nRmvL
1rOG+FlX3vSQwWxvN50jd7q7jzP7dkBUcrgCOTjNlZvG2XCspN6bs+qEbnFIxDAzz1WP/7rDidgQ
JGiE9w0SY+g4fgpPmhuSVxaITtpWmTshT6n4gDCaLbqCE2WDi1SEikToUSI01SCo67dRvhnOwvp0
0qbhhVzkYWrpq7jiUiqvv042CITzeJ4OjXq8iMlyV7RypmYdpARH7AWIyiR6Ul+OH1symGPYwCYo
JgO3BsYdkuApzpWnvgwP97JUGpHrdH4+3UOD3Q19Vo+bMDNM/Gedj6kGjL5lufgFyu4wxZvq0dty
ul4bF6MQciw11gd8H/fdg5Sr5NCWNs8ClirbPoDseUV/Dv1vxtJjZED4DY8duY0EZTaVghZbxJHD
Jv6J7oghOWfn0w+dUcPK1LD5+DWwKwUA+gxWmfqkjmRJJ5rcGHRwSL87QwG8vElSlKCq0kxA3sL8
ZZ7ItQs0v2W61f6rQVQN9MUki9pyFyI9VMr0vk1RWJ79HnwgzTjSGOtr94voG7K/fnJ/WGKhtS2b
tKDpemhyanaXLlRbOucDzw75HLTVpuxp5ctGgrxIDc0KXLc+jJTs7PXhiY6hvXHl9vSMjEiJ3W74
JrZiOq7RsC5Z9P05lci2flPjHb0FdvdAR4c0gRo410KZfjRO915fu591QULbcSYXTR+q8AsDrt2Z
LG5wqDJsN45VRGiDN09ceWg8O6F5RXrMiSa5PM+R81rxmZtnhGcR2itCfkhSl5vK0QYEH5kNKdf3
o22lNphDBelobvikOAEGRay1Sak62c2j3Hp8f4wss7wtdLX1oFJg+MKcEBqFkdkKIwy/Qd0BRuWF
FBcpmb7DCDXE4BvlVJwAjse8lAVT7+0sf4/vuQGuORyNVqfpXFtQkxAw5sitl81xvML23mrSwcUB
tAG6AE4kBSCQmi+9tZu1dtjlSo3zFJQRcq/2MvKHu6ZxOynj0Eo4kxJ3r1D056C//rj0aqpz89GU
QtgwC/5uV6ERx8VrREvuZ1wimvs0tU9Z71VJdFoIGsb9Q11JpWeyCRDqx0shKtqoPoh5T+30Kydj
yN77ZOD+ZzTdyg5SP5LMHi5oLuYeUw3yW02Ug0iJ3yfnHrcjWqpMiz+qnybKVMNHH+MBtp9JXf07
W3a98UUMwTHR00t061xDoe6roWC+SWmHvgzpzL501MduwTweykTR4oCr1ZU46t1L64UiXEpmoANS
kuLWw+VMr/N1fyCeSe1GGzwIF/uvji8ftIoiXqooV77nUBD0AA4lT1fGavBaGOnSDC6uTmll4FOg
yaaP4V8r0MexGsuo6zlhTiw9PL8CVQYV6AjEciaPihyyc/CUbYDI0NgqJTdTkUbN5VUVGW+ZeBf7
s8CcOLrQzwSLiLApQtWkCQ4+gac/gD+2kXtqea40l0b18qdyxpd1B3nVINGh1KF3YaDb6LgX1XW7
+farNJeqvPekCP5Tf55qJ1OrOsAAkjO2N/EDUBQFsIMbBEf5msvAJ7ERsVHW1jCyhcXNRuVnUiWg
KmB6hcnZZJRHvPJhdtV8SHx33IYM2ufWSkUFfWgv0A2EBUw7bc+7OnwnQhBUlJAKxlhf7PFYGivI
mMArO+ziLycxHS+4W0NGZAhM085/16ioEAsu/dV+nYSfOvb5SsKRzQqUvvEbKt88qmRpAT0ixa7a
73jlH0Y92YAkKvrHiAvxG1j1rg3zDbkhCNpdRyO3bDUK2eSIGmcqzMs9Mx1BLoZiAF/4oMUYjrqe
pbwkLMBL1wwLF4GsFIjUxqbFs2BvwRd1LlPIuScEQdWDJDo6mvAMMjVKSiGGoRNbzptyHa0QaM4r
kbQ1iig6ck+z7Yal8loRhsMHYxROwJujUX1usYedSgztzT9tLSf5dRIoPAi9re4Nmhes955xsMln
+u8HD8qY5H8KhdIGNHOBYC5IfLR/vGcpLqQ/ZrLEnOqb+V51nBmPs/Ysczw+0jUxD4d/xIhA6TDi
Nx+w3jVmQQtqO64juDj0JWA+B2mYChrSMlWUE8NQzk0N/RqdcNPHZIpKxPdyEYcEje1aFsktk7aH
627kn6XdEbVzFkXkLOqKjMvqGINZbzf8COjcpxDXg46ujUi8E/WBLhZq/KeL0I3iSRP7gw+wtw8p
Vj/RxTIseZU3R4rMMlT1ORmZC+vZwtOak3aCxqccLJQyLeXpLDga3pYfIb/RXJZCwlKJYu2zUVq4
FCUr5Fks+KkOyBwA5ykjNTgHkw4LoEUsrSQM6aZoipl6dybw7HLDpZGOJUU+ShMoPyhExWYDkAOc
4T2KeXDhDNtUhHgFObjhSv0h+ABfJQo0BmUM/WeYIK91YCndNSJ5zz9j5gyT1Zdi0Hmf+JsdGnhe
T93jaOIoRJ3rtJfYMVwrzeDuZd2Pc5j+XpqhJ86EqEzGrH5cd27SQpb7K96kpPNdGgsunMnFwA7W
zdFiRY085qQVxtu2XG+xoLNsMtvGjYA34v0r352amA6dHdjrrSdvojV2R5S6oGzXNe43nFG34mjD
VoEUsTFAcTednuP4QAwihQAIaHfXsheHejqDgqsmXpFtqul9PdnSDhdzk5dsIjXACOKBv5mX2vc4
4ZJbMVvDU50Yz7fDDbPyOkKA7xN9YTeNLZgEGAdmZhM/3ZTgdWW6NeCa+V0hNwYz61IgVF6SxoEj
Zo2XcYsDikQGRvtBx5XPbH/Phy2fxCv69Qh1txDcpIlJoqYdkiW+IZ2O3kzubiTebwKpYUgMD82z
uhW9d7ymmtDpo7VcPpAEkOw5jNH5rf7ootzoZyrqM5U0MQHEv3o9mM0VQYM8wlA1H823TLxYAT5v
FgnLgbzi9EOJXEvfvWYzlif7jIaKXPfP1UyLG9EfMvz6IiHI177x0rV9umGoT7YAz7+N7vbAV2AF
48q/T3icCsUVOJkuRiqUWaetmvYhPvLPdnSAeE7wMYcXJZxhHa7EEKfJrV8UOT8o0I0SE4JUFtLM
iTFRdiMJ2MDlGmle83GAaf/3B504FLfyrDQc1sjMY1Aj2Y1GaRU3fEt3WLGAMAx9Ayx3XLOrjNbh
auGsHagVPiwcxhgdbm3Fy5f3j0VmMI7JWWDh381nx+bWepXlL+a9C0Mpm+0Yqnk3S1FirvH8mjOb
x8hTqqFUG3g8OPzOqGBFNzvyhlB4FVouL+3biyTTf0KBkGFLRd99R0YrVXR83WpYNk+KshuzyXq9
nWjL5ftBfTTOwWsPxoUuCmZaEZZTcxK8mITIOxD73YuEQTdjlx19tEXtdlVNOnWaLl9VTpb8o9vT
4eMcVxfW4ravj22NKmLRx0Mnd9Y4Ki3cBRGjMTY9r3hbVAWTvUAZo9cbNgKGt0Wrn47Rs/pdYJAZ
zA9HIdfIyHZUEhUmuKoDcn5cHkSOEti4XHkQsM8mB3OeAQAG1CohgYQ/BFINKGCald2GtQVY2pq6
VfX89mkjEkRCU86inWIJ5PI9/1ArB4AcM6vndp02cVrIcRICR6B7RCPNNs1xTHqgoWEfS+vA/1j9
ju3PAuMFJrUtMR/87nJJ6ihIjKX2Xj/kmfp/Uga40XgLuxr/9lYJG9u0gPyG0G2FW2KtG/yP8ryZ
bLV4AfVh1Ph359krFR9sXwmTlrSjrEBfBaub2/lIr4g+LcOEli/mNX+vMCn68Ua2BjZJTQsuhPVH
jmY+uAdfeU8O8UbPtOjobu/fkuugMZRKH4s97hLMgMrQxra7zkIogjPe0oQYxGhsPlgW7K7PVG7k
zAcJk47TaQeA+2zz6E/3thA9r9sOTLDITTA06tfcN9u7CqyG65P4sj8NJW1MEgM/5AktgMKdrsJB
HNRCgZFJsFl6MViNtoRnjFV++VRK+PYYWP3P/UPgQDHH2oCgO5+RXh7GKFE+QVR/Pa7ZKOeqeUhq
Dk3DdYR/pdKkbJlIkvEAdku3wuoqgRIR1jpSXcXroXWDHRUvTI/xYfFhbJCxf8WTUaysg2k98zRF
hSejjryFYwMZ5L+xf5giAxpHenBn+1qq8Uo54ZwXNni6PqkGEfljK+w5jnWbVPwPuigXWGyPn8m0
s1OrpGcp0Ojkdx+XXLxhjK/hmYYPB2eZDhsBDVXiG6cmlm+oDLGjtdLUTaXccP6UMUQ/lxD6PqyZ
Z7AwM7T0zol4iNSthLl/nffd23CGz/53Sqvx0xdRd9vKIUe5QRHR8tVi6lTrugfZvr5/3qARdRlZ
4ItyEjOT4bO1NoiV9Q+EgE4e446MVuA6NItJgr1rCNrn7VMFRe2GK9hwit5M+S6Zvho6vSsUDLQ3
HoSjuohnQQBufAvmaTCtUr6ABfQifsbSMMRYwa4Mqqw+x+G2kmALTKUFsxprtQ0EuRLTR2v+xJkt
kfWQtUhsVmTbL8skWw/WZNSyZZHKf3T0ADP+jWRcvA+FCZskEEzFXfSNQ3UlTvxC5K9aXA44aoeg
JXcToqkjrxM4BPB+fK5lrcS4VzNkMv8zNY7G1iZntX629m25/umQ6bllnjpwIgMp55/wRWLlQzxr
R9IFWCAHjZ4xhtYiHmCa4/EwsrSaCwQm/7bu9zELetfValiplIay8DmHU+YHaGz9/jY9GkDwKyb8
QA49YKBqGW8wyWy7v5spmfLCKuSXKRHFYKCuYcfMN3Jk8V7xNbUFKx5VYQQ0/J+3xU1Ik0IYabja
afZlfoq0qDf1Vg7d2hZDKR46AuHZ2OT/hcIK3Z8WQj59fN++CvwlzUI3vUuGGXrwz0EE+snmw/jN
bASwW4eZlBi/M6jknrJNHFZvhmC4CcP63bHCDIoPBdS782WdxVQd4M07X7Y+yt/lmg4vtIrcvfhf
npOrCYlmMN3WlLsyPq+IsBpzuuJGzOu0lqq+dnpUQd2zm791Ew03rRZJLIYuJLvwKC3Oi0CqwMKy
4Yuy5SaDRi6nZ3O241YYDUysb+yz30bS6Hdy4PtKc6KHU+F0cSdZkAbNqWhyUHSar9au5+qGI29U
+Hs5JVqPSxnoTyqYDjrFAvumVvBwrCAG6X2l1o7F4fDIcm5e4yiG6Qai7uqxKh7JDmBWkO2awXif
tA2E/IWxej+MJDMNGx+FGoQk3f7RpGEE8sMtMHL4XyJ32ao3k7IONkIYWgBeMOuYmqZz2PF8pJua
jLWEyZtSlM7VNbx8jewOuYJjWUR8Y+O6oaqNO23yzj0Cl0rsnpA62AUvZvQLDrTYFvPC41wdei3I
+oyPxwKAJztvSf7BPXJpoj7vvzz+t7166P/dso/O9CuLzOT3kRRcQzMkz2xiznmO3sz78y3CxaAa
/2tO6W1GKRunZn57II8tMrrcDoiVM3F3ONUi3vBWzeuLvlKkEOfKK7jbsEs0NZWHd4+g/c2nnHlg
jdyyEvBR0biB5jAAYj2N0VdlkOphzFNqD1AXRJacPKcBxS5WFCo17mGtXCaaqAvp9O/SFt+6Dd4k
l+sv5fIggSePIZvoY3pEYZr/an25wi2bDWyroh/Nz2s9LLDrdBSIykGOJJfhBZGjKaqVEWcHPJa0
8g7lON1LU/m9l8A3bBuL6EzSqnfAMP0nVy1DkpOKT9IVCcg7E3RNLc4o1q85JMnarh5tQV1yP+rm
uAD4NLLgL+uFUp6NflYM97CBKGdZFbjBoNFcsOudHaJnpoZkC0RfzZUqe30xWzu5lyXeataq7PJO
H6pBbPXW+E2GFdhdBJxDKcRplnEyG3x5u/bTFndnf/QMWFRU6T/zGYWrxuiiT3S6ZOYh60BjsYJZ
ykwknIHimvqoIVfEAC1YQbj7k+zewEEMPU0+DQACXQXSQdMn9f7jVP5ZjXrgLP13WI144Q894B3q
W6uWKFALf1B+gnzR9yhO2BhQssO3RHV6nV+UQ7PZdj9YrWPUV0joxkm/SoxnIgVB9K+bVWqm7G3J
UGhsiKlxBvzL+sHHx6Kj7m2MI65yg0LVjRywQwnh6+LZWpJrijVEoJyWN8KiDAcVrQ41Vx09aah5
ETZnjWFO9GZQ3iRLbFP9LSQ220OtWj+fJTessxWt8D9FAshAoMCOGsTga5w5a9kgYhWwWwZJFqyb
dJTHf3Dc0o/kXYtuaT8KMVb1nM+y5RvHgkuGecR1pmtkPK0dGmXFw1NFrkCtYalI+CiHWXwdp0JK
v1mmKTtrKRLggJrOauC2jEsQI+06CbEbaIvySuZ4A6GWZj7pMD6B78b4NZJlkSpVyptEyJWzxCLy
CTOMPGjEiLKZkLqkfWr+kNf9CU/KMxes4oN4mZ2RMu1NqFoMnbFtI2ik4WmG552RtXtil9hiBGth
gC2EIqzZt6RcWEtiQAVbHMTguxfBMWcV/MqVGSYF9EFzs5Ez2/FbsILzh2eONwXWNio7giKcf1ow
IQYhB+ATkkm9CQjIOqJrDD8GRix24N1HU/ZKped3aWDk0sqp2ArWnNSJnCX+InUNUYtRqQyop2/n
Lk94zbaorKqzxYWtIn/y+YkBzzG0P8dNfpN7DLEUC0JvkHPspZ91vXlpRwIFjk84UDsE9YvrmNRl
Zcu6A4wky7L+wkHHmmE7irv1PrSm+VoEBQuaXba7360souUIUr3x0owx2LQVgk6WxLMq71MsaUSK
6XEiA59l1BLxwxYM8CwTNniTcEsigxmPSAD7uT7bDr+8ecNtoJXhTowhZSOixoFIaBIZCQA+XGnM
AXxfCn+T8JjdxV2OqUu7WEGiiMIdyF9Ih+zZ/klQ8bbzOnIAUpoJEzw1JQuvVTgL3rvxEzGyIxut
h2tcW33ffkrKP5ZP6EGr2VA3VqY1Z9qtSLN4TziDfQ4YjiTsljL+KhC04VsR9Zjq5r2ynUgdLQdn
wxJftVdT8pFJXDCKCdYWcjlFgiZUOhcIAfz14trQKli21G2BhZHjOd7Yb2D7IQe5qaPoc4cDpDTd
ZsZzgyjAAUWIGwhFOPcV8fzlccP0Rgrgusjb4LeWZIbkZSg4IQ54UnxCxfmbrVx+krJubN9vStoz
91kpDwR+yi2s3yhfpdOFH+oSzToHV2auRwTLtHLBr2aE6xhZ/gkbqxQEecpez4d+ksqu8NJTbvT0
iuQmnYdNEyA9SdtpvSOw9jurp9GoCcOFB2LIMGe78AUqt2KwrplBHPUW11/I7/EKGmIz9jJanFFn
CjYC9gmKsPgwp8z7BSQ/OnPBlq4hT+zwBFJJ+gxLiKVFfCzPnUhlKbpOOXC8GEbmiC5bMpCFhJxc
3OhPk6+KrJUIphc2lfSySM/6gxpCzamHgkUkBBEvz42INpSvaslw0ucZkXrhk8wKujE9iaH4paQ1
Imm7Uo9Z8XZV1K8vcDI1AJuSedkFLlSx5e/m9pjHoNE68LPcC3lY8OMp7QNZ/QQKV4yzeeY24UuS
wCTWeLvBzIlPHsa5tHyupkoJPI/aSYW3pGfHgDFuLSxcAil2wQRgs/BYMHCXjJVPcohL8AVhn1yT
LJP2kG3C9w1TFzTwA5mD8l4KOtmX193wWpAu+JBL7tFPfFVcsmyGkIOTDFfdEpripXamtk2qqnKi
LSoVgutiE7ZFp5GUJav3p0UJvSY0HEXtRY/mxZr1lQtzvqbv6h3lJ8Ava8S+zbu4vzAu6iiGvYqN
kqNJ1GSSFRt3PRGiSmZrPOY8SAC+Sg7oOi3QCsykEiuiZcDw1i3Q+kFuBy+brex7Qn5Ogy8AQGyW
W6g3NjSavne/rQV0QrTACcgeubidSuZmmzk/JWhiqiHk9rrnMLw2KtbK10E+jiA7bVUqtFIH0BId
YgHFnEy81lu4aZSLa1TTclGq04NfYZ6ijXF2FgeGarRTA9gHWGEVbDBUqZJp11BqjJWhDEf7zivX
WCX7/zByQEKOR5xOx4rsO3rGuvduNfFkFJ6ZtQ7vrhwa5NErEGJCFhI1rGebHjVl87iWFAdyAVn7
dlkiX6esDWSDFfbsMKzVh33J9INvb/69yy1RXERbRosbxhVzKCTnvdLgm8+pIQKD3TA2lnOX9/2m
ZHKPwEdJtto5ebU8FILwl9fG60qGYI9dd+DL++j9upBOfS6ygGPD02JVNK6hZ+DH8PDkO593qLtg
djw9So2/0+rbygAIOhCXweWE7ki9ymaEqSO4J59bO24JOUF8bP/IYDKNVyW1Ssus2Z42qnuwheA0
LoA6FynvW3h7h3GPiRs3bF/WtHJV8hBYIlj/L7qlHjl9uf0TkreIPsini8B5Kk3RmHqz3AYvnFtz
zNy2s8X2R8R8G/FdcEuNSuOhzqPwqWBj73FW2y1g+hkBzqyRpnttOokX1GmBv+xqh75sl86lXHBM
iAPL4X+5w3DilutHMFAl2FlGishCMtNxs8K4K+RkjiyJSC3cJPibFxHi5udw8Ks/iSQ7eg1iBqju
fMZGhivCjwLezh5b7OHbBjsj/B1kI8ltLO4yTZYRpL1efZZ4a74S3eD0PdCqiyqh4DoP+i3E4AJz
XurzUyKZyFJDU8Wmx8TbPnctrz1NLZ0aj3FhKPm6hX8yZe1FMvnQuPqWQBlFK0XFkN0FGvrDVKpn
+0jPW3yrPJP/JnfRVgo0xXoLIpDpDj4Equ57NPWdrbV22V8dV01g0eGKK3Bkoj88vZJRgPVoP0aW
7dAjZvKaV+KXGKwqIGi4uhxuD9SMMIPfxa8hGjarmDTxqWYjyq0TcJJIwPfW73wBCsmshEgnJipX
kAG00y8QbXOfegikMbss8ozbFEUITPCvB8wOcchwrthGk+boQ57tRI2IqT1GMqo3K+3R2bRWs2fQ
Sz0rRufZHpUGfggKAms+bvBmz4xX6brG4jbTyi1uNOl9LcqhGfRLYmoSH5XRyQcDoLD8CcQZVPmV
kIdjAqFoBTyWcSmtIbUKVZXVoVQBY8edqSl0sPBJtwA7B/juFX0TwKzg2vnS3rqsNAb+AgzekYzj
WffTt7kptnV9tPwqEAckFJA/hQIES48BhG4hjceWq0vrem+LQvuXEXctN/ggbM+tS4p4XkTGMnQm
IM3+lYZspPKRlWOZ2oIdpxxdzEt/jsa0SxCxe+i9k+hG4w193zAOq0bH3rBAZcbyX/0nJIj2T7KE
prTUY8bLT6KBizXFajpE1XKsSDfz77csfvMPXKFYIH14QiXYHYBH36V09Je65ZF/cVydVLCX7lag
TL4Zf9Med9FzqpzYir75yI0BYHD3itFTkvQvi3BUV4c2+zgdVGDg/MDx3RLsV4SI6YTKG+0dFkcj
AGEd8qk6eq8CboqjdGt4HUJj+rKOZZuEUaYfw8i86U5jmCcvwPIqyFO03w8q9WdX2scx5lD/HdZh
+sGCMoJfl98QLyguHbNlFe06UM9nBfA+ZmF4+jUXElAh29L1xoMmKmaC2Px7yb0xQDhYP6zjffOi
EhQ+us5kPPd2/Lr7iwtps6IQDvO9OO/ADTrjHPtBPgnGrY4j6h22biuzx4yHB8CIIg0Gv3o+42vG
Dq0BEJwE+yGF7zyBYjAyGYpBJJzH5VecKHkM3GV0b4XpeUMhvA9NyE4419j+fhoKb6tlQCv3gAFv
PlnShMHCFeTyljmVAdV5oa4gXlymEdTaVUGGBe5dkKSB3Dr95Fe0/BBIL+gXohDxCyStanKsTk8O
MhWdAhdW4NZyYsYyF6ykYCLj37s3d3uYuZfh4A8qc0FJPMjuSfzXdEeyDqId3AMSeIaiH0CSmD48
6vs9pI6oTV8c9U5UXrv+HIwYUx39XMEb24gyIsCE5/1F6Z7YBF+zWNtv7pzvFoE4We6rHzKFIp05
Upuqs2CMIeRpEFgiWuPo51kWXF+HcSmx0yHeqNvMWtbnnqG0dhbD8qym3qu9M6fiiupkAFyWOW+R
BTGdBoxT4LwyQddhRAsAUjxhaNl253x7vHyOX93XyzEubN9R59HtGHFxHHY074h4vnprWTk3gk8Y
76Kj5PDAJjoDIejMnlHENjyhMHWbsdkXIfLq8e++7+/YoXymefaIkCBwS7qzXgF0c3LKIPyOscE9
+ueRZsdkYytyVHCahi4P3gTKNolAz5rbX8SuGbcNKBW2VIULTGcY6P61Bjz9HhQhA/UcDOHmvh11
w/2+q7ZNIPmjnAMyYTyM6m/TgKeOsGAYjrkBkiiyG/L+yurs+yQ2xYqzPodMGBEzJT9t6bW0lQ4E
6j/7W2N0t6gOfvruZmmucseya/SyXg+N5fVj9zD2PB1R7jyiZ+DH5QvS5Z1teVMdlJVAlar8l77w
JVIzShI/hqeg0UuwamE/H4P2BzfB3+wbJomhN8Q+qFWsf79f6Ko6UCdarq1gQb3pxIrfD/jR9I38
c+PBJ1lCMMoX4kELnbdx1H/WAj12plE6WllIZbH/3Xa8F+Gp7CBLbYLJtHeFkL5OWnt4ID0dxMi+
E2SimjPB7DH/hKcrGD9IEQSrt4i4WVgFcGNhAzeyE1q1Vt4UpnRXNM9OpC0FHaYR0A/PqicGQ99z
jRglyJ3x88h0k2JCA3zPhSnZT0FkN53J1MboexQc5Km2KRudUzAAFn9jA9OEHM2KRZF2YAXTWcWW
7XpVp4XWbmuHvpQZ7dlL4uxJFwslBG46iLLmIPk8CCFWYvsBw72SPd2uLQz/UAB0cnRPeT13ZyXt
o8zJjccNTVvV+jPCxyuTUDDHalKXZpllKr6sPOr0njKcdLHcfZVBzl/PsCve0DurYLAm0jTq+RZq
BR0bqlK+755dsMdP4zSQ9xAc9Nl2Tgfm5GoLd6hHPBRWnArnfowpOrF1aAg5Qxwz7z4lPxpcumrz
MNxW3VmBWIuSagldSEaY6SvSgviWyg75OcDH67glRd+dviC0DhbnBjvjHy++bqm9olRJZozRRcGE
MkvvDAYnClqijD5X8Vc7gp+DTxCvkUmFRA5UbpiIRi89KvslasjwO+BL+57oQu5u6QdIKRcKCK8s
uz4vrxtn+5KJEoPSeMIy/o1euCY4ddo/kVnbs9ZP7u7Acd3pjoqAgCZCv0felQ7+zP1W/SDqXcRk
9Orbm+oR9gYhycdsxGUnGYxjP9WdhrZ3oEmoL3nVeAgz6B9+lGrFI1Lvy3Omm7ueX9VAR5W0adfy
7h1wvSgKtjiNcZnmZR59u554ad5fFLWRQau8RZvYp+DmPcBg2jR7LIT3E4826yYbAj4LGFvYk/Xm
d7l4ZfYVZVfuLOJNiGzsdwcGLdgIH1Vcqm8paH6aq88Tm40ufhvefawzQ6CCZ//x4z16sAeW2FZF
OZtTzsHhwXnC6CzDgn5j9w0gC1oGSAf/geI7Dy+77KCuRx/zjXLlv4HQ8ukZIe8F4fohzApUC3sl
t+SXN1hVi37Jvmrf1q1ycT4cSuHc+mXgOraLKmLFgBvPEi45xeC/JtJsNg3o2HvY9hghV/iH49gk
XSSMx5MSi3xgUWrR50LmDyhdQ+pA1FNUMhJZxaz4xfE1C94ejpGsuTPXOSOeCoOMIqlST66eZ8YJ
Zu95Kv+VgNl0b5QocTP2+RUR/QfT/Asy2yNgVTUXkpY6zFRH0O4c+xUAcn0LBFVAiLZmo7g+LMus
a5dR137ifjqi34QRgY1Z6O+uH/8/Z8SAuAXxpMA0URdD/ILvRmGzsiJCJoFqyd7kGjbJZsuHbrY5
IR85Pmi6D5skgcKltdhUmxx0y+4h1MX8X9rsvg+LRmaJ6U4dABCG78Uf0to/HOSwF7ZpZRiN3/F2
I7jjg3mNaRXn8mxA1blb5IWxCkbTXpxZsBtSCQFqOSOdSSQ6o8SPunJD/rGXlNJ3HXJuHB2DxqVO
ftSb55OTB5DCMLHgzACizPNC4mpr+PNspMlaVBt61ChcTtXnyzREgkORLd3dbWPih+zGP4Y7yFDn
I+G2hYRDVANz0tEpSFXEs4j5zjou85cENNoe74xjyKvpC4JuvQJBPU161XKrULCFLhbuGj8X1I3U
O+0DmM+BkjBOo+eNaFQn5iNsLasOz0ddCK5FAkpEbvDF2X7ZTJRUonDoqshoYvX2hbqq24JM0LYD
rsK8tIQ4opFh10olDkVbo6UUuegPrV+dYqO+tbdxyEX2Sxc7EFYnF3LUt2Qw0BnfBfUsfHJ4oTuV
/Sx8tms45wi2ttWvmJT7GYqPKdZcwVdaqI97MkiXFLHPyRMJAUcv716aG6NbcCPG1PLVXeX2y0MS
VZCY7PZS4Ii1HPMsbHqj4RWcQBki0VS6Fit9RZEsGSOTtWGOFJTcDcQnkr/F01ld8D5fPRHS7xXX
7Buil69WhKzixQMReCQShP4tD7TBJmHJxlMgBJHw5C3MQ8Qoll5kCwqGTWcEkg6hsfvQcf0kVvp7
D1wbSN3Wu4+4oL8C1ndqEHkvOs4EpDYFBUxTQrF588s+EOWwZCT1upQZmTpdj+tFZe308OUcWBLs
fyjpZGNvHa4p/PSDcxvy0KMmz3tDmCYNO6TrXk25aYtA6Q1x2+GjLhvV038txCLg0y39RwN0TCvi
yKkOOINRwiQ2oNIf0Iep0ul/YOzDJGUn1JUt6CaY1c5RiCp7YtRtZyyGGHthJBw3o7KX3Icg+//8
M9sDSdH2YLwZLc2NHghnQoiM9y6HgKjcJISZOQk8MDVI0JKjtAwptvNiWzXkG7CS0OmdUh1pGgAG
wQ3mlSdtLQwkQeVtmWNUmpVxhIFXpJwu8JKaYm3fzUy8bRf5gMMhe7Drg8A5PHdDAExNeypuqbi0
XR2cIHo4nw6rBjVhOs9UVaAaBngSG3kzu89hxOiimuFbO/5rMs/VfHCKJXe4as35J0/EgSJayToE
j3gFS5Utuh+SDJBt+5NPrIgv8tVpb99uDzm7gfLpZ0d4o5Az/N8/RArzB8MkjCOmo3FJIuFVnqGS
HQW769XjFRCd+F44FJ1BfC2obUGJdvtqZMlaSC6mmQps8/tjc5kcMlAS91Ckx5mPeh/TJqv1ijVI
n+Nw30+0CmptZ0gdywdK13HNIHhIg8I29BUaPUEaDFMEeH0ReWUZKLnrFw3dwq1RcbvltFAUayl/
wmNjMzsvqPMbgOg2vXOGtlEvHS5ptFAI/7rL50A9CNp7Vc1GxXOIcOhkTCGV/9b7CLLJ5zV/gfp4
TV9WLrPsemTO7K9ydod6DZmiIyqJS85ReAVT+HhFg/llAb+w4xe0T1a/p2NsUDbKSttPyZliuSZV
7MNroL7WGrdl0QZscjBpJOUkSJyfFWQ7YkN8SvMKpIKvvi8uAmYB8oIUpP7SMkudIHeQNLMuw0Pm
r5y2fBojHeN5E7QAKWHgJfbplBFC/kE9xWSc9wIpms01JRHSBT0DNThA9646dynmG346UUNCk8E8
KTSW/f3/kWe4rV1b9W38+A/Mp1uYV5/YJmuNhwB16zIk1E/R7YyjB5fG4UXlTpHGbiKMNN1Sxfpd
YPmxZK8GsqidGSCTE/2pRCgyUDyURdMPXhpMoUPbtvOcvoAJldCGD+a3EHlS1n0uJy3YlEN/Dglq
rTu5XdRBomOTIyFR1mfSM/N8TFU+2GwZNiIAxOKYyVrivCfVpsrDREgHRIffErGPN+c1BZIjpBZH
W0GF4FqyIo8eliTj5VVbfeIO2fBEdQV3VGriSKds76dljvOU9wwEL6pC38OSoqSF9LdJV8xy8VdB
3K75gyd8HHB3nUFGibnKV3bO81itVV0mRGPXIlDCRuFgZXFGqYlpX8xvZ2N6mo81TwOLbx24ZJul
LVI794P4Jj5yAOMvRDvQ1sqweFLJxauIMx4QmZMQXRZlv6v6K8AE+n1IP4yc0b5m4CRF9kX0YWs6
q8CtXzGypAuYLQMcSq+h+nFYT0v91nWGDcCAEWCO11lnHLHnAwtAh32JxwOfvImoVRo8DeASVzZ2
oG091nX2edoT/Ftzhd0moNcpt3u9vyC21np0yZb4TL59Xg/FpcadDpQYHbiWOrEXzjNVPA+wsZiE
JY2t501dnHBVy8FEWF6ey0i1E3F814zd8ihXxaFQopUsxqrQzEZx4XOJrOyBD/EvY+HbnT6f2c3P
OJxQOFBMmnTVyXsmbN169demiSk4okPE3vN2bg6D8JdUusAm0hPJi67rXewLT4vRhRFoo273hTQT
sc2z2HIdEpZk5jScY52UBQJEVauo6mUY4W6YboJh5YvNhuXWKlLwjIINMCwiMn3PiJwCLl65DFQl
lgtiK4AUVE1MtotXnPH+TEuRSZBR3UcbvASaSMYcZJRsQ4V6Cve/mr2vLmsa+G4b4YPrihdSd9S2
+0I0KqSayLEIEEx3Xj1yICNSYL8NNyxm8ycSPR/mlWJi5at+DkfllSwT11LST9rcW1r0yNEB4+Cl
T+D4nW4lprS+DJhi9A5DZj8Fvv7oXjwLXEgvnwO9qhJPmKxViBzkO038fzsIk/3M0k3BNwK69aAl
zdd+2fYn2GZ5SD6r515hS9QcJZrC2MSjmM/XIOsVPq2o3aTFGRA3sC/zuV83Xga2mPLLt5eyAGEd
ibl002mi4e1UxdcKjkgbInPLGOsOJx7VdhrTiekZGS2FaUEbT4QU7/aMO7MYyPk+CfJFbsNQNzSs
I3aso9sHJo5ohLRm4dLxd2+suy8j6bUScPK3uFaIKmt9jL1CWW1ofXxHS49ea69mCjCwZBadr6rS
sTs/lFxrnKjTyLQz82VhR9C8xFXq448DdbrcmO4IJmvbEx02UwN4XhQkCcffnPAlGDGaEJXaNIUm
4tvmh3PwCdK197iIAf9nbWxRYIdUQ3PRIVpBqF4TCDq/bYmfEmKXZHpn5Ce8Q+X6+TVFp8B16jbI
0GeFszxDmnoZyuqsNQjgQtncL1VW4A33Lq/t/DA4hctQLJmY2EpEptdoUlZN/PPXFhhM3S9q1vOX
1vf1mWDf0Eb1NdOqFp9ezFQ/whQrvDFIH4eg51x00jnaq5Fbb//2uP1nVb345dfkNv1YGAZAxZ9f
i0HobLxsfcbUSx9AaXFwNDEBRCielyzULv8TjKUpIMXvUOYN7yU0rVB9jUhv0cA8lqKAPxr388EQ
/F3U6nVYBGmmhFF7C14nIqK0TsytJX82lOGkLEpIOMcTsrnv079OKZBzY9LELdZf9IidNIzJyMfo
E5QQ/9VRcbY+B+/bKE5Vy42GfbxQ8+f68h99Ev/r8uUQYytRuTHtU3LgYAAblzcyNTeL+9bnOHFS
LOpZAs+3kNjsRUsTBkLilgt+PU4ItCm2GqacxOw8AGlpZwj5GBrZPpulpUO5pI9YPgdiivROsGxh
bmq4csG7A4p60CkdOXeA5IacRgSb4c64SFl1st/O+ATuSSCOq5U36vi1fcJXtHf57YIwXrB3qr20
VWWbdBbfosCv7LvTwrIsgLL8aV8d/5UVIUky6rYnpI5fdT6LcRFUr0JvGBHaFqQVXQlDrR6RcnKZ
bZxviVts02Hcp71oyq3WkjTmR/40Y05XnMInpWaPcOIXnZ2QJBltstTzpy5GIWhrPtbWkQ/ERdzH
u8CmMl1mkz/pRHLZRnivf6f2aOneCwEprwzZT3yxEZ/llvIUTWuvfPc1U3S8nBvWOrmuymlvhMMu
7yQRfiy6izAA6wtuFiS919GEN2lwqLPRBEUvjBqJJvyYdMAxpZ3t/3FOPY3YeedgFMOoGIxMBFeR
ck5MdSdPH4d8zYc6s3u8wzkHxZAbjb1iItkouDuTcdTrdCiGkLDq71ECngekz0BjslK3woMnDgTZ
kyp2K1bKQCCOQuCnzIOE/4IdSRcDpzKtbsskVJOm2qfhSSstb51wTLed+1azq65r6n0i4Jy8LqpQ
NbydaHYgrbwhU3lTQeMZpc5jKuobYO3kaIOEwLQEMNrCwunZIJEjVSNHrZDg8tRRNUkpkUDpsl9a
vQM10nnNfAdKNuD5d35Dv2cmQLwfs3RjiaSJDiaRS/tEU4fFW4vpp0gsoJJORFKLj9phNKnmCo76
laCF6sD7lWQEkrj3CI34ziELWWkIkwxJXFSQ+VjW3p9aeJvG3i0ungJqQbtyKYNTkCOtH5+eTbDB
8wT/nfZoaY7JGiagj9Jqw/r1psrkpgLVkIaXzuImn/bcjhMt2kblpfA4ov/Vo9HG/s4sJ9j3SXmp
PnVKVRfc+ek036GJ1bEBHUJysmupNv0meONMYzJnI5M/HVxrp3cbxCsCqf/A47CClA1TmwTWIOVf
V7LMMz7YNGOlhCdZ2BYTQMko/wHioZB6Bow36Sx1DXvJkkp9myW+fPKif5654lFmnv5okyrkyzxL
VzH9xiPGnp4iDAWwk2urIXeKFJZ1Ft2kSz7IpcANj8kUSIefxI7Z60a+QF1bbVPYrXaRwg7uebn0
Kn9xB53r8DDE+6yjhKE2ZsHiVUJfQEhlbjTv16P3Ei9EczBLAcwklFfCMOsTC9PBWJ6AmUY3V2EW
kNvWtwsyslDmh9v1aBcip3SU3dNAVL+obnEgZGC8w8qbDH2mM6gdr3CuTyZElmhZ0VrkqBH3pg7W
P4XZMpXCoyhBieDPScyFpbhDzo1Yvvsqjaouo6qpQ/JI58f4VRPfkC6H+6WXz2UlGd8adD7OPNKj
ifjTUt1va8sNrXjWq5nuoUCuFlqt0XNRNy4uv60Zoz2P+q6Y9aan+Hm1YuJZtZv5JGGhDey5ENlW
qLNj0dogUA7TFoPAHm+GMtEZCLkHgvJBouTi9zsVK2s701Ptn0BXDD8AiKah2BxcK39puxNm5MPt
AfPQqtmxMikfkmcvT5aZYvkUYcwInSur6Olhr/ehhYn0FnoxW2l7Knk+8WLc7EjCDdPFLaRWVwrV
ruyTIiZLGagSL958QsImQDvOHfzWXgPIqQJ2fjOlf9H7rlbKyE8D8P1CfxuJ9W2E8NsXQc4c10a/
dJN9jIMVbPDvNEOmxS+fGlP35wLh46rGbQ+aJZsx5YLiM1oj9KwTRrDkbVCD+Vw6JUNAh2D7bfZ4
ro4xZqKeNYQIT9ktIgEK+7ujsgseEsHImVz8xwxuv1Y9F7ZDWMjPzAvY1yDaoM8sWLzZS/mCIhpU
u6s4MqOA2Ohyd6OUiZIIP/35tArZTiRyTBO3N7ZLxcPOTPGUonCj5b+3C7Ba1VJaepSpmJF4PK8u
uIo+com/H4EqigMcOLowUbFEAtNmIOQTkar1YoyHPzZuhUkHd5u/IrM1N7W3HvZutQYC/Pctw2RD
oqrrmIfSuB59Fzs/cGGd59G+oQY4dlTcp7bC/uJ/vEpLwUXBq3zkwDi+tSnLRJqfkFUqUHzXIUeo
j5DttrTETx5GVNqrTVxRKGw9wMxgNGL9sy4nuo7QVwBhZkVgZe6qyEMOSGlCCSA41Pq6xgjtt8qE
myTz10LVi5A2SnXyuy2X7rTM2HP5CyFaqKO7hRRc7vrElwRseg5hiKbu3DBUIkl6xAGLbECcy9Vt
0jdh3UTh9orreikTuxwR3rEJupQxKKQ/FQ19QVtDNua9rQZ5pSrDPf1Uwsx/+201YBcecX/SaAq/
WemyEJ6vTBiyxAl/Ox7UDDd+cLdkxQ2dLfdP2QWRCPySJ2NoOGhQXA98FDgDzwNx4q5kaFTHUW7q
JEi9J2aSDGR/t0BnCe485QDTxpZtPB90M5GT96HYZAMSQIsaING85xBh5Z6/gnGrc5VLMEI6S8+s
W61tbhByxdy4MBzkEw11STnWrgim3U94f4VC8HHekh0sBIl7nWoA7EEL4VQomD8fB5D1V3az6muc
+3TRjgmtZb6f/3N41YZWljjlm7KH/54nT3hCkmr9Sm3qX573nPvryvRjWHWJCYaPU9S9g303Yw60
ESOan1YFIjHbCWFeP+LkDkjcy8pBSWjrLRZpch1f1ebNiDjAd4nFJKg+NqzoOYE/Jae/hhrX28l0
p3THDlkTAnXSQj500mHN9YdtiCrL53zWjb9SOT5oQYgV/k2AZVbIrsENf36t8FKna5paBwlmyQmh
n5qTHx31f/63zHaLLmv/KYhcdJOGJV9Zu+3h2DTt+8a6IG5e/f7xdKWl/hhk1c24ZNNZi1duHCRK
qCqywgfrbeUrFwvZyxeqZ1gK+pcYCXlJlVHS0jjOAFXTvTNKKUKY96VfC1ebla6JSTHyAKH6hHZm
a0gaEJPU+y60iGWzh6+T19g5kjYxmUrxlU7I7xBU5cD1csiQuJIOChXjKg3o0NZYG1MDcxYARouH
NA0TYY1OXM0iJKAMGteKMJUlf57yoX3dH2+b27Jg0rJaQ1IbIQnv4tbxOouQd4xlP2oyr5z4nTCJ
fkHPzj2s3+wzsCs4wg9+IVfp6tbN38aN8QEmMm6mvRE25+pUvzSZrNnkljEKpIUyzIAjC6weW/Pi
PLH889+hDJIwqeC9qTWY/LgS4V5J7fBVDJ7KWeHoemJsVaIuzmRyo/s+BHjfr0MBvVcvy8EwecdE
kKbQK2qDR10kq8Lc61FeDGhIwSlyiZt35/B6XJz+vo9FZ3iV6svWj6qxToWiRLQv2Ec/3lr9hE4f
YK+OYaItvM7OLjzUQlsXgouq25j67juCsDFeBbhjLKrdEIbLqMhA/WgzoDKMdCz/w/qNWNdX13mW
JJl4PDqbNCLiATSJxWVW31WrJFmARBN9JnhV2lZbBnVOrqODBGg3cZ8tAhwX9lvaOsgT3iMjY601
KkNmqbV5F0sDLPuxwCG6PUgMJg2uN09Suk5+FDDC1nxWLNtscgJk5aPvXSfhvw0lmtw8YU73i3k5
1g0IiiDBN5eQEgYunwei7u3izFrQhbYb6J2xosvgoeYQbt59c5UuZo4B+Pbp6EU0S9YrqnWrcJJM
1qaCVcD5Gh4HBC2q+MFAIiewZybV9ZgkZfABM8jbXU7QgFVwv/3zZwxVxb5IBjYjYLMOBa637P2K
euhpTi6zQeAGZOHJfQCPB8SBr5zxyONAZmjvqVGf+Oi/qlL/ULT+Vk557m/oMYAspqWEqsAvVQLS
DZKqJjCG/Fr1T75w+1hau3TQnMQa4J9kkauDD1JoFw+8wO+XBDen6U1RwLsOGVVfvvYRdE5lOkxK
2xM5+KgYgaL3LcD73LorMnUurB4AdBRZwN5o7rt/Q2eBU6rViJoyg4l5NYbE8THzpob+mPbBUtlo
G4Pjc5VZhHGJPGOARunZo+XI2ce1/mvJj94aAGeSNwxotdDIV2M6bpiJlhQOvflJtfDqmzNl+H42
6N3XpaRuYzWA8sTnUvgPIB4IsAsjLUptclv23c0/0iylOGclaRZjFBVXh7ox/0MhWPPWebr536FZ
Kev3w/zc59WOcaNRkl6gtJN2MS7gqmTUpoUFTVE+F/RSXRZVJ1mwtKz2C+ohzeSRPTb01BgfpVX7
6qjwNIs6s/ln0MHCHUolm57jzP9c724ZE8cPj5DoPv8VU/obabYbpNMKu/cJHogVPE1hlATt+ze2
pqFdvmvxgTr6NoCr/aN0bE/+FGYiHRC4Mmk1tR2ARoIB+B3I+eCMGa40mKUs4VZhN2KaQSm134eE
lYsNPpcUdgwFch3dzqsRnZU2gPq2Bq61SpySoMKFPvoy3lEtaxKx/f6eIkNyizXZs1xDPQbmW/Py
+1V+14B0cuEV9TjFOQng6isFgiMYdyoZFZpiiQlhFf6Qq1Ck2Z25Qj/PwEZvYHo+O/g4BLV5XxPV
kkfGutBHanSVE97TM5ZFiDYNEJ6Am94cIXX0fraNyPy4gA3bd/Uk4XOH2lVmvjDz9ZNdh1cPyMRq
z8i0Hc+bcyj7ZuIgMaUfRG7lSOZR59dfx/zqS2B+r2lkeEVoJtmglRo/oGsyu7Xtlc0C3MbNLC/i
JJomyJKsAqeTks9dsdddpF8Er3kZoT7ko4+UTUtmTUZjX6sFDlkFQNkuk8jHH/4sL4Jsi0XWUnQD
D4pdpThEwRpiGtVti0uzeBGAZ7yC+YxPzhTOzE5zSLLzF9WgjFPrnNKWwg8SELWItJwmIHxvCuNM
t9fSMpdhQ3IK+o9204QYj4NPTEaRvQQvKV4RVUDsx7IUKilQ+ZY7ywrl+69OzG/ooeVGsXn1ZEjQ
uQVanFbJVGfG6YsSQ+hbxrjUvipOQMgpsgwPq0fimpYDrEiN6uaJ7ujXn6IBdht7+RYHGN9dLEZ0
T302SWlov+9ryZhcqSjx2hXBeKF83ddfdUvmjKN5v4AwgIc/Cl/54bTGAEm9mYX+w5daoUP1B20o
PuKdewCRhtbqJtI6K+JtKZmOaUYo5WWhX5ARVT3PtDBFvDTcUoHAL4d7p59vVd7WVeFRMSuFdZ21
UN4T6eGjF9pXhAwUgarb3Epdu6wjyUnG6OiSqg7CL7fS7oixcyyYcxX3rlLjqbWXMHMjGGVt+H5Z
pRnMmjIcmBBqSsiDsUBp+ilyScSDX0wYE6sFDbrghlzsmjqYOcxf319RrZCpuzjs7W6KE1wAJcuX
ScqqNbNyNPrTERRunPnwkxeybfkccmXzMwIf449J4bZ1yFHvQjXo12XHps+jxzqmEHK8xsMqfcil
i9pkv+1+lqkQvbwepXZ7+4NssCwTLp5zP3eBJHZohm5mCQhWYWHL6shJ+kEfGO/xk2QlQ0RAQVN9
y85YijTNhPx2NjvzndSH83a3gpjIUVMMONha/DwvkxQGoS7iEIdf7eSHkDLgsVuFCMTjsbMB7lTx
cjXfYYeZlaIcVIAux26yQvwHZn5mJk8yYzDJiGph4/4L1GzSd2xZD0PV962CO+41mT5HvLfXeTUa
GoKmMPpsuPrPxrRcc731/9xJtunVRqe42wtD/QbreTOpssFUrTZRzpEQQFMROxPX8cbUIBt+IgsP
kJZF07aLohJ2HWBrDgYQfs9b24c4Fmv6eXEGFdfF1PKN3RgkAQS6d+skkbeewI5Pv0xc/X5SUNHV
Bn/h3WgAC9/OnRkqSxvIG7SkXgygK/XyQLPEd6eY7Ew7879hI87Lk4PD7OemoiqJXCCdbZ8ojfnn
UcwYPY0P5vrYnBi4MQM8fGeloVFss+b7ny93Jyne2KXdtS+Xs77XWWND5dJiEnITKKIcRcwXoqmc
CANKcZdvZX2cyj+6YvxaOzQca+HIZ/92zkE7ZMG9TO1Az9IF6q8hMaqAQweY1viaFf6w0UC6y+OX
xM8BC/TYb6nizoW+phb0Wd/JKiLxeCfidwdKNmdBN1e8PqT9hgn594HL8p2I0t1KJl9TwD1Rj4le
Xwq8Q9wu54+IGzTK0opFS0xMaFrrMwO3AIM3RJj3auZkyUBY1zj7gUx7av7tJ2zU/w237h5GemHp
Z3R0bkvGu4ieMVuxbQBmNqnwI5xJORC872gJt2cpeEx/JgrnOOscw6bEkLGh5ynncSRB8ftyl1HP
O5qRuwgQ2cTSxyfnKm/EIgYDX785kuPpbdKhgguI0WECKwRD0+vBlaEWmKc7WMbEs68/0GtXkuR9
YZNWPldsF3pp+BmzDtA4ZbqhKKk7QILzX7ValQgqoTo4wulVfwSDSEGI9TpzYIrQjiEC/JSst+Sm
qC8PR1OZoxWJmExAnFMPcZDjssryXiN0rtrgM588+6gMYHoPC2cl/lFXXHglBikxLjcrJyUUkpyW
ysnPdsoyLKvstWGMxwJ2lzc7UYycZB8V5T7KXa9PS1Nox3yIfYLfaQ3hvpxZDSLABQdkB2tU7NKV
M2Esfs7KP05xMAoStuvOB/QMv9SK0DfN7lniyjh3JUs1YPPYvUNNWwVx4g0UL0yyJH546NFJ5OTJ
p/rqd2V7GtHvrBpKwl7KHt1w0a3hrSuZNfGjrp+HqxsquBFAeK7Ac0/LE8EOSLwjNZ0vPJYh2ZGN
KjoQ/+urFE+B63yDrh4Es9/r2t3Bhv2nLZbAkO0ZTiex7sPnvbofA/EYw+jYoRzdxmQZjNtCis9K
6cEAr/ppF5bx+kFFifEASovv3vlGiHMPyhNA3IT/Ypcvve2j/G5cuhTrVGs45V92iFdL9EztFqhe
IFTsoAzPMuqwC1ANmLVhVDxZQIGymroQFBcTM3CgO+34o1noJ6gsE3ZgjO3uPcTibQbpGnmjxm/j
9fZQdU6RObLq/Q2BreyvL7bp4uyrT/N8fQwdxHr327xd13+OAPQ0Jm4XwpC0S09DQ8cmmxUFAPUl
zB2QW8rZtfkEDqvfoYWvmLdDp5ctpw4jo671Ow5U/OupLXHbhY+RUZfBJMQC6PhPb4oCCWFcK0tX
GPN0OKEFAxmpNLaZwGWlxBSWgA423GquMxQidWSjmUa1wTqKVy6nLrCGE15ULwDGuOSVQ+uo74Ax
7+2daAoPpeeuMhhlTaomeVzo+eyAYg9cuVUIZJcmiaPQeeR9I0+ZCbEZKt4ZlQi1YIJsrkdhyYgd
gH1TXzmk1yuh10bNAwuuoeYZPiwwgraejuMP4Um1Po6O3giYLpHakj/HWkjNIG50KdtfkaqaIdg5
1Z+aKqM1wH0eB41lRaV5V6j0+jG054HC6HD6Lw2j9FlN5uT69xuix/GLgDkKDLHU0WqNo4z9aPZf
jkNlYm87lAfFWmfSeXZMWO+UX5a68xyWh4xY769zkPG7ftDRz1BZBxCgr3F2qC+JiYtJZ5/pwYkj
oX/M0s+ICnsQnDnk3B/cmDsu2oOE4EwflE8ETj3XQEF/+aCzpLoQhWYp9/K76o/uoGnrvZ0mSdc7
TSc5wUOyuR0EULya0udgB4ALBi0ovyaX7hQQaKQhqgA3NyexnwbqzVsPjC1jwZGKg0+aPAHKMvEF
MtDzkb9EIt+VwHBQ65opd1QeVro9xYobxEwjiofRhcKMCw6+CNtaPpiQ1AQjuTPLtgvVSd24mBD9
dCzmYL7s3dmDJtA6vYUw5dLrrWfIsyop1kbqz+htZJ551B9SDXF+ZKd09e2EjJvATauw/lUN+tdL
O0uPTyVt+FlWtiMRM5EVWmsDQy4N5zhERPobzn6QYKVjSrh0UPzdeRN6zLVzlrK30zA+AL4DJTdl
ipBeBd1xCweDs2A4rLJ0es6/Ot4/i4vRw/gFz7/E43dwAdYaMkKT+2mwcXjn4nWiRUVyzE/eI9+U
XKrmott2NDh4ZWgsYQJ7y5nUfROUHXn8ACDLB8jMjJ50+YUl0Y1M1/QVS3G+0H7bZL+Udpv03mGC
xtnMbJdp2J1O2ns8EuOEc+Q6mtQMZJiyVJCoF2gMWubawa2YRwMIhO3yTARwZBz9GJ82rklQIdcg
V7hDDz5bBVwp9nB9QU72IvKPySRB+3i/2FYl8sA6kuGXxTt0vu/evpdiSKezcRRX/UHlD17nhSIG
Q53A/cvavWh1lRV3fr4fFzjRlXC7fHeMSoO2Soi66mtObfAuekPm3EqpzWlReBnpJpp00IXnpucu
thC3QmSymyGAaTRp4GepfXuING6EWshrZYoMoO+7g+g70ZA/oeadJf4cS96xJOpkWkdnFLtDaDCp
PdoNQ6kGxDqR4DwPxBf7lhQoQ34aTDIX4vusE18K+H2NmJklQvXmglQZGo1TBWJKlMb7RghLV2p1
OHzOdmdPA/JiQgd2/09++8PSOh93zRDjb5k14nJV1bGqcKW48nz4Dxdwo9XNjjpSKcNWVg8zE3CV
k5iABpZdToQjBiFa8Q+erfC9kb63alR+zJTySFLD3GB06KfY6RJtNUlRMo8y9qxnlX1uunnq5mio
+oW+Noo/VNC2izp0uuRPUuG5OktwKij9ZX7PERD3sbusxxtquTJyTyFjw3bgYH7ZjE+XSmRbk7bi
PQeOl958O4MqDwrFrbAZcM34SZI4yS7DT9SF49UKbxTwk2ydr7/p/DKJ+kfbTuUFR9oPjM0jl7Hv
5zRKPI32mMgc5Jz0DypVkJ1clzmDSSWp2/7p63Uh52wDVu8PORzDdDbFK595YDErKBsSVkmoY0Uf
8pQ/3qnY/Pqa724AZ0My5SysXgEkIL5+J4NIDXjrG9ADouO/1Tjp5HQjarK7nlDIiQOpGjlYgtSq
krCvwLwHaPZ6ypP8epMGNxUFodjczPvTG/UalmO7+H9ZGKcYwgh58KJIj5uAXulpROjmRGyuL8ym
pmYLNeX9XanMM0SyJEW4EW3PMjtQbg3OriqlcB523uXgllU1RycOekoTnGdBgkZ2h1jewAcjKEpI
qpomol0/1QKgTwI2TyjGtTvHV8y0AtXlAs/ngHFbBrjPA141sYMoHPgOLVgK8utI3i30dvkyp0nB
pEgM7T02WiqOZI/PsiYX8Z+4biqi843cSw21GFRd3xi95G3bzDv1LONkNeh0FJDw1bWJuAvgfp0S
wrYbwUOvMfOe7LfR34IU/8Y8HYwjMCxB6jsarNXnv1tY6b4JlT0Af9867L8ySUcVVpbea+Y4+lDL
pDY+eJe3+OJO/Kj8m/eWubIxCu0qQMjMyzdPDQNUbmQyZtS19fxwDhemGoCkdWuyl8ima5Ah+U5J
4ywCb7AL4faSLOy4N2awh7fDzMmsTatk1TAf4Bd2czvzXlYXShPGX4QpFmcvTLcNubxwOC4bQQeI
1quMt5vZv970zuEIPRqV9WzhgX3BOU4IC4R8znLJfTNnFPHJvGNqaA8fexD1XHFQjNmch6GS/1W5
8if2WE/+CtcfumK4AU1GI9zHzfn8RY83cusLis3aq1+28jyhwYEJcGuK0hfMtRkGR4BhnInIubFx
APr7skR/JIJA0xPQpe8dWngeZIpaccxzmuMVhxfHZFoj/SaTqdh5A5Ywrj/MhhU/OEHUeq5Bs9Vs
zYbTVCFGPI3IlUTD3KOX8HvBa8HnHNSLF5R8h1szb+XbA/XVlSbo156mO34hsOPl2JaJNk/FlisN
HRbO6Z/KUNp0rB/2HrFoDbfVuDZF8X2wj+aVZWUDTtUG/+D3x9T6TGdVogKH+zDaWz9emrLzr+3N
EHjgIGxTOX1awlUTEWrLOOPUEnybq93PbPJQmsL30bj+PoGvwPXSvhtoQXKUCxFe6KyPfbNqKwJm
dyIRQbh8SK9PrWheAdMc7K0UFhK0dsumJYwN12GkkN26osaJo4SBSzEa0mKeIbreYszYo/XYmL91
G32M4ePSnwlo+Qclig5mojURwlNsGcxPSjO74niONDvGvTPPenIgA3EsFbjtU5qUtz6U8LwUo3Or
ov79c9Qe6gVJ5klAlUzr5hrM6E8yGyu2Hr/YOMXB1L7CqLREOcRvAHhZeIn54SHOfKftN7zMpDJ2
ShzoUJRH/dEzf1Fsr/tui6Dcumx2S9HJVYKzCguCuVMPaMhECEjYbf/ew0a4j9/byxlHiybyfhbz
gIeflUBwVyMZ+N5p/EbcH3EmGzjoq/xKsaMw6X0WCZNdnFVwzzU646dZNYcQvQp48Ps3qoyicGmH
F/E61Z9snU3Yq0iEKmP196s867xwCtob9nW6LI9Cx7wH9xHEZRHnGbC5XMprqlYsyo6E+GAd9u39
vIcUFHSMS3kjQN95W1sfuBxPsVhrBOZEPi6t6U5PJEygymqLrxJI23CUu5oEyfy5mqjE89Ohl3OJ
1POiXZmJDmKM1J3/PwIJZelY0CrYUR51QgESE2W/u3CY9kZNK4R7wGhySn2ryA0VH/XzEJPWwiDX
rGHjRdUAof6wmi32u3Fk+nSx5x52jN7Z9mSFHPyOuAWxAQvWQ+FcYTji6oir2zW+eICMrezovXyz
IRLbp+c6RAXV+pgWDBDqVYJOdNHF5dB6Sahlb5Oh9N1G0Q01IPpHHLyVmD/AnoIzbZ/FGILyBBcm
mKpmISQrmLeXBKbjR/USwPGuT1Zy3T0srVQk5MxBO3Do11NbwoPvyJbgmjvcZaJ9oZ0zPT34k7z1
UcTLVp7bxbeKo+JvAA1m3NAhjEzMz4gUEhBw080VgctwtL7F9WKBjAKKspnsMKWW9efnZ2N91jCi
tcbYsh/kTKmMjTHCH3XTx3hiZUyJKrorToSv5uel2QuZptsuci004rUrCzUKwYnMN4Ng4Lmci6PC
FBPKO8qr73RqCBl7jHoUzZkROnAGaFTTuUxdbIjzq1owoyFdU/PZ45FAbRM7Qw8cP1Km8s8aesNq
Km9XLLDVZj4h2U6drvadaQfhWaxCvrpEkWO/6yh87RjzLyHcyQzzGAX6gze+Pa2FGxp6l25PU/JT
kSeGe7cTrAagrZGvGAdb6SPUxNkrSD/Advfplk9lLsI/rbKGjmLi3jlvxPEjWYmF1igL5JtCd7t1
3N+5Z6DkVG01HemFEPvO2KkuCiRJIc41G+/KFy+nAjhWrWLGZJitCjE7WIb39TXj8g9nNt+t9nSY
SGN2Y99z9ocfChbldnj8OuUcPDY09zu9THg7Yz+asgoRkEPJ1fCSyqgimPeCIEiHZ9Of0zrgsN7c
W1+2q0+tzbP+eEpqvtJABsj3naswcBr0eVxV9RPAp5LOWPxA0Gvy/t2GuIqdz9HWEu217pOdrd1F
ugiXgLxvKTRBADTqE2dwJYTzPjPIOhjoQEmWHIG95DV8YPXh9xf7iXoWKNaLWzAYAyliWQuymApT
Vf3BeNMqlhevVCZlGBE4EWvdwb+xYlIkCbMGA0KUJs3gL+v/qQCtLYWTQao5d8/Uc1mUP0PGzyaP
qB9hcuvVaNiZeJ1i9QEe49kGrYHe5h3mIiUMSmQZtIgX6nkYgq0502y8VL215xM1gDLcEqLMscI5
TXdZ/HWn3x9RA7eITA5sUCD0CJRRYDESRVyOBaqYcpJkqgiFnJ3Ax+wSCcAB0EM4UylsH5xEN5B0
Fd4ft7CbZ2rvx5kPus9thD8I9Qv+3qCzpUMfPovPxnolZZYfIRrtEKNpKLr2oLVQ5HkHjDsY15TO
Tdv77jDih48m8+7aps6kI8sH6nPFIojaixjK9oUFTAWEtz3SC6qIl2+crn+VKG+hd7AbKZSw3Cc8
o8bwC7I0aUmfQBBT5G0oLkd0X1vPe3BZtwkH1krJBy39/WTUmFkBnomavkDlahqsz2c71ZrinW32
EswHldaQNGr5foUBeuXyn2ZpW+0CW20NaG//xHd7TegdcAjiC+uLn4mvzh8grErlFgd8gFM9MRll
UdDbV750PZZr+kMO1zGk1DDkat1MMKLp3VrnovKK+c9BFuVjRsE7pN+eOtNrXGe1SD/nJOuhHutd
nK1gWMYtKrbNkVeuDSHwGDidNZofH81yLCwL+t/1qJRV/gTQB4LF+Guph9xeuh4G8f0i8OCgVsWS
8B2LTgU9STQYGdIBqUg/+zexV6wOsMwslRul5GpLfvS3oAUSdCE+a8N0aSmHnEInObcRXORWG0b3
hH1nVXCA+zGADsY6ELueHBLm/2/ltAG1cloHEozOBrIkqtJKXpVWwk/DvsEMBTmpxiS4WymaINYH
AgLxmdYB+vTUMLWsXtuEZR2lx5bjgasd6wlvgfvnoMtzLbA0A0a6FHIvLtgG1xMVdqMiw556l8xU
s8HTWVkpUE3ieBTqqisXEUfkud1cWBW3wBF1i0SoDEXunhaEV+5/chOITYX5+8M+Ky7vvrVNPIpC
lh8Y+H45/0MvtVLdereUhs60y01/brflNHtlOLYRmlgF6TtB3HGAVlo/aZQFXI/YXClYfsMBlqNC
bq9g7MFMGAdqSqdB+PxUx140mfD+gD7374KZhtqlH/9VUX98QQmwW3XOmyCFnxRYSyqoS3srmNOA
fnr9Xuf6OAQBwOOkH5FzAs/+Kzpi7qLgsYjZORw/UBL329XtuiQ96fnaEdGatFWrW/HYJIIMyLVU
faISshv4GCe2wrSmzFa9xd/9tebp1B5rJhU5dyMSogAby8zovYB2pvtfgNWHFhExwUaWa064kW1X
si+GVSeg2RteTvyv0cQgvwgrUf9iAa/hJcBhRjR/WXJpE/RBfIHDX1vJe4sQvWVFnQJzanlnQ3gF
9+FMgpDngMrpNvGSvnJfWmzRLGm+ZHbctmpcBhz0dxTlrpSIOf67TczyQh0WEKnw4dx5DVrTxxpB
+sik8ukJlbb/SVxPPUe2fuVSRT34QxhUyjaN4+6TOpa3iz1oIeNHWceI04Vtuwd8ezFy8TT6eHJO
BmUj2kY5iMVaRtEJRUU2knM/P17Z4BJohwPCeiGZv6TTfWpgwWQ8lZe5uf8PzJ3pH9TMVzeYKgHo
K7aVuSAQda+LbREFq0kvrbnwmpNm/WfeCRrYbEYDZo/9l6TWfiZjh00HMhZabfVur/FFn2gzsPJM
HG3mjfR+PlrAT2xFDkQq5REYvoD+mIX4YGl6NO8R7rn4+TLBY1VO1j4DBAsAI7g5972/tVtyXDmA
g7Ehh2DAkLgNFLZL9dIooRiZrb0QU7kPlSis72WPbXuWEEnI9qBocDBhKVm+2/TeRo7aqBo3frg4
CJpxJgDQ/RrpZ7Q5YQSXEzjBpofZWfkofibj9C+HRHI3BCJti8L6B/VBTUdTBBqjmDgVQjNkyrzu
sJg+633tj1oWir9rATkauqgrXRp4j6jdgQmh39DebeYRrZbq4VO1F2A9bMXwKIGL6kA91GF3x1Hv
tVr4iGaeVxp3bF752yobUMf7TqNPbagdZu7AsM5RtQPq0kvtaP1XrhQoUQwFnaDL9d7dwieiXzqh
xSbpbqfKZnRm3WrO5QMIfn3qrjCTAUIHm6Z0bWHyE9ng7mzw8ti5sWeX9du2uNDQB/Ts0TouPDs9
8BcOgGmY6b8EN9UbarhllZMHlekEiMKCdsg8d9zpJfS3ZDNRbC+bT0PCIvGk1l2/MdjCHcs1gGbW
EWe5MYNeHOhaJ4bqi+8Wm4HeDJu43fSclcOQml0Gg8/f/O3YiEg6/6gs0GW1wE1d4+0Yh1w7lfNu
E2ZJQkwV7VS9rT/CWGzmzGsOzmx0OGiU64gm6Sd3BGhboVTyc7f3XXmvBUtXBAYFAZvcP1h+bIrx
xW/0Ty80C79R6yxs/bG9nYX7Yhdb6z/5+0o28aASdBNOcKUzoY3airVW4GOAhJOAPi2EQMp+oHZS
GgSSfbRou8nHljyYcqY4+76a1uW+1kgTNKSyWPNUadH/l+nmgOdjFZB6IVH7Hxq0mN4sB3DNpoRi
aiHFsL1bImnVfZc1yTIWvhDJn7zMmMCOtmBWx2ccjFRsGRGwW5MzSfyNSawXow3GgV9Hp3p4i1Pz
MgGyxC2TXrb50PSPnLCDRnXHx0EWMvNU8z/Sp0x6KamdeEX4EI8/4p7OlOE4StXue6x1LtXFcApT
bvc+c58PACTpQ5CPjqB9DJKMBRayRKhyYDRqrEPPZT6rbSUxesUJQvqgjDYtnFK1LS6kyO2OhPy/
2v/5wGKrXRdkFJvt5CGOuH2EY5OLcZ+A2aU/1EfVKJKMbui9uaryp8NDUu/Awl6DtnE4THm+c+cV
rdUNzzsSBPX0i7lw1mCcrgnXYTNw6q1nL4isyt8bFwIYenRdZmPnbiAXpzl90swgRMiJzINqeLiO
tS8+fvUzj2ZwY8KzqvxN3ZT/DN/cAbsxi9g3WRHk7m5s/s3vHMkc1e+m++a9WEv/VvORBKkijA6C
o4ZeyLfXtqKjMLvCBHsUS/IhSQfIE0++zew/A7ttzUyREhlnzP+a3UH6F9itjH/VJ7Bvtzmt4IIZ
esgoc6XeSH9b67EqZqjr8ylOPn/f2rGZhmJEcdY5c4xg+g5jMo6kHTgkK9plfSP97xOFHTukYoes
vs60bU7pyqgdLiR3n+XYBJNt59ebMkQYLbJ5HoW0eHQzaHAdZLVHsMDjLEjgqq+GoWw3TWN1rOWQ
qy0mdbCmTAlVCZS3LWuPa+VncBkmz0vDZN1qN5ls5DSTs0LMJpWHlhxoKhZUlXjlCkfquEGDyPU4
rraoYQZRFVQWLSoPjRAxKailGhSj1Vh2bWdy3xXSQiNah7jZtYovXNePmkuK7nsdWfTO/blRD/Wm
LEfaqNJhku9LbTS/mWLTxJOhxvbyxgJa4S+3bbD+QSYK40FfKGT3ar1/Cskmt02nHx7LtTpkrmy4
RvIUwe5jLWO8DcJSdlJ5+lv4Kd84ZJHBA3L8bjeq74jhnL19zqLcoigBZqnP9Wg1j2Ov2c7b6eDU
pdJcwAUoFkg9ypJu1tWDVLu0wJUHlkkz8TK0tfUETZ/NjTb1YfiClMCkjVqs4qok82dbNBMWBOyR
8JW/GmGZdS2h+FqJcjdfVfXQrFqWTdt29FAumqhCQwX946No/R9D8B0nl4k12FwEWFPjs77M/HiO
ssiqSdjOU/L5ZQdgDA+NMZBRLqs4KGvMd9B21BRe6cSnDaG/gBxoCgt06pWTvt4prFmyE16KHgev
Eb1l0VAlNmJfZRysCyeLT9I+LvkCcum05QNNxrwEu0sg6D5y8cY+f8qCoRHIAoSC2EXKdW1I39NO
qp3ZK/NWmIwQHadaCeOCJY+tR/sAB6h+WXJK0T47yEcpjEfPpRFCXGI1gAEK1yJ7cG36I+ecc1Vw
R7D9txuiAq4BaAyDqz6qlsl18MV+xyGdMmpAxo/UFzSDzF5/To0+YgY+pFoQfI3loJ2QHyNYJrJG
kHCEHTvacs9fJQ99kOOGCp/w+OF/V+Jsdjm1LjVTpZ3SjdhpcCQNd4mdku+hNDvlrBEesn+vi+yV
5u/Q6PHVoVX7NrERG1TKSCEuI93BB+ruOj96Gklk65Hlf0NYMSAFlIu+1CGmMQqkVg7LpAOpWHk/
i4VmTEhc1OICli6ovnKAEc6XnIPkm+8KvWzXKNqB4fTNYeVLKaoPlkAbekuQMU350Qm22CXuCBIV
3bf1C5ydguc2PHMgUR8QWFVLaUcUSARb8xqZG+nOcRyLgfzsQsoZcerdT/rlHMiYw5faEIK+c+95
w3FoSaHa1QT/445QvJNfD5hClo9seU5uTuoTViyNUqaEmH4f13SszUbuM+ZAtMSETnXPnbk8WaK+
gd+FXveAB+3ayVWR5eMF0KCuNVjkiRqPaERTJnwejYKHiyrxkpU/Inpt8M2b5bZ2IIWK/AvXhh84
t04OHmyUdC+lVibiQiehNs/fbiPjmbRSwoTcfTeO3mucBznfdB9ulFcI0T2LnD7N00Gx20IZ226K
DNeJGhLtymwHWymG9wt1dTezEsW90iqR2nm8ixvK7e/Ca7/hBaTxxL2PBA6srJWA01apGw89NMf4
CwmH1omLBA99G6aTid8BNXhM5lulU64FxIvN4v5RT+OCV+w2YcaX08WoWNF9EzFnhmiKW1pyQ+ZC
r4OuETucEJIIy/M27nIjEtxMGGnalH+1vSJ8CcWdpMhxFu2yVXeXryeMzO/Hr8rnrYNkXkl7/9T4
50Odx0dA/PxDVUcrO0VlhoZBDxK9d11Iu97L2dl/LJi9rxdpaNDQHMSqCjWlgJMFSYWaliIrUy4O
Oo0+xGgmU+P9wyn0bRDWliRBT7ODaUE6mH5m4tryVv/6SpnorQNr+eELhPVJVcIXQQgmuxwEkgtU
0jIOW0bERSaspS8d2yb1awZ0hatBKP4qxwC2dnJ02PGSC1R/AOwtQE1KMySDqNx4DUG7are3eoZf
UwlYlVtEB3DdfkbTBS+faYLivT74SLbDFJOb1AaD8At6bHYe7OH8/7UpohpUIL/q3OYyBdxfhxO5
/IqNDFaGqFenlofp2SoM6WooH9+2LnLwknVrdQ4Te8ymDJGFrqAkaZB1vp2wLmcn4K+b5LgfGaWf
Sh9eZCRfugYg5FyijyHMEGC71TBGq3/kOns5wpHfsZ6CGUkHsq0Wjqu8VEK97Ip8ksV05VgtT1Ia
mEl6/6gb+jVvs9Ifdh9eqvXqLZinlEBd+bz+72yOPP1n6Q6nD6LqrYCYx5RzITaOkIwc1ZHKshFM
xzKf1vE/ZKDHS+XssASKN5/pwG5stiVFgBwQMGs1TP13Zni+3FIyEWtn4NMZIwjLWaohF9/Fw3Cd
jniAg5vhHgcj4zvXBtBO+trZNWi6MN6bqN9DgrdrbNr/iA0yF7qqSRNiG3HQQm58oaJHp++OWy3y
XuiE03cW79gaw8a78YClfh9KevMhCzAuNFCY2k6mf9TmK7kSIeCCgGTth8UTgyPjqWIPmg1bIXM8
38EGbIrdArId2DvVoIRBQTBfp6qjTenhi1IGiMIgYUfh39Eoy48K19F3gUDGmZNJ1VF1WZquBa3/
kC6kZhPjzZAsNzPOiziyl/el7BqQsFAKBuSEldqe5f/BsZmOjZGBM2kRSQo83Xt70Pt1wI9pNf51
yjmh60+mupqvfTpu8ts1hhutUG17UdlUKsT00Lb5cxBXhpfOcHm+2XolQaYuArdI9IB/Qi74WznC
M4OY1LXpY8SZbdIJPym/tsUUEG4Mu0VOQvS/xM/Kq11AsiyhJHg8PwkptQdtJDvFIsP3c+wKAOyS
a3Yid4SGREzrrgRtimJANGjPZtAK4d6eS8c79Axekx5ZGeyGSp73O51zMczcqtRtHdRE6t2XddGB
bcZlUnGkhIiG5UWFa76ACF56UDmM6AmAsq6Dwj6J3egGo6PTsDadXJLBP1P38NOKiWjxtyjx+nxt
MvwGsYz9Aha3Y9lpIHehz2OPCCb+yfDhN6L6RXVUfdrOxdhLdYD604HnPt+rn22PPdTEVMy+/Hnn
71JDbVkscJV50Nb74yq2sc3HbbyLVWjCvp7J7T3hI/7jmkKeRZ77GDHKEkZar4RVpiuy96RMsi+z
gadTaPYz9V2lPPOTCYItdP5PZPqJHH/cN994KDiE1eqSOJygzhkw5xLKhPc14z6XbGIsLCyyTf7n
SzacIbi/93oB41tk3rAEi5do6Hb5A5OR9qHLrCrObW16/Jp+eyiJYBaKw8yCWRqyyypJRusmoqPh
p1cXGVisLZq3KTL++7Ysw9IUDu99gQGml/DbnPCgm9tlWUxGNNPNJE0O/78Hu9Hf7ORS1aeuTvEF
m61UEyhp6x0AbfLFnkfbLAavdQw6XWV9LiRvVs32TfROsR1lPL5gEZYSkkbHraD0GmQPcFItgyvE
n8Gl/1I553pYtD/tsU9Xki4Y434p+yM9sH7PTLQtAJMxd86PZFUQ2AsIiDHIZ2ckDoIzp7RzFilU
jBcXraeKeDxJ3ngAygibjYXwWKzLvG0wQPc692nD/1v5JPm4jOU3IZ4NLKnWl5IVxjZto0jhrt0K
fqVLEVIzXGPGPZpQbu99GjQer24B+ALBhGPHOSJXC3Ae3dzo1b9pD0pDtmnmROh3XUujHu7yHIRZ
tcdGBR0Ew85y2MGVzDEu3PVIWO/GA0M6YjTENaUhzNW29jtyd2TRBUjyKZYpEFhGAV50YGOBsxGR
x3qd1k5UMVdV8ml9bN0Mxlkevbq4DBZqaotfTk98hmQDQhQEV03KDyB/VS08I5EEOpee24SKylxF
IJSYlbJqvJacu/gBCVfiKREkyaUVr6x/NvKTIYpXy3fMdyXTp+2IQKn1jgbK/pmgaDyrbIIgqaiv
0O/+Rd+kMCUX2UbVxcQyDOtsCYL6PEc1nIsqB8Flf7MpaG6lF07nrIhbcfgVAZuyEQbihYsGBrGw
wYltYkqxQaW3OFdqAQ+cdiLAWYrioOl01vuhR182mkmvNlr0/LDxaLYt+iPctkXyoTXVF0IhRSw7
T3yYLerbIz/a3FtMgdbyTdtmq56dDYRIpoiq+uMzQOkadxck4XbdjmyV1/oQtIk09nZ+zYN507XN
bhOLuNZ9fgyeytxtN4u+iwbr1tTwYBDxywP+XAlWzfdXGjjJLNO6YsD6QO0LCgFEpPsIl45zA9NY
gLxD5GEqT3gPzFsysBRSBfT0DggXL11UKAV5um0BC440UZ5m4Bg1krlX8DhmMGKa5OtrFGRySwA7
saqLFHcZcUijdSJgcfaIPnR/9yH0OQ/kAQG4EanoQMxXkqZunXy3k/coBqiqdgLBwDjTtAu/5FFB
iRyxPMMA0VvQ/m4AErDSrMZg3KUCvHZSSrCJIlvtoaxNnehw/HpF8rRqFhC8855KcolTdZinugov
cnO1d8tAMfAkSbi3hrIrVMxj4KcQeQAjMK8kBjl7jBG8NfsEuAdlAP/hsTRHunKYGByroD8hr4dG
2qk/u03uaCuoyVN+OEELB+D8W/c8TsyEQVeSIgWMsDup1AxnYnvBZhsfhJiTOSIoj1M2ZrTGkDBo
Sl+ItrqK9VUZNBr0/13f2yy3IdQibo9MDccOteYJwBAgw5eUd9vjBvs6SlvGs6zQyeXeEPjyT55C
UPSM0brCyCi7UdaR2lP9KlPAP/7i7MncMUPoJW1smBLyNPcvaHhh06KVhuXh+jDJgAqrw80KK7+C
mSgB+7DDBNc4Pp1i80zmuHOdcad5L7Oeho8NAe/hUiOKI4bs38BFR6zhbMAHBbU2FRTaqy0YPk4z
1UrZffLsuBb/YPksJbMHOeKZjxPcCSAr8EgDz9Nt4yXTWuMUrHpFSeRCeNtbCmY9I71pP9QCuuR8
pQtbsv9RmhcgSsrLBqhZ1dwOgQWiKLmUrZyDxC8Je2z9YoJt7YWIjByVFH2o1EV6Atqrfrv/zQfJ
e3a0AtVxMnjK8PPYhWMsU5PZ/QTDva1/uNmeXXwYmkTOs5l7Ufehv0M8Teg/vT+APbW1Z//4604X
9sactaMJnBF5VguavqRxcZWbPj5cxHU/6N0o484HFs/Zp2LUeX2XExoSbVs5yMhnnF3ZUYjz1PWI
xE61z5DLWXgtpATkEhy/O3tSwWxz76qVshM2FrxQTtcwz0nVlJdu9ZzZ83zIQXNIhqSHZvr03oAK
pYVX/vhN2BRT2wW/K/EZY7gzobmY6bNPLpCTCdEDtP6I6Onju0wTeuoZqgyfJCetX+K7W9kSx0tW
t98yr+edpGrxaHo27KHjvaQoY/7K1BnL8o/Rg8e4hWMO3MQj8BgzQkCWtNS984mGbURLQq83mWX/
WiyZBXitZoo1MPQO7gMC/q06Mwy2MAV/U7F6TMZcvwj2h3UoEX3Fjj9YAqLjDP0r2kw/HDIx0Sn1
2EVr6E5a0tWVjAaXzlHKkZriIlDo6JigD/Cg7o8qdyoFZrcCKBLgmypR1r10ARGUoWhdw0l9Agea
ED2DOzYmq+GfxZ4Nhum/WHkaXSLNQyW0VZQX1pPjj9tHHUiyFVFXVJngkG1J7OFwPt3RVtzsPnEu
tNRvxNAptD1vXDMk6/oigFT/pzUGodb5lHmmmc9TF+RTOTYwFKY3gI6LQqg7j7KGbr2V5RVgciwD
ImuboEjgAtQ9BtoadSBtAo3pEFCHgg1CD66WE+dRfO3x8ZoRexhQXFCXA85UkkDCUJoqvtS4sTAB
52b6ot2e4tsveOtCuX8AxeQqnYpVaHVt78977CsKq30GDesPgq+YDNrdzCWJS7i9Vto5BodXdfPq
hCIWMCjQzLqn1rBxfgAD5j1fLMT4Gu/x1XvXEvxLXDFfxaEg4Fam6jdPuUBtaMQ4+tDGrZA9xFo2
I6ZWDYANDuO2n6d8ECAuCFKmO2rSANvps2EnyMe6HIvRhKUZPDZFvS9Kijql5T50qX1WoSay8R3G
pMhhn+48UpeK/kMe7WbEMZYL+poTQDGZ9bT4uwmF9CiBg8z7vaYwU6QX/3/8+9tUElhQmm2b6q8q
GTInuZoneBKq2dR99tJKsFCXupo67Rmghmc2M6n4+EsofSDZtD4mXS2Q6vhdsyOo8GdkJyHSg1ZS
9J2KFcGrimRZsola7Juq2qdJbwKrwmWbtkJ4NmDWJ6eAP8ZkymHM2CZdGnkycBGjNgfgGztHkrfc
w4E2u/lM3f2udwQXx5Yl2jnS4KJoGQGFGzzb3mO7KGr67ayaffmN1ywgacyXUMzzWw1ah82jHFyP
aCPIUsDyTPxhCJQNwO3iG5JWNGqqtVdoeutNYa1+NxBl4exMwuYoQMGv/Pk2moFjdYkdNBuV8yzs
1UxZxIZCaFWP3ferZJ7CvV/t/b+SUlpTaNYCnRYnBymYwB8vWzQNucbmgatL/lkSZRUwv8sQbVPx
tDrgzhlSudBsIt6HvvHeTAAquzs9IovW+L4LtLKpGWqEb7XlzTOjLzwqsrLhIIaTS6lCd0dcdhME
eTeZGdrZhFNHfMbaUMq/X/SXkFwOuuogJ8CkToe0CWkicpUui71sVvvrNIb5fzMFb6a+vUXTfOy7
EvTA2RnYxqAVXu1jREBAX8PiIrHEjWJ3BBsyLAZIk4KndNnO66kEssXW2p3rFNmCJdNph1pBInAo
DpiEgsb2Bx+uNmcP5TrQr+0T8IgJgv/fQ7tuokmQ+6nubTdZbpNjv/on9tRSn8tfohIHUJqqf5hp
iLrsJFVg1MzVFs5UxG3gl2UwHtNWSaNvTeUMcXRcAtXREIyh2bNElvmZo/WBRlDXQ7d+5L4Y8Rjb
JjquKVAq1qEK4C88H509hLHbAX226tqWAlKdxijPOr+nf6ujf5mZ7bbj48Y4rp/FI4F//if3/Bdy
HzFBjnkIvr7yXFKFqrUJ10YUwIhvyCLmQMo61TOyA3+7ute9DUXonStZinhrIgA6GWm8CT2TsI4F
QgLkmBNSM6Fba+63m//ZKtTVMighaCMze/PM9wSUM8ykdebbhOgvSZki72BfZtXFn4vlKMtarzlz
1RWILijHV8/8cCRikbBu85335AGZiOw7vkSi65IR6SmAlhaiKZdPtHbQVm9CJTR5qm3Ii8kbPAts
29JNl7NflcR/qIABjtmTm/jGh6GW+9DGVfdf/7gnW95Fq9gZ9Ym4g022O3MeRbDj3nDHY0hOP1nV
r0mRH+A0WqAGhY+9nNcgZQR2D0GxpdnbDi2YfaSbtlZysXoKJEjXIqlN1H24cz39ymfNHlYDUCPO
Y5He4qIwU9GwfgbdkQg7BixO6EVRUk7/+nDtXVljxVKmTnQwBrrEb914kiXG0b2SJJSJ6RFXDgzT
7A7hmEV15k7vtx4lueUvQym2NJxOCk9Whexw3bgzfA+RExYNGWpgS02V+JaYwnDTY6YUZ27e8TGR
QiOkswSCHtS4pZwAzin7SZZ/B4Iv1zx5LCWJLHMlbTXpQNXXLnjNtOeZchH+ZTbwKPsr6U/U56H5
MSiTJ/fANFs7JuesDxRMQ3CXWBxoZgNLebcwUDPIDGIc7nEHDdtlzsh8PlFUs95vdzQF8OZJbPa+
Bhxcg8aco1fscKiMrCx6dD8iTEyOj1hh/KK1B3pN/wrPXyZirAIJ3xvrq6Aa/ZBG/UIBWjp2a9jl
FJFSIyHN98DgV+ou2UgkLlFY3kCYCjG6ZoYtmvqUTtemN/mKPEpANUtSi6/ea46qzvmgGTVVZ4dy
TfVIdw6MJSo9tmQY5r5C9q635Eo6oIKLDGnhnF2Eqv9GyUnL+vIEJ5laqOARZb7Q6JjkEGkuuuYl
mbRefV9uCXm4YSk0iQ2yTOUrHOufmng8WjmGcIit9YtHJUgpro4TrbOQP34/P0G0dce+VqE+Ugb1
2kwG3d5I5LEdXCxcr5pe0YClDWmRBMhSXuIUjVSL7ecEMf4iT/HYy4q1izGemNZJRzFvQoTrWJ2O
pB085ttMzrNSnUmnsAt5Jp5wrdQSVLpCfcA9yZuzzmA/LadMo8t7RrzBPUX1gjaKRsJ5HirhItcC
Y3pMJrZ1bCO08FFjasaUhOV6Dq8ZSP8qYKFzpCvg77URpaUZF/kuRJYgt3MfG8Q7QYx5on10E7Cn
E/VYxU/4jz1zojWpEG88NZcnXhNxlG9nqO1BsVhchLFFhYCBrAV8zVbEtGKhPByRyRKwKNZtZL8n
4BRqgk5mqxHDKeobOsbq8E1nuINDCuMVlP+CM5sh1IJTu5kgsmscOs+rHxdTaa6sP9KFMYNRmlci
EubTp1dJZOqxyCABaY4O/7pZ7ZYmasSLSfb2hN6IQn3sYx73ZJ02qCH7XEeh95OmRdWTKeJHqRrG
by9CFkHS1B50yF1Q8J2dH2TJsnjm/K3zNyPR5fwTOWCuKffnxBqCJPC/GmDIVKDZagHQJNZ5AM9+
ibNk1KjIxq+j6E8QqbrJ1cl+/Clf4vh7LDg+pxm5jmv63judFeOyDP0hXCghkHQHpfB7nWChxqcm
TlpaOvHRdYH/4vodsShcf+gAFIFUnWXifGcC2MnIrcoINqP29Ssph4y5IVSJ4WZLZAWX32aej0no
qmo21UxYh5fU4sI74UPps5qa8bCAWhwPzbfGS6gflzDEwoCkDUW/BzIMJ4KuSjZ1VE0vzQT6LAv8
calV7vXpNEH4FdOhS/7mhPJoN4mGoaQ+OMSvexm6W2vbfmPXqrV3R6tTlOkg5O991gTQ9+cDKo13
Fj683rsxB6dIWL53tL9R0Uqs3tAsaPKLpUzQk8rVx6tFLMY0YuRXOx8ndbSZ12qY+J/prlRbY9N2
4GodxA6HoZ7YiAi9krWpceKYHQG3H/UuQgDm4nRBEthwl2VdvPsXuZSGSzqfRxLgZPf6fcM1fOsQ
Z2y/dPebH48INvCnbhOwtbIQlQ3HJ7/8dphYLb2B/1wHxywGr0ZUp2JAQPnWlIGdOVLMNZxy8XAq
B/efejYH9a+Gw3O/30Mk+ZcMViFbiyTwcPDqlR/NvHTbdREWfsmeRtqI/ZaofsEdaEmTqIEsWh07
07lAMUeDABsmmzYfguce0/d4l+xjFDCqvnh2taaUEzABHeQHsoDxKyU3r18RQ4IWpMP8wKA8Tnhm
cgyjZghmDwKtxdEczzXBAosKGr3n80CB8ULy0ysuMVWNRip/KV/Uqew4m4HwsKdbghyzB2ajIrC1
1IUvXryI6+Pi9ewms9D8bkbh42AV5B+8gFilr2spxSjVk+5eZyOkL5fj5vKolHkVD7j/P5HD+8KC
yaURCL3HMa6WqMJ8nKE1leKLbAa/6NZraXABFjKNNRJITGNI8j+XL70vSQrbfKx6e9kEJ25PrImR
QUEQZjrHDMbW6XnTrhCoeU7C59u2GFJg0fFnojr5hfJI2ogEbtghz4D+hWFEQf35xXyNuXEKYJ95
5JYX+JQxN8/vhVuKrHer6x/WH3HYBbWeFW6wnbnPCg5DpXDq/6drjihiw4jqtyEH3L5gFGPdjnAb
mZl7gs9TGJxM0XLT13zfQsvwEjQ1q3KyoI0WRu/+RAxxgaU7pl8Af5xPUqD+iTnzCU2/QvVNcaEv
gE15CtO1mJJg0J3WEl6FKe1ra7MnviG25Byhpu6UQ8Dx1TwyjjB0OZaS9+Po19pF1ExHyzQN06Ow
Lmmy9meg+A6/SnAzYPdgJJdOCDQyd9J469WWEXOZpsOzlH2fHTSOEoq3PHfbkxhaWLHuT/y0dhxG
gqCLd+ZOG3kuPCgv2bnTuXx3q2/vz6NtVJpLLLFCgNCR0Q0skdYXERKaNmyCyDk6A2FA6tHuEUPA
Xs2tLQA334kEdFgWDB50GrrlucY8PZxbR/H0qAWvD/Bh6caUmEu7Fy0z0LJYUMYzvMT3De9MDUtZ
u6ywCTbpkUF1j+cVxXr1ne8iylI17QLHPnCw+ZM5V50A3LwKMF6YUs68jkuVWVSSiIEAttwbecIX
OO912cBkClj/PZuQbJwSvaBrz+QCm3ibAZAGmusgswBwAKjh8z9YyRSz48tADhDgvqJuREnSuZxT
gln2vVBj8fsVq9Uzh8dFbOfTxXe+yX8CCdjkO0VHJCPNW0XntNiYjXYbhxHtL3vZc7QYQz2aCk9R
KOsGJRPs+hQaSxbj8TW3E2pwU3SxHUsNqzVXlFtR2xYkvxGB4C2AWha2Jst1lGSdFHsgPvLg9Dw3
CWooWi/8pawAzosVp2nLV8RQVk/1S4xXuu3wR3S7CSVEo16z8K0nN4oj/WOMflGPQy7PehdtneHC
aZZiQdxHvP2X3RgLbC9BwdZ2/p2A/iGMgUEIsXrlE8abzBJmuzJFtgq+WanwnjjvIwlmy/7du3dT
lZotgTo69N0aYc8urrkFSi6Xi7Whr2JIVz+TLK20CnABsXHuHXJ5uOOBkhX37XP1OwdVQR+3uko1
rV4viy1iOnbT8NGYZpyMz45+Z3lyV1+9S12K6uptdr4gFW+ekb+u0V6tXGYQa0ki4BPfSAGVW9uJ
+JiiGpe31vtKkkLQ03sPTGoAh4pryrEiSJqNkeBAYXYLgAnWNowQJDvrJ0pEI8NzCLduUU7PyFKT
c1tZ9nNdBCeOlckz2RDevXeuc7406pAEKFaB/t2w6sCW07ZpoWjm8HgIquqV4MisUbUC2ypWdeSt
f/GI0NoVfJhUz2stOtBQ34Hqo5cyUnFbbQlFS/pGC47RQC7t2I4gSzmX8DSrs8aOAHGQI2YjNSqT
Of3e1qUziJqt5NRWA4HTMiRCQ1MCiDqRaPCJe3AD050GvXclizE5ytJEpnTmb8Z9+rLHODmH4rZD
Hg5BvtI1zzdPoStNEQPNsuOFMivOU4HHlytD5t37I32dal/4zBRVOKkPvGI3ZprIOZcL3hh3O71b
LfM1AVaVPP37NMB+6qmD57T/0/knNt1gDJHhCfD947Jyk1D5HnhDb6SRzyRg2IOlFpWk4uaTQo3E
q8JLpjLL6mvuGR5OAWcm2dZEvJ9MyfF/lawIfE8MG6l0AgfmlUG8U5ydUIgnPwUqg6zK+HMQnRa0
RJFCR+LoOxA95QtAluOHoSBbCYAY2gNBYWgqXPXpgTuTrnvUO0kuO9Rd2IIrNLcdNN7TTRv7Dudc
FEb6N3Nfw3gh8n62dGXfDARajmJAs6plwUar8cDrs8x136YDpo/xaEXUqyxGUF4ytAWMlQufUE0O
Qi7hsZ5xPTiHDuIzpxLZo4VudEPcxxy2NTXxq38lFLr4KvZ+fGXFs3pUU7AwWlmxXn5V39cmbmnr
TTKnfWLhy8/zxBQ7CehnSUWggHaNh7Dm1/fCVLl62wAWoqxGlsAW5muptej2v+WvINWOWwkUkZdl
fFV5ok0nebM2ei1ZHKqI0WxzAbtB5SGQtjsxVvGiQLcUioB4C4Swq2+uI0oa8wNPJUexnBypWbPZ
BwVV9QxMmiuxrHZONySbcoiwoCYBLHsoGu9zjdGHL66CuvhFwRqCHa5fpLdv6dYtbZaTxW+k6q8c
xOAS6pC13Zp0qhdG9fnuSUYytGKsEOzVHYj8zvvasQZQ/exHwQur7CCwVLyG7a+ibnOMVy5vO93G
OfnCcSk4+gNj7iU8jRHz2RM2W4ioOFiJKFKj7ET5Ci3QQajxmsHAPJPMwxEuVugRV2VQxLKcaG28
tT7CIfGQmFhO9+dJd0be74La12WNmHBfblhc55kKGGrvQKI4WEAwRdUXt4kGJ/jB9fJ+RjKVzsvG
+jmFP2mdLGvsDBYmxYuZD+JOT/gPCtODsYd1OpBSOnJNmwY7GoW0fXgPtqhV1NfEY0HwOSHAZhFD
WoD2ZtNwerYfwWHPZ6keBPN83rlRwzkIuFJnWYxXDWpzIOvcX0l+FlvRd6bpiDSlZz7LHs1UOdW6
TIOlv9iDcSyMwqUvB0kyVlZejabrgP+yICIMj2c8qvnvuHkYFMH9BmhZx2P5d1mnbg0O8wv3yZmS
EcWbPbVwSrSQ8WhG2XElNjodnxJK/G0APkko2V6M1VNZqG7aSw76b+f36hNTtMBbHOYfieatURX4
Ms6um4RHZXhVb/pungnG9jUP90i+OSKz+JggvOmYcgTThcM3dEBduFpS8OgyJ7cSlPsRlbCw0T+Q
CQeu+KCeNwFBoO2M0cL2MdpUbsF/J6xDomELrUVMh15Kj34OKzP5C6iBofhzhslWUkpu2Jlxf0A3
z+znb1/lCUPsdJD/zNqXb6svSq6A7o5b7yIO7pFfTK7Y+roPjPKP4ZSjYgiBd5txdxC3zRGLGLuv
nXa1n524c0wPsUV7OQcRaI5ud541LwX6AN2L0HZW6qhE0m7wZQToG0EqnVB288Zpe/m3yLlZQKlJ
jr6JPxI15+V04gHCW15WLCTjOLgGGAdjNx/lploFZcDqzOsGGVT4y2idNxjWczutj/wiZsycgopD
hd/4T58B3KZ3yO7Lew2fXDTrLHEt99DBXeKmoGmxWR4xkPliaTWYPYD3p6riOBjCm6afp6Lp83os
X1+doXjvvctvKplk0FZU07GTt/38IEJZGAovRQtJhZfLAs6UGpd7j9PCo6LRIdQQUBZhjylMpiNJ
iqkYeyfKjpfHttCwTSBa4Yzt3qRXoiP0ORCblf/te/2Gr1P28Yg023HC//AjAbIIwRnduUGOVJGS
UeNU5GOBTCnzPwFkqPSJL+v3epDUD81lpJVqrPDsKi/3dsqBZNRASZT9Smz9gJZRGGPT+/zJ6u6i
xr4leLTInij+yGvSS7HiGYBjKXbRcRVVwb4e6AHDvtoOOpYQHRsuSChp9wJd0D6dIBDraC6b5zea
Fp/1OLQDMiPa5wectnXfhy/pwG7enBu8/p2WJZ02cGaTENxIGyJ7W0pYpgpy9gkoe1527c5ZYU05
6bvAUvqRD6uQJXnwGW1vPrkvzYsibpmkoLIVLQMcSJ7gyBwaw0SxhvG+1xLvva4cGCn5iX3nUrhH
F7xdK1Q3dj6G+VVt7zJ+BbJo+h7q1jwIQfOC2jWStMl5jNyCLUiTRThWo0gszEUZig8ewXexPJ2G
yisynQktOGOVq8FYAxkRwr0rs2lKvtVW0llOtuJt8+jReF/nwen8biH5ZGjGBKN+6Tr/GLC/9BW9
TtVUTQiVlqCrbtEByXmx795oUYAxws3uzS4cAtwpFFBjxJnOJwltAjdWB5z/u3kJDEzU321n6K/a
/eJGCNwPpDTvO0ZeawrZm5BastXa+IQBfkrQjbdjha6NPmZ5Xirpfkewp1xDKwGlvQGj6AL7h5wj
KsGbH161567EI/ks7y7lcjhcT6LnPKVJF4UnhIEcf0fONtz2SwQS2UUv4W9RtACmM4TMOxQYye7i
JzCCgPw38laDGMmGSMRWvyfZbSi1cXf86Jau0kvONA7nAlzxE2oqJml9HsCU2Syy7LtTKw9OnmUE
MtN51sfEVBsThpYhBPYHwzwadA71HndebVXdUip/aDCB5fx1XZUJ76bMoHeW3iYQMv2urHdW4dl1
pCsXC0iE6kKNZfeWGjJN+RcqPLomQKde9aHDokyB+Q6lVw4CNAFgK/iy1vX8VjXjOIEg45gCXxQ4
kqXJCLjk467/OsLCuBX2Z/hJ9BsRTDL77Uf3FQgbpRr4Y/JmEqHG7vXnf6dDPreplHtAVUjpJOKI
K/4u54ZT2JJ8f7x2zVHIH07PLLIxxVuDIltA2S+zVQAW5obpoJt5casUK5mcSkpQw0x3RJJwBmFc
DrSb7BxX6GwAXY1/lQCQhqi8/5oCoEWoCe2dvO2S4unkqGvrwNjGMZCthpr5DUqR0V4J80GPL5rV
/4JCTW0azDAEXGtqM5qKVCzDTR/2zNkkgx55ynMH3l+q3mC00KvQ2hxHn5ZIoZ+z9O65Thmp33ec
iM5HlBq0UQg1HZRK8AjEIy/KAaYJU3ER+1y9NCFufzR0pwzsSVzlR56Y7EgLFOl0WgjmwSvNBN+6
/suWf5pKcdlNaVzjd0FtEf+KBRj48Y4sNxXFT8qkJdFy6J4StHPLGT0Y8uBXOVb6AnVoR/msGkVO
Zuao2V67P6fqeM3mGixjWItZYCGyZi0z2dp2x98b+kZkYKl91RV/EEsIF81PdAEvkatsMkZqEHZu
j9kWelXR6i+0u7nfIR76umyNlxWEEGpqkc8rQI2ScjBGl+hcDSo9aqGYJVYGQlqKVaYhoYOV722W
530HMHMp26zW9sq8E4RFavZlfUAdjMN5z7Brzi5aVKlpcCVRrr0obQjrNfiBuppO67rnaoOJqmkQ
H8z/0NglVrunobUX9WIz6mGChb03uNxZg9moikYrRCbquLT7ufs/ZfPCvenczYr00mNWjb5hatDC
/UVWoH8qh5U4j6snsswEfjuAvQdamCgdRLPblJIjJmiNoL0B/8K/2oSUUuZssG+TGzNzPUu47Up2
gZQQsr5JCePU9FUy4jrO2t73qlsIB7/Helr/nsWotNIozZu88ulolsxw9FS+xwBJJuOduhzyUHXd
rFFy7Vby/wpHmaoU42qecoDkViCx9q//RHq53G8OMAwmyKSgG4o6DUqrmaW5VP6FuyWTtmNBup1m
GEQ6uG/MPDNl1ZWdUfDz/ewcrABb+r+zWSgOB3GFLPtrrJ1TLduiwC7zZZOWFiXJEaGKudC/Sw06
+/D67Ix1VlcPUX6RJfYzNgZGPygfs6/7njmVuX22veKmifaJKHE2yRHmA8naQXtn5FpLcSAd0Aw3
jiNcFZ65zo0dGKOApIHbylOmjJq49iM3aeHVsSGBlhcGb/9l9LmIZ8mA6Ah9/RnNaQdzOI998VgN
CNAMZT6HsloBuMTWQSJNr8OUSTp9CZOWWLiXuYTnbkplNq+CJrHhPBU5mLXZxzxFNf0BPeX9+72H
m6RG8yRgYQSKEP7MZM9PC6wGF1MZV0CIl4xdTDKPw6AW8pHpoRLnMD5Uy9PtR+HBIodrq9DfVJKe
LZHx5xcKCuKzDNkvtb6K7DomQWNrR8qdh5DlJ5tKiF8tG7+FhAo+AIk8R3UOXT2nfZI4p63H3eKF
mz+wnSJRdqnNrJ9Fnrr32trCYxrDa9X/f01OgCNI
`protect end_protected
